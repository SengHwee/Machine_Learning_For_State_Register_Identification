
module siphash(clk, reset_n, cs, we, \addr[0] , \addr[1] , \addr[2] , \addr[3] , \addr[4] , \addr[5] , \addr[6] , \addr[7] , \write_data[0] , \write_data[1] , \write_data[2] , \write_data[3] , \write_data[4] , \write_data[5] , \write_data[6] , \write_data[7] , \write_data[8] , \write_data[9] , \write_data[10] , \write_data[11] , \write_data[12] , \write_data[13] , \write_data[14] , \write_data[15] , \write_data[16] , \write_data[17] , \write_data[18] , \write_data[19] , \write_data[20] , \write_data[21] , \write_data[22] , \write_data[23] , \write_data[24] , \write_data[25] , \write_data[26] , \write_data[27] , \write_data[28] , \write_data[29] , \write_data[30] , \write_data[31] , \read_data[0] , \read_data[1] , \read_data[2] , \read_data[3] , \read_data[4] , \read_data[5] , \read_data[6] , \read_data[7] , \read_data[8] , \read_data[9] , \read_data[10] , \read_data[11] , \read_data[12] , \read_data[13] , \read_data[14] , \read_data[15] , \read_data[16] , \read_data[17] , \read_data[18] , \read_data[19] , \read_data[20] , \read_data[21] , \read_data[22] , \read_data[23] , \read_data[24] , \read_data[25] , \read_data[26] , \read_data[27] , \read_data[28] , \read_data[29] , \read_data[30] , \read_data[31] );
  wire _abc_19068_n1000_1;
  wire _abc_19068_n1001;
  wire _abc_19068_n1002_1;
  wire _abc_19068_n1003_1;
  wire _abc_19068_n1005_1;
  wire _abc_19068_n1006_1;
  wire _abc_19068_n1007;
  wire _abc_19068_n1008_1;
  wire _abc_19068_n1009_1;
  wire _abc_19068_n1010;
  wire _abc_19068_n1011_1;
  wire _abc_19068_n1012_1;
  wire _abc_19068_n1013;
  wire _abc_19068_n1014_1;
  wire _abc_19068_n1015_1;
  wire _abc_19068_n1016;
  wire _abc_19068_n1017_1;
  wire _abc_19068_n1018_1;
  wire _abc_19068_n1019;
  wire _abc_19068_n1020_1;
  wire _abc_19068_n1021_1;
  wire _abc_19068_n1022;
  wire _abc_19068_n1023_1;
  wire _abc_19068_n1024_1;
  wire _abc_19068_n1025;
  wire _abc_19068_n1026_1;
  wire _abc_19068_n1028;
  wire _abc_19068_n1029_1;
  wire _abc_19068_n1030_1;
  wire _abc_19068_n1031;
  wire _abc_19068_n1032_1;
  wire _abc_19068_n1033_1;
  wire _abc_19068_n1034;
  wire _abc_19068_n1035_1;
  wire _abc_19068_n1036_1;
  wire _abc_19068_n1037;
  wire _abc_19068_n1038_1;
  wire _abc_19068_n1039_1;
  wire _abc_19068_n1040;
  wire _abc_19068_n1041_1;
  wire _abc_19068_n1042_1;
  wire _abc_19068_n1043;
  wire _abc_19068_n1044_1;
  wire _abc_19068_n1045_1;
  wire _abc_19068_n1046;
  wire _abc_19068_n1047_1;
  wire _abc_19068_n1048_1;
  wire _abc_19068_n1049;
  wire _abc_19068_n1050_1;
  wire _abc_19068_n1052;
  wire _abc_19068_n1053_1;
  wire _abc_19068_n1054_1;
  wire _abc_19068_n1055;
  wire _abc_19068_n1056_1;
  wire _abc_19068_n1057_1;
  wire _abc_19068_n1058;
  wire _abc_19068_n1059_1;
  wire _abc_19068_n1060_1;
  wire _abc_19068_n1061;
  wire _abc_19068_n1062_1;
  wire _abc_19068_n1063_1;
  wire _abc_19068_n1064;
  wire _abc_19068_n1065_1;
  wire _abc_19068_n1066_1;
  wire _abc_19068_n1067;
  wire _abc_19068_n1068_1;
  wire _abc_19068_n1069_1;
  wire _abc_19068_n1070;
  wire _abc_19068_n1071_1;
  wire _abc_19068_n1072_1;
  wire _abc_19068_n1073;
  wire _abc_19068_n1075_1;
  wire _abc_19068_n1076;
  wire _abc_19068_n1077_1;
  wire _abc_19068_n1078_1;
  wire _abc_19068_n1079;
  wire _abc_19068_n1080_1;
  wire _abc_19068_n1081_1;
  wire _abc_19068_n1082;
  wire _abc_19068_n1083_1;
  wire _abc_19068_n1084_1;
  wire _abc_19068_n1085;
  wire _abc_19068_n1086_1;
  wire _abc_19068_n1087_1;
  wire _abc_19068_n1088;
  wire _abc_19068_n1089_1;
  wire _abc_19068_n1090_1;
  wire _abc_19068_n1091;
  wire _abc_19068_n1092_1;
  wire _abc_19068_n1093_1;
  wire _abc_19068_n1094;
  wire _abc_19068_n1095_1;
  wire _abc_19068_n1096_1;
  wire _abc_19068_n1098_1;
  wire _abc_19068_n1099_1;
  wire _abc_19068_n1100;
  wire _abc_19068_n1101_1;
  wire _abc_19068_n1102_1;
  wire _abc_19068_n1103;
  wire _abc_19068_n1104_1;
  wire _abc_19068_n1105_1;
  wire _abc_19068_n1106;
  wire _abc_19068_n1107_1;
  wire _abc_19068_n1108_1;
  wire _abc_19068_n1109;
  wire _abc_19068_n1110_1;
  wire _abc_19068_n1111_1;
  wire _abc_19068_n1112;
  wire _abc_19068_n1113_1;
  wire _abc_19068_n1114_1;
  wire _abc_19068_n1115;
  wire _abc_19068_n1116_1;
  wire _abc_19068_n1117_1;
  wire _abc_19068_n1118;
  wire _abc_19068_n1120_1;
  wire _abc_19068_n1121;
  wire _abc_19068_n1122_1;
  wire _abc_19068_n1123_1;
  wire _abc_19068_n1124;
  wire _abc_19068_n1125_1;
  wire _abc_19068_n1126_1;
  wire _abc_19068_n1127;
  wire _abc_19068_n1128_1;
  wire _abc_19068_n1129_1;
  wire _abc_19068_n1130;
  wire _abc_19068_n1131_1;
  wire _abc_19068_n1132;
  wire _abc_19068_n1133;
  wire _abc_19068_n1134_1;
  wire _abc_19068_n1135;
  wire _abc_19068_n1136_1;
  wire _abc_19068_n1137_1;
  wire _abc_19068_n1138;
  wire _abc_19068_n1140_1;
  wire _abc_19068_n1141;
  wire _abc_19068_n1142_1;
  wire _abc_19068_n1143;
  wire _abc_19068_n1144_1;
  wire _abc_19068_n1145;
  wire _abc_19068_n1146_1;
  wire _abc_19068_n1147_1;
  wire _abc_19068_n1148;
  wire _abc_19068_n1149_1;
  wire _abc_19068_n1150_1;
  wire _abc_19068_n1151;
  wire _abc_19068_n1152_1;
  wire _abc_19068_n1153_1;
  wire _abc_19068_n1154;
  wire _abc_19068_n1155_1;
  wire _abc_19068_n1156_1;
  wire _abc_19068_n1157;
  wire _abc_19068_n1158_1;
  wire _abc_19068_n1160;
  wire _abc_19068_n1161_1;
  wire _abc_19068_n1162_1;
  wire _abc_19068_n1163;
  wire _abc_19068_n1164_1;
  wire _abc_19068_n1165_1;
  wire _abc_19068_n1166;
  wire _abc_19068_n1167_1;
  wire _abc_19068_n1168_1;
  wire _abc_19068_n1169;
  wire _abc_19068_n1170_1;
  wire _abc_19068_n1171_1;
  wire _abc_19068_n1172;
  wire _abc_19068_n1173_1;
  wire _abc_19068_n1174_1;
  wire _abc_19068_n1175;
  wire _abc_19068_n1176_1;
  wire _abc_19068_n1177_1;
  wire _abc_19068_n1178;
  wire _abc_19068_n1180_1;
  wire _abc_19068_n1181;
  wire _abc_19068_n1182_1;
  wire _abc_19068_n1183_1;
  wire _abc_19068_n1184;
  wire _abc_19068_n1185_1;
  wire _abc_19068_n1186_1;
  wire _abc_19068_n1187;
  wire _abc_19068_n1188_1;
  wire _abc_19068_n1189_1;
  wire _abc_19068_n1190;
  wire _abc_19068_n1191_1;
  wire _abc_19068_n1192_1;
  wire _abc_19068_n1193;
  wire _abc_19068_n1194_1;
  wire _abc_19068_n1195_1;
  wire _abc_19068_n1196;
  wire _abc_19068_n1197_1;
  wire _abc_19068_n1198_1;
  wire _abc_19068_n1199;
  wire _abc_19068_n1200_1;
  wire _abc_19068_n1202;
  wire _abc_19068_n1203_1;
  wire _abc_19068_n1204_1;
  wire _abc_19068_n1205;
  wire _abc_19068_n1206_1;
  wire _abc_19068_n1207_1;
  wire _abc_19068_n1208;
  wire _abc_19068_n1209_1;
  wire _abc_19068_n1210_1;
  wire _abc_19068_n1211;
  wire _abc_19068_n1212_1;
  wire _abc_19068_n1213_1;
  wire _abc_19068_n1214;
  wire _abc_19068_n1215_1;
  wire _abc_19068_n1216_1;
  wire _abc_19068_n1217;
  wire _abc_19068_n1218_1;
  wire _abc_19068_n1219_1;
  wire _abc_19068_n1220;
  wire _abc_19068_n1221_1;
  wire _abc_19068_n1222_1;
  wire _abc_19068_n1224_1;
  wire _abc_19068_n1225_1;
  wire _abc_19068_n1226;
  wire _abc_19068_n1227_1;
  wire _abc_19068_n1228_1;
  wire _abc_19068_n1229;
  wire _abc_19068_n1230_1;
  wire _abc_19068_n1231;
  wire _abc_19068_n1232;
  wire _abc_19068_n1233_1;
  wire _abc_19068_n1234;
  wire _abc_19068_n1235_1;
  wire _abc_19068_n1236;
  wire _abc_19068_n1237_1;
  wire _abc_19068_n1238;
  wire _abc_19068_n1239_1;
  wire _abc_19068_n1240;
  wire _abc_19068_n1241_1;
  wire _abc_19068_n1242;
  wire _abc_19068_n1243_1;
  wire _abc_19068_n1245_1;
  wire _abc_19068_n1246;
  wire _abc_19068_n1247_1;
  wire _abc_19068_n1248;
  wire _abc_19068_n1249_1;
  wire _abc_19068_n1250;
  wire _abc_19068_n1251_1;
  wire _abc_19068_n1252;
  wire _abc_19068_n1253_1;
  wire _abc_19068_n1254;
  wire _abc_19068_n1255_1;
  wire _abc_19068_n1256;
  wire _abc_19068_n1257_1;
  wire _abc_19068_n1258;
  wire _abc_19068_n1259_1;
  wire _abc_19068_n1260;
  wire _abc_19068_n1261_1;
  wire _abc_19068_n1262;
  wire _abc_19068_n1263_1;
  wire _abc_19068_n1264;
  wire _abc_19068_n1265_1;
  wire _abc_19068_n1267_1;
  wire _abc_19068_n1268;
  wire _abc_19068_n1269_1;
  wire _abc_19068_n1270;
  wire _abc_19068_n1271_1;
  wire _abc_19068_n1272;
  wire _abc_19068_n1273_1;
  wire _abc_19068_n1274;
  wire _abc_19068_n1275_1;
  wire _abc_19068_n1276;
  wire _abc_19068_n1277_1;
  wire _abc_19068_n1278;
  wire _abc_19068_n1279_1;
  wire _abc_19068_n1280;
  wire _abc_19068_n1281_1;
  wire _abc_19068_n1282;
  wire _abc_19068_n1283_1;
  wire _abc_19068_n1284;
  wire _abc_19068_n1285_1;
  wire _abc_19068_n1287_1;
  wire _abc_19068_n1288;
  wire _abc_19068_n1289_1;
  wire _abc_19068_n1290;
  wire _abc_19068_n1291_1;
  wire _abc_19068_n1292;
  wire _abc_19068_n1293_1;
  wire _abc_19068_n1294;
  wire _abc_19068_n1295_1;
  wire _abc_19068_n1296;
  wire _abc_19068_n1297;
  wire _abc_19068_n1298_1;
  wire _abc_19068_n1299;
  wire _abc_19068_n1300_1;
  wire _abc_19068_n1301;
  wire _abc_19068_n1302_1;
  wire _abc_19068_n1303;
  wire _abc_19068_n1304_1;
  wire _abc_19068_n1305;
  wire _abc_19068_n1306_1;
  wire _abc_19068_n1308_1;
  wire _abc_19068_n1309;
  wire _abc_19068_n1310_1;
  wire _abc_19068_n1311;
  wire _abc_19068_n1312_1;
  wire _abc_19068_n1313;
  wire _abc_19068_n1314_1;
  wire _abc_19068_n1315;
  wire _abc_19068_n1316_1;
  wire _abc_19068_n1317;
  wire _abc_19068_n1318_1;
  wire _abc_19068_n1319;
  wire _abc_19068_n1320_1;
  wire _abc_19068_n1321;
  wire _abc_19068_n1322_1;
  wire _abc_19068_n1323;
  wire _abc_19068_n1324_1;
  wire _abc_19068_n1325;
  wire _abc_19068_n1326_1;
  wire _abc_19068_n1327;
  wire _abc_19068_n1329;
  wire _abc_19068_n1330_1;
  wire _abc_19068_n1331;
  wire _abc_19068_n1332_1;
  wire _abc_19068_n1333;
  wire _abc_19068_n1334_1;
  wire _abc_19068_n1335;
  wire _abc_19068_n1336_1;
  wire _abc_19068_n1337;
  wire _abc_19068_n1338_1;
  wire _abc_19068_n1339;
  wire _abc_19068_n1340_1;
  wire _abc_19068_n1341;
  wire _abc_19068_n1342_1;
  wire _abc_19068_n1343;
  wire _abc_19068_n1344_1;
  wire _abc_19068_n1345;
  wire _abc_19068_n1346_1;
  wire _abc_19068_n1347;
  wire _abc_19068_n1348_1;
  wire _abc_19068_n1350_1;
  wire _abc_19068_n1351;
  wire _abc_19068_n1352_1;
  wire _abc_19068_n1353;
  wire _abc_19068_n1354_1;
  wire _abc_19068_n1355;
  wire _abc_19068_n1356_1;
  wire _abc_19068_n1357;
  wire _abc_19068_n1358_1;
  wire _abc_19068_n1359;
  wire _abc_19068_n1360_1;
  wire _abc_19068_n1361;
  wire _abc_19068_n1362;
  wire _abc_19068_n1363_1;
  wire _abc_19068_n1364;
  wire _abc_19068_n1365_1;
  wire _abc_19068_n1366;
  wire _abc_19068_n1367_1;
  wire _abc_19068_n1368;
  wire _abc_19068_n1369_1;
  wire _abc_19068_n1371_1;
  wire _abc_19068_n1372;
  wire _abc_19068_n1373_1;
  wire _abc_19068_n1374;
  wire _abc_19068_n1375_1;
  wire _abc_19068_n1376;
  wire _abc_19068_n1377_1;
  wire _abc_19068_n1378;
  wire _abc_19068_n1379_1;
  wire _abc_19068_n1380;
  wire _abc_19068_n1381_1;
  wire _abc_19068_n1382;
  wire _abc_19068_n1383_1;
  wire _abc_19068_n1384;
  wire _abc_19068_n1385_1;
  wire _abc_19068_n1386;
  wire _abc_19068_n1387_1;
  wire _abc_19068_n1388;
  wire _abc_19068_n1389_1;
  wire _abc_19068_n1390;
  wire _abc_19068_n1392;
  wire _abc_19068_n1393_1;
  wire _abc_19068_n1394;
  wire _abc_19068_n1395_1;
  wire _abc_19068_n1396;
  wire _abc_19068_n1397_1;
  wire _abc_19068_n1398;
  wire _abc_19068_n1399_1;
  wire _abc_19068_n1400;
  wire _abc_19068_n1401_1;
  wire _abc_19068_n1402;
  wire _abc_19068_n1403_1;
  wire _abc_19068_n1404;
  wire _abc_19068_n1405_1;
  wire _abc_19068_n1406;
  wire _abc_19068_n1407_1;
  wire _abc_19068_n1408;
  wire _abc_19068_n1409_1;
  wire _abc_19068_n1410;
  wire _abc_19068_n1411_1;
  wire _abc_19068_n1413_1;
  wire _abc_19068_n1414;
  wire _abc_19068_n1415_1;
  wire _abc_19068_n1416;
  wire _abc_19068_n1417_1;
  wire _abc_19068_n1418;
  wire _abc_19068_n1419_1;
  wire _abc_19068_n1420;
  wire _abc_19068_n1421_1;
  wire _abc_19068_n1422;
  wire _abc_19068_n1423_1;
  wire _abc_19068_n1424;
  wire _abc_19068_n1425_1;
  wire _abc_19068_n1426;
  wire _abc_19068_n1427;
  wire _abc_19068_n1428_1;
  wire _abc_19068_n1429;
  wire _abc_19068_n1430_1;
  wire _abc_19068_n1431;
  wire _abc_19068_n1432_1;
  wire _abc_19068_n1434_1;
  wire _abc_19068_n1435;
  wire _abc_19068_n1436_1;
  wire _abc_19068_n1437;
  wire _abc_19068_n1438_1;
  wire _abc_19068_n1439;
  wire _abc_19068_n1440_1;
  wire _abc_19068_n1441;
  wire _abc_19068_n1442_1;
  wire _abc_19068_n1443;
  wire _abc_19068_n1444_1;
  wire _abc_19068_n1445;
  wire _abc_19068_n1446_1;
  wire _abc_19068_n1447;
  wire _abc_19068_n1448_1;
  wire _abc_19068_n1449;
  wire _abc_19068_n1450_1;
  wire _abc_19068_n1451;
  wire _abc_19068_n1452_1;
  wire _abc_19068_n1454_1;
  wire _abc_19068_n1455;
  wire _abc_19068_n1456_1;
  wire _abc_19068_n1457;
  wire _abc_19068_n1458_1;
  wire _abc_19068_n1459;
  wire _abc_19068_n1460_1;
  wire _abc_19068_n1461;
  wire _abc_19068_n1462_1;
  wire _abc_19068_n1463;
  wire _abc_19068_n1464_1;
  wire _abc_19068_n1465;
  wire _abc_19068_n1466_1;
  wire _abc_19068_n1467;
  wire _abc_19068_n1468_1;
  wire _abc_19068_n1469;
  wire _abc_19068_n1470_1;
  wire _abc_19068_n1471;
  wire _abc_19068_n1472_1;
  wire _abc_19068_n1473;
  wire _abc_19068_n1475;
  wire _abc_19068_n1476_1;
  wire _abc_19068_n1477;
  wire _abc_19068_n1478_1;
  wire _abc_19068_n1479;
  wire _abc_19068_n1480_1;
  wire _abc_19068_n1481;
  wire _abc_19068_n1482_1;
  wire _abc_19068_n1483;
  wire _abc_19068_n1484_1;
  wire _abc_19068_n1485;
  wire _abc_19068_n1486_1;
  wire _abc_19068_n1487;
  wire _abc_19068_n1488_1;
  wire _abc_19068_n1489;
  wire _abc_19068_n1490_1;
  wire _abc_19068_n1491;
  wire _abc_19068_n1492;
  wire _abc_19068_n1493_1;
  wire _abc_19068_n1494;
  wire _abc_19068_n1496;
  wire _abc_19068_n1497_1;
  wire _abc_19068_n1498;
  wire _abc_19068_n1499_1;
  wire _abc_19068_n1500;
  wire _abc_19068_n1501_1;
  wire _abc_19068_n1502;
  wire _abc_19068_n1503_1;
  wire _abc_19068_n1504;
  wire _abc_19068_n1505_1;
  wire _abc_19068_n1506;
  wire _abc_19068_n1507_1;
  wire _abc_19068_n1508;
  wire _abc_19068_n1509_1;
  wire _abc_19068_n1510;
  wire _abc_19068_n1511_1;
  wire _abc_19068_n1512;
  wire _abc_19068_n1513_1;
  wire _abc_19068_n1514;
  wire _abc_19068_n1516;
  wire _abc_19068_n1517_1;
  wire _abc_19068_n1518;
  wire _abc_19068_n1519_1;
  wire _abc_19068_n1520;
  wire _abc_19068_n1521_1;
  wire _abc_19068_n1522;
  wire _abc_19068_n1523_1;
  wire _abc_19068_n1524;
  wire _abc_19068_n1525_1;
  wire _abc_19068_n1526;
  wire _abc_19068_n1527_1;
  wire _abc_19068_n1528;
  wire _abc_19068_n1529_1;
  wire _abc_19068_n1530;
  wire _abc_19068_n1531_1;
  wire _abc_19068_n1532;
  wire _abc_19068_n1533_1;
  wire _abc_19068_n1534;
  wire _abc_19068_n1536;
  wire _abc_19068_n1537_1;
  wire _abc_19068_n1538;
  wire _abc_19068_n1539_1;
  wire _abc_19068_n1540;
  wire _abc_19068_n1541_1;
  wire _abc_19068_n1542;
  wire _abc_19068_n1543_1;
  wire _abc_19068_n1544;
  wire _abc_19068_n1545_1;
  wire _abc_19068_n1546;
  wire _abc_19068_n1547_1;
  wire _abc_19068_n1548;
  wire _abc_19068_n1549_1;
  wire _abc_19068_n1550;
  wire _abc_19068_n1551_1;
  wire _abc_19068_n1552;
  wire _abc_19068_n1553_1;
  wire _abc_19068_n1554;
  wire _abc_19068_n1555_1;
  wire _abc_19068_n1557;
  wire _abc_19068_n1558_1;
  wire _abc_19068_n1559;
  wire _abc_19068_n1560;
  wire _abc_19068_n1561_1;
  wire _abc_19068_n1562;
  wire _abc_19068_n1563_1;
  wire _abc_19068_n1564;
  wire _abc_19068_n1565_1;
  wire _abc_19068_n1566;
  wire _abc_19068_n1567_1;
  wire _abc_19068_n1568;
  wire _abc_19068_n1569_1;
  wire _abc_19068_n1570;
  wire _abc_19068_n1571_1;
  wire _abc_19068_n1572;
  wire _abc_19068_n1573_1;
  wire _abc_19068_n1574;
  wire _abc_19068_n1575;
  wire _abc_19068_n1576;
  wire _abc_19068_n1578;
  wire _abc_19068_n1579;
  wire _abc_19068_n1580_1;
  wire _abc_19068_n1581;
  wire _abc_19068_n1582;
  wire _abc_19068_n1583_1;
  wire _abc_19068_n1584;
  wire _abc_19068_n1585;
  wire _abc_19068_n1586;
  wire _abc_19068_n1587_1;
  wire _abc_19068_n1588;
  wire _abc_19068_n1589_1;
  wire _abc_19068_n1590;
  wire _abc_19068_n1591;
  wire _abc_19068_n1592;
  wire _abc_19068_n1593;
  wire _abc_19068_n1594;
  wire _abc_19068_n1595;
  wire _abc_19068_n1596;
  wire _abc_19068_n1597;
  wire _abc_19068_n1599;
  wire _abc_19068_n1600;
  wire _abc_19068_n1601;
  wire _abc_19068_n1602;
  wire _abc_19068_n1603;
  wire _abc_19068_n1604;
  wire _abc_19068_n1605;
  wire _abc_19068_n1606;
  wire _abc_19068_n1607;
  wire _abc_19068_n1608;
  wire _abc_19068_n1609;
  wire _abc_19068_n1610;
  wire _abc_19068_n1611;
  wire _abc_19068_n1612;
  wire _abc_19068_n1613;
  wire _abc_19068_n1614;
  wire _abc_19068_n1615;
  wire _abc_19068_n1616;
  wire _abc_19068_n1617;
  wire _abc_19068_n1619;
  wire _abc_19068_n1620;
  wire _abc_19068_n1620_bF_buf0;
  wire _abc_19068_n1620_bF_buf1;
  wire _abc_19068_n1620_bF_buf10;
  wire _abc_19068_n1620_bF_buf2;
  wire _abc_19068_n1620_bF_buf3;
  wire _abc_19068_n1620_bF_buf4;
  wire _abc_19068_n1620_bF_buf5;
  wire _abc_19068_n1620_bF_buf6;
  wire _abc_19068_n1620_bF_buf7;
  wire _abc_19068_n1620_bF_buf8;
  wire _abc_19068_n1620_bF_buf9;
  wire _abc_19068_n1621;
  wire _abc_19068_n1622;
  wire _abc_19068_n1624;
  wire _abc_19068_n1625;
  wire _abc_19068_n1626;
  wire _abc_19068_n1628;
  wire _abc_19068_n1629;
  wire _abc_19068_n1630;
  wire _abc_19068_n1632;
  wire _abc_19068_n1633;
  wire _abc_19068_n1634;
  wire _abc_19068_n1636;
  wire _abc_19068_n1637;
  wire _abc_19068_n1638;
  wire _abc_19068_n1640;
  wire _abc_19068_n1641;
  wire _abc_19068_n1642;
  wire _abc_19068_n1644;
  wire _abc_19068_n1645;
  wire _abc_19068_n1646;
  wire _abc_19068_n1648;
  wire _abc_19068_n1649;
  wire _abc_19068_n1650;
  wire _abc_19068_n1652;
  wire _abc_19068_n1653;
  wire _abc_19068_n1654;
  wire _abc_19068_n1656;
  wire _abc_19068_n1657;
  wire _abc_19068_n1658;
  wire _abc_19068_n1660;
  wire _abc_19068_n1661;
  wire _abc_19068_n1662;
  wire _abc_19068_n1664;
  wire _abc_19068_n1665;
  wire _abc_19068_n1666;
  wire _abc_19068_n1668;
  wire _abc_19068_n1669;
  wire _abc_19068_n1670;
  wire _abc_19068_n1672;
  wire _abc_19068_n1673;
  wire _abc_19068_n1674;
  wire _abc_19068_n1676;
  wire _abc_19068_n1677;
  wire _abc_19068_n1678;
  wire _abc_19068_n1680;
  wire _abc_19068_n1681;
  wire _abc_19068_n1682;
  wire _abc_19068_n1684;
  wire _abc_19068_n1685;
  wire _abc_19068_n1686;
  wire _abc_19068_n1688;
  wire _abc_19068_n1689;
  wire _abc_19068_n1690;
  wire _abc_19068_n1692;
  wire _abc_19068_n1693;
  wire _abc_19068_n1694;
  wire _abc_19068_n1696;
  wire _abc_19068_n1697;
  wire _abc_19068_n1698;
  wire _abc_19068_n1700;
  wire _abc_19068_n1701;
  wire _abc_19068_n1702;
  wire _abc_19068_n1704;
  wire _abc_19068_n1705;
  wire _abc_19068_n1706;
  wire _abc_19068_n1708;
  wire _abc_19068_n1709;
  wire _abc_19068_n1710;
  wire _abc_19068_n1712;
  wire _abc_19068_n1713;
  wire _abc_19068_n1714;
  wire _abc_19068_n1716;
  wire _abc_19068_n1717;
  wire _abc_19068_n1718;
  wire _abc_19068_n1720;
  wire _abc_19068_n1721;
  wire _abc_19068_n1722;
  wire _abc_19068_n1724;
  wire _abc_19068_n1725;
  wire _abc_19068_n1726;
  wire _abc_19068_n1728;
  wire _abc_19068_n1729;
  wire _abc_19068_n1730;
  wire _abc_19068_n1732;
  wire _abc_19068_n1733;
  wire _abc_19068_n1734;
  wire _abc_19068_n1736;
  wire _abc_19068_n1737;
  wire _abc_19068_n1738;
  wire _abc_19068_n1740;
  wire _abc_19068_n1741;
  wire _abc_19068_n1742;
  wire _abc_19068_n1744;
  wire _abc_19068_n1745;
  wire _abc_19068_n1746;
  wire _abc_19068_n1748;
  wire _abc_19068_n1749;
  wire _abc_19068_n1750;
  wire _abc_19068_n1752;
  wire _abc_19068_n1753;
  wire _abc_19068_n1754;
  wire _abc_19068_n1756;
  wire _abc_19068_n1757;
  wire _abc_19068_n1758;
  wire _abc_19068_n1760;
  wire _abc_19068_n1761;
  wire _abc_19068_n1762;
  wire _abc_19068_n1764;
  wire _abc_19068_n1765;
  wire _abc_19068_n1766;
  wire _abc_19068_n1768;
  wire _abc_19068_n1769;
  wire _abc_19068_n1770;
  wire _abc_19068_n1772;
  wire _abc_19068_n1773;
  wire _abc_19068_n1774;
  wire _abc_19068_n1776;
  wire _abc_19068_n1777;
  wire _abc_19068_n1778;
  wire _abc_19068_n1780;
  wire _abc_19068_n1781;
  wire _abc_19068_n1782;
  wire _abc_19068_n1784;
  wire _abc_19068_n1785;
  wire _abc_19068_n1786;
  wire _abc_19068_n1788;
  wire _abc_19068_n1789;
  wire _abc_19068_n1790;
  wire _abc_19068_n1792;
  wire _abc_19068_n1793;
  wire _abc_19068_n1794;
  wire _abc_19068_n1796;
  wire _abc_19068_n1797;
  wire _abc_19068_n1798;
  wire _abc_19068_n1800;
  wire _abc_19068_n1801;
  wire _abc_19068_n1802;
  wire _abc_19068_n1804;
  wire _abc_19068_n1805;
  wire _abc_19068_n1806;
  wire _abc_19068_n1808;
  wire _abc_19068_n1809;
  wire _abc_19068_n1810;
  wire _abc_19068_n1812;
  wire _abc_19068_n1813;
  wire _abc_19068_n1814;
  wire _abc_19068_n1816;
  wire _abc_19068_n1817;
  wire _abc_19068_n1818;
  wire _abc_19068_n1820;
  wire _abc_19068_n1821;
  wire _abc_19068_n1822;
  wire _abc_19068_n1824;
  wire _abc_19068_n1825;
  wire _abc_19068_n1826;
  wire _abc_19068_n1828;
  wire _abc_19068_n1829;
  wire _abc_19068_n1830;
  wire _abc_19068_n1832;
  wire _abc_19068_n1833;
  wire _abc_19068_n1834;
  wire _abc_19068_n1836;
  wire _abc_19068_n1837;
  wire _abc_19068_n1838;
  wire _abc_19068_n1840;
  wire _abc_19068_n1841;
  wire _abc_19068_n1842;
  wire _abc_19068_n1844;
  wire _abc_19068_n1845;
  wire _abc_19068_n1846;
  wire _abc_19068_n1848;
  wire _abc_19068_n1849;
  wire _abc_19068_n1850;
  wire _abc_19068_n1852;
  wire _abc_19068_n1853;
  wire _abc_19068_n1854;
  wire _abc_19068_n1856;
  wire _abc_19068_n1857;
  wire _abc_19068_n1858;
  wire _abc_19068_n1860;
  wire _abc_19068_n1861;
  wire _abc_19068_n1862;
  wire _abc_19068_n1864;
  wire _abc_19068_n1865;
  wire _abc_19068_n1866;
  wire _abc_19068_n1868;
  wire _abc_19068_n1869;
  wire _abc_19068_n1870;
  wire _abc_19068_n1872;
  wire _abc_19068_n1873;
  wire _abc_19068_n1874;
  wire _abc_19068_n1876;
  wire _abc_19068_n1877;
  wire _abc_19068_n1878;
  wire _abc_19068_n1880;
  wire _abc_19068_n1881;
  wire _abc_19068_n1882;
  wire _abc_19068_n1884;
  wire _abc_19068_n1885;
  wire _abc_19068_n1886;
  wire _abc_19068_n1888;
  wire _abc_19068_n1889;
  wire _abc_19068_n1890;
  wire _abc_19068_n1892;
  wire _abc_19068_n1893;
  wire _abc_19068_n1894;
  wire _abc_19068_n1896;
  wire _abc_19068_n1897;
  wire _abc_19068_n1898;
  wire _abc_19068_n1900;
  wire _abc_19068_n1901;
  wire _abc_19068_n1902;
  wire _abc_19068_n1904;
  wire _abc_19068_n1905;
  wire _abc_19068_n1906;
  wire _abc_19068_n1908;
  wire _abc_19068_n1909;
  wire _abc_19068_n1910;
  wire _abc_19068_n1912;
  wire _abc_19068_n1913;
  wire _abc_19068_n1914;
  wire _abc_19068_n1916;
  wire _abc_19068_n1917;
  wire _abc_19068_n1918;
  wire _abc_19068_n1920;
  wire _abc_19068_n1921;
  wire _abc_19068_n1922;
  wire _abc_19068_n1924;
  wire _abc_19068_n1925;
  wire _abc_19068_n1926;
  wire _abc_19068_n1928;
  wire _abc_19068_n1929;
  wire _abc_19068_n1930;
  wire _abc_19068_n1932;
  wire _abc_19068_n1933;
  wire _abc_19068_n1934;
  wire _abc_19068_n1936;
  wire _abc_19068_n1937;
  wire _abc_19068_n1938;
  wire _abc_19068_n1940;
  wire _abc_19068_n1941;
  wire _abc_19068_n1942;
  wire _abc_19068_n1944;
  wire _abc_19068_n1945;
  wire _abc_19068_n1946;
  wire _abc_19068_n1948;
  wire _abc_19068_n1949;
  wire _abc_19068_n1950;
  wire _abc_19068_n1952;
  wire _abc_19068_n1953;
  wire _abc_19068_n1954;
  wire _abc_19068_n1956;
  wire _abc_19068_n1957;
  wire _abc_19068_n1958;
  wire _abc_19068_n1960;
  wire _abc_19068_n1961;
  wire _abc_19068_n1962;
  wire _abc_19068_n1964;
  wire _abc_19068_n1965;
  wire _abc_19068_n1966;
  wire _abc_19068_n1968;
  wire _abc_19068_n1969;
  wire _abc_19068_n1970;
  wire _abc_19068_n1972;
  wire _abc_19068_n1973;
  wire _abc_19068_n1974;
  wire _abc_19068_n1976;
  wire _abc_19068_n1977;
  wire _abc_19068_n1978;
  wire _abc_19068_n1980;
  wire _abc_19068_n1981;
  wire _abc_19068_n1982;
  wire _abc_19068_n1984;
  wire _abc_19068_n1985;
  wire _abc_19068_n1986;
  wire _abc_19068_n1988;
  wire _abc_19068_n1989;
  wire _abc_19068_n1990;
  wire _abc_19068_n1992;
  wire _abc_19068_n1993;
  wire _abc_19068_n1994;
  wire _abc_19068_n1996;
  wire _abc_19068_n1997;
  wire _abc_19068_n1998;
  wire _abc_19068_n2000;
  wire _abc_19068_n2001;
  wire _abc_19068_n2002;
  wire _abc_19068_n2004;
  wire _abc_19068_n2005;
  wire _abc_19068_n2006;
  wire _abc_19068_n2008;
  wire _abc_19068_n2009;
  wire _abc_19068_n2010;
  wire _abc_19068_n2012;
  wire _abc_19068_n2013;
  wire _abc_19068_n2014;
  wire _abc_19068_n2016;
  wire _abc_19068_n2017;
  wire _abc_19068_n2018;
  wire _abc_19068_n2020;
  wire _abc_19068_n2021;
  wire _abc_19068_n2022;
  wire _abc_19068_n2024;
  wire _abc_19068_n2025;
  wire _abc_19068_n2026;
  wire _abc_19068_n2028;
  wire _abc_19068_n2029;
  wire _abc_19068_n2030;
  wire _abc_19068_n2032;
  wire _abc_19068_n2033;
  wire _abc_19068_n2034;
  wire _abc_19068_n2036;
  wire _abc_19068_n2037;
  wire _abc_19068_n2038;
  wire _abc_19068_n2040;
  wire _abc_19068_n2041;
  wire _abc_19068_n2042;
  wire _abc_19068_n2044;
  wire _abc_19068_n2045;
  wire _abc_19068_n2046;
  wire _abc_19068_n2048;
  wire _abc_19068_n2049;
  wire _abc_19068_n2050;
  wire _abc_19068_n2052;
  wire _abc_19068_n2053;
  wire _abc_19068_n2054;
  wire _abc_19068_n2056;
  wire _abc_19068_n2057;
  wire _abc_19068_n2058;
  wire _abc_19068_n2060;
  wire _abc_19068_n2061;
  wire _abc_19068_n2062;
  wire _abc_19068_n2064;
  wire _abc_19068_n2065;
  wire _abc_19068_n2066;
  wire _abc_19068_n2068;
  wire _abc_19068_n2069;
  wire _abc_19068_n2070;
  wire _abc_19068_n2072;
  wire _abc_19068_n2073;
  wire _abc_19068_n2074;
  wire _abc_19068_n2076;
  wire _abc_19068_n2077;
  wire _abc_19068_n2078;
  wire _abc_19068_n2080;
  wire _abc_19068_n2081;
  wire _abc_19068_n2082;
  wire _abc_19068_n2084;
  wire _abc_19068_n2085;
  wire _abc_19068_n2086;
  wire _abc_19068_n2088;
  wire _abc_19068_n2089;
  wire _abc_19068_n2090;
  wire _abc_19068_n2092;
  wire _abc_19068_n2093;
  wire _abc_19068_n2094;
  wire _abc_19068_n2096;
  wire _abc_19068_n2097;
  wire _abc_19068_n2098;
  wire _abc_19068_n2100;
  wire _abc_19068_n2101;
  wire _abc_19068_n2102;
  wire _abc_19068_n2104;
  wire _abc_19068_n2105;
  wire _abc_19068_n2106;
  wire _abc_19068_n2108;
  wire _abc_19068_n2109;
  wire _abc_19068_n2110;
  wire _abc_19068_n2112;
  wire _abc_19068_n2113;
  wire _abc_19068_n2114;
  wire _abc_19068_n2116;
  wire _abc_19068_n2117;
  wire _abc_19068_n2118;
  wire _abc_19068_n2120;
  wire _abc_19068_n2121;
  wire _abc_19068_n2122;
  wire _abc_19068_n2124;
  wire _abc_19068_n2125;
  wire _abc_19068_n2126;
  wire _abc_19068_n2128;
  wire _abc_19068_n2129;
  wire _abc_19068_n2130;
  wire _abc_19068_n2132;
  wire _abc_19068_n2133;
  wire _abc_19068_n2133_bF_buf0;
  wire _abc_19068_n2133_bF_buf1;
  wire _abc_19068_n2133_bF_buf2;
  wire _abc_19068_n2133_bF_buf3;
  wire _abc_19068_n2133_bF_buf4;
  wire _abc_19068_n2133_bF_buf5;
  wire _abc_19068_n2133_bF_buf6;
  wire _abc_19068_n2133_bF_buf7;
  wire _abc_19068_n2134;
  wire _abc_19068_n2135;
  wire _abc_19068_n2136;
  wire _abc_19068_n2137;
  wire _abc_19068_n2138;
  wire _abc_19068_n2140;
  wire _abc_19068_n2141;
  wire _abc_19068_n2142;
  wire _abc_19068_n2143;
  wire _abc_19068_n2144;
  wire _abc_19068_n2146;
  wire _abc_19068_n2147;
  wire _abc_19068_n2148;
  wire _abc_19068_n2149;
  wire _abc_19068_n2150;
  wire _abc_19068_n2152;
  wire _abc_19068_n2153;
  wire _abc_19068_n2154;
  wire _abc_19068_n2155;
  wire _abc_19068_n2156;
  wire _abc_19068_n2158;
  wire _abc_19068_n2159;
  wire _abc_19068_n2160;
  wire _abc_19068_n2161;
  wire _abc_19068_n2162;
  wire _abc_19068_n2164;
  wire _abc_19068_n2165;
  wire _abc_19068_n2166;
  wire _abc_19068_n2167;
  wire _abc_19068_n2168;
  wire _abc_19068_n2170;
  wire _abc_19068_n2171;
  wire _abc_19068_n2172;
  wire _abc_19068_n2173;
  wire _abc_19068_n2174;
  wire _abc_19068_n2176;
  wire _abc_19068_n2177;
  wire _abc_19068_n2178;
  wire _abc_19068_n2179;
  wire _abc_19068_n2180;
  wire _abc_19068_n2182;
  wire _abc_19068_n2183;
  wire _abc_19068_n2184;
  wire _abc_19068_n2185;
  wire _abc_19068_n2186;
  wire _abc_19068_n2188;
  wire _abc_19068_n2189;
  wire _abc_19068_n2190;
  wire _abc_19068_n2191;
  wire _abc_19068_n2192;
  wire _abc_19068_n2194;
  wire _abc_19068_n2195;
  wire _abc_19068_n2196;
  wire _abc_19068_n2197;
  wire _abc_19068_n2198;
  wire _abc_19068_n2200;
  wire _abc_19068_n2201;
  wire _abc_19068_n2202;
  wire _abc_19068_n2203;
  wire _abc_19068_n2204;
  wire _abc_19068_n2206;
  wire _abc_19068_n2207;
  wire _abc_19068_n2208;
  wire _abc_19068_n2209;
  wire _abc_19068_n2210;
  wire _abc_19068_n2212;
  wire _abc_19068_n2213;
  wire _abc_19068_n2214;
  wire _abc_19068_n2215;
  wire _abc_19068_n2216;
  wire _abc_19068_n2218;
  wire _abc_19068_n2219;
  wire _abc_19068_n2220;
  wire _abc_19068_n2221;
  wire _abc_19068_n2222;
  wire _abc_19068_n2224;
  wire _abc_19068_n2225;
  wire _abc_19068_n2226;
  wire _abc_19068_n2227;
  wire _abc_19068_n2228;
  wire _abc_19068_n2230;
  wire _abc_19068_n2231;
  wire _abc_19068_n2232;
  wire _abc_19068_n2233;
  wire _abc_19068_n2234;
  wire _abc_19068_n2236;
  wire _abc_19068_n2237;
  wire _abc_19068_n2238;
  wire _abc_19068_n2239;
  wire _abc_19068_n2240;
  wire _abc_19068_n2242;
  wire _abc_19068_n2243;
  wire _abc_19068_n2244;
  wire _abc_19068_n2245;
  wire _abc_19068_n2246;
  wire _abc_19068_n2248;
  wire _abc_19068_n2249;
  wire _abc_19068_n2250;
  wire _abc_19068_n2251;
  wire _abc_19068_n2252;
  wire _abc_19068_n2254;
  wire _abc_19068_n2255;
  wire _abc_19068_n2256;
  wire _abc_19068_n2257;
  wire _abc_19068_n2258;
  wire _abc_19068_n2260;
  wire _abc_19068_n2261;
  wire _abc_19068_n2262;
  wire _abc_19068_n2263;
  wire _abc_19068_n2264;
  wire _abc_19068_n2266;
  wire _abc_19068_n2267;
  wire _abc_19068_n2268;
  wire _abc_19068_n2269;
  wire _abc_19068_n2270;
  wire _abc_19068_n2272;
  wire _abc_19068_n2273;
  wire _abc_19068_n2274;
  wire _abc_19068_n2275;
  wire _abc_19068_n2276;
  wire _abc_19068_n2278;
  wire _abc_19068_n2279;
  wire _abc_19068_n2280;
  wire _abc_19068_n2281;
  wire _abc_19068_n2282;
  wire _abc_19068_n2284;
  wire _abc_19068_n2285;
  wire _abc_19068_n2286;
  wire _abc_19068_n2287;
  wire _abc_19068_n2288;
  wire _abc_19068_n2290;
  wire _abc_19068_n2291;
  wire _abc_19068_n2292;
  wire _abc_19068_n2293;
  wire _abc_19068_n2294;
  wire _abc_19068_n2296;
  wire _abc_19068_n2297;
  wire _abc_19068_n2298;
  wire _abc_19068_n2299;
  wire _abc_19068_n2300;
  wire _abc_19068_n2302;
  wire _abc_19068_n2303;
  wire _abc_19068_n2304;
  wire _abc_19068_n2305;
  wire _abc_19068_n2306;
  wire _abc_19068_n2308;
  wire _abc_19068_n2309;
  wire _abc_19068_n2310;
  wire _abc_19068_n2311;
  wire _abc_19068_n2312;
  wire _abc_19068_n2314;
  wire _abc_19068_n2315;
  wire _abc_19068_n2316;
  wire _abc_19068_n2317;
  wire _abc_19068_n2318;
  wire _abc_19068_n2320;
  wire _abc_19068_n2321;
  wire _abc_19068_n2322;
  wire _abc_19068_n2323;
  wire _abc_19068_n2324;
  wire _abc_19068_n2326;
  wire _abc_19068_n2326_bF_buf0;
  wire _abc_19068_n2326_bF_buf1;
  wire _abc_19068_n2326_bF_buf2;
  wire _abc_19068_n2326_bF_buf3;
  wire _abc_19068_n2326_bF_buf4;
  wire _abc_19068_n2326_bF_buf5;
  wire _abc_19068_n2326_bF_buf6;
  wire _abc_19068_n2326_bF_buf7;
  wire _abc_19068_n2327;
  wire _abc_19068_n2328;
  wire _abc_19068_n2329;
  wire _abc_19068_n2330;
  wire _abc_19068_n2332;
  wire _abc_19068_n2333;
  wire _abc_19068_n2334;
  wire _abc_19068_n2335;
  wire _abc_19068_n2337;
  wire _abc_19068_n2338;
  wire _abc_19068_n2339;
  wire _abc_19068_n2340;
  wire _abc_19068_n2342;
  wire _abc_19068_n2343;
  wire _abc_19068_n2344;
  wire _abc_19068_n2345;
  wire _abc_19068_n2347;
  wire _abc_19068_n2348;
  wire _abc_19068_n2349;
  wire _abc_19068_n2350;
  wire _abc_19068_n2352;
  wire _abc_19068_n2353;
  wire _abc_19068_n2354;
  wire _abc_19068_n2355;
  wire _abc_19068_n2357;
  wire _abc_19068_n2358;
  wire _abc_19068_n2359;
  wire _abc_19068_n2360;
  wire _abc_19068_n2362;
  wire _abc_19068_n2363;
  wire _abc_19068_n2364;
  wire _abc_19068_n2365;
  wire _abc_19068_n2367;
  wire _abc_19068_n2368;
  wire _abc_19068_n2369;
  wire _abc_19068_n2370;
  wire _abc_19068_n2372;
  wire _abc_19068_n2373;
  wire _abc_19068_n2374;
  wire _abc_19068_n2375;
  wire _abc_19068_n2377;
  wire _abc_19068_n2378;
  wire _abc_19068_n2379;
  wire _abc_19068_n2380;
  wire _abc_19068_n2382;
  wire _abc_19068_n2383;
  wire _abc_19068_n2384;
  wire _abc_19068_n2385;
  wire _abc_19068_n2387;
  wire _abc_19068_n2388;
  wire _abc_19068_n2389;
  wire _abc_19068_n2390;
  wire _abc_19068_n2392;
  wire _abc_19068_n2393;
  wire _abc_19068_n2394;
  wire _abc_19068_n2395;
  wire _abc_19068_n2397;
  wire _abc_19068_n2398;
  wire _abc_19068_n2399;
  wire _abc_19068_n2400;
  wire _abc_19068_n2402;
  wire _abc_19068_n2403;
  wire _abc_19068_n2404;
  wire _abc_19068_n2405;
  wire _abc_19068_n2407;
  wire _abc_19068_n2408;
  wire _abc_19068_n2409;
  wire _abc_19068_n2410;
  wire _abc_19068_n2412;
  wire _abc_19068_n2413;
  wire _abc_19068_n2414;
  wire _abc_19068_n2415;
  wire _abc_19068_n2417;
  wire _abc_19068_n2418;
  wire _abc_19068_n2419;
  wire _abc_19068_n2420;
  wire _abc_19068_n2422;
  wire _abc_19068_n2423;
  wire _abc_19068_n2424;
  wire _abc_19068_n2425;
  wire _abc_19068_n2427;
  wire _abc_19068_n2428;
  wire _abc_19068_n2429;
  wire _abc_19068_n2430;
  wire _abc_19068_n2432;
  wire _abc_19068_n2433;
  wire _abc_19068_n2434;
  wire _abc_19068_n2435;
  wire _abc_19068_n2437;
  wire _abc_19068_n2438;
  wire _abc_19068_n2439;
  wire _abc_19068_n2440;
  wire _abc_19068_n2442;
  wire _abc_19068_n2443;
  wire _abc_19068_n2444;
  wire _abc_19068_n2445;
  wire _abc_19068_n2447;
  wire _abc_19068_n2448;
  wire _abc_19068_n2449;
  wire _abc_19068_n2450;
  wire _abc_19068_n2452;
  wire _abc_19068_n2453;
  wire _abc_19068_n2454;
  wire _abc_19068_n2455;
  wire _abc_19068_n2457;
  wire _abc_19068_n2458;
  wire _abc_19068_n2459;
  wire _abc_19068_n2460;
  wire _abc_19068_n2462;
  wire _abc_19068_n2463;
  wire _abc_19068_n2464;
  wire _abc_19068_n2465;
  wire _abc_19068_n2467;
  wire _abc_19068_n2468;
  wire _abc_19068_n2469;
  wire _abc_19068_n2470;
  wire _abc_19068_n2472;
  wire _abc_19068_n2473;
  wire _abc_19068_n2474;
  wire _abc_19068_n2475;
  wire _abc_19068_n2477;
  wire _abc_19068_n2478;
  wire _abc_19068_n2479;
  wire _abc_19068_n2480;
  wire _abc_19068_n2482;
  wire _abc_19068_n2483;
  wire _abc_19068_n2484;
  wire _abc_19068_n2485;
  wire _abc_19068_n2487;
  wire _abc_19068_n2487_bF_buf0;
  wire _abc_19068_n2487_bF_buf1;
  wire _abc_19068_n2487_bF_buf2;
  wire _abc_19068_n2487_bF_buf3;
  wire _abc_19068_n2487_bF_buf4;
  wire _abc_19068_n2487_bF_buf5;
  wire _abc_19068_n2487_bF_buf6;
  wire _abc_19068_n2487_bF_buf7;
  wire _abc_19068_n2488;
  wire _abc_19068_n2489;
  wire _abc_19068_n2490;
  wire _abc_19068_n2491;
  wire _abc_19068_n2493;
  wire _abc_19068_n2494;
  wire _abc_19068_n2495;
  wire _abc_19068_n2496;
  wire _abc_19068_n2498;
  wire _abc_19068_n2499;
  wire _abc_19068_n2500;
  wire _abc_19068_n2501;
  wire _abc_19068_n2503;
  wire _abc_19068_n2504;
  wire _abc_19068_n2505;
  wire _abc_19068_n2506;
  wire _abc_19068_n2508;
  wire _abc_19068_n2509;
  wire _abc_19068_n2510;
  wire _abc_19068_n2511;
  wire _abc_19068_n2513;
  wire _abc_19068_n2514;
  wire _abc_19068_n2515;
  wire _abc_19068_n2516;
  wire _abc_19068_n2518;
  wire _abc_19068_n2519;
  wire _abc_19068_n2520;
  wire _abc_19068_n2521;
  wire _abc_19068_n2523;
  wire _abc_19068_n2524;
  wire _abc_19068_n2525;
  wire _abc_19068_n2526;
  wire _abc_19068_n2528;
  wire _abc_19068_n2529;
  wire _abc_19068_n2530;
  wire _abc_19068_n2531;
  wire _abc_19068_n2533;
  wire _abc_19068_n2534;
  wire _abc_19068_n2535;
  wire _abc_19068_n2536;
  wire _abc_19068_n2538;
  wire _abc_19068_n2539;
  wire _abc_19068_n2540;
  wire _abc_19068_n2541;
  wire _abc_19068_n2543;
  wire _abc_19068_n2544;
  wire _abc_19068_n2545;
  wire _abc_19068_n2546;
  wire _abc_19068_n2548;
  wire _abc_19068_n2549;
  wire _abc_19068_n2550;
  wire _abc_19068_n2551;
  wire _abc_19068_n2553;
  wire _abc_19068_n2554;
  wire _abc_19068_n2555;
  wire _abc_19068_n2556;
  wire _abc_19068_n2558;
  wire _abc_19068_n2559;
  wire _abc_19068_n2560;
  wire _abc_19068_n2561;
  wire _abc_19068_n2563;
  wire _abc_19068_n2564;
  wire _abc_19068_n2565;
  wire _abc_19068_n2566;
  wire _abc_19068_n2568;
  wire _abc_19068_n2569;
  wire _abc_19068_n2570;
  wire _abc_19068_n2571;
  wire _abc_19068_n2573;
  wire _abc_19068_n2574;
  wire _abc_19068_n2575;
  wire _abc_19068_n2576;
  wire _abc_19068_n2578;
  wire _abc_19068_n2579;
  wire _abc_19068_n2580;
  wire _abc_19068_n2581;
  wire _abc_19068_n2583;
  wire _abc_19068_n2584;
  wire _abc_19068_n2585;
  wire _abc_19068_n2586;
  wire _abc_19068_n2588;
  wire _abc_19068_n2589;
  wire _abc_19068_n2590;
  wire _abc_19068_n2591;
  wire _abc_19068_n2593;
  wire _abc_19068_n2594;
  wire _abc_19068_n2595;
  wire _abc_19068_n2596;
  wire _abc_19068_n2598;
  wire _abc_19068_n2599;
  wire _abc_19068_n2600;
  wire _abc_19068_n2601;
  wire _abc_19068_n2603;
  wire _abc_19068_n2604;
  wire _abc_19068_n2605;
  wire _abc_19068_n2606;
  wire _abc_19068_n2608;
  wire _abc_19068_n2609;
  wire _abc_19068_n2610;
  wire _abc_19068_n2611;
  wire _abc_19068_n2613;
  wire _abc_19068_n2614;
  wire _abc_19068_n2615;
  wire _abc_19068_n2616;
  wire _abc_19068_n2618;
  wire _abc_19068_n2619;
  wire _abc_19068_n2620;
  wire _abc_19068_n2621;
  wire _abc_19068_n2623;
  wire _abc_19068_n2624;
  wire _abc_19068_n2625;
  wire _abc_19068_n2626;
  wire _abc_19068_n2628;
  wire _abc_19068_n2629;
  wire _abc_19068_n2630;
  wire _abc_19068_n2631;
  wire _abc_19068_n2633;
  wire _abc_19068_n2634;
  wire _abc_19068_n2635;
  wire _abc_19068_n2636;
  wire _abc_19068_n2638;
  wire _abc_19068_n2639;
  wire _abc_19068_n2640;
  wire _abc_19068_n2641;
  wire _abc_19068_n2643;
  wire _abc_19068_n2644;
  wire _abc_19068_n2645;
  wire _abc_19068_n2646;
  wire _abc_19068_n2648;
  wire _abc_19068_n2648_bF_buf0;
  wire _abc_19068_n2648_bF_buf1;
  wire _abc_19068_n2648_bF_buf2;
  wire _abc_19068_n2648_bF_buf3;
  wire _abc_19068_n2648_bF_buf4;
  wire _abc_19068_n2648_bF_buf5;
  wire _abc_19068_n2648_bF_buf6;
  wire _abc_19068_n2648_bF_buf7;
  wire _abc_19068_n2649;
  wire _abc_19068_n2650;
  wire _abc_19068_n2651;
  wire _abc_19068_n2652;
  wire _abc_19068_n2654;
  wire _abc_19068_n2655;
  wire _abc_19068_n2656;
  wire _abc_19068_n2657;
  wire _abc_19068_n2659;
  wire _abc_19068_n2660;
  wire _abc_19068_n2661;
  wire _abc_19068_n2662;
  wire _abc_19068_n2664;
  wire _abc_19068_n2665;
  wire _abc_19068_n2666;
  wire _abc_19068_n2667;
  wire _abc_19068_n2669;
  wire _abc_19068_n2670;
  wire _abc_19068_n2671;
  wire _abc_19068_n2672;
  wire _abc_19068_n2674;
  wire _abc_19068_n2675;
  wire _abc_19068_n2676;
  wire _abc_19068_n2677;
  wire _abc_19068_n2679;
  wire _abc_19068_n2680;
  wire _abc_19068_n2681;
  wire _abc_19068_n2682;
  wire _abc_19068_n2684;
  wire _abc_19068_n2685;
  wire _abc_19068_n2686;
  wire _abc_19068_n2687;
  wire _abc_19068_n2689;
  wire _abc_19068_n2690;
  wire _abc_19068_n2691;
  wire _abc_19068_n2692;
  wire _abc_19068_n2694;
  wire _abc_19068_n2695;
  wire _abc_19068_n2696;
  wire _abc_19068_n2697;
  wire _abc_19068_n2699;
  wire _abc_19068_n2700;
  wire _abc_19068_n2701;
  wire _abc_19068_n2702;
  wire _abc_19068_n2704;
  wire _abc_19068_n2705;
  wire _abc_19068_n2706;
  wire _abc_19068_n2707;
  wire _abc_19068_n2709;
  wire _abc_19068_n2710;
  wire _abc_19068_n2711;
  wire _abc_19068_n2712;
  wire _abc_19068_n2714;
  wire _abc_19068_n2715;
  wire _abc_19068_n2716;
  wire _abc_19068_n2717;
  wire _abc_19068_n2719;
  wire _abc_19068_n2720;
  wire _abc_19068_n2721;
  wire _abc_19068_n2722;
  wire _abc_19068_n2724;
  wire _abc_19068_n2725;
  wire _abc_19068_n2726;
  wire _abc_19068_n2727;
  wire _abc_19068_n2729;
  wire _abc_19068_n2730;
  wire _abc_19068_n2731;
  wire _abc_19068_n2732;
  wire _abc_19068_n2734;
  wire _abc_19068_n2735;
  wire _abc_19068_n2736;
  wire _abc_19068_n2737;
  wire _abc_19068_n2739;
  wire _abc_19068_n2740;
  wire _abc_19068_n2741;
  wire _abc_19068_n2742;
  wire _abc_19068_n2744;
  wire _abc_19068_n2745;
  wire _abc_19068_n2746;
  wire _abc_19068_n2747;
  wire _abc_19068_n2749;
  wire _abc_19068_n2750;
  wire _abc_19068_n2751;
  wire _abc_19068_n2752;
  wire _abc_19068_n2754;
  wire _abc_19068_n2755;
  wire _abc_19068_n2756;
  wire _abc_19068_n2757;
  wire _abc_19068_n2759;
  wire _abc_19068_n2760;
  wire _abc_19068_n2761;
  wire _abc_19068_n2762;
  wire _abc_19068_n2764;
  wire _abc_19068_n2765;
  wire _abc_19068_n2766;
  wire _abc_19068_n2767;
  wire _abc_19068_n2769;
  wire _abc_19068_n2770;
  wire _abc_19068_n2771;
  wire _abc_19068_n2772;
  wire _abc_19068_n2774;
  wire _abc_19068_n2775;
  wire _abc_19068_n2776;
  wire _abc_19068_n2777;
  wire _abc_19068_n2779;
  wire _abc_19068_n2780;
  wire _abc_19068_n2781;
  wire _abc_19068_n2782;
  wire _abc_19068_n2784;
  wire _abc_19068_n2785;
  wire _abc_19068_n2786;
  wire _abc_19068_n2787;
  wire _abc_19068_n2789;
  wire _abc_19068_n2790;
  wire _abc_19068_n2791;
  wire _abc_19068_n2792;
  wire _abc_19068_n2794;
  wire _abc_19068_n2795;
  wire _abc_19068_n2796;
  wire _abc_19068_n2797;
  wire _abc_19068_n2799;
  wire _abc_19068_n2800;
  wire _abc_19068_n2801;
  wire _abc_19068_n2802;
  wire _abc_19068_n2804;
  wire _abc_19068_n2805;
  wire _abc_19068_n2806;
  wire _abc_19068_n2807;
  wire _abc_19068_n2809;
  wire _abc_19068_n2809_bF_buf0;
  wire _abc_19068_n2809_bF_buf1;
  wire _abc_19068_n2809_bF_buf2;
  wire _abc_19068_n2809_bF_buf3;
  wire _abc_19068_n2809_bF_buf4;
  wire _abc_19068_n2809_bF_buf5;
  wire _abc_19068_n2809_bF_buf6;
  wire _abc_19068_n2809_bF_buf7;
  wire _abc_19068_n2810;
  wire _abc_19068_n2811;
  wire _abc_19068_n2812;
  wire _abc_19068_n2813;
  wire _abc_19068_n2815;
  wire _abc_19068_n2816;
  wire _abc_19068_n2817;
  wire _abc_19068_n2818;
  wire _abc_19068_n2820;
  wire _abc_19068_n2821;
  wire _abc_19068_n2822;
  wire _abc_19068_n2823;
  wire _abc_19068_n2825;
  wire _abc_19068_n2826;
  wire _abc_19068_n2827;
  wire _abc_19068_n2828;
  wire _abc_19068_n2830;
  wire _abc_19068_n2831;
  wire _abc_19068_n2832;
  wire _abc_19068_n2833;
  wire _abc_19068_n2835;
  wire _abc_19068_n2836;
  wire _abc_19068_n2837;
  wire _abc_19068_n2838;
  wire _abc_19068_n2840;
  wire _abc_19068_n2841;
  wire _abc_19068_n2842;
  wire _abc_19068_n2843;
  wire _abc_19068_n2845;
  wire _abc_19068_n2846;
  wire _abc_19068_n2847;
  wire _abc_19068_n2848;
  wire _abc_19068_n2850;
  wire _abc_19068_n2851;
  wire _abc_19068_n2852;
  wire _abc_19068_n2853;
  wire _abc_19068_n2855;
  wire _abc_19068_n2856;
  wire _abc_19068_n2857;
  wire _abc_19068_n2858;
  wire _abc_19068_n2860;
  wire _abc_19068_n2861;
  wire _abc_19068_n2862;
  wire _abc_19068_n2863;
  wire _abc_19068_n2865;
  wire _abc_19068_n2866;
  wire _abc_19068_n2867;
  wire _abc_19068_n2868;
  wire _abc_19068_n2870;
  wire _abc_19068_n2871;
  wire _abc_19068_n2872;
  wire _abc_19068_n2873;
  wire _abc_19068_n2875;
  wire _abc_19068_n2876;
  wire _abc_19068_n2877;
  wire _abc_19068_n2878;
  wire _abc_19068_n2880;
  wire _abc_19068_n2881;
  wire _abc_19068_n2882;
  wire _abc_19068_n2883;
  wire _abc_19068_n2885;
  wire _abc_19068_n2886;
  wire _abc_19068_n2887;
  wire _abc_19068_n2888;
  wire _abc_19068_n2890;
  wire _abc_19068_n2891;
  wire _abc_19068_n2892;
  wire _abc_19068_n2893;
  wire _abc_19068_n2895;
  wire _abc_19068_n2896;
  wire _abc_19068_n2897;
  wire _abc_19068_n2898;
  wire _abc_19068_n2900;
  wire _abc_19068_n2901;
  wire _abc_19068_n2902;
  wire _abc_19068_n2903;
  wire _abc_19068_n2905;
  wire _abc_19068_n2906;
  wire _abc_19068_n2907;
  wire _abc_19068_n2908;
  wire _abc_19068_n2910;
  wire _abc_19068_n2911;
  wire _abc_19068_n2912;
  wire _abc_19068_n2913;
  wire _abc_19068_n2915;
  wire _abc_19068_n2916;
  wire _abc_19068_n2917;
  wire _abc_19068_n2918;
  wire _abc_19068_n2920;
  wire _abc_19068_n2921;
  wire _abc_19068_n2922;
  wire _abc_19068_n2923;
  wire _abc_19068_n2925;
  wire _abc_19068_n2926;
  wire _abc_19068_n2927;
  wire _abc_19068_n2928;
  wire _abc_19068_n2930;
  wire _abc_19068_n2931;
  wire _abc_19068_n2932;
  wire _abc_19068_n2933;
  wire _abc_19068_n2935;
  wire _abc_19068_n2936;
  wire _abc_19068_n2937;
  wire _abc_19068_n2938;
  wire _abc_19068_n2940;
  wire _abc_19068_n2941;
  wire _abc_19068_n2942;
  wire _abc_19068_n2943;
  wire _abc_19068_n2945;
  wire _abc_19068_n2946;
  wire _abc_19068_n2947;
  wire _abc_19068_n2948;
  wire _abc_19068_n2950;
  wire _abc_19068_n2951;
  wire _abc_19068_n2952;
  wire _abc_19068_n2953;
  wire _abc_19068_n2955;
  wire _abc_19068_n2956;
  wire _abc_19068_n2957;
  wire _abc_19068_n2958;
  wire _abc_19068_n2960;
  wire _abc_19068_n2961;
  wire _abc_19068_n2962;
  wire _abc_19068_n2963;
  wire _abc_19068_n2965;
  wire _abc_19068_n2966;
  wire _abc_19068_n2967;
  wire _abc_19068_n2968;
  wire _abc_19068_n2970;
  wire _abc_19068_n2970_bF_buf0;
  wire _abc_19068_n2970_bF_buf1;
  wire _abc_19068_n2970_bF_buf2;
  wire _abc_19068_n2970_bF_buf3;
  wire _abc_19068_n2970_bF_buf4;
  wire _abc_19068_n2970_bF_buf5;
  wire _abc_19068_n2970_bF_buf6;
  wire _abc_19068_n2970_bF_buf7;
  wire _abc_19068_n2971;
  wire _abc_19068_n2972;
  wire _abc_19068_n2973;
  wire _abc_19068_n2974;
  wire _abc_19068_n2976;
  wire _abc_19068_n2977;
  wire _abc_19068_n2978;
  wire _abc_19068_n2979;
  wire _abc_19068_n2981;
  wire _abc_19068_n2982;
  wire _abc_19068_n2983;
  wire _abc_19068_n2984;
  wire _abc_19068_n2986;
  wire _abc_19068_n2987;
  wire _abc_19068_n2988;
  wire _abc_19068_n2989;
  wire _abc_19068_n2991;
  wire _abc_19068_n2992;
  wire _abc_19068_n2993;
  wire _abc_19068_n2994;
  wire _abc_19068_n2996;
  wire _abc_19068_n2997;
  wire _abc_19068_n2998;
  wire _abc_19068_n2999;
  wire _abc_19068_n3001;
  wire _abc_19068_n3002;
  wire _abc_19068_n3003;
  wire _abc_19068_n3004;
  wire _abc_19068_n3006;
  wire _abc_19068_n3007;
  wire _abc_19068_n3008;
  wire _abc_19068_n3009;
  wire _abc_19068_n3011;
  wire _abc_19068_n3012;
  wire _abc_19068_n3013;
  wire _abc_19068_n3014;
  wire _abc_19068_n3016;
  wire _abc_19068_n3017;
  wire _abc_19068_n3018;
  wire _abc_19068_n3019;
  wire _abc_19068_n3021;
  wire _abc_19068_n3022;
  wire _abc_19068_n3023;
  wire _abc_19068_n3024;
  wire _abc_19068_n3026;
  wire _abc_19068_n3027;
  wire _abc_19068_n3028;
  wire _abc_19068_n3029;
  wire _abc_19068_n3031;
  wire _abc_19068_n3032;
  wire _abc_19068_n3033;
  wire _abc_19068_n3034;
  wire _abc_19068_n3036;
  wire _abc_19068_n3037;
  wire _abc_19068_n3038;
  wire _abc_19068_n3039;
  wire _abc_19068_n3041;
  wire _abc_19068_n3042;
  wire _abc_19068_n3043;
  wire _abc_19068_n3044;
  wire _abc_19068_n3046;
  wire _abc_19068_n3047;
  wire _abc_19068_n3048;
  wire _abc_19068_n3049;
  wire _abc_19068_n3051;
  wire _abc_19068_n3052;
  wire _abc_19068_n3053;
  wire _abc_19068_n3054;
  wire _abc_19068_n3056;
  wire _abc_19068_n3057;
  wire _abc_19068_n3058;
  wire _abc_19068_n3059;
  wire _abc_19068_n3061;
  wire _abc_19068_n3062;
  wire _abc_19068_n3063;
  wire _abc_19068_n3064;
  wire _abc_19068_n3066;
  wire _abc_19068_n3067;
  wire _abc_19068_n3068;
  wire _abc_19068_n3069;
  wire _abc_19068_n3071;
  wire _abc_19068_n3072;
  wire _abc_19068_n3073;
  wire _abc_19068_n3074;
  wire _abc_19068_n3076;
  wire _abc_19068_n3077;
  wire _abc_19068_n3078;
  wire _abc_19068_n3079;
  wire _abc_19068_n3081;
  wire _abc_19068_n3082;
  wire _abc_19068_n3083;
  wire _abc_19068_n3084;
  wire _abc_19068_n3086;
  wire _abc_19068_n3087;
  wire _abc_19068_n3088;
  wire _abc_19068_n3089;
  wire _abc_19068_n3091;
  wire _abc_19068_n3092;
  wire _abc_19068_n3093;
  wire _abc_19068_n3094;
  wire _abc_19068_n3096;
  wire _abc_19068_n3097;
  wire _abc_19068_n3098;
  wire _abc_19068_n3099;
  wire _abc_19068_n3101;
  wire _abc_19068_n3102;
  wire _abc_19068_n3103;
  wire _abc_19068_n3104;
  wire _abc_19068_n3106;
  wire _abc_19068_n3107;
  wire _abc_19068_n3108;
  wire _abc_19068_n3109;
  wire _abc_19068_n3111;
  wire _abc_19068_n3112;
  wire _abc_19068_n3113;
  wire _abc_19068_n3114;
  wire _abc_19068_n3116;
  wire _abc_19068_n3117;
  wire _abc_19068_n3118;
  wire _abc_19068_n3119;
  wire _abc_19068_n3121;
  wire _abc_19068_n3122;
  wire _abc_19068_n3123;
  wire _abc_19068_n3124;
  wire _abc_19068_n3126;
  wire _abc_19068_n3127;
  wire _abc_19068_n3128;
  wire _abc_19068_n3129;
  wire _abc_19068_n3131;
  wire _abc_19068_n3132;
  wire _abc_19068_n3133;
  wire _abc_19068_n3134;
  wire _abc_19068_n3135;
  wire _abc_19068_n3137;
  wire _abc_19068_n3138;
  wire _abc_19068_n3139;
  wire _abc_19068_n3140;
  wire _abc_19068_n3142;
  wire _abc_19068_n3143;
  wire _abc_19068_n3144;
  wire _abc_19068_n3146;
  wire _abc_19068_n3147;
  wire _abc_19068_n3148;
  wire _abc_19068_n3150;
  wire _abc_19068_n3151;
  wire _abc_19068_n3152;
  wire _abc_19068_n3154;
  wire _abc_19068_n3155;
  wire _abc_19068_n3156;
  wire _abc_19068_n3158;
  wire _abc_19068_n3159;
  wire _abc_19068_n3160;
  wire _abc_19068_n3162;
  wire _abc_19068_n3163;
  wire _abc_19068_n3164;
  wire _abc_19068_n3166;
  wire _abc_19068_n3167;
  wire _abc_19068_n3169;
  wire _abc_19068_n3171;
  wire _abc_19068_n3173;
  wire _abc_19068_n3174;
  wire _abc_19068_n3175;
  wire _abc_19068_n3176;
  wire _abc_19068_n3177;
  wire _abc_19068_n3178;
  wire _abc_19068_n3179;
  wire _abc_19068_n870_1;
  wire _abc_19068_n871_1;
  wire _abc_19068_n872;
  wire _abc_19068_n873_1;
  wire _abc_19068_n874_1;
  wire _abc_19068_n875;
  wire _abc_19068_n876_1;
  wire _abc_19068_n877_1;
  wire _abc_19068_n878;
  wire _abc_19068_n879_1;
  wire _abc_19068_n880_1;
  wire _abc_19068_n881;
  wire _abc_19068_n882_1;
  wire _abc_19068_n883_1;
  wire _abc_19068_n884;
  wire _abc_19068_n885_1;
  wire _abc_19068_n886_1;
  wire _abc_19068_n887;
  wire _abc_19068_n888_1;
  wire _abc_19068_n889_1;
  wire _abc_19068_n890;
  wire _abc_19068_n891_1;
  wire _abc_19068_n892_1;
  wire _abc_19068_n893;
  wire _abc_19068_n894_1;
  wire _abc_19068_n895_1;
  wire _abc_19068_n896;
  wire _abc_19068_n897_1;
  wire _abc_19068_n897_1_bF_buf0;
  wire _abc_19068_n897_1_bF_buf1;
  wire _abc_19068_n897_1_bF_buf2;
  wire _abc_19068_n897_1_bF_buf3;
  wire _abc_19068_n897_1_bF_buf4;
  wire _abc_19068_n898_1;
  wire _abc_19068_n899;
  wire _abc_19068_n899_bF_buf0;
  wire _abc_19068_n899_bF_buf1;
  wire _abc_19068_n899_bF_buf2;
  wire _abc_19068_n899_bF_buf3;
  wire _abc_19068_n899_bF_buf4;
  wire _abc_19068_n900_1;
  wire _abc_19068_n901_1;
  wire _abc_19068_n902;
  wire _abc_19068_n902_bF_buf0;
  wire _abc_19068_n902_bF_buf1;
  wire _abc_19068_n902_bF_buf2;
  wire _abc_19068_n902_bF_buf3;
  wire _abc_19068_n902_bF_buf4;
  wire _abc_19068_n903_1;
  wire _abc_19068_n904_1;
  wire _abc_19068_n905;
  wire _abc_19068_n906_1;
  wire _abc_19068_n907_1;
  wire _abc_19068_n908;
  wire _abc_19068_n909_1;
  wire _abc_19068_n910_1;
  wire _abc_19068_n911;
  wire _abc_19068_n912_1;
  wire _abc_19068_n913_1;
  wire _abc_19068_n914;
  wire _abc_19068_n915_1;
  wire _abc_19068_n915_1_bF_buf0;
  wire _abc_19068_n915_1_bF_buf1;
  wire _abc_19068_n915_1_bF_buf2;
  wire _abc_19068_n915_1_bF_buf3;
  wire _abc_19068_n915_1_bF_buf4;
  wire _abc_19068_n916_1;
  wire _abc_19068_n916_1_bF_buf0;
  wire _abc_19068_n916_1_bF_buf1;
  wire _abc_19068_n916_1_bF_buf2;
  wire _abc_19068_n916_1_bF_buf3;
  wire _abc_19068_n916_1_bF_buf4;
  wire _abc_19068_n917;
  wire _abc_19068_n918_1;
  wire _abc_19068_n919_1;
  wire _abc_19068_n920;
  wire _abc_19068_n921_1;
  wire _abc_19068_n922_1;
  wire _abc_19068_n923;
  wire _abc_19068_n923_bF_buf0;
  wire _abc_19068_n923_bF_buf1;
  wire _abc_19068_n923_bF_buf2;
  wire _abc_19068_n923_bF_buf3;
  wire _abc_19068_n923_bF_buf4;
  wire _abc_19068_n924_1;
  wire _abc_19068_n924_1_bF_buf0;
  wire _abc_19068_n924_1_bF_buf1;
  wire _abc_19068_n924_1_bF_buf2;
  wire _abc_19068_n924_1_bF_buf3;
  wire _abc_19068_n924_1_bF_buf4;
  wire _abc_19068_n925_1;
  wire _abc_19068_n926;
  wire _abc_19068_n926_bF_buf0;
  wire _abc_19068_n926_bF_buf1;
  wire _abc_19068_n926_bF_buf2;
  wire _abc_19068_n926_bF_buf3;
  wire _abc_19068_n926_bF_buf4;
  wire _abc_19068_n927_1;
  wire _abc_19068_n928_1;
  wire _abc_19068_n929;
  wire _abc_19068_n930_1;
  wire _abc_19068_n931_1;
  wire _abc_19068_n932;
  wire _abc_19068_n933_1;
  wire _abc_19068_n934_1;
  wire _abc_19068_n935;
  wire _abc_19068_n936_1;
  wire _abc_19068_n937_1;
  wire _abc_19068_n938;
  wire _abc_19068_n939_1;
  wire _abc_19068_n939_1_bF_buf0;
  wire _abc_19068_n939_1_bF_buf1;
  wire _abc_19068_n939_1_bF_buf2;
  wire _abc_19068_n939_1_bF_buf3;
  wire _abc_19068_n939_1_bF_buf4;
  wire _abc_19068_n940_1;
  wire _abc_19068_n941;
  wire _abc_19068_n941_bF_buf0;
  wire _abc_19068_n941_bF_buf1;
  wire _abc_19068_n941_bF_buf2;
  wire _abc_19068_n941_bF_buf3;
  wire _abc_19068_n941_bF_buf4;
  wire _abc_19068_n942_1;
  wire _abc_19068_n943_1;
  wire _abc_19068_n944;
  wire _abc_19068_n945_1;
  wire _abc_19068_n945_1_bF_buf0;
  wire _abc_19068_n945_1_bF_buf1;
  wire _abc_19068_n945_1_bF_buf2;
  wire _abc_19068_n945_1_bF_buf3;
  wire _abc_19068_n945_1_bF_buf4;
  wire _abc_19068_n946_1;
  wire _abc_19068_n947;
  wire _abc_19068_n948_1;
  wire _abc_19068_n949_1;
  wire _abc_19068_n950;
  wire _abc_19068_n951_1;
  wire _abc_19068_n952_1;
  wire _abc_19068_n953;
  wire _abc_19068_n955_1;
  wire _abc_19068_n956;
  wire _abc_19068_n957_1;
  wire _abc_19068_n958_1;
  wire _abc_19068_n959;
  wire _abc_19068_n960_1;
  wire _abc_19068_n961_1;
  wire _abc_19068_n962;
  wire _abc_19068_n963_1;
  wire _abc_19068_n964_1;
  wire _abc_19068_n965;
  wire _abc_19068_n966_1;
  wire _abc_19068_n967_1;
  wire _abc_19068_n968;
  wire _abc_19068_n969_1;
  wire _abc_19068_n970_1;
  wire _abc_19068_n971;
  wire _abc_19068_n972_1;
  wire _abc_19068_n973_1;
  wire _abc_19068_n974;
  wire _abc_19068_n975_1;
  wire _abc_19068_n976_1;
  wire _abc_19068_n977;
  wire _abc_19068_n978_1;
  wire _abc_19068_n979_1;
  wire _abc_19068_n981_1;
  wire _abc_19068_n982_1;
  wire _abc_19068_n983;
  wire _abc_19068_n984_1;
  wire _abc_19068_n985_1;
  wire _abc_19068_n986;
  wire _abc_19068_n987_1;
  wire _abc_19068_n988_1;
  wire _abc_19068_n989;
  wire _abc_19068_n990_1;
  wire _abc_19068_n991_1;
  wire _abc_19068_n992;
  wire _abc_19068_n993_1;
  wire _abc_19068_n994_1;
  wire _abc_19068_n995;
  wire _abc_19068_n996_1;
  wire _abc_19068_n997_1;
  wire _abc_19068_n998;
  wire _abc_19068_n999_1;
  wire _auto_iopadmap_cc_313_execute_30317_0_;
  wire _auto_iopadmap_cc_313_execute_30317_10_;
  wire _auto_iopadmap_cc_313_execute_30317_11_;
  wire _auto_iopadmap_cc_313_execute_30317_12_;
  wire _auto_iopadmap_cc_313_execute_30317_13_;
  wire _auto_iopadmap_cc_313_execute_30317_14_;
  wire _auto_iopadmap_cc_313_execute_30317_15_;
  wire _auto_iopadmap_cc_313_execute_30317_16_;
  wire _auto_iopadmap_cc_313_execute_30317_17_;
  wire _auto_iopadmap_cc_313_execute_30317_18_;
  wire _auto_iopadmap_cc_313_execute_30317_19_;
  wire _auto_iopadmap_cc_313_execute_30317_1_;
  wire _auto_iopadmap_cc_313_execute_30317_20_;
  wire _auto_iopadmap_cc_313_execute_30317_21_;
  wire _auto_iopadmap_cc_313_execute_30317_22_;
  wire _auto_iopadmap_cc_313_execute_30317_23_;
  wire _auto_iopadmap_cc_313_execute_30317_24_;
  wire _auto_iopadmap_cc_313_execute_30317_25_;
  wire _auto_iopadmap_cc_313_execute_30317_26_;
  wire _auto_iopadmap_cc_313_execute_30317_27_;
  wire _auto_iopadmap_cc_313_execute_30317_28_;
  wire _auto_iopadmap_cc_313_execute_30317_29_;
  wire _auto_iopadmap_cc_313_execute_30317_2_;
  wire _auto_iopadmap_cc_313_execute_30317_30_;
  wire _auto_iopadmap_cc_313_execute_30317_31_;
  wire _auto_iopadmap_cc_313_execute_30317_3_;
  wire _auto_iopadmap_cc_313_execute_30317_4_;
  wire _auto_iopadmap_cc_313_execute_30317_5_;
  wire _auto_iopadmap_cc_313_execute_30317_6_;
  wire _auto_iopadmap_cc_313_execute_30317_7_;
  wire _auto_iopadmap_cc_313_execute_30317_8_;
  wire _auto_iopadmap_cc_313_execute_30317_9_;
  input \addr[0] ;
  input \addr[1] ;
  input \addr[2] ;
  input \addr[3] ;
  input \addr[4] ;
  input \addr[5] ;
  input \addr[6] ;
  input \addr[7] ;
  input clk;
  wire clk_bF_buf0;
  wire clk_bF_buf1;
  wire clk_bF_buf10;
  wire clk_bF_buf11;
  wire clk_bF_buf12;
  wire clk_bF_buf13;
  wire clk_bF_buf14;
  wire clk_bF_buf15;
  wire clk_bF_buf16;
  wire clk_bF_buf17;
  wire clk_bF_buf18;
  wire clk_bF_buf19;
  wire clk_bF_buf2;
  wire clk_bF_buf20;
  wire clk_bF_buf21;
  wire clk_bF_buf22;
  wire clk_bF_buf23;
  wire clk_bF_buf24;
  wire clk_bF_buf25;
  wire clk_bF_buf26;
  wire clk_bF_buf27;
  wire clk_bF_buf28;
  wire clk_bF_buf29;
  wire clk_bF_buf3;
  wire clk_bF_buf30;
  wire clk_bF_buf31;
  wire clk_bF_buf32;
  wire clk_bF_buf33;
  wire clk_bF_buf34;
  wire clk_bF_buf35;
  wire clk_bF_buf36;
  wire clk_bF_buf37;
  wire clk_bF_buf38;
  wire clk_bF_buf39;
  wire clk_bF_buf4;
  wire clk_bF_buf40;
  wire clk_bF_buf41;
  wire clk_bF_buf42;
  wire clk_bF_buf43;
  wire clk_bF_buf44;
  wire clk_bF_buf45;
  wire clk_bF_buf46;
  wire clk_bF_buf47;
  wire clk_bF_buf48;
  wire clk_bF_buf49;
  wire clk_bF_buf5;
  wire clk_bF_buf50;
  wire clk_bF_buf51;
  wire clk_bF_buf52;
  wire clk_bF_buf53;
  wire clk_bF_buf54;
  wire clk_bF_buf55;
  wire clk_bF_buf56;
  wire clk_bF_buf57;
  wire clk_bF_buf58;
  wire clk_bF_buf59;
  wire clk_bF_buf6;
  wire clk_bF_buf60;
  wire clk_bF_buf61;
  wire clk_bF_buf62;
  wire clk_bF_buf63;
  wire clk_bF_buf64;
  wire clk_bF_buf65;
  wire clk_bF_buf66;
  wire clk_bF_buf67;
  wire clk_bF_buf68;
  wire clk_bF_buf69;
  wire clk_bF_buf7;
  wire clk_bF_buf70;
  wire clk_bF_buf71;
  wire clk_bF_buf72;
  wire clk_bF_buf73;
  wire clk_bF_buf74;
  wire clk_bF_buf75;
  wire clk_bF_buf76;
  wire clk_bF_buf77;
  wire clk_bF_buf78;
  wire clk_bF_buf79;
  wire clk_bF_buf8;
  wire clk_bF_buf80;
  wire clk_bF_buf81;
  wire clk_bF_buf82;
  wire clk_bF_buf83;
  wire clk_bF_buf84;
  wire clk_bF_buf9;
  wire clk_hier0_bF_buf0;
  wire clk_hier0_bF_buf1;
  wire clk_hier0_bF_buf2;
  wire clk_hier0_bF_buf3;
  wire clk_hier0_bF_buf4;
  wire clk_hier0_bF_buf5;
  wire clk_hier0_bF_buf6;
  wire clk_hier0_bF_buf7;
  wire clk_hier0_bF_buf8;
  wire core__abc_14829_n1285;
  wire core__abc_14829_n1310;
  wire core__abc_14829_n1316;
  wire core__abc_14829_n1330;
  wire core__abc_14829_n6021;
  wire core__abc_14829_n6022;
  wire core__abc_14829_n6023;
  wire core__abc_14829_n6024;
  wire core__abc_21380_n10000;
  wire core__abc_21380_n10001;
  wire core__abc_21380_n10002;
  wire core__abc_21380_n10004;
  wire core__abc_21380_n10005;
  wire core__abc_21380_n10006;
  wire core__abc_21380_n10007;
  wire core__abc_21380_n10008;
  wire core__abc_21380_n10009;
  wire core__abc_21380_n10010;
  wire core__abc_21380_n10011;
  wire core__abc_21380_n10012;
  wire core__abc_21380_n10013;
  wire core__abc_21380_n10014;
  wire core__abc_21380_n10015;
  wire core__abc_21380_n10016;
  wire core__abc_21380_n10018;
  wire core__abc_21380_n10019;
  wire core__abc_21380_n10020;
  wire core__abc_21380_n10021;
  wire core__abc_21380_n10022;
  wire core__abc_21380_n10023;
  wire core__abc_21380_n10024;
  wire core__abc_21380_n10025;
  wire core__abc_21380_n10026;
  wire core__abc_21380_n10027;
  wire core__abc_21380_n10028;
  wire core__abc_21380_n10030;
  wire core__abc_21380_n10031;
  wire core__abc_21380_n10032;
  wire core__abc_21380_n10033;
  wire core__abc_21380_n10034;
  wire core__abc_21380_n10035;
  wire core__abc_21380_n10036;
  wire core__abc_21380_n10037;
  wire core__abc_21380_n10038;
  wire core__abc_21380_n10039;
  wire core__abc_21380_n10040;
  wire core__abc_21380_n10042;
  wire core__abc_21380_n10043;
  wire core__abc_21380_n10044;
  wire core__abc_21380_n10045;
  wire core__abc_21380_n10046;
  wire core__abc_21380_n10047;
  wire core__abc_21380_n10048;
  wire core__abc_21380_n10049;
  wire core__abc_21380_n10050;
  wire core__abc_21380_n10051;
  wire core__abc_21380_n10052;
  wire core__abc_21380_n10054;
  wire core__abc_21380_n10055;
  wire core__abc_21380_n10056;
  wire core__abc_21380_n10061;
  wire core__abc_21380_n10062;
  wire core__abc_21380_n10063;
  wire core__abc_21380_n10064;
  wire core__abc_21380_n1130_1;
  wire core__abc_21380_n1131;
  wire core__abc_21380_n1132_1;
  wire core__abc_21380_n1133_1;
  wire core__abc_21380_n1134_1;
  wire core__abc_21380_n1134_1_bF_buf0;
  wire core__abc_21380_n1134_1_bF_buf1;
  wire core__abc_21380_n1134_1_bF_buf2;
  wire core__abc_21380_n1134_1_bF_buf3;
  wire core__abc_21380_n1134_1_bF_buf4;
  wire core__abc_21380_n1134_1_bF_buf5;
  wire core__abc_21380_n1134_1_bF_buf6;
  wire core__abc_21380_n1134_1_bF_buf7;
  wire core__abc_21380_n1135;
  wire core__abc_21380_n1136_1;
  wire core__abc_21380_n1137_1;
  wire core__abc_21380_n1138_1;
  wire core__abc_21380_n1139;
  wire core__abc_21380_n1140_1;
  wire core__abc_21380_n1141_1;
  wire core__abc_21380_n1142_1;
  wire core__abc_21380_n1143;
  wire core__abc_21380_n1144_1;
  wire core__abc_21380_n1145_1;
  wire core__abc_21380_n1146_1;
  wire core__abc_21380_n1147;
  wire core__abc_21380_n1148_1;
  wire core__abc_21380_n1149_1;
  wire core__abc_21380_n1150_1;
  wire core__abc_21380_n1151;
  wire core__abc_21380_n1152_1;
  wire core__abc_21380_n1153_1;
  wire core__abc_21380_n1154_1;
  wire core__abc_21380_n1155;
  wire core__abc_21380_n1156_1;
  wire core__abc_21380_n1157_1;
  wire core__abc_21380_n1158_1;
  wire core__abc_21380_n1159;
  wire core__abc_21380_n1160_1;
  wire core__abc_21380_n1161_1;
  wire core__abc_21380_n1162_1;
  wire core__abc_21380_n1163;
  wire core__abc_21380_n1164_1;
  wire core__abc_21380_n1165_1;
  wire core__abc_21380_n1166_1;
  wire core__abc_21380_n1167;
  wire core__abc_21380_n1168_1;
  wire core__abc_21380_n1169_1;
  wire core__abc_21380_n1170_1;
  wire core__abc_21380_n1171;
  wire core__abc_21380_n1172_1;
  wire core__abc_21380_n1173_1;
  wire core__abc_21380_n1174_1;
  wire core__abc_21380_n1175;
  wire core__abc_21380_n1176_1;
  wire core__abc_21380_n1177_1;
  wire core__abc_21380_n1178_1;
  wire core__abc_21380_n1179;
  wire core__abc_21380_n1180_1;
  wire core__abc_21380_n1181_1;
  wire core__abc_21380_n1182_1;
  wire core__abc_21380_n1183;
  wire core__abc_21380_n1184_1;
  wire core__abc_21380_n1185_1;
  wire core__abc_21380_n1186_1;
  wire core__abc_21380_n1187;
  wire core__abc_21380_n1188_1;
  wire core__abc_21380_n1189_1;
  wire core__abc_21380_n1190_1;
  wire core__abc_21380_n1191;
  wire core__abc_21380_n1192_1;
  wire core__abc_21380_n1193_1;
  wire core__abc_21380_n1194_1;
  wire core__abc_21380_n1195;
  wire core__abc_21380_n1196_1;
  wire core__abc_21380_n1197_1;
  wire core__abc_21380_n1198_1;
  wire core__abc_21380_n1199;
  wire core__abc_21380_n1200_1;
  wire core__abc_21380_n1201_1;
  wire core__abc_21380_n1202_1;
  wire core__abc_21380_n1203;
  wire core__abc_21380_n1204_1;
  wire core__abc_21380_n1205_1;
  wire core__abc_21380_n1206_1;
  wire core__abc_21380_n1207;
  wire core__abc_21380_n1208_1;
  wire core__abc_21380_n1209_1;
  wire core__abc_21380_n1210_1;
  wire core__abc_21380_n1211;
  wire core__abc_21380_n1212_1;
  wire core__abc_21380_n1213_1;
  wire core__abc_21380_n1214_1;
  wire core__abc_21380_n1215;
  wire core__abc_21380_n1216_1;
  wire core__abc_21380_n1217_1;
  wire core__abc_21380_n1218_1;
  wire core__abc_21380_n1219;
  wire core__abc_21380_n1220_1;
  wire core__abc_21380_n1221_1;
  wire core__abc_21380_n1222_1;
  wire core__abc_21380_n1223;
  wire core__abc_21380_n1224_1;
  wire core__abc_21380_n1225_1;
  wire core__abc_21380_n1226_1;
  wire core__abc_21380_n1227;
  wire core__abc_21380_n1228_1;
  wire core__abc_21380_n1229_1;
  wire core__abc_21380_n1230_1;
  wire core__abc_21380_n1231;
  wire core__abc_21380_n1232_1;
  wire core__abc_21380_n1233_1;
  wire core__abc_21380_n1234_1;
  wire core__abc_21380_n1235;
  wire core__abc_21380_n1236_1;
  wire core__abc_21380_n1237_1;
  wire core__abc_21380_n1238_1;
  wire core__abc_21380_n1239;
  wire core__abc_21380_n1240_1;
  wire core__abc_21380_n1241_1;
  wire core__abc_21380_n1242_1;
  wire core__abc_21380_n1243;
  wire core__abc_21380_n1244_1;
  wire core__abc_21380_n1245_1;
  wire core__abc_21380_n1246_1;
  wire core__abc_21380_n1248_1;
  wire core__abc_21380_n1249_1;
  wire core__abc_21380_n1250_1;
  wire core__abc_21380_n1252_1;
  wire core__abc_21380_n1253_1;
  wire core__abc_21380_n1255;
  wire core__abc_21380_n1256_1;
  wire core__abc_21380_n1257_1;
  wire core__abc_21380_n1259;
  wire core__abc_21380_n1260_1;
  wire core__abc_21380_n1261_1;
  wire core__abc_21380_n1262_1;
  wire core__abc_21380_n1263;
  wire core__abc_21380_n1264_1;
  wire core__abc_21380_n1265_1;
  wire core__abc_21380_n1266_1;
  wire core__abc_21380_n1267;
  wire core__abc_21380_n1268_1;
  wire core__abc_21380_n1269_1;
  wire core__abc_21380_n1270_1;
  wire core__abc_21380_n1271;
  wire core__abc_21380_n1272_1;
  wire core__abc_21380_n1273_1;
  wire core__abc_21380_n1274_1;
  wire core__abc_21380_n1275;
  wire core__abc_21380_n1277_1;
  wire core__abc_21380_n1278_1;
  wire core__abc_21380_n1279;
  wire core__abc_21380_n1280_1;
  wire core__abc_21380_n1281_1;
  wire core__abc_21380_n1282_1;
  wire core__abc_21380_n1283;
  wire core__abc_21380_n1284_1;
  wire core__abc_21380_n1285_1;
  wire core__abc_21380_n1286_1;
  wire core__abc_21380_n1287;
  wire core__abc_21380_n1288_1;
  wire core__abc_21380_n1289;
  wire core__abc_21380_n1290;
  wire core__abc_21380_n1291;
  wire core__abc_21380_n1292;
  wire core__abc_21380_n1293;
  wire core__abc_21380_n1294;
  wire core__abc_21380_n1295;
  wire core__abc_21380_n1296;
  wire core__abc_21380_n1298;
  wire core__abc_21380_n1299;
  wire core__abc_21380_n1300;
  wire core__abc_21380_n1301;
  wire core__abc_21380_n1302;
  wire core__abc_21380_n1303;
  wire core__abc_21380_n1304;
  wire core__abc_21380_n1305;
  wire core__abc_21380_n1306;
  wire core__abc_21380_n1307;
  wire core__abc_21380_n1308;
  wire core__abc_21380_n1309;
  wire core__abc_21380_n1310;
  wire core__abc_21380_n1311;
  wire core__abc_21380_n1312;
  wire core__abc_21380_n1313;
  wire core__abc_21380_n1314;
  wire core__abc_21380_n1315;
  wire core__abc_21380_n1317;
  wire core__abc_21380_n1318;
  wire core__abc_21380_n1319;
  wire core__abc_21380_n1320;
  wire core__abc_21380_n1321;
  wire core__abc_21380_n1322;
  wire core__abc_21380_n1323;
  wire core__abc_21380_n1324;
  wire core__abc_21380_n1325;
  wire core__abc_21380_n1326;
  wire core__abc_21380_n1327;
  wire core__abc_21380_n1328;
  wire core__abc_21380_n1329;
  wire core__abc_21380_n1330;
  wire core__abc_21380_n1331;
  wire core__abc_21380_n1332;
  wire core__abc_21380_n1333;
  wire core__abc_21380_n1334;
  wire core__abc_21380_n1336;
  wire core__abc_21380_n1337;
  wire core__abc_21380_n1338;
  wire core__abc_21380_n1339;
  wire core__abc_21380_n1340;
  wire core__abc_21380_n1341;
  wire core__abc_21380_n1342;
  wire core__abc_21380_n1343;
  wire core__abc_21380_n1344;
  wire core__abc_21380_n1345;
  wire core__abc_21380_n1346;
  wire core__abc_21380_n1347;
  wire core__abc_21380_n1348;
  wire core__abc_21380_n1349;
  wire core__abc_21380_n1350;
  wire core__abc_21380_n1351;
  wire core__abc_21380_n1352;
  wire core__abc_21380_n1354;
  wire core__abc_21380_n1355;
  wire core__abc_21380_n1356;
  wire core__abc_21380_n1357;
  wire core__abc_21380_n1358;
  wire core__abc_21380_n1359;
  wire core__abc_21380_n1360;
  wire core__abc_21380_n1361;
  wire core__abc_21380_n1362;
  wire core__abc_21380_n1363;
  wire core__abc_21380_n1364;
  wire core__abc_21380_n1365;
  wire core__abc_21380_n1366;
  wire core__abc_21380_n1367;
  wire core__abc_21380_n1368;
  wire core__abc_21380_n1369;
  wire core__abc_21380_n1370;
  wire core__abc_21380_n1371;
  wire core__abc_21380_n1373;
  wire core__abc_21380_n1374;
  wire core__abc_21380_n1375;
  wire core__abc_21380_n1376;
  wire core__abc_21380_n1377;
  wire core__abc_21380_n1378;
  wire core__abc_21380_n1379;
  wire core__abc_21380_n1380;
  wire core__abc_21380_n1381;
  wire core__abc_21380_n1382;
  wire core__abc_21380_n1383;
  wire core__abc_21380_n1384;
  wire core__abc_21380_n1385;
  wire core__abc_21380_n1386;
  wire core__abc_21380_n1387;
  wire core__abc_21380_n1388;
  wire core__abc_21380_n1389;
  wire core__abc_21380_n1390;
  wire core__abc_21380_n1392;
  wire core__abc_21380_n1393;
  wire core__abc_21380_n1394;
  wire core__abc_21380_n1395;
  wire core__abc_21380_n1396;
  wire core__abc_21380_n1397;
  wire core__abc_21380_n1398;
  wire core__abc_21380_n1399;
  wire core__abc_21380_n1400;
  wire core__abc_21380_n1401;
  wire core__abc_21380_n1402;
  wire core__abc_21380_n1403;
  wire core__abc_21380_n1404;
  wire core__abc_21380_n1405;
  wire core__abc_21380_n1406;
  wire core__abc_21380_n1407;
  wire core__abc_21380_n1408;
  wire core__abc_21380_n1409;
  wire core__abc_21380_n1411;
  wire core__abc_21380_n1412;
  wire core__abc_21380_n1413;
  wire core__abc_21380_n1414;
  wire core__abc_21380_n1415;
  wire core__abc_21380_n1416;
  wire core__abc_21380_n1417;
  wire core__abc_21380_n1418;
  wire core__abc_21380_n1419;
  wire core__abc_21380_n1420;
  wire core__abc_21380_n1421;
  wire core__abc_21380_n1422;
  wire core__abc_21380_n1423;
  wire core__abc_21380_n1424;
  wire core__abc_21380_n1425;
  wire core__abc_21380_n1426;
  wire core__abc_21380_n1428;
  wire core__abc_21380_n1429;
  wire core__abc_21380_n1430;
  wire core__abc_21380_n1431;
  wire core__abc_21380_n1432;
  wire core__abc_21380_n1433;
  wire core__abc_21380_n1434;
  wire core__abc_21380_n1435;
  wire core__abc_21380_n1436;
  wire core__abc_21380_n1437;
  wire core__abc_21380_n1438;
  wire core__abc_21380_n1439;
  wire core__abc_21380_n1440;
  wire core__abc_21380_n1441;
  wire core__abc_21380_n1442;
  wire core__abc_21380_n1443;
  wire core__abc_21380_n1444;
  wire core__abc_21380_n1445;
  wire core__abc_21380_n1446;
  wire core__abc_21380_n1448;
  wire core__abc_21380_n1449;
  wire core__abc_21380_n1450;
  wire core__abc_21380_n1451;
  wire core__abc_21380_n1452;
  wire core__abc_21380_n1453;
  wire core__abc_21380_n1454;
  wire core__abc_21380_n1455;
  wire core__abc_21380_n1456;
  wire core__abc_21380_n1457;
  wire core__abc_21380_n1458;
  wire core__abc_21380_n1459;
  wire core__abc_21380_n1460;
  wire core__abc_21380_n1461;
  wire core__abc_21380_n1462;
  wire core__abc_21380_n1463;
  wire core__abc_21380_n1465;
  wire core__abc_21380_n1466;
  wire core__abc_21380_n1467;
  wire core__abc_21380_n1468;
  wire core__abc_21380_n1469;
  wire core__abc_21380_n1470;
  wire core__abc_21380_n1471;
  wire core__abc_21380_n1472;
  wire core__abc_21380_n1473;
  wire core__abc_21380_n1474;
  wire core__abc_21380_n1475;
  wire core__abc_21380_n1476;
  wire core__abc_21380_n1477;
  wire core__abc_21380_n1478;
  wire core__abc_21380_n1479;
  wire core__abc_21380_n1480;
  wire core__abc_21380_n1482;
  wire core__abc_21380_n1483;
  wire core__abc_21380_n1484;
  wire core__abc_21380_n1485;
  wire core__abc_21380_n1486;
  wire core__abc_21380_n1487;
  wire core__abc_21380_n1488;
  wire core__abc_21380_n1489;
  wire core__abc_21380_n1490;
  wire core__abc_21380_n1491;
  wire core__abc_21380_n1492;
  wire core__abc_21380_n1493;
  wire core__abc_21380_n1494;
  wire core__abc_21380_n1495;
  wire core__abc_21380_n1496;
  wire core__abc_21380_n1497;
  wire core__abc_21380_n1498;
  wire core__abc_21380_n1500;
  wire core__abc_21380_n1501;
  wire core__abc_21380_n1502;
  wire core__abc_21380_n1503;
  wire core__abc_21380_n1504;
  wire core__abc_21380_n1505;
  wire core__abc_21380_n1506;
  wire core__abc_21380_n1507;
  wire core__abc_21380_n1508;
  wire core__abc_21380_n1509;
  wire core__abc_21380_n1510;
  wire core__abc_21380_n1511;
  wire core__abc_21380_n1512;
  wire core__abc_21380_n1513;
  wire core__abc_21380_n1514;
  wire core__abc_21380_n1515;
  wire core__abc_21380_n1516;
  wire core__abc_21380_n1518;
  wire core__abc_21380_n1519;
  wire core__abc_21380_n1520;
  wire core__abc_21380_n1521;
  wire core__abc_21380_n1522;
  wire core__abc_21380_n1523;
  wire core__abc_21380_n1524;
  wire core__abc_21380_n1525;
  wire core__abc_21380_n1526;
  wire core__abc_21380_n1527;
  wire core__abc_21380_n1528;
  wire core__abc_21380_n1529;
  wire core__abc_21380_n1530;
  wire core__abc_21380_n1531;
  wire core__abc_21380_n1532;
  wire core__abc_21380_n1533;
  wire core__abc_21380_n1534;
  wire core__abc_21380_n1536;
  wire core__abc_21380_n1537;
  wire core__abc_21380_n1538;
  wire core__abc_21380_n1539;
  wire core__abc_21380_n1540;
  wire core__abc_21380_n1541;
  wire core__abc_21380_n1542;
  wire core__abc_21380_n1543;
  wire core__abc_21380_n1544;
  wire core__abc_21380_n1545;
  wire core__abc_21380_n1546;
  wire core__abc_21380_n1547;
  wire core__abc_21380_n1548;
  wire core__abc_21380_n1549;
  wire core__abc_21380_n1550;
  wire core__abc_21380_n1551;
  wire core__abc_21380_n1552;
  wire core__abc_21380_n1553;
  wire core__abc_21380_n1554;
  wire core__abc_21380_n1556;
  wire core__abc_21380_n1557;
  wire core__abc_21380_n1558;
  wire core__abc_21380_n1559;
  wire core__abc_21380_n1560;
  wire core__abc_21380_n1561;
  wire core__abc_21380_n1562;
  wire core__abc_21380_n1563;
  wire core__abc_21380_n1564;
  wire core__abc_21380_n1565;
  wire core__abc_21380_n1566;
  wire core__abc_21380_n1567;
  wire core__abc_21380_n1568;
  wire core__abc_21380_n1569;
  wire core__abc_21380_n1570;
  wire core__abc_21380_n1571;
  wire core__abc_21380_n1572;
  wire core__abc_21380_n1574;
  wire core__abc_21380_n1575;
  wire core__abc_21380_n1576;
  wire core__abc_21380_n1577;
  wire core__abc_21380_n1578;
  wire core__abc_21380_n1579;
  wire core__abc_21380_n1580;
  wire core__abc_21380_n1581;
  wire core__abc_21380_n1582;
  wire core__abc_21380_n1583;
  wire core__abc_21380_n1584;
  wire core__abc_21380_n1585;
  wire core__abc_21380_n1586;
  wire core__abc_21380_n1587;
  wire core__abc_21380_n1588;
  wire core__abc_21380_n1589;
  wire core__abc_21380_n1590;
  wire core__abc_21380_n1591;
  wire core__abc_21380_n1592;
  wire core__abc_21380_n1594;
  wire core__abc_21380_n1595;
  wire core__abc_21380_n1596;
  wire core__abc_21380_n1597;
  wire core__abc_21380_n1598;
  wire core__abc_21380_n1599;
  wire core__abc_21380_n1600;
  wire core__abc_21380_n1601;
  wire core__abc_21380_n1602;
  wire core__abc_21380_n1603;
  wire core__abc_21380_n1604;
  wire core__abc_21380_n1605;
  wire core__abc_21380_n1606;
  wire core__abc_21380_n1607;
  wire core__abc_21380_n1608;
  wire core__abc_21380_n1609;
  wire core__abc_21380_n1611;
  wire core__abc_21380_n1612;
  wire core__abc_21380_n1613;
  wire core__abc_21380_n1614;
  wire core__abc_21380_n1615;
  wire core__abc_21380_n1616;
  wire core__abc_21380_n1617;
  wire core__abc_21380_n1618;
  wire core__abc_21380_n1619;
  wire core__abc_21380_n1620;
  wire core__abc_21380_n1621;
  wire core__abc_21380_n1622;
  wire core__abc_21380_n1623;
  wire core__abc_21380_n1624;
  wire core__abc_21380_n1625;
  wire core__abc_21380_n1626;
  wire core__abc_21380_n1628;
  wire core__abc_21380_n1629;
  wire core__abc_21380_n1630;
  wire core__abc_21380_n1631;
  wire core__abc_21380_n1632;
  wire core__abc_21380_n1633;
  wire core__abc_21380_n1634;
  wire core__abc_21380_n1635;
  wire core__abc_21380_n1636;
  wire core__abc_21380_n1637;
  wire core__abc_21380_n1638;
  wire core__abc_21380_n1639;
  wire core__abc_21380_n1640;
  wire core__abc_21380_n1641;
  wire core__abc_21380_n1642;
  wire core__abc_21380_n1643;
  wire core__abc_21380_n1644;
  wire core__abc_21380_n1646;
  wire core__abc_21380_n1647;
  wire core__abc_21380_n1648;
  wire core__abc_21380_n1649_1;
  wire core__abc_21380_n1650;
  wire core__abc_21380_n1651;
  wire core__abc_21380_n1652;
  wire core__abc_21380_n1653;
  wire core__abc_21380_n1654;
  wire core__abc_21380_n1655_1;
  wire core__abc_21380_n1656;
  wire core__abc_21380_n1657;
  wire core__abc_21380_n1658;
  wire core__abc_21380_n1659;
  wire core__abc_21380_n1660;
  wire core__abc_21380_n1661;
  wire core__abc_21380_n1662;
  wire core__abc_21380_n1664;
  wire core__abc_21380_n1665;
  wire core__abc_21380_n1666;
  wire core__abc_21380_n1667;
  wire core__abc_21380_n1668;
  wire core__abc_21380_n1669;
  wire core__abc_21380_n1670;
  wire core__abc_21380_n1671;
  wire core__abc_21380_n1672;
  wire core__abc_21380_n1673;
  wire core__abc_21380_n1674;
  wire core__abc_21380_n1675;
  wire core__abc_21380_n1676;
  wire core__abc_21380_n1677;
  wire core__abc_21380_n1678;
  wire core__abc_21380_n1679;
  wire core__abc_21380_n1680;
  wire core__abc_21380_n1682;
  wire core__abc_21380_n1683;
  wire core__abc_21380_n1684;
  wire core__abc_21380_n1685;
  wire core__abc_21380_n1686;
  wire core__abc_21380_n1687;
  wire core__abc_21380_n1688;
  wire core__abc_21380_n1689;
  wire core__abc_21380_n1690;
  wire core__abc_21380_n1691;
  wire core__abc_21380_n1692;
  wire core__abc_21380_n1693;
  wire core__abc_21380_n1694;
  wire core__abc_21380_n1695;
  wire core__abc_21380_n1696;
  wire core__abc_21380_n1697;
  wire core__abc_21380_n1698;
  wire core__abc_21380_n1699;
  wire core__abc_21380_n1700;
  wire core__abc_21380_n1702;
  wire core__abc_21380_n1703;
  wire core__abc_21380_n1704;
  wire core__abc_21380_n1705;
  wire core__abc_21380_n1706;
  wire core__abc_21380_n1707;
  wire core__abc_21380_n1708;
  wire core__abc_21380_n1709;
  wire core__abc_21380_n1710;
  wire core__abc_21380_n1711;
  wire core__abc_21380_n1712;
  wire core__abc_21380_n1713;
  wire core__abc_21380_n1714;
  wire core__abc_21380_n1715;
  wire core__abc_21380_n1716;
  wire core__abc_21380_n1717;
  wire core__abc_21380_n1718;
  wire core__abc_21380_n1720;
  wire core__abc_21380_n1721;
  wire core__abc_21380_n1722;
  wire core__abc_21380_n1723;
  wire core__abc_21380_n1724;
  wire core__abc_21380_n1725;
  wire core__abc_21380_n1726;
  wire core__abc_21380_n1727;
  wire core__abc_21380_n1728;
  wire core__abc_21380_n1729;
  wire core__abc_21380_n1730;
  wire core__abc_21380_n1731;
  wire core__abc_21380_n1732;
  wire core__abc_21380_n1733;
  wire core__abc_21380_n1734;
  wire core__abc_21380_n1735;
  wire core__abc_21380_n1736;
  wire core__abc_21380_n1737;
  wire core__abc_21380_n1738;
  wire core__abc_21380_n1740;
  wire core__abc_21380_n1741;
  wire core__abc_21380_n1742;
  wire core__abc_21380_n1743;
  wire core__abc_21380_n1744;
  wire core__abc_21380_n1745;
  wire core__abc_21380_n1746;
  wire core__abc_21380_n1747;
  wire core__abc_21380_n1748;
  wire core__abc_21380_n1749;
  wire core__abc_21380_n1750;
  wire core__abc_21380_n1751;
  wire core__abc_21380_n1752;
  wire core__abc_21380_n1753;
  wire core__abc_21380_n1754_1;
  wire core__abc_21380_n1755;
  wire core__abc_21380_n1757;
  wire core__abc_21380_n1758;
  wire core__abc_21380_n1759;
  wire core__abc_21380_n1760_1;
  wire core__abc_21380_n1761;
  wire core__abc_21380_n1762;
  wire core__abc_21380_n1763;
  wire core__abc_21380_n1764;
  wire core__abc_21380_n1765;
  wire core__abc_21380_n1766;
  wire core__abc_21380_n1767;
  wire core__abc_21380_n1768;
  wire core__abc_21380_n1769;
  wire core__abc_21380_n1770;
  wire core__abc_21380_n1771;
  wire core__abc_21380_n1772;
  wire core__abc_21380_n1773;
  wire core__abc_21380_n1774;
  wire core__abc_21380_n1775;
  wire core__abc_21380_n1777;
  wire core__abc_21380_n1778;
  wire core__abc_21380_n1779;
  wire core__abc_21380_n1780;
  wire core__abc_21380_n1781;
  wire core__abc_21380_n1782_1;
  wire core__abc_21380_n1783;
  wire core__abc_21380_n1784;
  wire core__abc_21380_n1785;
  wire core__abc_21380_n1786_1;
  wire core__abc_21380_n1787;
  wire core__abc_21380_n1788;
  wire core__abc_21380_n1789;
  wire core__abc_21380_n1790;
  wire core__abc_21380_n1791;
  wire core__abc_21380_n1792;
  wire core__abc_21380_n1793;
  wire core__abc_21380_n1795;
  wire core__abc_21380_n1796;
  wire core__abc_21380_n1797;
  wire core__abc_21380_n1798;
  wire core__abc_21380_n1799;
  wire core__abc_21380_n1800;
  wire core__abc_21380_n1801;
  wire core__abc_21380_n1802;
  wire core__abc_21380_n1803;
  wire core__abc_21380_n1804;
  wire core__abc_21380_n1805;
  wire core__abc_21380_n1806;
  wire core__abc_21380_n1807;
  wire core__abc_21380_n1808;
  wire core__abc_21380_n1809;
  wire core__abc_21380_n1810;
  wire core__abc_21380_n1811;
  wire core__abc_21380_n1812_1;
  wire core__abc_21380_n1813;
  wire core__abc_21380_n1815;
  wire core__abc_21380_n1816_1;
  wire core__abc_21380_n1817;
  wire core__abc_21380_n1818;
  wire core__abc_21380_n1819;
  wire core__abc_21380_n1820;
  wire core__abc_21380_n1821;
  wire core__abc_21380_n1822;
  wire core__abc_21380_n1823;
  wire core__abc_21380_n1824;
  wire core__abc_21380_n1825;
  wire core__abc_21380_n1826;
  wire core__abc_21380_n1827;
  wire core__abc_21380_n1828;
  wire core__abc_21380_n1829;
  wire core__abc_21380_n1830;
  wire core__abc_21380_n1831;
  wire core__abc_21380_n1833;
  wire core__abc_21380_n1834;
  wire core__abc_21380_n1835;
  wire core__abc_21380_n1836;
  wire core__abc_21380_n1837;
  wire core__abc_21380_n1838;
  wire core__abc_21380_n1839;
  wire core__abc_21380_n1840;
  wire core__abc_21380_n1841;
  wire core__abc_21380_n1842;
  wire core__abc_21380_n1843;
  wire core__abc_21380_n1844;
  wire core__abc_21380_n1845;
  wire core__abc_21380_n1846_1;
  wire core__abc_21380_n1847;
  wire core__abc_21380_n1848;
  wire core__abc_21380_n1849;
  wire core__abc_21380_n1850;
  wire core__abc_21380_n1851;
  wire core__abc_21380_n1853;
  wire core__abc_21380_n1854;
  wire core__abc_21380_n1855;
  wire core__abc_21380_n1856;
  wire core__abc_21380_n1857;
  wire core__abc_21380_n1858;
  wire core__abc_21380_n1859;
  wire core__abc_21380_n1860;
  wire core__abc_21380_n1861;
  wire core__abc_21380_n1862;
  wire core__abc_21380_n1863;
  wire core__abc_21380_n1864;
  wire core__abc_21380_n1865;
  wire core__abc_21380_n1866;
  wire core__abc_21380_n1867;
  wire core__abc_21380_n1868;
  wire core__abc_21380_n1869;
  wire core__abc_21380_n1871;
  wire core__abc_21380_n1872;
  wire core__abc_21380_n1873;
  wire core__abc_21380_n1874;
  wire core__abc_21380_n1875;
  wire core__abc_21380_n1876;
  wire core__abc_21380_n1877;
  wire core__abc_21380_n1878;
  wire core__abc_21380_n1879;
  wire core__abc_21380_n1880;
  wire core__abc_21380_n1881;
  wire core__abc_21380_n1882;
  wire core__abc_21380_n1883;
  wire core__abc_21380_n1884;
  wire core__abc_21380_n1885;
  wire core__abc_21380_n1886;
  wire core__abc_21380_n1887;
  wire core__abc_21380_n1889;
  wire core__abc_21380_n1890;
  wire core__abc_21380_n1891;
  wire core__abc_21380_n1892;
  wire core__abc_21380_n1893;
  wire core__abc_21380_n1894_1;
  wire core__abc_21380_n1895;
  wire core__abc_21380_n1896;
  wire core__abc_21380_n1897;
  wire core__abc_21380_n1898;
  wire core__abc_21380_n1899;
  wire core__abc_21380_n1900;
  wire core__abc_21380_n1901;
  wire core__abc_21380_n1902;
  wire core__abc_21380_n1903;
  wire core__abc_21380_n1904;
  wire core__abc_21380_n1905;
  wire core__abc_21380_n1907;
  wire core__abc_21380_n1908;
  wire core__abc_21380_n1909;
  wire core__abc_21380_n1910;
  wire core__abc_21380_n1911;
  wire core__abc_21380_n1912;
  wire core__abc_21380_n1913;
  wire core__abc_21380_n1914;
  wire core__abc_21380_n1915;
  wire core__abc_21380_n1916;
  wire core__abc_21380_n1917;
  wire core__abc_21380_n1918;
  wire core__abc_21380_n1919;
  wire core__abc_21380_n1920;
  wire core__abc_21380_n1921;
  wire core__abc_21380_n1922;
  wire core__abc_21380_n1923;
  wire core__abc_21380_n1924;
  wire core__abc_21380_n1925;
  wire core__abc_21380_n1927;
  wire core__abc_21380_n1928_1;
  wire core__abc_21380_n1929;
  wire core__abc_21380_n1930;
  wire core__abc_21380_n1931;
  wire core__abc_21380_n1932;
  wire core__abc_21380_n1933;
  wire core__abc_21380_n1934_1;
  wire core__abc_21380_n1935;
  wire core__abc_21380_n1936;
  wire core__abc_21380_n1937;
  wire core__abc_21380_n1938;
  wire core__abc_21380_n1939;
  wire core__abc_21380_n1940;
  wire core__abc_21380_n1941;
  wire core__abc_21380_n1942;
  wire core__abc_21380_n1943;
  wire core__abc_21380_n1945;
  wire core__abc_21380_n1946;
  wire core__abc_21380_n1947;
  wire core__abc_21380_n1948;
  wire core__abc_21380_n1949;
  wire core__abc_21380_n1950;
  wire core__abc_21380_n1951;
  wire core__abc_21380_n1952;
  wire core__abc_21380_n1953;
  wire core__abc_21380_n1954;
  wire core__abc_21380_n1955;
  wire core__abc_21380_n1956;
  wire core__abc_21380_n1957;
  wire core__abc_21380_n1958;
  wire core__abc_21380_n1959;
  wire core__abc_21380_n1960;
  wire core__abc_21380_n1961_1;
  wire core__abc_21380_n1962;
  wire core__abc_21380_n1963;
  wire core__abc_21380_n1965_1;
  wire core__abc_21380_n1966;
  wire core__abc_21380_n1967;
  wire core__abc_21380_n1968;
  wire core__abc_21380_n1969;
  wire core__abc_21380_n1970;
  wire core__abc_21380_n1971;
  wire core__abc_21380_n1972;
  wire core__abc_21380_n1973;
  wire core__abc_21380_n1974;
  wire core__abc_21380_n1975;
  wire core__abc_21380_n1976;
  wire core__abc_21380_n1977;
  wire core__abc_21380_n1978;
  wire core__abc_21380_n1979;
  wire core__abc_21380_n1980;
  wire core__abc_21380_n1981;
  wire core__abc_21380_n1983;
  wire core__abc_21380_n1984;
  wire core__abc_21380_n1985;
  wire core__abc_21380_n1986;
  wire core__abc_21380_n1987;
  wire core__abc_21380_n1988;
  wire core__abc_21380_n1989;
  wire core__abc_21380_n1990;
  wire core__abc_21380_n1991;
  wire core__abc_21380_n1992;
  wire core__abc_21380_n1993;
  wire core__abc_21380_n1994;
  wire core__abc_21380_n1995_1;
  wire core__abc_21380_n1996;
  wire core__abc_21380_n1997;
  wire core__abc_21380_n1998;
  wire core__abc_21380_n1999;
  wire core__abc_21380_n2000;
  wire core__abc_21380_n2001_1;
  wire core__abc_21380_n2003;
  wire core__abc_21380_n2004;
  wire core__abc_21380_n2005;
  wire core__abc_21380_n2006;
  wire core__abc_21380_n2007;
  wire core__abc_21380_n2008;
  wire core__abc_21380_n2009;
  wire core__abc_21380_n2010;
  wire core__abc_21380_n2011;
  wire core__abc_21380_n2012;
  wire core__abc_21380_n2013;
  wire core__abc_21380_n2014;
  wire core__abc_21380_n2015;
  wire core__abc_21380_n2016;
  wire core__abc_21380_n2017;
  wire core__abc_21380_n2018;
  wire core__abc_21380_n2019;
  wire core__abc_21380_n2021;
  wire core__abc_21380_n2022;
  wire core__abc_21380_n2023;
  wire core__abc_21380_n2024;
  wire core__abc_21380_n2025;
  wire core__abc_21380_n2026;
  wire core__abc_21380_n2027;
  wire core__abc_21380_n2028;
  wire core__abc_21380_n2029;
  wire core__abc_21380_n2030;
  wire core__abc_21380_n2031;
  wire core__abc_21380_n2032;
  wire core__abc_21380_n2033;
  wire core__abc_21380_n2034;
  wire core__abc_21380_n2035_1;
  wire core__abc_21380_n2036;
  wire core__abc_21380_n2037;
  wire core__abc_21380_n2039_1;
  wire core__abc_21380_n2040;
  wire core__abc_21380_n2041;
  wire core__abc_21380_n2042;
  wire core__abc_21380_n2043;
  wire core__abc_21380_n2044;
  wire core__abc_21380_n2045;
  wire core__abc_21380_n2046;
  wire core__abc_21380_n2047;
  wire core__abc_21380_n2048;
  wire core__abc_21380_n2049;
  wire core__abc_21380_n2050;
  wire core__abc_21380_n2051;
  wire core__abc_21380_n2052;
  wire core__abc_21380_n2053;
  wire core__abc_21380_n2054;
  wire core__abc_21380_n2055;
  wire core__abc_21380_n2057;
  wire core__abc_21380_n2058;
  wire core__abc_21380_n2059;
  wire core__abc_21380_n2060;
  wire core__abc_21380_n2061;
  wire core__abc_21380_n2062;
  wire core__abc_21380_n2063;
  wire core__abc_21380_n2064;
  wire core__abc_21380_n2065;
  wire core__abc_21380_n2066;
  wire core__abc_21380_n2067_1;
  wire core__abc_21380_n2068;
  wire core__abc_21380_n2069;
  wire core__abc_21380_n2070;
  wire core__abc_21380_n2071;
  wire core__abc_21380_n2072;
  wire core__abc_21380_n2073_1;
  wire core__abc_21380_n2074;
  wire core__abc_21380_n2075;
  wire core__abc_21380_n2077;
  wire core__abc_21380_n2078;
  wire core__abc_21380_n2079;
  wire core__abc_21380_n2080;
  wire core__abc_21380_n2081;
  wire core__abc_21380_n2082;
  wire core__abc_21380_n2083;
  wire core__abc_21380_n2084;
  wire core__abc_21380_n2085;
  wire core__abc_21380_n2086;
  wire core__abc_21380_n2087;
  wire core__abc_21380_n2088;
  wire core__abc_21380_n2089;
  wire core__abc_21380_n2090;
  wire core__abc_21380_n2091;
  wire core__abc_21380_n2092;
  wire core__abc_21380_n2093;
  wire core__abc_21380_n2095;
  wire core__abc_21380_n2096;
  wire core__abc_21380_n2097;
  wire core__abc_21380_n2098;
  wire core__abc_21380_n2099_1;
  wire core__abc_21380_n2100;
  wire core__abc_21380_n2101;
  wire core__abc_21380_n2102;
  wire core__abc_21380_n2103_1;
  wire core__abc_21380_n2104;
  wire core__abc_21380_n2105;
  wire core__abc_21380_n2106;
  wire core__abc_21380_n2107;
  wire core__abc_21380_n2108;
  wire core__abc_21380_n2109;
  wire core__abc_21380_n2110;
  wire core__abc_21380_n2111;
  wire core__abc_21380_n2112;
  wire core__abc_21380_n2113;
  wire core__abc_21380_n2115;
  wire core__abc_21380_n2116;
  wire core__abc_21380_n2117;
  wire core__abc_21380_n2118;
  wire core__abc_21380_n2119;
  wire core__abc_21380_n2120;
  wire core__abc_21380_n2121;
  wire core__abc_21380_n2122;
  wire core__abc_21380_n2123;
  wire core__abc_21380_n2124;
  wire core__abc_21380_n2125;
  wire core__abc_21380_n2126;
  wire core__abc_21380_n2127;
  wire core__abc_21380_n2128;
  wire core__abc_21380_n2129;
  wire core__abc_21380_n2130;
  wire core__abc_21380_n2131;
  wire core__abc_21380_n2133;
  wire core__abc_21380_n2134;
  wire core__abc_21380_n2135;
  wire core__abc_21380_n2136;
  wire core__abc_21380_n2137;
  wire core__abc_21380_n2138;
  wire core__abc_21380_n2139_1;
  wire core__abc_21380_n2140;
  wire core__abc_21380_n2141;
  wire core__abc_21380_n2142;
  wire core__abc_21380_n2143_1;
  wire core__abc_21380_n2144;
  wire core__abc_21380_n2145;
  wire core__abc_21380_n2146;
  wire core__abc_21380_n2147;
  wire core__abc_21380_n2148;
  wire core__abc_21380_n2149;
  wire core__abc_21380_n2150;
  wire core__abc_21380_n2151;
  wire core__abc_21380_n2153;
  wire core__abc_21380_n2154;
  wire core__abc_21380_n2155;
  wire core__abc_21380_n2156;
  wire core__abc_21380_n2157;
  wire core__abc_21380_n2158;
  wire core__abc_21380_n2159;
  wire core__abc_21380_n2160;
  wire core__abc_21380_n2161;
  wire core__abc_21380_n2162;
  wire core__abc_21380_n2163;
  wire core__abc_21380_n2164;
  wire core__abc_21380_n2165;
  wire core__abc_21380_n2166;
  wire core__abc_21380_n2167;
  wire core__abc_21380_n2168;
  wire core__abc_21380_n2169;
  wire core__abc_21380_n2171;
  wire core__abc_21380_n2172;
  wire core__abc_21380_n2173;
  wire core__abc_21380_n2174;
  wire core__abc_21380_n2175;
  wire core__abc_21380_n2176;
  wire core__abc_21380_n2177;
  wire core__abc_21380_n2178;
  wire core__abc_21380_n2179_1;
  wire core__abc_21380_n2180;
  wire core__abc_21380_n2181;
  wire core__abc_21380_n2182;
  wire core__abc_21380_n2183;
  wire core__abc_21380_n2184;
  wire core__abc_21380_n2185_1;
  wire core__abc_21380_n2186;
  wire core__abc_21380_n2187;
  wire core__abc_21380_n2189;
  wire core__abc_21380_n2190;
  wire core__abc_21380_n2191;
  wire core__abc_21380_n2192;
  wire core__abc_21380_n2193;
  wire core__abc_21380_n2194;
  wire core__abc_21380_n2195;
  wire core__abc_21380_n2196;
  wire core__abc_21380_n2197;
  wire core__abc_21380_n2198;
  wire core__abc_21380_n2199;
  wire core__abc_21380_n2200;
  wire core__abc_21380_n2201;
  wire core__abc_21380_n2202;
  wire core__abc_21380_n2203;
  wire core__abc_21380_n2204;
  wire core__abc_21380_n2205;
  wire core__abc_21380_n2207;
  wire core__abc_21380_n2208;
  wire core__abc_21380_n2209;
  wire core__abc_21380_n2210;
  wire core__abc_21380_n2211;
  wire core__abc_21380_n2212;
  wire core__abc_21380_n2213_1;
  wire core__abc_21380_n2214;
  wire core__abc_21380_n2215;
  wire core__abc_21380_n2216;
  wire core__abc_21380_n2217;
  wire core__abc_21380_n2218;
  wire core__abc_21380_n2219_1;
  wire core__abc_21380_n2220;
  wire core__abc_21380_n2221;
  wire core__abc_21380_n2222;
  wire core__abc_21380_n2223;
  wire core__abc_21380_n2224;
  wire core__abc_21380_n2225;
  wire core__abc_21380_n2227;
  wire core__abc_21380_n2228;
  wire core__abc_21380_n2229;
  wire core__abc_21380_n2230;
  wire core__abc_21380_n2231;
  wire core__abc_21380_n2232;
  wire core__abc_21380_n2233;
  wire core__abc_21380_n2234;
  wire core__abc_21380_n2235;
  wire core__abc_21380_n2236;
  wire core__abc_21380_n2237;
  wire core__abc_21380_n2238;
  wire core__abc_21380_n2239;
  wire core__abc_21380_n2240;
  wire core__abc_21380_n2241;
  wire core__abc_21380_n2242;
  wire core__abc_21380_n2244;
  wire core__abc_21380_n2245;
  wire core__abc_21380_n2246;
  wire core__abc_21380_n2247_1;
  wire core__abc_21380_n2248;
  wire core__abc_21380_n2249;
  wire core__abc_21380_n2250;
  wire core__abc_21380_n2251;
  wire core__abc_21380_n2252;
  wire core__abc_21380_n2253;
  wire core__abc_21380_n2254;
  wire core__abc_21380_n2255;
  wire core__abc_21380_n2256;
  wire core__abc_21380_n2257;
  wire core__abc_21380_n2258;
  wire core__abc_21380_n2259;
  wire core__abc_21380_n2260;
  wire core__abc_21380_n2261;
  wire core__abc_21380_n2262;
  wire core__abc_21380_n2264;
  wire core__abc_21380_n2265;
  wire core__abc_21380_n2266;
  wire core__abc_21380_n2267;
  wire core__abc_21380_n2268;
  wire core__abc_21380_n2269;
  wire core__abc_21380_n2270;
  wire core__abc_21380_n2271;
  wire core__abc_21380_n2272;
  wire core__abc_21380_n2273;
  wire core__abc_21380_n2274;
  wire core__abc_21380_n2275;
  wire core__abc_21380_n2276;
  wire core__abc_21380_n2277;
  wire core__abc_21380_n2278;
  wire core__abc_21380_n2279;
  wire core__abc_21380_n2280;
  wire core__abc_21380_n2282;
  wire core__abc_21380_n2283;
  wire core__abc_21380_n2284;
  wire core__abc_21380_n2285;
  wire core__abc_21380_n2286;
  wire core__abc_21380_n2287;
  wire core__abc_21380_n2288;
  wire core__abc_21380_n2289;
  wire core__abc_21380_n2290;
  wire core__abc_21380_n2291;
  wire core__abc_21380_n2292;
  wire core__abc_21380_n2293;
  wire core__abc_21380_n2294_1;
  wire core__abc_21380_n2295;
  wire core__abc_21380_n2296;
  wire core__abc_21380_n2297;
  wire core__abc_21380_n2298_1;
  wire core__abc_21380_n2299;
  wire core__abc_21380_n2300;
  wire core__abc_21380_n2302;
  wire core__abc_21380_n2303;
  wire core__abc_21380_n2304;
  wire core__abc_21380_n2305;
  wire core__abc_21380_n2306;
  wire core__abc_21380_n2307;
  wire core__abc_21380_n2308;
  wire core__abc_21380_n2309;
  wire core__abc_21380_n2310;
  wire core__abc_21380_n2311;
  wire core__abc_21380_n2312;
  wire core__abc_21380_n2313;
  wire core__abc_21380_n2314;
  wire core__abc_21380_n2315;
  wire core__abc_21380_n2316;
  wire core__abc_21380_n2317;
  wire core__abc_21380_n2318;
  wire core__abc_21380_n2320;
  wire core__abc_21380_n2321;
  wire core__abc_21380_n2322;
  wire core__abc_21380_n2323;
  wire core__abc_21380_n2324;
  wire core__abc_21380_n2325;
  wire core__abc_21380_n2326;
  wire core__abc_21380_n2327;
  wire core__abc_21380_n2328_1;
  wire core__abc_21380_n2329;
  wire core__abc_21380_n2330;
  wire core__abc_21380_n2331;
  wire core__abc_21380_n2332_1;
  wire core__abc_21380_n2333;
  wire core__abc_21380_n2334;
  wire core__abc_21380_n2335;
  wire core__abc_21380_n2336;
  wire core__abc_21380_n2338;
  wire core__abc_21380_n2339;
  wire core__abc_21380_n2340;
  wire core__abc_21380_n2341;
  wire core__abc_21380_n2342;
  wire core__abc_21380_n2343;
  wire core__abc_21380_n2344;
  wire core__abc_21380_n2345;
  wire core__abc_21380_n2346;
  wire core__abc_21380_n2347;
  wire core__abc_21380_n2348;
  wire core__abc_21380_n2349;
  wire core__abc_21380_n2350;
  wire core__abc_21380_n2351;
  wire core__abc_21380_n2352;
  wire core__abc_21380_n2353;
  wire core__abc_21380_n2354;
  wire core__abc_21380_n2356;
  wire core__abc_21380_n2357;
  wire core__abc_21380_n2358;
  wire core__abc_21380_n2359;
  wire core__abc_21380_n2360;
  wire core__abc_21380_n2361;
  wire core__abc_21380_n2362;
  wire core__abc_21380_n2363_1;
  wire core__abc_21380_n2364;
  wire core__abc_21380_n2365;
  wire core__abc_21380_n2366;
  wire core__abc_21380_n2367;
  wire core__abc_21380_n2368;
  wire core__abc_21380_n2369_1;
  wire core__abc_21380_n2370;
  wire core__abc_21380_n2371;
  wire core__abc_21380_n2372;
  wire core__abc_21380_n2373;
  wire core__abc_21380_n2374;
  wire core__abc_21380_n2376;
  wire core__abc_21380_n2377;
  wire core__abc_21380_n2378;
  wire core__abc_21380_n2379;
  wire core__abc_21380_n2380;
  wire core__abc_21380_n2381;
  wire core__abc_21380_n2382;
  wire core__abc_21380_n2383;
  wire core__abc_21380_n2384;
  wire core__abc_21380_n2385;
  wire core__abc_21380_n2386;
  wire core__abc_21380_n2387;
  wire core__abc_21380_n2388;
  wire core__abc_21380_n2389;
  wire core__abc_21380_n2390;
  wire core__abc_21380_n2391_1;
  wire core__abc_21380_n2392;
  wire core__abc_21380_n2394;
  wire core__abc_21380_n2395_1;
  wire core__abc_21380_n2396;
  wire core__abc_21380_n2397;
  wire core__abc_21380_n2398;
  wire core__abc_21380_n2399;
  wire core__abc_21380_n2400;
  wire core__abc_21380_n2401;
  wire core__abc_21380_n2402;
  wire core__abc_21380_n2403;
  wire core__abc_21380_n2404;
  wire core__abc_21380_n2405;
  wire core__abc_21380_n2406;
  wire core__abc_21380_n2407;
  wire core__abc_21380_n2408;
  wire core__abc_21380_n2409;
  wire core__abc_21380_n2410;
  wire core__abc_21380_n2412;
  wire core__abc_21380_n2413;
  wire core__abc_21380_n2414;
  wire core__abc_21380_n2415;
  wire core__abc_21380_n2416;
  wire core__abc_21380_n2417;
  wire core__abc_21380_n2418;
  wire core__abc_21380_n2419;
  wire core__abc_21380_n2420;
  wire core__abc_21380_n2421;
  wire core__abc_21380_n2422;
  wire core__abc_21380_n2423;
  wire core__abc_21380_n2424_1;
  wire core__abc_21380_n2425;
  wire core__abc_21380_n2426;
  wire core__abc_21380_n2427;
  wire core__abc_21380_n2428;
  wire core__abc_21380_n2430_1;
  wire core__abc_21380_n2431;
  wire core__abc_21380_n2432;
  wire core__abc_21380_n2433;
  wire core__abc_21380_n2434;
  wire core__abc_21380_n2435;
  wire core__abc_21380_n2436;
  wire core__abc_21380_n2437;
  wire core__abc_21380_n2438;
  wire core__abc_21380_n2439;
  wire core__abc_21380_n2440;
  wire core__abc_21380_n2441;
  wire core__abc_21380_n2442;
  wire core__abc_21380_n2443;
  wire core__abc_21380_n2444;
  wire core__abc_21380_n2445_1;
  wire core__abc_21380_n2446;
  wire core__abc_21380_n2448;
  wire core__abc_21380_n2449;
  wire core__abc_21380_n2450;
  wire core__abc_21380_n2451_1;
  wire core__abc_21380_n2451_1_bF_buf0;
  wire core__abc_21380_n2451_1_bF_buf1;
  wire core__abc_21380_n2451_1_bF_buf2;
  wire core__abc_21380_n2451_1_bF_buf3;
  wire core__abc_21380_n2451_1_bF_buf4;
  wire core__abc_21380_n2451_1_bF_buf5;
  wire core__abc_21380_n2451_1_bF_buf6;
  wire core__abc_21380_n2451_1_bF_buf7;
  wire core__abc_21380_n2452;
  wire core__abc_21380_n2452_bF_buf0;
  wire core__abc_21380_n2452_bF_buf1;
  wire core__abc_21380_n2452_bF_buf2;
  wire core__abc_21380_n2452_bF_buf3;
  wire core__abc_21380_n2452_bF_buf4;
  wire core__abc_21380_n2452_bF_buf5;
  wire core__abc_21380_n2452_bF_buf6;
  wire core__abc_21380_n2452_bF_buf7;
  wire core__abc_21380_n2453;
  wire core__abc_21380_n2454;
  wire core__abc_21380_n2455;
  wire core__abc_21380_n2457;
  wire core__abc_21380_n2458;
  wire core__abc_21380_n2459;
  wire core__abc_21380_n2461;
  wire core__abc_21380_n2462;
  wire core__abc_21380_n2463;
  wire core__abc_21380_n2465;
  wire core__abc_21380_n2466;
  wire core__abc_21380_n2467;
  wire core__abc_21380_n2469;
  wire core__abc_21380_n2470;
  wire core__abc_21380_n2471_1;
  wire core__abc_21380_n2473;
  wire core__abc_21380_n2474;
  wire core__abc_21380_n2475;
  wire core__abc_21380_n2477_1;
  wire core__abc_21380_n2478;
  wire core__abc_21380_n2479;
  wire core__abc_21380_n2481;
  wire core__abc_21380_n2482;
  wire core__abc_21380_n2483;
  wire core__abc_21380_n2485;
  wire core__abc_21380_n2486;
  wire core__abc_21380_n2487;
  wire core__abc_21380_n2489;
  wire core__abc_21380_n2490;
  wire core__abc_21380_n2491;
  wire core__abc_21380_n2493_1;
  wire core__abc_21380_n2494;
  wire core__abc_21380_n2495;
  wire core__abc_21380_n2497_1;
  wire core__abc_21380_n2498;
  wire core__abc_21380_n2499;
  wire core__abc_21380_n2501;
  wire core__abc_21380_n2502;
  wire core__abc_21380_n2503;
  wire core__abc_21380_n2505;
  wire core__abc_21380_n2506;
  wire core__abc_21380_n2507;
  wire core__abc_21380_n2509;
  wire core__abc_21380_n2510;
  wire core__abc_21380_n2511;
  wire core__abc_21380_n2513;
  wire core__abc_21380_n2514;
  wire core__abc_21380_n2515;
  wire core__abc_21380_n2517;
  wire core__abc_21380_n2518;
  wire core__abc_21380_n2519;
  wire core__abc_21380_n2521;
  wire core__abc_21380_n2522;
  wire core__abc_21380_n2523;
  wire core__abc_21380_n2525;
  wire core__abc_21380_n2526;
  wire core__abc_21380_n2527;
  wire core__abc_21380_n2529;
  wire core__abc_21380_n2530;
  wire core__abc_21380_n2531;
  wire core__abc_21380_n2533;
  wire core__abc_21380_n2534_1;
  wire core__abc_21380_n2535;
  wire core__abc_21380_n2537;
  wire core__abc_21380_n2538;
  wire core__abc_21380_n2539;
  wire core__abc_21380_n2541;
  wire core__abc_21380_n2542;
  wire core__abc_21380_n2543;
  wire core__abc_21380_n2545;
  wire core__abc_21380_n2546;
  wire core__abc_21380_n2547;
  wire core__abc_21380_n2549;
  wire core__abc_21380_n2550;
  wire core__abc_21380_n2551_1;
  wire core__abc_21380_n2553;
  wire core__abc_21380_n2554;
  wire core__abc_21380_n2555_1;
  wire core__abc_21380_n2557;
  wire core__abc_21380_n2558;
  wire core__abc_21380_n2559;
  wire core__abc_21380_n2561;
  wire core__abc_21380_n2562;
  wire core__abc_21380_n2563;
  wire core__abc_21380_n2565;
  wire core__abc_21380_n2566;
  wire core__abc_21380_n2567;
  wire core__abc_21380_n2569;
  wire core__abc_21380_n2570;
  wire core__abc_21380_n2571;
  wire core__abc_21380_n2573;
  wire core__abc_21380_n2574;
  wire core__abc_21380_n2575;
  wire core__abc_21380_n2577;
  wire core__abc_21380_n2578_1;
  wire core__abc_21380_n2579;
  wire core__abc_21380_n2581;
  wire core__abc_21380_n2582_1;
  wire core__abc_21380_n2583;
  wire core__abc_21380_n2585;
  wire core__abc_21380_n2586;
  wire core__abc_21380_n2587;
  wire core__abc_21380_n2589;
  wire core__abc_21380_n2590;
  wire core__abc_21380_n2591;
  wire core__abc_21380_n2593;
  wire core__abc_21380_n2594;
  wire core__abc_21380_n2595;
  wire core__abc_21380_n2597_1;
  wire core__abc_21380_n2598;
  wire core__abc_21380_n2599;
  wire core__abc_21380_n2601;
  wire core__abc_21380_n2602;
  wire core__abc_21380_n2603_1;
  wire core__abc_21380_n2605;
  wire core__abc_21380_n2606;
  wire core__abc_21380_n2607;
  wire core__abc_21380_n2609;
  wire core__abc_21380_n2610;
  wire core__abc_21380_n2611;
  wire core__abc_21380_n2613;
  wire core__abc_21380_n2614;
  wire core__abc_21380_n2615;
  wire core__abc_21380_n2617;
  wire core__abc_21380_n2618;
  wire core__abc_21380_n2619;
  wire core__abc_21380_n2621;
  wire core__abc_21380_n2622;
  wire core__abc_21380_n2623;
  wire core__abc_21380_n2625;
  wire core__abc_21380_n2626;
  wire core__abc_21380_n2627_1;
  wire core__abc_21380_n2629;
  wire core__abc_21380_n2630;
  wire core__abc_21380_n2631;
  wire core__abc_21380_n2633_1;
  wire core__abc_21380_n2634;
  wire core__abc_21380_n2635;
  wire core__abc_21380_n2637;
  wire core__abc_21380_n2638;
  wire core__abc_21380_n2639;
  wire core__abc_21380_n2641;
  wire core__abc_21380_n2642;
  wire core__abc_21380_n2643;
  wire core__abc_21380_n2645;
  wire core__abc_21380_n2646;
  wire core__abc_21380_n2647;
  wire core__abc_21380_n2649;
  wire core__abc_21380_n2650;
  wire core__abc_21380_n2651;
  wire core__abc_21380_n2653;
  wire core__abc_21380_n2654_1;
  wire core__abc_21380_n2655;
  wire core__abc_21380_n2657;
  wire core__abc_21380_n2658;
  wire core__abc_21380_n2659;
  wire core__abc_21380_n2661;
  wire core__abc_21380_n2662;
  wire core__abc_21380_n2663;
  wire core__abc_21380_n2665;
  wire core__abc_21380_n2666;
  wire core__abc_21380_n2667;
  wire core__abc_21380_n2669;
  wire core__abc_21380_n2670;
  wire core__abc_21380_n2671;
  wire core__abc_21380_n2673;
  wire core__abc_21380_n2674;
  wire core__abc_21380_n2675;
  wire core__abc_21380_n2677;
  wire core__abc_21380_n2678;
  wire core__abc_21380_n2679;
  wire core__abc_21380_n2681;
  wire core__abc_21380_n2682_1;
  wire core__abc_21380_n2683;
  wire core__abc_21380_n2685;
  wire core__abc_21380_n2686;
  wire core__abc_21380_n2687;
  wire core__abc_21380_n2689;
  wire core__abc_21380_n2690;
  wire core__abc_21380_n2691;
  wire core__abc_21380_n2693;
  wire core__abc_21380_n2694;
  wire core__abc_21380_n2695;
  wire core__abc_21380_n2697;
  wire core__abc_21380_n2698;
  wire core__abc_21380_n2699;
  wire core__abc_21380_n2701;
  wire core__abc_21380_n2702;
  wire core__abc_21380_n2703;
  wire core__abc_21380_n2705;
  wire core__abc_21380_n2706;
  wire core__abc_21380_n2707;
  wire core__abc_21380_n2709;
  wire core__abc_21380_n2710;
  wire core__abc_21380_n2711;
  wire core__abc_21380_n2712;
  wire core__abc_21380_n2713;
  wire core__abc_21380_n2715;
  wire core__abc_21380_n2716;
  wire core__abc_21380_n2717;
  wire core__abc_21380_n2718;
  wire core__abc_21380_n2719;
  wire core__abc_21380_n2720;
  wire core__abc_21380_n2721;
  wire core__abc_21380_n2722;
  wire core__abc_21380_n2724_1;
  wire core__abc_21380_n2725;
  wire core__abc_21380_n2726;
  wire core__abc_21380_n2727;
  wire core__abc_21380_n2728_1;
  wire core__abc_21380_n2729;
  wire core__abc_21380_n2730;
  wire core__abc_21380_n2732;
  wire core__abc_21380_n2733;
  wire core__abc_21380_n2734;
  wire core__abc_21380_n2735;
  wire core__abc_21380_n2736;
  wire core__abc_21380_n2737;
  wire core__abc_21380_n2738;
  wire core__abc_21380_n2740;
  wire core__abc_21380_n2741;
  wire core__abc_21380_n2742;
  wire core__abc_21380_n2743;
  wire core__abc_21380_n2744;
  wire core__abc_21380_n2746;
  wire core__abc_21380_n2747;
  wire core__abc_21380_n2748;
  wire core__abc_21380_n2749;
  wire core__abc_21380_n2749_bF_buf0;
  wire core__abc_21380_n2749_bF_buf1;
  wire core__abc_21380_n2749_bF_buf10;
  wire core__abc_21380_n2749_bF_buf2;
  wire core__abc_21380_n2749_bF_buf3;
  wire core__abc_21380_n2749_bF_buf4;
  wire core__abc_21380_n2749_bF_buf5;
  wire core__abc_21380_n2749_bF_buf6;
  wire core__abc_21380_n2749_bF_buf7;
  wire core__abc_21380_n2749_bF_buf8;
  wire core__abc_21380_n2749_bF_buf9;
  wire core__abc_21380_n2750;
  wire core__abc_21380_n2750_bF_buf0;
  wire core__abc_21380_n2750_bF_buf1;
  wire core__abc_21380_n2750_bF_buf2;
  wire core__abc_21380_n2750_bF_buf3;
  wire core__abc_21380_n2750_bF_buf4;
  wire core__abc_21380_n2750_bF_buf5;
  wire core__abc_21380_n2750_bF_buf6;
  wire core__abc_21380_n2750_bF_buf7;
  wire core__abc_21380_n2751;
  wire core__abc_21380_n2752;
  wire core__abc_21380_n2753;
  wire core__abc_21380_n2755;
  wire core__abc_21380_n2756;
  wire core__abc_21380_n2757;
  wire core__abc_21380_n2759;
  wire core__abc_21380_n2760;
  wire core__abc_21380_n2761;
  wire core__abc_21380_n2763;
  wire core__abc_21380_n2764;
  wire core__abc_21380_n2765;
  wire core__abc_21380_n2767;
  wire core__abc_21380_n2768;
  wire core__abc_21380_n2769;
  wire core__abc_21380_n2771;
  wire core__abc_21380_n2772;
  wire core__abc_21380_n2773;
  wire core__abc_21380_n2775;
  wire core__abc_21380_n2776;
  wire core__abc_21380_n2777;
  wire core__abc_21380_n2779;
  wire core__abc_21380_n2780;
  wire core__abc_21380_n2781;
  wire core__abc_21380_n2783;
  wire core__abc_21380_n2784;
  wire core__abc_21380_n2785;
  wire core__abc_21380_n2787;
  wire core__abc_21380_n2788;
  wire core__abc_21380_n2789;
  wire core__abc_21380_n2791;
  wire core__abc_21380_n2792;
  wire core__abc_21380_n2793;
  wire core__abc_21380_n2795;
  wire core__abc_21380_n2796;
  wire core__abc_21380_n2797;
  wire core__abc_21380_n2799;
  wire core__abc_21380_n2800_1;
  wire core__abc_21380_n2801;
  wire core__abc_21380_n2803;
  wire core__abc_21380_n2804_1;
  wire core__abc_21380_n2805;
  wire core__abc_21380_n2807;
  wire core__abc_21380_n2808;
  wire core__abc_21380_n2809;
  wire core__abc_21380_n2811;
  wire core__abc_21380_n2812;
  wire core__abc_21380_n2813;
  wire core__abc_21380_n2815;
  wire core__abc_21380_n2816;
  wire core__abc_21380_n2817_1;
  wire core__abc_21380_n2819;
  wire core__abc_21380_n2820;
  wire core__abc_21380_n2821;
  wire core__abc_21380_n2823_1;
  wire core__abc_21380_n2824;
  wire core__abc_21380_n2825;
  wire core__abc_21380_n2827;
  wire core__abc_21380_n2828;
  wire core__abc_21380_n2829;
  wire core__abc_21380_n2831;
  wire core__abc_21380_n2832;
  wire core__abc_21380_n2833;
  wire core__abc_21380_n2835;
  wire core__abc_21380_n2836;
  wire core__abc_21380_n2837;
  wire core__abc_21380_n2839_1;
  wire core__abc_21380_n2840;
  wire core__abc_21380_n2841;
  wire core__abc_21380_n2843;
  wire core__abc_21380_n2844;
  wire core__abc_21380_n2845_1;
  wire core__abc_21380_n2847;
  wire core__abc_21380_n2848;
  wire core__abc_21380_n2849;
  wire core__abc_21380_n2851;
  wire core__abc_21380_n2852;
  wire core__abc_21380_n2853;
  wire core__abc_21380_n2855;
  wire core__abc_21380_n2856;
  wire core__abc_21380_n2857;
  wire core__abc_21380_n2859;
  wire core__abc_21380_n2860_1;
  wire core__abc_21380_n2861;
  wire core__abc_21380_n2863;
  wire core__abc_21380_n2864_1;
  wire core__abc_21380_n2865;
  wire core__abc_21380_n2867;
  wire core__abc_21380_n2868;
  wire core__abc_21380_n2869;
  wire core__abc_21380_n2871;
  wire core__abc_21380_n2872;
  wire core__abc_21380_n2873;
  wire core__abc_21380_n2875;
  wire core__abc_21380_n2876;
  wire core__abc_21380_n2877;
  wire core__abc_21380_n2879;
  wire core__abc_21380_n2880;
  wire core__abc_21380_n2881_1;
  wire core__abc_21380_n2883;
  wire core__abc_21380_n2884;
  wire core__abc_21380_n2885_1;
  wire core__abc_21380_n2887;
  wire core__abc_21380_n2888;
  wire core__abc_21380_n2889;
  wire core__abc_21380_n2891;
  wire core__abc_21380_n2892;
  wire core__abc_21380_n2893;
  wire core__abc_21380_n2895;
  wire core__abc_21380_n2896;
  wire core__abc_21380_n2897;
  wire core__abc_21380_n2899;
  wire core__abc_21380_n2900_1;
  wire core__abc_21380_n2901;
  wire core__abc_21380_n2903;
  wire core__abc_21380_n2904_1;
  wire core__abc_21380_n2905;
  wire core__abc_21380_n2907;
  wire core__abc_21380_n2908;
  wire core__abc_21380_n2909;
  wire core__abc_21380_n2911;
  wire core__abc_21380_n2912;
  wire core__abc_21380_n2913;
  wire core__abc_21380_n2915;
  wire core__abc_21380_n2916_1;
  wire core__abc_21380_n2917;
  wire core__abc_21380_n2919;
  wire core__abc_21380_n2920;
  wire core__abc_21380_n2921;
  wire core__abc_21380_n2923;
  wire core__abc_21380_n2924;
  wire core__abc_21380_n2925;
  wire core__abc_21380_n2927;
  wire core__abc_21380_n2928;
  wire core__abc_21380_n2929;
  wire core__abc_21380_n2931;
  wire core__abc_21380_n2932;
  wire core__abc_21380_n2933;
  wire core__abc_21380_n2935;
  wire core__abc_21380_n2936;
  wire core__abc_21380_n2937;
  wire core__abc_21380_n2939;
  wire core__abc_21380_n2940;
  wire core__abc_21380_n2941;
  wire core__abc_21380_n2943;
  wire core__abc_21380_n2944;
  wire core__abc_21380_n2945;
  wire core__abc_21380_n2947;
  wire core__abc_21380_n2948;
  wire core__abc_21380_n2949;
  wire core__abc_21380_n2951;
  wire core__abc_21380_n2952_1;
  wire core__abc_21380_n2953;
  wire core__abc_21380_n2955;
  wire core__abc_21380_n2956_1;
  wire core__abc_21380_n2957;
  wire core__abc_21380_n2959;
  wire core__abc_21380_n2960;
  wire core__abc_21380_n2961;
  wire core__abc_21380_n2963;
  wire core__abc_21380_n2964;
  wire core__abc_21380_n2965_1;
  wire core__abc_21380_n2967;
  wire core__abc_21380_n2968;
  wire core__abc_21380_n2969;
  wire core__abc_21380_n2971_1;
  wire core__abc_21380_n2972;
  wire core__abc_21380_n2973;
  wire core__abc_21380_n2975;
  wire core__abc_21380_n2976;
  wire core__abc_21380_n2977;
  wire core__abc_21380_n2979;
  wire core__abc_21380_n2980;
  wire core__abc_21380_n2981;
  wire core__abc_21380_n2983;
  wire core__abc_21380_n2984;
  wire core__abc_21380_n2985;
  wire core__abc_21380_n2987;
  wire core__abc_21380_n2988_1;
  wire core__abc_21380_n2989;
  wire core__abc_21380_n2991;
  wire core__abc_21380_n2992;
  wire core__abc_21380_n2993;
  wire core__abc_21380_n2995;
  wire core__abc_21380_n2996;
  wire core__abc_21380_n2997;
  wire core__abc_21380_n2999;
  wire core__abc_21380_n3000;
  wire core__abc_21380_n3001_1;
  wire core__abc_21380_n3003;
  wire core__abc_21380_n3004;
  wire core__abc_21380_n3005_1;
  wire core__abc_21380_n3007;
  wire core__abc_21380_n3008;
  wire core__abc_21380_n3009;
  wire core__abc_21380_n3010;
  wire core__abc_21380_n3011;
  wire core__abc_21380_n3012;
  wire core__abc_21380_n3013;
  wire core__abc_21380_n3014;
  wire core__abc_21380_n3015;
  wire core__abc_21380_n3016;
  wire core__abc_21380_n3017;
  wire core__abc_21380_n3018;
  wire core__abc_21380_n3019;
  wire core__abc_21380_n3020;
  wire core__abc_21380_n3021;
  wire core__abc_21380_n3022;
  wire core__abc_21380_n3023;
  wire core__abc_21380_n3024_1;
  wire core__abc_21380_n3025;
  wire core__abc_21380_n3026;
  wire core__abc_21380_n3027;
  wire core__abc_21380_n3028;
  wire core__abc_21380_n3029;
  wire core__abc_21380_n3030_1;
  wire core__abc_21380_n3031;
  wire core__abc_21380_n3032;
  wire core__abc_21380_n3033;
  wire core__abc_21380_n3034;
  wire core__abc_21380_n3035;
  wire core__abc_21380_n3036;
  wire core__abc_21380_n3037;
  wire core__abc_21380_n3038;
  wire core__abc_21380_n3039;
  wire core__abc_21380_n3040_1;
  wire core__abc_21380_n3041;
  wire core__abc_21380_n3042;
  wire core__abc_21380_n3043;
  wire core__abc_21380_n3044_1;
  wire core__abc_21380_n3045;
  wire core__abc_21380_n3046;
  wire core__abc_21380_n3047;
  wire core__abc_21380_n3048;
  wire core__abc_21380_n3049;
  wire core__abc_21380_n3050;
  wire core__abc_21380_n3051;
  wire core__abc_21380_n3052;
  wire core__abc_21380_n3053;
  wire core__abc_21380_n3054;
  wire core__abc_21380_n3055_1;
  wire core__abc_21380_n3056;
  wire core__abc_21380_n3057;
  wire core__abc_21380_n3058;
  wire core__abc_21380_n3059;
  wire core__abc_21380_n3060;
  wire core__abc_21380_n3061_1;
  wire core__abc_21380_n3062;
  wire core__abc_21380_n3063;
  wire core__abc_21380_n3064;
  wire core__abc_21380_n3065;
  wire core__abc_21380_n3066;
  wire core__abc_21380_n3067;
  wire core__abc_21380_n3068;
  wire core__abc_21380_n3069;
  wire core__abc_21380_n3070;
  wire core__abc_21380_n3071;
  wire core__abc_21380_n3072;
  wire core__abc_21380_n3073_1;
  wire core__abc_21380_n3074;
  wire core__abc_21380_n3075;
  wire core__abc_21380_n3076;
  wire core__abc_21380_n3077_1;
  wire core__abc_21380_n3078;
  wire core__abc_21380_n3079;
  wire core__abc_21380_n3080;
  wire core__abc_21380_n3081;
  wire core__abc_21380_n3082;
  wire core__abc_21380_n3083;
  wire core__abc_21380_n3084;
  wire core__abc_21380_n3085;
  wire core__abc_21380_n3086;
  wire core__abc_21380_n3087;
  wire core__abc_21380_n3088;
  wire core__abc_21380_n3089;
  wire core__abc_21380_n3090;
  wire core__abc_21380_n3091_1;
  wire core__abc_21380_n3092;
  wire core__abc_21380_n3093;
  wire core__abc_21380_n3094;
  wire core__abc_21380_n3095_1;
  wire core__abc_21380_n3096;
  wire core__abc_21380_n3097;
  wire core__abc_21380_n3098;
  wire core__abc_21380_n3099;
  wire core__abc_21380_n3100;
  wire core__abc_21380_n3101;
  wire core__abc_21380_n3102;
  wire core__abc_21380_n3103;
  wire core__abc_21380_n3104_1;
  wire core__abc_21380_n3105;
  wire core__abc_21380_n3106;
  wire core__abc_21380_n3107;
  wire core__abc_21380_n3108;
  wire core__abc_21380_n3109;
  wire core__abc_21380_n3110_1;
  wire core__abc_21380_n3111;
  wire core__abc_21380_n3112;
  wire core__abc_21380_n3113;
  wire core__abc_21380_n3114;
  wire core__abc_21380_n3115;
  wire core__abc_21380_n3116;
  wire core__abc_21380_n3117;
  wire core__abc_21380_n3118;
  wire core__abc_21380_n3119;
  wire core__abc_21380_n3120;
  wire core__abc_21380_n3121;
  wire core__abc_21380_n3122_1;
  wire core__abc_21380_n3123;
  wire core__abc_21380_n3124;
  wire core__abc_21380_n3125;
  wire core__abc_21380_n3126;
  wire core__abc_21380_n3127;
  wire core__abc_21380_n3128_1;
  wire core__abc_21380_n3129;
  wire core__abc_21380_n3130;
  wire core__abc_21380_n3131;
  wire core__abc_21380_n3132;
  wire core__abc_21380_n3133;
  wire core__abc_21380_n3134;
  wire core__abc_21380_n3135;
  wire core__abc_21380_n3136;
  wire core__abc_21380_n3137;
  wire core__abc_21380_n3138;
  wire core__abc_21380_n3139;
  wire core__abc_21380_n3140;
  wire core__abc_21380_n3141_1;
  wire core__abc_21380_n3142;
  wire core__abc_21380_n3143;
  wire core__abc_21380_n3144;
  wire core__abc_21380_n3145_1;
  wire core__abc_21380_n3146;
  wire core__abc_21380_n3147;
  wire core__abc_21380_n3148;
  wire core__abc_21380_n3149;
  wire core__abc_21380_n3150;
  wire core__abc_21380_n3151;
  wire core__abc_21380_n3152;
  wire core__abc_21380_n3153;
  wire core__abc_21380_n3154;
  wire core__abc_21380_n3155;
  wire core__abc_21380_n3156;
  wire core__abc_21380_n3157;
  wire core__abc_21380_n3158;
  wire core__abc_21380_n3159;
  wire core__abc_21380_n3160;
  wire core__abc_21380_n3161;
  wire core__abc_21380_n3162;
  wire core__abc_21380_n3163_1;
  wire core__abc_21380_n3163_1_bF_buf0;
  wire core__abc_21380_n3163_1_bF_buf1;
  wire core__abc_21380_n3163_1_bF_buf2;
  wire core__abc_21380_n3163_1_bF_buf3;
  wire core__abc_21380_n3163_1_bF_buf4;
  wire core__abc_21380_n3163_1_bF_buf5;
  wire core__abc_21380_n3163_1_bF_buf6;
  wire core__abc_21380_n3164;
  wire core__abc_21380_n3165;
  wire core__abc_21380_n3166;
  wire core__abc_21380_n3167_1;
  wire core__abc_21380_n3167_1_bF_buf0;
  wire core__abc_21380_n3167_1_bF_buf1;
  wire core__abc_21380_n3167_1_bF_buf10;
  wire core__abc_21380_n3167_1_bF_buf11;
  wire core__abc_21380_n3167_1_bF_buf12;
  wire core__abc_21380_n3167_1_bF_buf13;
  wire core__abc_21380_n3167_1_bF_buf14;
  wire core__abc_21380_n3167_1_bF_buf14_bF_buf0;
  wire core__abc_21380_n3167_1_bF_buf14_bF_buf1;
  wire core__abc_21380_n3167_1_bF_buf14_bF_buf2;
  wire core__abc_21380_n3167_1_bF_buf14_bF_buf3;
  wire core__abc_21380_n3167_1_bF_buf15;
  wire core__abc_21380_n3167_1_bF_buf15_bF_buf0;
  wire core__abc_21380_n3167_1_bF_buf15_bF_buf1;
  wire core__abc_21380_n3167_1_bF_buf15_bF_buf2;
  wire core__abc_21380_n3167_1_bF_buf15_bF_buf3;
  wire core__abc_21380_n3167_1_bF_buf2;
  wire core__abc_21380_n3167_1_bF_buf3;
  wire core__abc_21380_n3167_1_bF_buf4;
  wire core__abc_21380_n3167_1_bF_buf5;
  wire core__abc_21380_n3167_1_bF_buf6;
  wire core__abc_21380_n3167_1_bF_buf7;
  wire core__abc_21380_n3167_1_bF_buf8;
  wire core__abc_21380_n3167_1_bF_buf9;
  wire core__abc_21380_n3168;
  wire core__abc_21380_n3169;
  wire core__abc_21380_n3170;
  wire core__abc_21380_n3171;
  wire core__abc_21380_n3172;
  wire core__abc_21380_n3173;
  wire core__abc_21380_n3174;
  wire core__abc_21380_n3175;
  wire core__abc_21380_n3176;
  wire core__abc_21380_n3177_1;
  wire core__abc_21380_n3178;
  wire core__abc_21380_n3179;
  wire core__abc_21380_n3180;
  wire core__abc_21380_n3181_1;
  wire core__abc_21380_n3182;
  wire core__abc_21380_n3183;
  wire core__abc_21380_n3184;
  wire core__abc_21380_n3185;
  wire core__abc_21380_n3186;
  wire core__abc_21380_n3187;
  wire core__abc_21380_n3188;
  wire core__abc_21380_n3189;
  wire core__abc_21380_n3190;
  wire core__abc_21380_n3191;
  wire core__abc_21380_n3192;
  wire core__abc_21380_n3193;
  wire core__abc_21380_n3194_1;
  wire core__abc_21380_n3195;
  wire core__abc_21380_n3196;
  wire core__abc_21380_n3197;
  wire core__abc_21380_n3198;
  wire core__abc_21380_n3199;
  wire core__abc_21380_n3200_1;
  wire core__abc_21380_n3201;
  wire core__abc_21380_n3202;
  wire core__abc_21380_n3203;
  wire core__abc_21380_n3204;
  wire core__abc_21380_n3205;
  wire core__abc_21380_n3206;
  wire core__abc_21380_n3207;
  wire core__abc_21380_n3208;
  wire core__abc_21380_n3209;
  wire core__abc_21380_n3210;
  wire core__abc_21380_n3211_1;
  wire core__abc_21380_n3212;
  wire core__abc_21380_n3213;
  wire core__abc_21380_n3214;
  wire core__abc_21380_n3215_1;
  wire core__abc_21380_n3216;
  wire core__abc_21380_n3217;
  wire core__abc_21380_n3218;
  wire core__abc_21380_n3219;
  wire core__abc_21380_n3220;
  wire core__abc_21380_n3221;
  wire core__abc_21380_n3222;
  wire core__abc_21380_n3223;
  wire core__abc_21380_n3224;
  wire core__abc_21380_n3225;
  wire core__abc_21380_n3226;
  wire core__abc_21380_n3227;
  wire core__abc_21380_n3228;
  wire core__abc_21380_n3229;
  wire core__abc_21380_n3230_1;
  wire core__abc_21380_n3231;
  wire core__abc_21380_n3232;
  wire core__abc_21380_n3233;
  wire core__abc_21380_n3234;
  wire core__abc_21380_n3235;
  wire core__abc_21380_n3236_1;
  wire core__abc_21380_n3237;
  wire core__abc_21380_n3238;
  wire core__abc_21380_n3239;
  wire core__abc_21380_n3240;
  wire core__abc_21380_n3241;
  wire core__abc_21380_n3242;
  wire core__abc_21380_n3243;
  wire core__abc_21380_n3244;
  wire core__abc_21380_n3245_1;
  wire core__abc_21380_n3246;
  wire core__abc_21380_n3247;
  wire core__abc_21380_n3248;
  wire core__abc_21380_n3249;
  wire core__abc_21380_n3250;
  wire core__abc_21380_n3251_1;
  wire core__abc_21380_n3252;
  wire core__abc_21380_n3253;
  wire core__abc_21380_n3254;
  wire core__abc_21380_n3255;
  wire core__abc_21380_n3256;
  wire core__abc_21380_n3257;
  wire core__abc_21380_n3258;
  wire core__abc_21380_n3259;
  wire core__abc_21380_n3260;
  wire core__abc_21380_n3261;
  wire core__abc_21380_n3262_1;
  wire core__abc_21380_n3263;
  wire core__abc_21380_n3264;
  wire core__abc_21380_n3265;
  wire core__abc_21380_n3266;
  wire core__abc_21380_n3267;
  wire core__abc_21380_n3268_1;
  wire core__abc_21380_n3269;
  wire core__abc_21380_n3270;
  wire core__abc_21380_n3271;
  wire core__abc_21380_n3272;
  wire core__abc_21380_n3273;
  wire core__abc_21380_n3274;
  wire core__abc_21380_n3275;
  wire core__abc_21380_n3276;
  wire core__abc_21380_n3277_1;
  wire core__abc_21380_n3278;
  wire core__abc_21380_n3279;
  wire core__abc_21380_n3280;
  wire core__abc_21380_n3281_1;
  wire core__abc_21380_n3282;
  wire core__abc_21380_n3283;
  wire core__abc_21380_n3284;
  wire core__abc_21380_n3285;
  wire core__abc_21380_n3286;
  wire core__abc_21380_n3287;
  wire core__abc_21380_n3288;
  wire core__abc_21380_n3289;
  wire core__abc_21380_n3290;
  wire core__abc_21380_n3291;
  wire core__abc_21380_n3292;
  wire core__abc_21380_n3293;
  wire core__abc_21380_n3294;
  wire core__abc_21380_n3295;
  wire core__abc_21380_n3296;
  wire core__abc_21380_n3297;
  wire core__abc_21380_n3298;
  wire core__abc_21380_n3299;
  wire core__abc_21380_n3300;
  wire core__abc_21380_n3301;
  wire core__abc_21380_n3302;
  wire core__abc_21380_n3303;
  wire core__abc_21380_n3304;
  wire core__abc_21380_n3305;
  wire core__abc_21380_n3306;
  wire core__abc_21380_n3307;
  wire core__abc_21380_n3308;
  wire core__abc_21380_n3309;
  wire core__abc_21380_n3310;
  wire core__abc_21380_n3311;
  wire core__abc_21380_n3312;
  wire core__abc_21380_n3313;
  wire core__abc_21380_n3313_bF_buf0;
  wire core__abc_21380_n3313_bF_buf1;
  wire core__abc_21380_n3313_bF_buf10;
  wire core__abc_21380_n3313_bF_buf11;
  wire core__abc_21380_n3313_bF_buf12;
  wire core__abc_21380_n3313_bF_buf2;
  wire core__abc_21380_n3313_bF_buf3;
  wire core__abc_21380_n3313_bF_buf4;
  wire core__abc_21380_n3313_bF_buf5;
  wire core__abc_21380_n3313_bF_buf6;
  wire core__abc_21380_n3313_bF_buf7;
  wire core__abc_21380_n3313_bF_buf8;
  wire core__abc_21380_n3313_bF_buf9;
  wire core__abc_21380_n3314;
  wire core__abc_21380_n3315;
  wire core__abc_21380_n3316;
  wire core__abc_21380_n3317;
  wire core__abc_21380_n3317_bF_buf0;
  wire core__abc_21380_n3317_bF_buf1;
  wire core__abc_21380_n3317_bF_buf2;
  wire core__abc_21380_n3317_bF_buf3;
  wire core__abc_21380_n3317_bF_buf4;
  wire core__abc_21380_n3317_bF_buf5;
  wire core__abc_21380_n3317_bF_buf6;
  wire core__abc_21380_n3317_bF_buf7;
  wire core__abc_21380_n3318;
  wire core__abc_21380_n3319;
  wire core__abc_21380_n3320;
  wire core__abc_21380_n3321;
  wire core__abc_21380_n3322;
  wire core__abc_21380_n3323;
  wire core__abc_21380_n3324;
  wire core__abc_21380_n3325;
  wire core__abc_21380_n3326;
  wire core__abc_21380_n3327;
  wire core__abc_21380_n3328;
  wire core__abc_21380_n3328_bF_buf0;
  wire core__abc_21380_n3328_bF_buf1;
  wire core__abc_21380_n3328_bF_buf2;
  wire core__abc_21380_n3328_bF_buf3;
  wire core__abc_21380_n3328_bF_buf4;
  wire core__abc_21380_n3328_bF_buf5;
  wire core__abc_21380_n3328_bF_buf6;
  wire core__abc_21380_n3328_bF_buf7;
  wire core__abc_21380_n3329;
  wire core__abc_21380_n3330;
  wire core__abc_21380_n3332;
  wire core__abc_21380_n3333;
  wire core__abc_21380_n3334;
  wire core__abc_21380_n3335;
  wire core__abc_21380_n3336;
  wire core__abc_21380_n3337;
  wire core__abc_21380_n3338;
  wire core__abc_21380_n3339;
  wire core__abc_21380_n3340;
  wire core__abc_21380_n3341;
  wire core__abc_21380_n3342;
  wire core__abc_21380_n3343;
  wire core__abc_21380_n3344;
  wire core__abc_21380_n3345;
  wire core__abc_21380_n3346;
  wire core__abc_21380_n3347;
  wire core__abc_21380_n3348;
  wire core__abc_21380_n3349;
  wire core__abc_21380_n3350;
  wire core__abc_21380_n3351;
  wire core__abc_21380_n3352;
  wire core__abc_21380_n3353;
  wire core__abc_21380_n3354;
  wire core__abc_21380_n3355;
  wire core__abc_21380_n3356;
  wire core__abc_21380_n3357;
  wire core__abc_21380_n3358;
  wire core__abc_21380_n3359;
  wire core__abc_21380_n3360;
  wire core__abc_21380_n3361;
  wire core__abc_21380_n3362;
  wire core__abc_21380_n3363;
  wire core__abc_21380_n3364;
  wire core__abc_21380_n3365;
  wire core__abc_21380_n3366;
  wire core__abc_21380_n3367;
  wire core__abc_21380_n3368;
  wire core__abc_21380_n3369;
  wire core__abc_21380_n3370;
  wire core__abc_21380_n3371;
  wire core__abc_21380_n3372;
  wire core__abc_21380_n3373;
  wire core__abc_21380_n3374;
  wire core__abc_21380_n3375;
  wire core__abc_21380_n3376;
  wire core__abc_21380_n3377;
  wire core__abc_21380_n3378;
  wire core__abc_21380_n3379;
  wire core__abc_21380_n3380;
  wire core__abc_21380_n3381;
  wire core__abc_21380_n3382;
  wire core__abc_21380_n3383;
  wire core__abc_21380_n3384;
  wire core__abc_21380_n3385;
  wire core__abc_21380_n3386;
  wire core__abc_21380_n3387;
  wire core__abc_21380_n3388;
  wire core__abc_21380_n3389;
  wire core__abc_21380_n3390;
  wire core__abc_21380_n3391;
  wire core__abc_21380_n3392;
  wire core__abc_21380_n3393;
  wire core__abc_21380_n3394;
  wire core__abc_21380_n3395;
  wire core__abc_21380_n3396;
  wire core__abc_21380_n3397;
  wire core__abc_21380_n3398;
  wire core__abc_21380_n3399;
  wire core__abc_21380_n3400;
  wire core__abc_21380_n3402;
  wire core__abc_21380_n3403;
  wire core__abc_21380_n3404;
  wire core__abc_21380_n3405;
  wire core__abc_21380_n3406;
  wire core__abc_21380_n3407;
  wire core__abc_21380_n3408;
  wire core__abc_21380_n3409;
  wire core__abc_21380_n3410;
  wire core__abc_21380_n3411;
  wire core__abc_21380_n3412;
  wire core__abc_21380_n3413;
  wire core__abc_21380_n3414;
  wire core__abc_21380_n3415;
  wire core__abc_21380_n3416;
  wire core__abc_21380_n3417;
  wire core__abc_21380_n3418;
  wire core__abc_21380_n3419;
  wire core__abc_21380_n3420;
  wire core__abc_21380_n3421;
  wire core__abc_21380_n3422;
  wire core__abc_21380_n3423;
  wire core__abc_21380_n3424;
  wire core__abc_21380_n3425;
  wire core__abc_21380_n3426;
  wire core__abc_21380_n3427;
  wire core__abc_21380_n3428;
  wire core__abc_21380_n3429;
  wire core__abc_21380_n3430;
  wire core__abc_21380_n3431;
  wire core__abc_21380_n3432;
  wire core__abc_21380_n3433;
  wire core__abc_21380_n3434;
  wire core__abc_21380_n3435;
  wire core__abc_21380_n3436;
  wire core__abc_21380_n3437;
  wire core__abc_21380_n3438;
  wire core__abc_21380_n3439;
  wire core__abc_21380_n3440;
  wire core__abc_21380_n3441;
  wire core__abc_21380_n3442;
  wire core__abc_21380_n3443;
  wire core__abc_21380_n3444;
  wire core__abc_21380_n3445;
  wire core__abc_21380_n3446;
  wire core__abc_21380_n3447;
  wire core__abc_21380_n3448;
  wire core__abc_21380_n3449;
  wire core__abc_21380_n3450;
  wire core__abc_21380_n3451;
  wire core__abc_21380_n3452;
  wire core__abc_21380_n3453;
  wire core__abc_21380_n3454;
  wire core__abc_21380_n3455;
  wire core__abc_21380_n3456;
  wire core__abc_21380_n3457;
  wire core__abc_21380_n3459;
  wire core__abc_21380_n3460;
  wire core__abc_21380_n3461;
  wire core__abc_21380_n3462;
  wire core__abc_21380_n3463;
  wire core__abc_21380_n3464;
  wire core__abc_21380_n3465;
  wire core__abc_21380_n3466;
  wire core__abc_21380_n3467;
  wire core__abc_21380_n3468;
  wire core__abc_21380_n3469;
  wire core__abc_21380_n3470;
  wire core__abc_21380_n3471;
  wire core__abc_21380_n3472;
  wire core__abc_21380_n3473;
  wire core__abc_21380_n3474;
  wire core__abc_21380_n3475;
  wire core__abc_21380_n3476;
  wire core__abc_21380_n3477;
  wire core__abc_21380_n3478;
  wire core__abc_21380_n3479;
  wire core__abc_21380_n3480;
  wire core__abc_21380_n3481;
  wire core__abc_21380_n3482;
  wire core__abc_21380_n3483_1;
  wire core__abc_21380_n3484;
  wire core__abc_21380_n3485_1;
  wire core__abc_21380_n3486;
  wire core__abc_21380_n3487;
  wire core__abc_21380_n3488;
  wire core__abc_21380_n3489;
  wire core__abc_21380_n3490_1;
  wire core__abc_21380_n3491;
  wire core__abc_21380_n3492;
  wire core__abc_21380_n3493;
  wire core__abc_21380_n3494;
  wire core__abc_21380_n3495;
  wire core__abc_21380_n3496;
  wire core__abc_21380_n3497;
  wire core__abc_21380_n3498;
  wire core__abc_21380_n3499;
  wire core__abc_21380_n3500;
  wire core__abc_21380_n3501_1;
  wire core__abc_21380_n3502;
  wire core__abc_21380_n3503;
  wire core__abc_21380_n3504;
  wire core__abc_21380_n3505_1;
  wire core__abc_21380_n3506;
  wire core__abc_21380_n3507;
  wire core__abc_21380_n3508;
  wire core__abc_21380_n3509;
  wire core__abc_21380_n3510;
  wire core__abc_21380_n3511;
  wire core__abc_21380_n3512;
  wire core__abc_21380_n3513;
  wire core__abc_21380_n3514;
  wire core__abc_21380_n3515;
  wire core__abc_21380_n3516;
  wire core__abc_21380_n3517;
  wire core__abc_21380_n3518_1;
  wire core__abc_21380_n3519;
  wire core__abc_21380_n3520;
  wire core__abc_21380_n3521;
  wire core__abc_21380_n3523;
  wire core__abc_21380_n3524;
  wire core__abc_21380_n3525;
  wire core__abc_21380_n3526;
  wire core__abc_21380_n3527;
  wire core__abc_21380_n3528;
  wire core__abc_21380_n3529;
  wire core__abc_21380_n3530;
  wire core__abc_21380_n3531_1;
  wire core__abc_21380_n3532;
  wire core__abc_21380_n3533;
  wire core__abc_21380_n3534;
  wire core__abc_21380_n3535_1;
  wire core__abc_21380_n3536;
  wire core__abc_21380_n3537;
  wire core__abc_21380_n3538;
  wire core__abc_21380_n3539;
  wire core__abc_21380_n3540;
  wire core__abc_21380_n3541;
  wire core__abc_21380_n3542;
  wire core__abc_21380_n3543;
  wire core__abc_21380_n3544;
  wire core__abc_21380_n3545;
  wire core__abc_21380_n3546;
  wire core__abc_21380_n3547;
  wire core__abc_21380_n3548_1;
  wire core__abc_21380_n3549;
  wire core__abc_21380_n3550;
  wire core__abc_21380_n3551;
  wire core__abc_21380_n3552_1;
  wire core__abc_21380_n3553;
  wire core__abc_21380_n3554;
  wire core__abc_21380_n3555;
  wire core__abc_21380_n3556;
  wire core__abc_21380_n3557;
  wire core__abc_21380_n3558;
  wire core__abc_21380_n3559;
  wire core__abc_21380_n3560;
  wire core__abc_21380_n3561_1;
  wire core__abc_21380_n3562;
  wire core__abc_21380_n3563;
  wire core__abc_21380_n3564;
  wire core__abc_21380_n3565;
  wire core__abc_21380_n3566;
  wire core__abc_21380_n3567;
  wire core__abc_21380_n3568;
  wire core__abc_21380_n3569_1;
  wire core__abc_21380_n3570;
  wire core__abc_21380_n3571;
  wire core__abc_21380_n3572;
  wire core__abc_21380_n3573;
  wire core__abc_21380_n3574;
  wire core__abc_21380_n3575;
  wire core__abc_21380_n3576;
  wire core__abc_21380_n3577;
  wire core__abc_21380_n3578;
  wire core__abc_21380_n3579;
  wire core__abc_21380_n3580;
  wire core__abc_21380_n3581_1;
  wire core__abc_21380_n3582;
  wire core__abc_21380_n3583;
  wire core__abc_21380_n3584;
  wire core__abc_21380_n3585;
  wire core__abc_21380_n3586;
  wire core__abc_21380_n3587;
  wire core__abc_21380_n3588;
  wire core__abc_21380_n3589_1;
  wire core__abc_21380_n3590;
  wire core__abc_21380_n3591;
  wire core__abc_21380_n3592;
  wire core__abc_21380_n3593;
  wire core__abc_21380_n3594;
  wire core__abc_21380_n3595;
  wire core__abc_21380_n3597;
  wire core__abc_21380_n3598;
  wire core__abc_21380_n3599;
  wire core__abc_21380_n3600_1;
  wire core__abc_21380_n3601;
  wire core__abc_21380_n3602;
  wire core__abc_21380_n3603;
  wire core__abc_21380_n3604_1;
  wire core__abc_21380_n3605;
  wire core__abc_21380_n3606;
  wire core__abc_21380_n3607;
  wire core__abc_21380_n3608;
  wire core__abc_21380_n3609;
  wire core__abc_21380_n3610;
  wire core__abc_21380_n3611;
  wire core__abc_21380_n3612;
  wire core__abc_21380_n3613;
  wire core__abc_21380_n3614;
  wire core__abc_21380_n3615;
  wire core__abc_21380_n3616;
  wire core__abc_21380_n3617;
  wire core__abc_21380_n3618;
  wire core__abc_21380_n3619_1;
  wire core__abc_21380_n3620;
  wire core__abc_21380_n3621;
  wire core__abc_21380_n3622;
  wire core__abc_21380_n3623_1;
  wire core__abc_21380_n3624;
  wire core__abc_21380_n3625;
  wire core__abc_21380_n3626;
  wire core__abc_21380_n3627;
  wire core__abc_21380_n3628;
  wire core__abc_21380_n3629;
  wire core__abc_21380_n3630;
  wire core__abc_21380_n3631_1;
  wire core__abc_21380_n3632;
  wire core__abc_21380_n3633;
  wire core__abc_21380_n3634;
  wire core__abc_21380_n3635;
  wire core__abc_21380_n3636_1;
  wire core__abc_21380_n3637;
  wire core__abc_21380_n3638;
  wire core__abc_21380_n3639;
  wire core__abc_21380_n3640;
  wire core__abc_21380_n3641;
  wire core__abc_21380_n3642;
  wire core__abc_21380_n3643;
  wire core__abc_21380_n3644;
  wire core__abc_21380_n3645;
  wire core__abc_21380_n3646;
  wire core__abc_21380_n3647_1;
  wire core__abc_21380_n3648;
  wire core__abc_21380_n3649;
  wire core__abc_21380_n3650;
  wire core__abc_21380_n3651_1;
  wire core__abc_21380_n3652;
  wire core__abc_21380_n3653;
  wire core__abc_21380_n3654;
  wire core__abc_21380_n3655;
  wire core__abc_21380_n3656;
  wire core__abc_21380_n3657;
  wire core__abc_21380_n3658;
  wire core__abc_21380_n3659_1;
  wire core__abc_21380_n3660;
  wire core__abc_21380_n3661;
  wire core__abc_21380_n3662;
  wire core__abc_21380_n3663_1;
  wire core__abc_21380_n3664;
  wire core__abc_21380_n3666;
  wire core__abc_21380_n3667;
  wire core__abc_21380_n3668;
  wire core__abc_21380_n3669;
  wire core__abc_21380_n3670;
  wire core__abc_21380_n3671;
  wire core__abc_21380_n3672;
  wire core__abc_21380_n3673;
  wire core__abc_21380_n3674;
  wire core__abc_21380_n3675;
  wire core__abc_21380_n3676_1;
  wire core__abc_21380_n3677;
  wire core__abc_21380_n3678;
  wire core__abc_21380_n3679;
  wire core__abc_21380_n3680;
  wire core__abc_21380_n3681_1;
  wire core__abc_21380_n3682;
  wire core__abc_21380_n3683;
  wire core__abc_21380_n3684;
  wire core__abc_21380_n3685;
  wire core__abc_21380_n3686;
  wire core__abc_21380_n3687;
  wire core__abc_21380_n3688_1;
  wire core__abc_21380_n3689;
  wire core__abc_21380_n3690;
  wire core__abc_21380_n3691;
  wire core__abc_21380_n3692;
  wire core__abc_21380_n3693_1;
  wire core__abc_21380_n3694;
  wire core__abc_21380_n3695;
  wire core__abc_21380_n3696;
  wire core__abc_21380_n3697;
  wire core__abc_21380_n3698;
  wire core__abc_21380_n3699;
  wire core__abc_21380_n3700;
  wire core__abc_21380_n3701;
  wire core__abc_21380_n3702;
  wire core__abc_21380_n3703_1;
  wire core__abc_21380_n3704;
  wire core__abc_21380_n3705;
  wire core__abc_21380_n3706;
  wire core__abc_21380_n3707;
  wire core__abc_21380_n3708_1;
  wire core__abc_21380_n3709;
  wire core__abc_21380_n3710;
  wire core__abc_21380_n3711;
  wire core__abc_21380_n3712;
  wire core__abc_21380_n3713;
  wire core__abc_21380_n3714;
  wire core__abc_21380_n3715;
  wire core__abc_21380_n3716_1;
  wire core__abc_21380_n3717;
  wire core__abc_21380_n3718;
  wire core__abc_21380_n3719;
  wire core__abc_21380_n3720_1;
  wire core__abc_21380_n3721;
  wire core__abc_21380_n3722;
  wire core__abc_21380_n3723;
  wire core__abc_21380_n3724;
  wire core__abc_21380_n3725;
  wire core__abc_21380_n3726;
  wire core__abc_21380_n3727;
  wire core__abc_21380_n3728;
  wire core__abc_21380_n3729;
  wire core__abc_21380_n3730;
  wire core__abc_21380_n3731;
  wire core__abc_21380_n3732;
  wire core__abc_21380_n3733;
  wire core__abc_21380_n3734;
  wire core__abc_21380_n3735;
  wire core__abc_21380_n3736;
  wire core__abc_21380_n3738;
  wire core__abc_21380_n3739;
  wire core__abc_21380_n3740_1;
  wire core__abc_21380_n3741;
  wire core__abc_21380_n3742;
  wire core__abc_21380_n3743;
  wire core__abc_21380_n3744;
  wire core__abc_21380_n3745_1;
  wire core__abc_21380_n3746;
  wire core__abc_21380_n3747;
  wire core__abc_21380_n3748;
  wire core__abc_21380_n3749;
  wire core__abc_21380_n3750;
  wire core__abc_21380_n3751;
  wire core__abc_21380_n3752_1;
  wire core__abc_21380_n3753;
  wire core__abc_21380_n3754;
  wire core__abc_21380_n3755;
  wire core__abc_21380_n3756_1;
  wire core__abc_21380_n3757;
  wire core__abc_21380_n3758;
  wire core__abc_21380_n3759;
  wire core__abc_21380_n3760;
  wire core__abc_21380_n3761;
  wire core__abc_21380_n3762;
  wire core__abc_21380_n3763;
  wire core__abc_21380_n3764;
  wire core__abc_21380_n3765;
  wire core__abc_21380_n3766;
  wire core__abc_21380_n3767_1;
  wire core__abc_21380_n3768;
  wire core__abc_21380_n3769;
  wire core__abc_21380_n3770;
  wire core__abc_21380_n3771;
  wire core__abc_21380_n3772_1;
  wire core__abc_21380_n3773;
  wire core__abc_21380_n3774;
  wire core__abc_21380_n3775;
  wire core__abc_21380_n3776;
  wire core__abc_21380_n3777;
  wire core__abc_21380_n3778;
  wire core__abc_21380_n3779_1;
  wire core__abc_21380_n3780;
  wire core__abc_21380_n3781;
  wire core__abc_21380_n3782;
  wire core__abc_21380_n3783_1;
  wire core__abc_21380_n3784;
  wire core__abc_21380_n3785;
  wire core__abc_21380_n3786;
  wire core__abc_21380_n3787;
  wire core__abc_21380_n3788;
  wire core__abc_21380_n3789;
  wire core__abc_21380_n3790;
  wire core__abc_21380_n3791;
  wire core__abc_21380_n3792;
  wire core__abc_21380_n3793;
  wire core__abc_21380_n3794;
  wire core__abc_21380_n3795;
  wire core__abc_21380_n3797_1;
  wire core__abc_21380_n3798;
  wire core__abc_21380_n3799;
  wire core__abc_21380_n3800;
  wire core__abc_21380_n3801_1;
  wire core__abc_21380_n3802;
  wire core__abc_21380_n3803;
  wire core__abc_21380_n3804;
  wire core__abc_21380_n3805;
  wire core__abc_21380_n3806;
  wire core__abc_21380_n3807;
  wire core__abc_21380_n3808;
  wire core__abc_21380_n3809_1;
  wire core__abc_21380_n3810;
  wire core__abc_21380_n3811;
  wire core__abc_21380_n3812;
  wire core__abc_21380_n3813;
  wire core__abc_21380_n3814_1;
  wire core__abc_21380_n3815;
  wire core__abc_21380_n3816;
  wire core__abc_21380_n3817;
  wire core__abc_21380_n3818;
  wire core__abc_21380_n3819;
  wire core__abc_21380_n3820;
  wire core__abc_21380_n3821;
  wire core__abc_21380_n3822;
  wire core__abc_21380_n3823_1;
  wire core__abc_21380_n3824;
  wire core__abc_21380_n3825;
  wire core__abc_21380_n3826;
  wire core__abc_21380_n3827;
  wire core__abc_21380_n3828_1;
  wire core__abc_21380_n3829;
  wire core__abc_21380_n3830;
  wire core__abc_21380_n3831;
  wire core__abc_21380_n3832;
  wire core__abc_21380_n3833;
  wire core__abc_21380_n3834_1;
  wire core__abc_21380_n3835;
  wire core__abc_21380_n3836;
  wire core__abc_21380_n3837;
  wire core__abc_21380_n3838_1;
  wire core__abc_21380_n3839;
  wire core__abc_21380_n3840;
  wire core__abc_21380_n3841;
  wire core__abc_21380_n3842;
  wire core__abc_21380_n3843;
  wire core__abc_21380_n3844;
  wire core__abc_21380_n3845;
  wire core__abc_21380_n3846;
  wire core__abc_21380_n3847;
  wire core__abc_21380_n3848;
  wire core__abc_21380_n3849;
  wire core__abc_21380_n3850;
  wire core__abc_21380_n3851;
  wire core__abc_21380_n3852;
  wire core__abc_21380_n3853_1;
  wire core__abc_21380_n3854;
  wire core__abc_21380_n3855;
  wire core__abc_21380_n3856;
  wire core__abc_21380_n3857_1;
  wire core__abc_21380_n3858;
  wire core__abc_21380_n3859;
  wire core__abc_21380_n3860;
  wire core__abc_21380_n3861;
  wire core__abc_21380_n3862;
  wire core__abc_21380_n3863;
  wire core__abc_21380_n3864_1;
  wire core__abc_21380_n3865;
  wire core__abc_21380_n3866;
  wire core__abc_21380_n3867;
  wire core__abc_21380_n3868;
  wire core__abc_21380_n3869_1;
  wire core__abc_21380_n3870;
  wire core__abc_21380_n3871;
  wire core__abc_21380_n3872;
  wire core__abc_21380_n3873;
  wire core__abc_21380_n3874;
  wire core__abc_21380_n3875;
  wire core__abc_21380_n3876;
  wire core__abc_21380_n3877;
  wire core__abc_21380_n3879;
  wire core__abc_21380_n3880;
  wire core__abc_21380_n3881_1;
  wire core__abc_21380_n3882;
  wire core__abc_21380_n3883;
  wire core__abc_21380_n3884;
  wire core__abc_21380_n3885;
  wire core__abc_21380_n3886_1;
  wire core__abc_21380_n3887;
  wire core__abc_21380_n3888;
  wire core__abc_21380_n3889;
  wire core__abc_21380_n3890;
  wire core__abc_21380_n3891;
  wire core__abc_21380_n3892;
  wire core__abc_21380_n3893_1;
  wire core__abc_21380_n3894;
  wire core__abc_21380_n3895;
  wire core__abc_21380_n3896;
  wire core__abc_21380_n3897;
  wire core__abc_21380_n3898_1;
  wire core__abc_21380_n3899;
  wire core__abc_21380_n3900;
  wire core__abc_21380_n3901;
  wire core__abc_21380_n3902;
  wire core__abc_21380_n3903;
  wire core__abc_21380_n3904;
  wire core__abc_21380_n3905;
  wire core__abc_21380_n3906;
  wire core__abc_21380_n3907;
  wire core__abc_21380_n3908;
  wire core__abc_21380_n3909;
  wire core__abc_21380_n3910_1;
  wire core__abc_21380_n3911;
  wire core__abc_21380_n3912;
  wire core__abc_21380_n3913;
  wire core__abc_21380_n3914_1;
  wire core__abc_21380_n3915;
  wire core__abc_21380_n3916;
  wire core__abc_21380_n3917;
  wire core__abc_21380_n3918;
  wire core__abc_21380_n3919;
  wire core__abc_21380_n3920;
  wire core__abc_21380_n3921;
  wire core__abc_21380_n3922_1;
  wire core__abc_21380_n3923;
  wire core__abc_21380_n3924;
  wire core__abc_21380_n3925;
  wire core__abc_21380_n3926;
  wire core__abc_21380_n3927_1;
  wire core__abc_21380_n3928;
  wire core__abc_21380_n3929;
  wire core__abc_21380_n3930;
  wire core__abc_21380_n3931;
  wire core__abc_21380_n3932;
  wire core__abc_21380_n3933;
  wire core__abc_21380_n3934;
  wire core__abc_21380_n3935;
  wire core__abc_21380_n3936;
  wire core__abc_21380_n3937_1;
  wire core__abc_21380_n3938;
  wire core__abc_21380_n3939;
  wire core__abc_21380_n3940;
  wire core__abc_21380_n3941;
  wire core__abc_21380_n3942_1;
  wire core__abc_21380_n3943;
  wire core__abc_21380_n3944;
  wire core__abc_21380_n3946;
  wire core__abc_21380_n3947;
  wire core__abc_21380_n3948_1;
  wire core__abc_21380_n3949;
  wire core__abc_21380_n3950;
  wire core__abc_21380_n3951;
  wire core__abc_21380_n3952_1;
  wire core__abc_21380_n3953;
  wire core__abc_21380_n3954;
  wire core__abc_21380_n3955_1;
  wire core__abc_21380_n3956;
  wire core__abc_21380_n3957;
  wire core__abc_21380_n3958;
  wire core__abc_21380_n3959;
  wire core__abc_21380_n3960;
  wire core__abc_21380_n3961_1;
  wire core__abc_21380_n3962;
  wire core__abc_21380_n3963;
  wire core__abc_21380_n3964;
  wire core__abc_21380_n3965_1;
  wire core__abc_21380_n3966;
  wire core__abc_21380_n3967;
  wire core__abc_21380_n3968;
  wire core__abc_21380_n3969_1;
  wire core__abc_21380_n3970;
  wire core__abc_21380_n3971;
  wire core__abc_21380_n3972;
  wire core__abc_21380_n3973;
  wire core__abc_21380_n3974_1;
  wire core__abc_21380_n3975;
  wire core__abc_21380_n3976;
  wire core__abc_21380_n3977;
  wire core__abc_21380_n3978;
  wire core__abc_21380_n3979_1;
  wire core__abc_21380_n3980;
  wire core__abc_21380_n3981;
  wire core__abc_21380_n3982_1;
  wire core__abc_21380_n3983;
  wire core__abc_21380_n3984;
  wire core__abc_21380_n3985;
  wire core__abc_21380_n3986_1;
  wire core__abc_21380_n3987;
  wire core__abc_21380_n3988_1;
  wire core__abc_21380_n3989;
  wire core__abc_21380_n3990;
  wire core__abc_21380_n3991;
  wire core__abc_21380_n3992_1;
  wire core__abc_21380_n3993;
  wire core__abc_21380_n3994;
  wire core__abc_21380_n3995_1;
  wire core__abc_21380_n3996;
  wire core__abc_21380_n3997;
  wire core__abc_21380_n3998;
  wire core__abc_21380_n3999;
  wire core__abc_21380_n4000_1;
  wire core__abc_21380_n4001;
  wire core__abc_21380_n4002;
  wire core__abc_21380_n4003_1;
  wire core__abc_21380_n4004;
  wire core__abc_21380_n4006;
  wire core__abc_21380_n4007;
  wire core__abc_21380_n4008_1;
  wire core__abc_21380_n4009;
  wire core__abc_21380_n4010;
  wire core__abc_21380_n4011;
  wire core__abc_21380_n4012_1;
  wire core__abc_21380_n4013;
  wire core__abc_21380_n4014;
  wire core__abc_21380_n4015;
  wire core__abc_21380_n4016_1;
  wire core__abc_21380_n4017;
  wire core__abc_21380_n4018_1;
  wire core__abc_21380_n4019;
  wire core__abc_21380_n4020;
  wire core__abc_21380_n4021;
  wire core__abc_21380_n4022;
  wire core__abc_21380_n4023_1;
  wire core__abc_21380_n4024;
  wire core__abc_21380_n4025;
  wire core__abc_21380_n4026_1;
  wire core__abc_21380_n4027;
  wire core__abc_21380_n4028;
  wire core__abc_21380_n4029;
  wire core__abc_21380_n4030;
  wire core__abc_21380_n4031_1;
  wire core__abc_21380_n4032;
  wire core__abc_21380_n4033;
  wire core__abc_21380_n4034_1;
  wire core__abc_21380_n4035;
  wire core__abc_21380_n4036;
  wire core__abc_21380_n4037;
  wire core__abc_21380_n4038;
  wire core__abc_21380_n4039_1;
  wire core__abc_21380_n4040;
  wire core__abc_21380_n4041;
  wire core__abc_21380_n4042;
  wire core__abc_21380_n4043_1;
  wire core__abc_21380_n4044;
  wire core__abc_21380_n4045;
  wire core__abc_21380_n4046;
  wire core__abc_21380_n4047_1;
  wire core__abc_21380_n4048;
  wire core__abc_21380_n4049;
  wire core__abc_21380_n4050_1;
  wire core__abc_21380_n4051;
  wire core__abc_21380_n4052;
  wire core__abc_21380_n4053;
  wire core__abc_21380_n4054_1;
  wire core__abc_21380_n4055;
  wire core__abc_21380_n4056;
  wire core__abc_21380_n4057_1;
  wire core__abc_21380_n4058;
  wire core__abc_21380_n4059;
  wire core__abc_21380_n4060;
  wire core__abc_21380_n4061;
  wire core__abc_21380_n4062_1;
  wire core__abc_21380_n4064;
  wire core__abc_21380_n4065;
  wire core__abc_21380_n4066;
  wire core__abc_21380_n4067_1;
  wire core__abc_21380_n4068;
  wire core__abc_21380_n4069;
  wire core__abc_21380_n4070;
  wire core__abc_21380_n4071;
  wire core__abc_21380_n4072_1;
  wire core__abc_21380_n4073;
  wire core__abc_21380_n4074;
  wire core__abc_21380_n4075;
  wire core__abc_21380_n4076_1;
  wire core__abc_21380_n4077;
  wire core__abc_21380_n4078;
  wire core__abc_21380_n4079;
  wire core__abc_21380_n4080_1;
  wire core__abc_21380_n4081;
  wire core__abc_21380_n4082_1;
  wire core__abc_21380_n4083;
  wire core__abc_21380_n4084;
  wire core__abc_21380_n4085;
  wire core__abc_21380_n4086;
  wire core__abc_21380_n4087_1;
  wire core__abc_21380_n4088;
  wire core__abc_21380_n4089;
  wire core__abc_21380_n4090;
  wire core__abc_21380_n4091_1;
  wire core__abc_21380_n4092;
  wire core__abc_21380_n4093;
  wire core__abc_21380_n4094;
  wire core__abc_21380_n4095_1;
  wire core__abc_21380_n4096;
  wire core__abc_21380_n4097;
  wire core__abc_21380_n4098_1;
  wire core__abc_21380_n4099;
  wire core__abc_21380_n4100;
  wire core__abc_21380_n4101;
  wire core__abc_21380_n4102_1;
  wire core__abc_21380_n4103;
  wire core__abc_21380_n4104;
  wire core__abc_21380_n4105;
  wire core__abc_21380_n4106_1;
  wire core__abc_21380_n4107;
  wire core__abc_21380_n4108;
  wire core__abc_21380_n4109;
  wire core__abc_21380_n4110;
  wire core__abc_21380_n4111_1;
  wire core__abc_21380_n4112;
  wire core__abc_21380_n4113;
  wire core__abc_21380_n4114;
  wire core__abc_21380_n4115_1;
  wire core__abc_21380_n4116;
  wire core__abc_21380_n4117;
  wire core__abc_21380_n4118;
  wire core__abc_21380_n4119;
  wire core__abc_21380_n4120_1;
  wire core__abc_21380_n4121;
  wire core__abc_21380_n4122;
  wire core__abc_21380_n4123;
  wire core__abc_21380_n4124_1;
  wire core__abc_21380_n4125;
  wire core__abc_21380_n4126;
  wire core__abc_21380_n4127;
  wire core__abc_21380_n4128;
  wire core__abc_21380_n4129_1;
  wire core__abc_21380_n4130;
  wire core__abc_21380_n4131;
  wire core__abc_21380_n4132;
  wire core__abc_21380_n4133_1;
  wire core__abc_21380_n4134;
  wire core__abc_21380_n4135;
  wire core__abc_21380_n4136;
  wire core__abc_21380_n4137;
  wire core__abc_21380_n4138_1;
  wire core__abc_21380_n4139;
  wire core__abc_21380_n4140;
  wire core__abc_21380_n4141_1;
  wire core__abc_21380_n4142;
  wire core__abc_21380_n4143;
  wire core__abc_21380_n4144;
  wire core__abc_21380_n4145_1;
  wire core__abc_21380_n4146;
  wire core__abc_21380_n4147;
  wire core__abc_21380_n4148;
  wire core__abc_21380_n4149_1;
  wire core__abc_21380_n4150;
  wire core__abc_21380_n4152;
  wire core__abc_21380_n4153_1;
  wire core__abc_21380_n4154;
  wire core__abc_21380_n4155;
  wire core__abc_21380_n4156;
  wire core__abc_21380_n4157_1;
  wire core__abc_21380_n4158;
  wire core__abc_21380_n4159;
  wire core__abc_21380_n4160;
  wire core__abc_21380_n4161_1;
  wire core__abc_21380_n4162;
  wire core__abc_21380_n4163;
  wire core__abc_21380_n4164;
  wire core__abc_21380_n4165_1;
  wire core__abc_21380_n4166;
  wire core__abc_21380_n4167;
  wire core__abc_21380_n4168;
  wire core__abc_21380_n4169;
  wire core__abc_21380_n4170_1;
  wire core__abc_21380_n4171;
  wire core__abc_21380_n4172;
  wire core__abc_21380_n4173_1;
  wire core__abc_21380_n4174;
  wire core__abc_21380_n4175;
  wire core__abc_21380_n4176;
  wire core__abc_21380_n4177;
  wire core__abc_21380_n4178_1;
  wire core__abc_21380_n4179;
  wire core__abc_21380_n4180;
  wire core__abc_21380_n4181;
  wire core__abc_21380_n4182_1;
  wire core__abc_21380_n4183;
  wire core__abc_21380_n4184;
  wire core__abc_21380_n4185;
  wire core__abc_21380_n4186_1;
  wire core__abc_21380_n4187;
  wire core__abc_21380_n4188;
  wire core__abc_21380_n4189_1;
  wire core__abc_21380_n4190;
  wire core__abc_21380_n4191;
  wire core__abc_21380_n4192;
  wire core__abc_21380_n4193;
  wire core__abc_21380_n4194_1;
  wire core__abc_21380_n4195;
  wire core__abc_21380_n4196;
  wire core__abc_21380_n4197;
  wire core__abc_21380_n4198_1;
  wire core__abc_21380_n4199;
  wire core__abc_21380_n4200;
  wire core__abc_21380_n4201;
  wire core__abc_21380_n4202;
  wire core__abc_21380_n4203_1;
  wire core__abc_21380_n4204;
  wire core__abc_21380_n4205;
  wire core__abc_21380_n4206_1;
  wire core__abc_21380_n4207;
  wire core__abc_21380_n4208;
  wire core__abc_21380_n4209;
  wire core__abc_21380_n4210_1;
  wire core__abc_21380_n4211;
  wire core__abc_21380_n4212;
  wire core__abc_21380_n4213;
  wire core__abc_21380_n4214;
  wire core__abc_21380_n4215;
  wire core__abc_21380_n4216;
  wire core__abc_21380_n4217;
  wire core__abc_21380_n4218_1;
  wire core__abc_21380_n4219;
  wire core__abc_21380_n4220;
  wire core__abc_21380_n4222;
  wire core__abc_21380_n4223;
  wire core__abc_21380_n4224_1;
  wire core__abc_21380_n4225;
  wire core__abc_21380_n4226;
  wire core__abc_21380_n4227;
  wire core__abc_21380_n4228;
  wire core__abc_21380_n4229;
  wire core__abc_21380_n4230_1;
  wire core__abc_21380_n4231;
  wire core__abc_21380_n4232;
  wire core__abc_21380_n4233;
  wire core__abc_21380_n4234;
  wire core__abc_21380_n4235;
  wire core__abc_21380_n4236;
  wire core__abc_21380_n4237_1;
  wire core__abc_21380_n4238;
  wire core__abc_21380_n4239;
  wire core__abc_21380_n4240;
  wire core__abc_21380_n4241;
  wire core__abc_21380_n4242;
  wire core__abc_21380_n4243_1;
  wire core__abc_21380_n4244;
  wire core__abc_21380_n4245;
  wire core__abc_21380_n4246;
  wire core__abc_21380_n4247;
  wire core__abc_21380_n4248;
  wire core__abc_21380_n4249_1;
  wire core__abc_21380_n4250;
  wire core__abc_21380_n4251;
  wire core__abc_21380_n4252;
  wire core__abc_21380_n4253;
  wire core__abc_21380_n4254;
  wire core__abc_21380_n4255_1;
  wire core__abc_21380_n4256;
  wire core__abc_21380_n4257;
  wire core__abc_21380_n4258;
  wire core__abc_21380_n4259;
  wire core__abc_21380_n4260;
  wire core__abc_21380_n4261;
  wire core__abc_21380_n4262_1;
  wire core__abc_21380_n4263;
  wire core__abc_21380_n4264;
  wire core__abc_21380_n4265;
  wire core__abc_21380_n4266;
  wire core__abc_21380_n4267_1;
  wire core__abc_21380_n4268;
  wire core__abc_21380_n4269;
  wire core__abc_21380_n4270;
  wire core__abc_21380_n4271;
  wire core__abc_21380_n4272;
  wire core__abc_21380_n4273_1;
  wire core__abc_21380_n4274;
  wire core__abc_21380_n4275;
  wire core__abc_21380_n4276;
  wire core__abc_21380_n4277;
  wire core__abc_21380_n4278_1;
  wire core__abc_21380_n4279;
  wire core__abc_21380_n4280;
  wire core__abc_21380_n4281;
  wire core__abc_21380_n4282;
  wire core__abc_21380_n4283;
  wire core__abc_21380_n4284_1;
  wire core__abc_21380_n4285;
  wire core__abc_21380_n4286;
  wire core__abc_21380_n4287;
  wire core__abc_21380_n4288;
  wire core__abc_21380_n4289_1;
  wire core__abc_21380_n4290;
  wire core__abc_21380_n4292;
  wire core__abc_21380_n4293;
  wire core__abc_21380_n4294_1;
  wire core__abc_21380_n4295;
  wire core__abc_21380_n4296;
  wire core__abc_21380_n4297;
  wire core__abc_21380_n4298;
  wire core__abc_21380_n4299_1;
  wire core__abc_21380_n4300;
  wire core__abc_21380_n4301;
  wire core__abc_21380_n4302;
  wire core__abc_21380_n4303;
  wire core__abc_21380_n4304_1;
  wire core__abc_21380_n4305;
  wire core__abc_21380_n4306;
  wire core__abc_21380_n4307;
  wire core__abc_21380_n4308;
  wire core__abc_21380_n4309_1;
  wire core__abc_21380_n4310;
  wire core__abc_21380_n4311;
  wire core__abc_21380_n4312;
  wire core__abc_21380_n4313;
  wire core__abc_21380_n4314_1;
  wire core__abc_21380_n4315;
  wire core__abc_21380_n4316;
  wire core__abc_21380_n4317;
  wire core__abc_21380_n4318;
  wire core__abc_21380_n4319_1;
  wire core__abc_21380_n4320;
  wire core__abc_21380_n4321;
  wire core__abc_21380_n4322;
  wire core__abc_21380_n4323;
  wire core__abc_21380_n4324_1;
  wire core__abc_21380_n4325;
  wire core__abc_21380_n4326;
  wire core__abc_21380_n4327;
  wire core__abc_21380_n4328;
  wire core__abc_21380_n4329_1;
  wire core__abc_21380_n4330;
  wire core__abc_21380_n4331;
  wire core__abc_21380_n4332;
  wire core__abc_21380_n4333;
  wire core__abc_21380_n4334_1;
  wire core__abc_21380_n4335;
  wire core__abc_21380_n4336;
  wire core__abc_21380_n4337;
  wire core__abc_21380_n4338;
  wire core__abc_21380_n4339_1;
  wire core__abc_21380_n4340;
  wire core__abc_21380_n4341;
  wire core__abc_21380_n4342;
  wire core__abc_21380_n4343;
  wire core__abc_21380_n4344_1;
  wire core__abc_21380_n4345;
  wire core__abc_21380_n4346;
  wire core__abc_21380_n4347;
  wire core__abc_21380_n4348;
  wire core__abc_21380_n4349_1;
  wire core__abc_21380_n4351;
  wire core__abc_21380_n4352;
  wire core__abc_21380_n4353;
  wire core__abc_21380_n4354;
  wire core__abc_21380_n4355_1;
  wire core__abc_21380_n4356;
  wire core__abc_21380_n4357;
  wire core__abc_21380_n4358;
  wire core__abc_21380_n4359;
  wire core__abc_21380_n4360;
  wire core__abc_21380_n4361_1;
  wire core__abc_21380_n4362;
  wire core__abc_21380_n4363;
  wire core__abc_21380_n4364;
  wire core__abc_21380_n4365;
  wire core__abc_21380_n4366_1;
  wire core__abc_21380_n4367;
  wire core__abc_21380_n4368;
  wire core__abc_21380_n4369;
  wire core__abc_21380_n4370;
  wire core__abc_21380_n4371_1;
  wire core__abc_21380_n4372;
  wire core__abc_21380_n4373;
  wire core__abc_21380_n4374;
  wire core__abc_21380_n4375;
  wire core__abc_21380_n4376_1;
  wire core__abc_21380_n4377;
  wire core__abc_21380_n4378;
  wire core__abc_21380_n4379;
  wire core__abc_21380_n4380;
  wire core__abc_21380_n4381_1;
  wire core__abc_21380_n4382;
  wire core__abc_21380_n4383;
  wire core__abc_21380_n4384;
  wire core__abc_21380_n4385;
  wire core__abc_21380_n4386_1;
  wire core__abc_21380_n4387;
  wire core__abc_21380_n4388;
  wire core__abc_21380_n4389;
  wire core__abc_21380_n4390;
  wire core__abc_21380_n4391;
  wire core__abc_21380_n4392_1;
  wire core__abc_21380_n4393;
  wire core__abc_21380_n4394;
  wire core__abc_21380_n4395;
  wire core__abc_21380_n4396;
  wire core__abc_21380_n4397_1;
  wire core__abc_21380_n4398;
  wire core__abc_21380_n4399;
  wire core__abc_21380_n4400;
  wire core__abc_21380_n4401;
  wire core__abc_21380_n4402_1;
  wire core__abc_21380_n4403;
  wire core__abc_21380_n4404;
  wire core__abc_21380_n4405;
  wire core__abc_21380_n4406;
  wire core__abc_21380_n4407_1;
  wire core__abc_21380_n4408;
  wire core__abc_21380_n4409;
  wire core__abc_21380_n4410;
  wire core__abc_21380_n4411;
  wire core__abc_21380_n4412_1;
  wire core__abc_21380_n4413;
  wire core__abc_21380_n4414;
  wire core__abc_21380_n4415;
  wire core__abc_21380_n4416;
  wire core__abc_21380_n4417_1;
  wire core__abc_21380_n4418;
  wire core__abc_21380_n4419;
  wire core__abc_21380_n4420;
  wire core__abc_21380_n4421;
  wire core__abc_21380_n4422_1;
  wire core__abc_21380_n4423;
  wire core__abc_21380_n4424;
  wire core__abc_21380_n4425;
  wire core__abc_21380_n4426;
  wire core__abc_21380_n4427_1;
  wire core__abc_21380_n4428;
  wire core__abc_21380_n4429;
  wire core__abc_21380_n4430;
  wire core__abc_21380_n4431;
  wire core__abc_21380_n4432_1;
  wire core__abc_21380_n4433;
  wire core__abc_21380_n4434;
  wire core__abc_21380_n4435;
  wire core__abc_21380_n4436;
  wire core__abc_21380_n4437;
  wire core__abc_21380_n4438_1;
  wire core__abc_21380_n4439;
  wire core__abc_21380_n4440;
  wire core__abc_21380_n4441;
  wire core__abc_21380_n4442;
  wire core__abc_21380_n4443_1;
  wire core__abc_21380_n4444;
  wire core__abc_21380_n4446;
  wire core__abc_21380_n4447;
  wire core__abc_21380_n4448_1;
  wire core__abc_21380_n4449;
  wire core__abc_21380_n4450;
  wire core__abc_21380_n4451;
  wire core__abc_21380_n4452;
  wire core__abc_21380_n4453;
  wire core__abc_21380_n4454_1;
  wire core__abc_21380_n4455;
  wire core__abc_21380_n4456;
  wire core__abc_21380_n4457;
  wire core__abc_21380_n4458;
  wire core__abc_21380_n4459_1;
  wire core__abc_21380_n4460;
  wire core__abc_21380_n4461;
  wire core__abc_21380_n4462;
  wire core__abc_21380_n4463;
  wire core__abc_21380_n4464_1;
  wire core__abc_21380_n4465;
  wire core__abc_21380_n4466;
  wire core__abc_21380_n4467;
  wire core__abc_21380_n4468;
  wire core__abc_21380_n4469_1;
  wire core__abc_21380_n4470;
  wire core__abc_21380_n4471;
  wire core__abc_21380_n4472;
  wire core__abc_21380_n4473;
  wire core__abc_21380_n4474_1;
  wire core__abc_21380_n4475;
  wire core__abc_21380_n4476;
  wire core__abc_21380_n4477;
  wire core__abc_21380_n4478;
  wire core__abc_21380_n4479;
  wire core__abc_21380_n4480_1;
  wire core__abc_21380_n4481;
  wire core__abc_21380_n4482;
  wire core__abc_21380_n4483;
  wire core__abc_21380_n4484;
  wire core__abc_21380_n4485_1;
  wire core__abc_21380_n4486;
  wire core__abc_21380_n4487;
  wire core__abc_21380_n4488;
  wire core__abc_21380_n4489;
  wire core__abc_21380_n4490;
  wire core__abc_21380_n4491_1;
  wire core__abc_21380_n4492;
  wire core__abc_21380_n4493;
  wire core__abc_21380_n4494;
  wire core__abc_21380_n4495;
  wire core__abc_21380_n4496_1;
  wire core__abc_21380_n4497;
  wire core__abc_21380_n4498;
  wire core__abc_21380_n4499;
  wire core__abc_21380_n4500;
  wire core__abc_21380_n4501_1;
  wire core__abc_21380_n4502;
  wire core__abc_21380_n4503;
  wire core__abc_21380_n4504;
  wire core__abc_21380_n4505;
  wire core__abc_21380_n4506_1;
  wire core__abc_21380_n4507;
  wire core__abc_21380_n4508;
  wire core__abc_21380_n4509;
  wire core__abc_21380_n4510;
  wire core__abc_21380_n4511_1;
  wire core__abc_21380_n4513;
  wire core__abc_21380_n4514;
  wire core__abc_21380_n4515;
  wire core__abc_21380_n4516_1;
  wire core__abc_21380_n4517;
  wire core__abc_21380_n4518;
  wire core__abc_21380_n4519;
  wire core__abc_21380_n4520;
  wire core__abc_21380_n4521;
  wire core__abc_21380_n4522_1;
  wire core__abc_21380_n4523;
  wire core__abc_21380_n4524;
  wire core__abc_21380_n4525;
  wire core__abc_21380_n4526;
  wire core__abc_21380_n4527_1;
  wire core__abc_21380_n4528;
  wire core__abc_21380_n4529;
  wire core__abc_21380_n4530;
  wire core__abc_21380_n4531;
  wire core__abc_21380_n4532_1;
  wire core__abc_21380_n4533;
  wire core__abc_21380_n4534;
  wire core__abc_21380_n4535;
  wire core__abc_21380_n4536;
  wire core__abc_21380_n4537_1;
  wire core__abc_21380_n4538;
  wire core__abc_21380_n4539;
  wire core__abc_21380_n4540;
  wire core__abc_21380_n4541;
  wire core__abc_21380_n4542_1;
  wire core__abc_21380_n4543;
  wire core__abc_21380_n4544;
  wire core__abc_21380_n4545;
  wire core__abc_21380_n4546;
  wire core__abc_21380_n4547_1;
  wire core__abc_21380_n4548;
  wire core__abc_21380_n4549;
  wire core__abc_21380_n4550;
  wire core__abc_21380_n4551;
  wire core__abc_21380_n4552_1;
  wire core__abc_21380_n4553;
  wire core__abc_21380_n4554;
  wire core__abc_21380_n4555;
  wire core__abc_21380_n4556;
  wire core__abc_21380_n4557;
  wire core__abc_21380_n4558;
  wire core__abc_21380_n4559;
  wire core__abc_21380_n4560_1;
  wire core__abc_21380_n4561;
  wire core__abc_21380_n4562;
  wire core__abc_21380_n4563;
  wire core__abc_21380_n4564;
  wire core__abc_21380_n4565_1;
  wire core__abc_21380_n4566;
  wire core__abc_21380_n4567;
  wire core__abc_21380_n4568;
  wire core__abc_21380_n4569;
  wire core__abc_21380_n4570;
  wire core__abc_21380_n4571_1;
  wire core__abc_21380_n4572;
  wire core__abc_21380_n4574;
  wire core__abc_21380_n4575;
  wire core__abc_21380_n4576_1;
  wire core__abc_21380_n4577;
  wire core__abc_21380_n4578;
  wire core__abc_21380_n4579;
  wire core__abc_21380_n4580;
  wire core__abc_21380_n4581;
  wire core__abc_21380_n4582_1;
  wire core__abc_21380_n4583;
  wire core__abc_21380_n4584;
  wire core__abc_21380_n4585;
  wire core__abc_21380_n4586;
  wire core__abc_21380_n4587_1;
  wire core__abc_21380_n4588;
  wire core__abc_21380_n4589;
  wire core__abc_21380_n4590;
  wire core__abc_21380_n4591;
  wire core__abc_21380_n4592_1;
  wire core__abc_21380_n4593;
  wire core__abc_21380_n4594;
  wire core__abc_21380_n4595;
  wire core__abc_21380_n4596;
  wire core__abc_21380_n4597_1;
  wire core__abc_21380_n4598;
  wire core__abc_21380_n4599;
  wire core__abc_21380_n4600;
  wire core__abc_21380_n4601;
  wire core__abc_21380_n4602;
  wire core__abc_21380_n4603_1;
  wire core__abc_21380_n4604;
  wire core__abc_21380_n4605;
  wire core__abc_21380_n4606;
  wire core__abc_21380_n4607;
  wire core__abc_21380_n4608_1;
  wire core__abc_21380_n4609;
  wire core__abc_21380_n4610;
  wire core__abc_21380_n4611;
  wire core__abc_21380_n4612;
  wire core__abc_21380_n4613;
  wire core__abc_21380_n4614_1;
  wire core__abc_21380_n4615;
  wire core__abc_21380_n4616;
  wire core__abc_21380_n4617;
  wire core__abc_21380_n4618;
  wire core__abc_21380_n4619_1;
  wire core__abc_21380_n4620;
  wire core__abc_21380_n4621;
  wire core__abc_21380_n4622;
  wire core__abc_21380_n4623;
  wire core__abc_21380_n4624_1;
  wire core__abc_21380_n4625;
  wire core__abc_21380_n4626;
  wire core__abc_21380_n4627;
  wire core__abc_21380_n4628;
  wire core__abc_21380_n4629_1;
  wire core__abc_21380_n4630;
  wire core__abc_21380_n4632;
  wire core__abc_21380_n4633;
  wire core__abc_21380_n4634_1;
  wire core__abc_21380_n4635;
  wire core__abc_21380_n4636;
  wire core__abc_21380_n4637;
  wire core__abc_21380_n4638;
  wire core__abc_21380_n4639_1;
  wire core__abc_21380_n4640;
  wire core__abc_21380_n4641;
  wire core__abc_21380_n4642;
  wire core__abc_21380_n4643;
  wire core__abc_21380_n4644_1;
  wire core__abc_21380_n4645;
  wire core__abc_21380_n4646;
  wire core__abc_21380_n4647;
  wire core__abc_21380_n4648;
  wire core__abc_21380_n4649;
  wire core__abc_21380_n4650_1;
  wire core__abc_21380_n4651;
  wire core__abc_21380_n4652;
  wire core__abc_21380_n4653;
  wire core__abc_21380_n4654;
  wire core__abc_21380_n4655_1;
  wire core__abc_21380_n4656;
  wire core__abc_21380_n4657;
  wire core__abc_21380_n4658;
  wire core__abc_21380_n4659;
  wire core__abc_21380_n4660_1;
  wire core__abc_21380_n4661;
  wire core__abc_21380_n4662;
  wire core__abc_21380_n4663;
  wire core__abc_21380_n4664;
  wire core__abc_21380_n4665;
  wire core__abc_21380_n4666_1;
  wire core__abc_21380_n4667;
  wire core__abc_21380_n4668;
  wire core__abc_21380_n4669;
  wire core__abc_21380_n4670;
  wire core__abc_21380_n4671_1;
  wire core__abc_21380_n4672;
  wire core__abc_21380_n4673;
  wire core__abc_21380_n4674;
  wire core__abc_21380_n4675;
  wire core__abc_21380_n4676_1;
  wire core__abc_21380_n4677;
  wire core__abc_21380_n4678;
  wire core__abc_21380_n4679;
  wire core__abc_21380_n4680;
  wire core__abc_21380_n4681_1;
  wire core__abc_21380_n4682;
  wire core__abc_21380_n4683;
  wire core__abc_21380_n4684;
  wire core__abc_21380_n4685;
  wire core__abc_21380_n4686_1;
  wire core__abc_21380_n4687;
  wire core__abc_21380_n4688;
  wire core__abc_21380_n4689;
  wire core__abc_21380_n4690;
  wire core__abc_21380_n4691_1;
  wire core__abc_21380_n4692;
  wire core__abc_21380_n4693;
  wire core__abc_21380_n4694;
  wire core__abc_21380_n4695;
  wire core__abc_21380_n4696_1;
  wire core__abc_21380_n4697;
  wire core__abc_21380_n4698;
  wire core__abc_21380_n4699;
  wire core__abc_21380_n4700;
  wire core__abc_21380_n4701_1;
  wire core__abc_21380_n4702;
  wire core__abc_21380_n4703;
  wire core__abc_21380_n4704;
  wire core__abc_21380_n4706;
  wire core__abc_21380_n4707_1;
  wire core__abc_21380_n4708;
  wire core__abc_21380_n4709;
  wire core__abc_21380_n4710;
  wire core__abc_21380_n4711;
  wire core__abc_21380_n4712_1;
  wire core__abc_21380_n4713;
  wire core__abc_21380_n4714;
  wire core__abc_21380_n4715;
  wire core__abc_21380_n4716;
  wire core__abc_21380_n4717_1;
  wire core__abc_21380_n4718;
  wire core__abc_21380_n4719;
  wire core__abc_21380_n4720;
  wire core__abc_21380_n4721;
  wire core__abc_21380_n4722_1;
  wire core__abc_21380_n4723;
  wire core__abc_21380_n4724;
  wire core__abc_21380_n4725;
  wire core__abc_21380_n4726;
  wire core__abc_21380_n4727_1;
  wire core__abc_21380_n4728;
  wire core__abc_21380_n4729;
  wire core__abc_21380_n4730;
  wire core__abc_21380_n4731;
  wire core__abc_21380_n4732_1;
  wire core__abc_21380_n4733;
  wire core__abc_21380_n4734;
  wire core__abc_21380_n4735;
  wire core__abc_21380_n4736;
  wire core__abc_21380_n4737_1;
  wire core__abc_21380_n4738;
  wire core__abc_21380_n4739;
  wire core__abc_21380_n4740;
  wire core__abc_21380_n4741;
  wire core__abc_21380_n4742_1;
  wire core__abc_21380_n4743;
  wire core__abc_21380_n4744;
  wire core__abc_21380_n4745;
  wire core__abc_21380_n4746;
  wire core__abc_21380_n4747_1;
  wire core__abc_21380_n4749;
  wire core__abc_21380_n4750;
  wire core__abc_21380_n4751;
  wire core__abc_21380_n4752_1;
  wire core__abc_21380_n4753;
  wire core__abc_21380_n4754;
  wire core__abc_21380_n4755;
  wire core__abc_21380_n4756;
  wire core__abc_21380_n4757_1;
  wire core__abc_21380_n4758;
  wire core__abc_21380_n4759;
  wire core__abc_21380_n4760;
  wire core__abc_21380_n4761;
  wire core__abc_21380_n4762_1;
  wire core__abc_21380_n4763;
  wire core__abc_21380_n4764;
  wire core__abc_21380_n4765;
  wire core__abc_21380_n4766;
  wire core__abc_21380_n4767_1;
  wire core__abc_21380_n4768;
  wire core__abc_21380_n4769;
  wire core__abc_21380_n4770;
  wire core__abc_21380_n4771;
  wire core__abc_21380_n4772_1;
  wire core__abc_21380_n4773;
  wire core__abc_21380_n4774;
  wire core__abc_21380_n4775;
  wire core__abc_21380_n4776;
  wire core__abc_21380_n4777_1;
  wire core__abc_21380_n4778;
  wire core__abc_21380_n4779;
  wire core__abc_21380_n4780;
  wire core__abc_21380_n4781;
  wire core__abc_21380_n4782;
  wire core__abc_21380_n4783_1;
  wire core__abc_21380_n4784;
  wire core__abc_21380_n4785;
  wire core__abc_21380_n4786;
  wire core__abc_21380_n4787;
  wire core__abc_21380_n4788_1;
  wire core__abc_21380_n4789;
  wire core__abc_21380_n4790;
  wire core__abc_21380_n4791;
  wire core__abc_21380_n4792;
  wire core__abc_21380_n4793_1;
  wire core__abc_21380_n4794;
  wire core__abc_21380_n4795;
  wire core__abc_21380_n4796;
  wire core__abc_21380_n4797;
  wire core__abc_21380_n4798_1;
  wire core__abc_21380_n4799;
  wire core__abc_21380_n4800;
  wire core__abc_21380_n4802;
  wire core__abc_21380_n4803_1;
  wire core__abc_21380_n4804;
  wire core__abc_21380_n4805;
  wire core__abc_21380_n4806;
  wire core__abc_21380_n4807;
  wire core__abc_21380_n4808_1;
  wire core__abc_21380_n4809;
  wire core__abc_21380_n4810;
  wire core__abc_21380_n4811;
  wire core__abc_21380_n4812;
  wire core__abc_21380_n4813;
  wire core__abc_21380_n4814_1;
  wire core__abc_21380_n4815;
  wire core__abc_21380_n4816;
  wire core__abc_21380_n4817;
  wire core__abc_21380_n4818;
  wire core__abc_21380_n4819;
  wire core__abc_21380_n4820_1;
  wire core__abc_21380_n4821;
  wire core__abc_21380_n4822;
  wire core__abc_21380_n4823;
  wire core__abc_21380_n4824;
  wire core__abc_21380_n4825_1;
  wire core__abc_21380_n4826;
  wire core__abc_21380_n4827;
  wire core__abc_21380_n4828;
  wire core__abc_21380_n4829;
  wire core__abc_21380_n4830_1;
  wire core__abc_21380_n4831;
  wire core__abc_21380_n4832;
  wire core__abc_21380_n4833;
  wire core__abc_21380_n4834;
  wire core__abc_21380_n4835_1;
  wire core__abc_21380_n4836;
  wire core__abc_21380_n4837;
  wire core__abc_21380_n4838;
  wire core__abc_21380_n4839;
  wire core__abc_21380_n4840_1;
  wire core__abc_21380_n4841;
  wire core__abc_21380_n4842;
  wire core__abc_21380_n4843;
  wire core__abc_21380_n4844;
  wire core__abc_21380_n4845_1;
  wire core__abc_21380_n4846;
  wire core__abc_21380_n4847;
  wire core__abc_21380_n4848;
  wire core__abc_21380_n4850;
  wire core__abc_21380_n4851_1;
  wire core__abc_21380_n4852;
  wire core__abc_21380_n4853;
  wire core__abc_21380_n4854;
  wire core__abc_21380_n4855;
  wire core__abc_21380_n4856;
  wire core__abc_21380_n4857_1;
  wire core__abc_21380_n4858;
  wire core__abc_21380_n4859;
  wire core__abc_21380_n4860;
  wire core__abc_21380_n4861;
  wire core__abc_21380_n4862_1;
  wire core__abc_21380_n4863;
  wire core__abc_21380_n4864;
  wire core__abc_21380_n4865;
  wire core__abc_21380_n4866;
  wire core__abc_21380_n4867_1;
  wire core__abc_21380_n4868;
  wire core__abc_21380_n4869;
  wire core__abc_21380_n4870;
  wire core__abc_21380_n4871;
  wire core__abc_21380_n4872;
  wire core__abc_21380_n4873_1;
  wire core__abc_21380_n4874;
  wire core__abc_21380_n4875;
  wire core__abc_21380_n4876;
  wire core__abc_21380_n4877;
  wire core__abc_21380_n4878_1;
  wire core__abc_21380_n4879;
  wire core__abc_21380_n4880;
  wire core__abc_21380_n4881;
  wire core__abc_21380_n4882;
  wire core__abc_21380_n4883_1;
  wire core__abc_21380_n4884;
  wire core__abc_21380_n4885;
  wire core__abc_21380_n4886;
  wire core__abc_21380_n4887;
  wire core__abc_21380_n4888_1;
  wire core__abc_21380_n4889;
  wire core__abc_21380_n4890;
  wire core__abc_21380_n4891;
  wire core__abc_21380_n4892_1;
  wire core__abc_21380_n4893_1;
  wire core__abc_21380_n4894;
  wire core__abc_21380_n4895;
  wire core__abc_21380_n4896_1;
  wire core__abc_21380_n4897;
  wire core__abc_21380_n4898_1;
  wire core__abc_21380_n4899;
  wire core__abc_21380_n4900_1;
  wire core__abc_21380_n4901;
  wire core__abc_21380_n4902_1;
  wire core__abc_21380_n4903;
  wire core__abc_21380_n4904;
  wire core__abc_21380_n4905;
  wire core__abc_21380_n4906;
  wire core__abc_21380_n4907;
  wire core__abc_21380_n4908;
  wire core__abc_21380_n4909;
  wire core__abc_21380_n4910;
  wire core__abc_21380_n4911;
  wire core__abc_21380_n4912;
  wire core__abc_21380_n4913;
  wire core__abc_21380_n4914;
  wire core__abc_21380_n4915;
  wire core__abc_21380_n4916;
  wire core__abc_21380_n4917;
  wire core__abc_21380_n4918;
  wire core__abc_21380_n4919;
  wire core__abc_21380_n4920;
  wire core__abc_21380_n4921;
  wire core__abc_21380_n4922;
  wire core__abc_21380_n4923;
  wire core__abc_21380_n4924;
  wire core__abc_21380_n4926;
  wire core__abc_21380_n4927;
  wire core__abc_21380_n4928;
  wire core__abc_21380_n4929;
  wire core__abc_21380_n4930;
  wire core__abc_21380_n4931;
  wire core__abc_21380_n4932;
  wire core__abc_21380_n4933;
  wire core__abc_21380_n4934;
  wire core__abc_21380_n4935;
  wire core__abc_21380_n4936;
  wire core__abc_21380_n4937;
  wire core__abc_21380_n4938;
  wire core__abc_21380_n4939;
  wire core__abc_21380_n4940;
  wire core__abc_21380_n4941;
  wire core__abc_21380_n4942;
  wire core__abc_21380_n4943;
  wire core__abc_21380_n4944;
  wire core__abc_21380_n4945;
  wire core__abc_21380_n4946;
  wire core__abc_21380_n4947;
  wire core__abc_21380_n4948;
  wire core__abc_21380_n4949;
  wire core__abc_21380_n4950;
  wire core__abc_21380_n4951;
  wire core__abc_21380_n4952;
  wire core__abc_21380_n4953;
  wire core__abc_21380_n4954;
  wire core__abc_21380_n4955;
  wire core__abc_21380_n4956;
  wire core__abc_21380_n4957;
  wire core__abc_21380_n4958;
  wire core__abc_21380_n4959;
  wire core__abc_21380_n4960;
  wire core__abc_21380_n4961;
  wire core__abc_21380_n4962;
  wire core__abc_21380_n4963;
  wire core__abc_21380_n4964;
  wire core__abc_21380_n4965;
  wire core__abc_21380_n4966;
  wire core__abc_21380_n4967;
  wire core__abc_21380_n4968;
  wire core__abc_21380_n4969;
  wire core__abc_21380_n4970;
  wire core__abc_21380_n4971;
  wire core__abc_21380_n4973;
  wire core__abc_21380_n4974;
  wire core__abc_21380_n4975;
  wire core__abc_21380_n4976;
  wire core__abc_21380_n4977;
  wire core__abc_21380_n4978;
  wire core__abc_21380_n4979;
  wire core__abc_21380_n4980;
  wire core__abc_21380_n4981;
  wire core__abc_21380_n4982;
  wire core__abc_21380_n4983;
  wire core__abc_21380_n4984;
  wire core__abc_21380_n4985;
  wire core__abc_21380_n4986;
  wire core__abc_21380_n4987;
  wire core__abc_21380_n4988;
  wire core__abc_21380_n4989;
  wire core__abc_21380_n4990;
  wire core__abc_21380_n4991;
  wire core__abc_21380_n4992;
  wire core__abc_21380_n4993;
  wire core__abc_21380_n4994;
  wire core__abc_21380_n4995;
  wire core__abc_21380_n4996;
  wire core__abc_21380_n4997;
  wire core__abc_21380_n4998;
  wire core__abc_21380_n4999;
  wire core__abc_21380_n5000;
  wire core__abc_21380_n5001;
  wire core__abc_21380_n5002;
  wire core__abc_21380_n5003;
  wire core__abc_21380_n5004;
  wire core__abc_21380_n5005;
  wire core__abc_21380_n5006;
  wire core__abc_21380_n5007;
  wire core__abc_21380_n5008;
  wire core__abc_21380_n5009;
  wire core__abc_21380_n5010;
  wire core__abc_21380_n5011;
  wire core__abc_21380_n5012;
  wire core__abc_21380_n5013;
  wire core__abc_21380_n5014;
  wire core__abc_21380_n5015;
  wire core__abc_21380_n5016;
  wire core__abc_21380_n5017;
  wire core__abc_21380_n5018;
  wire core__abc_21380_n5019;
  wire core__abc_21380_n5020;
  wire core__abc_21380_n5022;
  wire core__abc_21380_n5023;
  wire core__abc_21380_n5024;
  wire core__abc_21380_n5025;
  wire core__abc_21380_n5026;
  wire core__abc_21380_n5027;
  wire core__abc_21380_n5028;
  wire core__abc_21380_n5029;
  wire core__abc_21380_n5030;
  wire core__abc_21380_n5031;
  wire core__abc_21380_n5032;
  wire core__abc_21380_n5033;
  wire core__abc_21380_n5034;
  wire core__abc_21380_n5035;
  wire core__abc_21380_n5036;
  wire core__abc_21380_n5037;
  wire core__abc_21380_n5038;
  wire core__abc_21380_n5039;
  wire core__abc_21380_n5040;
  wire core__abc_21380_n5041;
  wire core__abc_21380_n5042;
  wire core__abc_21380_n5043;
  wire core__abc_21380_n5044;
  wire core__abc_21380_n5045;
  wire core__abc_21380_n5046;
  wire core__abc_21380_n5047;
  wire core__abc_21380_n5048;
  wire core__abc_21380_n5049;
  wire core__abc_21380_n5050;
  wire core__abc_21380_n5051;
  wire core__abc_21380_n5052;
  wire core__abc_21380_n5053;
  wire core__abc_21380_n5054;
  wire core__abc_21380_n5055;
  wire core__abc_21380_n5056;
  wire core__abc_21380_n5057;
  wire core__abc_21380_n5058;
  wire core__abc_21380_n5059;
  wire core__abc_21380_n5060;
  wire core__abc_21380_n5061;
  wire core__abc_21380_n5062;
  wire core__abc_21380_n5063;
  wire core__abc_21380_n5064;
  wire core__abc_21380_n5065;
  wire core__abc_21380_n5066;
  wire core__abc_21380_n5067;
  wire core__abc_21380_n5068;
  wire core__abc_21380_n5069;
  wire core__abc_21380_n5070;
  wire core__abc_21380_n5071;
  wire core__abc_21380_n5073;
  wire core__abc_21380_n5074;
  wire core__abc_21380_n5075;
  wire core__abc_21380_n5076;
  wire core__abc_21380_n5077;
  wire core__abc_21380_n5078;
  wire core__abc_21380_n5079;
  wire core__abc_21380_n5080;
  wire core__abc_21380_n5081;
  wire core__abc_21380_n5082;
  wire core__abc_21380_n5083;
  wire core__abc_21380_n5084;
  wire core__abc_21380_n5085;
  wire core__abc_21380_n5086;
  wire core__abc_21380_n5087;
  wire core__abc_21380_n5088;
  wire core__abc_21380_n5089;
  wire core__abc_21380_n5090;
  wire core__abc_21380_n5091;
  wire core__abc_21380_n5092;
  wire core__abc_21380_n5093;
  wire core__abc_21380_n5094;
  wire core__abc_21380_n5095;
  wire core__abc_21380_n5096;
  wire core__abc_21380_n5097;
  wire core__abc_21380_n5098;
  wire core__abc_21380_n5099;
  wire core__abc_21380_n5100;
  wire core__abc_21380_n5101;
  wire core__abc_21380_n5102;
  wire core__abc_21380_n5103;
  wire core__abc_21380_n5104;
  wire core__abc_21380_n5105;
  wire core__abc_21380_n5106;
  wire core__abc_21380_n5107;
  wire core__abc_21380_n5108;
  wire core__abc_21380_n5109;
  wire core__abc_21380_n5110;
  wire core__abc_21380_n5111;
  wire core__abc_21380_n5112;
  wire core__abc_21380_n5113;
  wire core__abc_21380_n5114;
  wire core__abc_21380_n5115;
  wire core__abc_21380_n5116;
  wire core__abc_21380_n5117;
  wire core__abc_21380_n5118;
  wire core__abc_21380_n5119;
  wire core__abc_21380_n5120;
  wire core__abc_21380_n5121;
  wire core__abc_21380_n5122;
  wire core__abc_21380_n5123;
  wire core__abc_21380_n5124;
  wire core__abc_21380_n5125;
  wire core__abc_21380_n5126;
  wire core__abc_21380_n5127;
  wire core__abc_21380_n5128;
  wire core__abc_21380_n5129;
  wire core__abc_21380_n5130;
  wire core__abc_21380_n5131;
  wire core__abc_21380_n5132;
  wire core__abc_21380_n5133;
  wire core__abc_21380_n5134;
  wire core__abc_21380_n5135;
  wire core__abc_21380_n5136;
  wire core__abc_21380_n5137;
  wire core__abc_21380_n5139;
  wire core__abc_21380_n5140;
  wire core__abc_21380_n5141;
  wire core__abc_21380_n5142;
  wire core__abc_21380_n5143;
  wire core__abc_21380_n5144;
  wire core__abc_21380_n5145;
  wire core__abc_21380_n5146;
  wire core__abc_21380_n5147;
  wire core__abc_21380_n5148;
  wire core__abc_21380_n5149;
  wire core__abc_21380_n5150;
  wire core__abc_21380_n5151;
  wire core__abc_21380_n5152;
  wire core__abc_21380_n5153;
  wire core__abc_21380_n5154;
  wire core__abc_21380_n5155;
  wire core__abc_21380_n5156;
  wire core__abc_21380_n5157;
  wire core__abc_21380_n5158;
  wire core__abc_21380_n5159;
  wire core__abc_21380_n5160;
  wire core__abc_21380_n5161;
  wire core__abc_21380_n5162;
  wire core__abc_21380_n5163;
  wire core__abc_21380_n5164;
  wire core__abc_21380_n5165;
  wire core__abc_21380_n5166;
  wire core__abc_21380_n5167;
  wire core__abc_21380_n5168;
  wire core__abc_21380_n5169;
  wire core__abc_21380_n5170;
  wire core__abc_21380_n5171;
  wire core__abc_21380_n5172;
  wire core__abc_21380_n5173;
  wire core__abc_21380_n5174;
  wire core__abc_21380_n5175;
  wire core__abc_21380_n5176;
  wire core__abc_21380_n5177;
  wire core__abc_21380_n5178;
  wire core__abc_21380_n5179;
  wire core__abc_21380_n5180;
  wire core__abc_21380_n5181;
  wire core__abc_21380_n5182;
  wire core__abc_21380_n5183;
  wire core__abc_21380_n5184;
  wire core__abc_21380_n5185;
  wire core__abc_21380_n5186;
  wire core__abc_21380_n5187;
  wire core__abc_21380_n5188;
  wire core__abc_21380_n5189;
  wire core__abc_21380_n5190;
  wire core__abc_21380_n5191;
  wire core__abc_21380_n5192;
  wire core__abc_21380_n5193;
  wire core__abc_21380_n5195;
  wire core__abc_21380_n5196;
  wire core__abc_21380_n5197;
  wire core__abc_21380_n5198;
  wire core__abc_21380_n5199;
  wire core__abc_21380_n5200;
  wire core__abc_21380_n5201;
  wire core__abc_21380_n5202;
  wire core__abc_21380_n5203;
  wire core__abc_21380_n5204;
  wire core__abc_21380_n5205;
  wire core__abc_21380_n5206;
  wire core__abc_21380_n5207;
  wire core__abc_21380_n5208;
  wire core__abc_21380_n5209;
  wire core__abc_21380_n5210;
  wire core__abc_21380_n5211;
  wire core__abc_21380_n5212;
  wire core__abc_21380_n5213;
  wire core__abc_21380_n5214;
  wire core__abc_21380_n5215;
  wire core__abc_21380_n5216;
  wire core__abc_21380_n5217;
  wire core__abc_21380_n5218;
  wire core__abc_21380_n5219;
  wire core__abc_21380_n5220;
  wire core__abc_21380_n5221;
  wire core__abc_21380_n5222;
  wire core__abc_21380_n5223;
  wire core__abc_21380_n5224;
  wire core__abc_21380_n5225;
  wire core__abc_21380_n5226;
  wire core__abc_21380_n5227;
  wire core__abc_21380_n5228;
  wire core__abc_21380_n5229;
  wire core__abc_21380_n5230;
  wire core__abc_21380_n5231;
  wire core__abc_21380_n5232;
  wire core__abc_21380_n5233;
  wire core__abc_21380_n5234;
  wire core__abc_21380_n5235;
  wire core__abc_21380_n5236;
  wire core__abc_21380_n5237;
  wire core__abc_21380_n5238;
  wire core__abc_21380_n5239;
  wire core__abc_21380_n5240;
  wire core__abc_21380_n5241;
  wire core__abc_21380_n5242;
  wire core__abc_21380_n5243;
  wire core__abc_21380_n5244;
  wire core__abc_21380_n5246;
  wire core__abc_21380_n5247;
  wire core__abc_21380_n5248;
  wire core__abc_21380_n5249;
  wire core__abc_21380_n5250;
  wire core__abc_21380_n5251;
  wire core__abc_21380_n5252;
  wire core__abc_21380_n5253;
  wire core__abc_21380_n5254;
  wire core__abc_21380_n5255;
  wire core__abc_21380_n5256;
  wire core__abc_21380_n5257;
  wire core__abc_21380_n5258;
  wire core__abc_21380_n5259;
  wire core__abc_21380_n5260;
  wire core__abc_21380_n5261;
  wire core__abc_21380_n5262;
  wire core__abc_21380_n5263;
  wire core__abc_21380_n5264;
  wire core__abc_21380_n5265;
  wire core__abc_21380_n5266;
  wire core__abc_21380_n5267;
  wire core__abc_21380_n5268;
  wire core__abc_21380_n5269;
  wire core__abc_21380_n5270;
  wire core__abc_21380_n5271;
  wire core__abc_21380_n5272;
  wire core__abc_21380_n5273;
  wire core__abc_21380_n5274;
  wire core__abc_21380_n5275;
  wire core__abc_21380_n5276;
  wire core__abc_21380_n5277;
  wire core__abc_21380_n5278;
  wire core__abc_21380_n5279;
  wire core__abc_21380_n5280;
  wire core__abc_21380_n5281;
  wire core__abc_21380_n5282;
  wire core__abc_21380_n5283;
  wire core__abc_21380_n5284;
  wire core__abc_21380_n5285;
  wire core__abc_21380_n5286;
  wire core__abc_21380_n5287;
  wire core__abc_21380_n5288;
  wire core__abc_21380_n5289;
  wire core__abc_21380_n5290;
  wire core__abc_21380_n5291;
  wire core__abc_21380_n5292;
  wire core__abc_21380_n5293;
  wire core__abc_21380_n5294;
  wire core__abc_21380_n5295;
  wire core__abc_21380_n5296;
  wire core__abc_21380_n5297;
  wire core__abc_21380_n5299;
  wire core__abc_21380_n5300;
  wire core__abc_21380_n5301;
  wire core__abc_21380_n5302;
  wire core__abc_21380_n5303;
  wire core__abc_21380_n5304;
  wire core__abc_21380_n5305;
  wire core__abc_21380_n5306;
  wire core__abc_21380_n5307;
  wire core__abc_21380_n5308;
  wire core__abc_21380_n5309;
  wire core__abc_21380_n5310;
  wire core__abc_21380_n5311;
  wire core__abc_21380_n5312;
  wire core__abc_21380_n5313;
  wire core__abc_21380_n5314;
  wire core__abc_21380_n5315;
  wire core__abc_21380_n5316;
  wire core__abc_21380_n5317;
  wire core__abc_21380_n5318;
  wire core__abc_21380_n5319;
  wire core__abc_21380_n5320;
  wire core__abc_21380_n5321;
  wire core__abc_21380_n5322;
  wire core__abc_21380_n5323;
  wire core__abc_21380_n5324;
  wire core__abc_21380_n5325;
  wire core__abc_21380_n5326;
  wire core__abc_21380_n5327;
  wire core__abc_21380_n5328;
  wire core__abc_21380_n5329;
  wire core__abc_21380_n5330;
  wire core__abc_21380_n5331;
  wire core__abc_21380_n5332;
  wire core__abc_21380_n5333;
  wire core__abc_21380_n5334;
  wire core__abc_21380_n5335;
  wire core__abc_21380_n5336;
  wire core__abc_21380_n5337;
  wire core__abc_21380_n5338;
  wire core__abc_21380_n5339;
  wire core__abc_21380_n5340;
  wire core__abc_21380_n5341;
  wire core__abc_21380_n5342;
  wire core__abc_21380_n5343;
  wire core__abc_21380_n5344;
  wire core__abc_21380_n5345;
  wire core__abc_21380_n5346;
  wire core__abc_21380_n5347;
  wire core__abc_21380_n5348;
  wire core__abc_21380_n5349;
  wire core__abc_21380_n5350;
  wire core__abc_21380_n5351;
  wire core__abc_21380_n5352;
  wire core__abc_21380_n5353;
  wire core__abc_21380_n5354;
  wire core__abc_21380_n5355;
  wire core__abc_21380_n5356;
  wire core__abc_21380_n5357;
  wire core__abc_21380_n5358;
  wire core__abc_21380_n5359;
  wire core__abc_21380_n5360;
  wire core__abc_21380_n5361;
  wire core__abc_21380_n5362;
  wire core__abc_21380_n5363;
  wire core__abc_21380_n5364;
  wire core__abc_21380_n5365;
  wire core__abc_21380_n5366;
  wire core__abc_21380_n5367;
  wire core__abc_21380_n5368;
  wire core__abc_21380_n5369;
  wire core__abc_21380_n5370;
  wire core__abc_21380_n5371;
  wire core__abc_21380_n5372;
  wire core__abc_21380_n5374;
  wire core__abc_21380_n5375;
  wire core__abc_21380_n5376;
  wire core__abc_21380_n5377;
  wire core__abc_21380_n5378;
  wire core__abc_21380_n5379;
  wire core__abc_21380_n5380;
  wire core__abc_21380_n5381;
  wire core__abc_21380_n5382;
  wire core__abc_21380_n5383;
  wire core__abc_21380_n5384;
  wire core__abc_21380_n5385;
  wire core__abc_21380_n5386;
  wire core__abc_21380_n5387;
  wire core__abc_21380_n5388;
  wire core__abc_21380_n5389;
  wire core__abc_21380_n5390;
  wire core__abc_21380_n5391;
  wire core__abc_21380_n5392;
  wire core__abc_21380_n5393;
  wire core__abc_21380_n5394;
  wire core__abc_21380_n5395;
  wire core__abc_21380_n5396;
  wire core__abc_21380_n5397;
  wire core__abc_21380_n5398;
  wire core__abc_21380_n5399;
  wire core__abc_21380_n5400;
  wire core__abc_21380_n5401;
  wire core__abc_21380_n5402;
  wire core__abc_21380_n5403;
  wire core__abc_21380_n5404;
  wire core__abc_21380_n5405;
  wire core__abc_21380_n5406;
  wire core__abc_21380_n5407;
  wire core__abc_21380_n5408;
  wire core__abc_21380_n5409;
  wire core__abc_21380_n5410;
  wire core__abc_21380_n5411;
  wire core__abc_21380_n5412;
  wire core__abc_21380_n5413;
  wire core__abc_21380_n5414;
  wire core__abc_21380_n5416;
  wire core__abc_21380_n5417;
  wire core__abc_21380_n5418;
  wire core__abc_21380_n5419;
  wire core__abc_21380_n5420;
  wire core__abc_21380_n5421;
  wire core__abc_21380_n5422;
  wire core__abc_21380_n5423;
  wire core__abc_21380_n5424;
  wire core__abc_21380_n5425;
  wire core__abc_21380_n5426;
  wire core__abc_21380_n5427;
  wire core__abc_21380_n5428;
  wire core__abc_21380_n5429;
  wire core__abc_21380_n5430;
  wire core__abc_21380_n5431;
  wire core__abc_21380_n5432;
  wire core__abc_21380_n5433;
  wire core__abc_21380_n5434;
  wire core__abc_21380_n5435;
  wire core__abc_21380_n5436;
  wire core__abc_21380_n5437;
  wire core__abc_21380_n5438;
  wire core__abc_21380_n5439;
  wire core__abc_21380_n5440;
  wire core__abc_21380_n5441;
  wire core__abc_21380_n5442;
  wire core__abc_21380_n5443;
  wire core__abc_21380_n5444;
  wire core__abc_21380_n5445;
  wire core__abc_21380_n5446;
  wire core__abc_21380_n5447;
  wire core__abc_21380_n5448;
  wire core__abc_21380_n5449;
  wire core__abc_21380_n5450;
  wire core__abc_21380_n5451;
  wire core__abc_21380_n5452;
  wire core__abc_21380_n5453;
  wire core__abc_21380_n5454;
  wire core__abc_21380_n5455;
  wire core__abc_21380_n5456;
  wire core__abc_21380_n5457;
  wire core__abc_21380_n5458;
  wire core__abc_21380_n5459;
  wire core__abc_21380_n5460;
  wire core__abc_21380_n5461;
  wire core__abc_21380_n5462;
  wire core__abc_21380_n5463;
  wire core__abc_21380_n5465;
  wire core__abc_21380_n5466;
  wire core__abc_21380_n5467;
  wire core__abc_21380_n5468;
  wire core__abc_21380_n5469;
  wire core__abc_21380_n5470;
  wire core__abc_21380_n5471;
  wire core__abc_21380_n5472;
  wire core__abc_21380_n5473;
  wire core__abc_21380_n5474;
  wire core__abc_21380_n5475;
  wire core__abc_21380_n5476;
  wire core__abc_21380_n5477;
  wire core__abc_21380_n5478;
  wire core__abc_21380_n5479;
  wire core__abc_21380_n5480;
  wire core__abc_21380_n5481;
  wire core__abc_21380_n5482;
  wire core__abc_21380_n5483;
  wire core__abc_21380_n5484;
  wire core__abc_21380_n5485;
  wire core__abc_21380_n5486;
  wire core__abc_21380_n5487;
  wire core__abc_21380_n5488;
  wire core__abc_21380_n5489;
  wire core__abc_21380_n5490;
  wire core__abc_21380_n5491;
  wire core__abc_21380_n5492;
  wire core__abc_21380_n5493;
  wire core__abc_21380_n5494;
  wire core__abc_21380_n5495;
  wire core__abc_21380_n5496;
  wire core__abc_21380_n5497;
  wire core__abc_21380_n5498;
  wire core__abc_21380_n5499;
  wire core__abc_21380_n5500;
  wire core__abc_21380_n5501;
  wire core__abc_21380_n5502;
  wire core__abc_21380_n5503;
  wire core__abc_21380_n5504;
  wire core__abc_21380_n5505;
  wire core__abc_21380_n5506;
  wire core__abc_21380_n5507;
  wire core__abc_21380_n5509;
  wire core__abc_21380_n5510;
  wire core__abc_21380_n5511;
  wire core__abc_21380_n5512;
  wire core__abc_21380_n5513;
  wire core__abc_21380_n5514;
  wire core__abc_21380_n5515;
  wire core__abc_21380_n5516;
  wire core__abc_21380_n5517;
  wire core__abc_21380_n5518;
  wire core__abc_21380_n5519;
  wire core__abc_21380_n5520;
  wire core__abc_21380_n5521;
  wire core__abc_21380_n5522;
  wire core__abc_21380_n5523;
  wire core__abc_21380_n5524;
  wire core__abc_21380_n5525;
  wire core__abc_21380_n5526;
  wire core__abc_21380_n5527;
  wire core__abc_21380_n5528;
  wire core__abc_21380_n5529;
  wire core__abc_21380_n5530;
  wire core__abc_21380_n5531;
  wire core__abc_21380_n5532;
  wire core__abc_21380_n5533;
  wire core__abc_21380_n5534;
  wire core__abc_21380_n5535;
  wire core__abc_21380_n5536;
  wire core__abc_21380_n5537;
  wire core__abc_21380_n5538;
  wire core__abc_21380_n5539;
  wire core__abc_21380_n5540;
  wire core__abc_21380_n5541;
  wire core__abc_21380_n5542;
  wire core__abc_21380_n5543;
  wire core__abc_21380_n5544;
  wire core__abc_21380_n5545;
  wire core__abc_21380_n5546;
  wire core__abc_21380_n5547;
  wire core__abc_21380_n5548;
  wire core__abc_21380_n5549;
  wire core__abc_21380_n5550;
  wire core__abc_21380_n5551;
  wire core__abc_21380_n5552;
  wire core__abc_21380_n5553;
  wire core__abc_21380_n5554;
  wire core__abc_21380_n5555;
  wire core__abc_21380_n5556;
  wire core__abc_21380_n5557;
  wire core__abc_21380_n5558;
  wire core__abc_21380_n5559;
  wire core__abc_21380_n5561;
  wire core__abc_21380_n5562;
  wire core__abc_21380_n5563;
  wire core__abc_21380_n5564;
  wire core__abc_21380_n5565;
  wire core__abc_21380_n5566;
  wire core__abc_21380_n5567;
  wire core__abc_21380_n5568;
  wire core__abc_21380_n5569;
  wire core__abc_21380_n5570;
  wire core__abc_21380_n5571;
  wire core__abc_21380_n5572;
  wire core__abc_21380_n5573;
  wire core__abc_21380_n5574;
  wire core__abc_21380_n5575;
  wire core__abc_21380_n5576;
  wire core__abc_21380_n5577;
  wire core__abc_21380_n5578;
  wire core__abc_21380_n5579;
  wire core__abc_21380_n5580;
  wire core__abc_21380_n5581;
  wire core__abc_21380_n5582;
  wire core__abc_21380_n5583;
  wire core__abc_21380_n5584;
  wire core__abc_21380_n5585;
  wire core__abc_21380_n5586;
  wire core__abc_21380_n5587;
  wire core__abc_21380_n5588;
  wire core__abc_21380_n5589;
  wire core__abc_21380_n5590;
  wire core__abc_21380_n5591;
  wire core__abc_21380_n5592;
  wire core__abc_21380_n5593;
  wire core__abc_21380_n5594;
  wire core__abc_21380_n5595;
  wire core__abc_21380_n5596;
  wire core__abc_21380_n5597;
  wire core__abc_21380_n5598;
  wire core__abc_21380_n5599;
  wire core__abc_21380_n5600;
  wire core__abc_21380_n5601;
  wire core__abc_21380_n5602;
  wire core__abc_21380_n5603;
  wire core__abc_21380_n5604;
  wire core__abc_21380_n5606;
  wire core__abc_21380_n5607;
  wire core__abc_21380_n5608;
  wire core__abc_21380_n5609;
  wire core__abc_21380_n5610;
  wire core__abc_21380_n5611;
  wire core__abc_21380_n5612;
  wire core__abc_21380_n5613;
  wire core__abc_21380_n5614;
  wire core__abc_21380_n5615;
  wire core__abc_21380_n5616;
  wire core__abc_21380_n5617;
  wire core__abc_21380_n5618;
  wire core__abc_21380_n5619;
  wire core__abc_21380_n5620;
  wire core__abc_21380_n5621;
  wire core__abc_21380_n5622;
  wire core__abc_21380_n5623;
  wire core__abc_21380_n5624;
  wire core__abc_21380_n5625;
  wire core__abc_21380_n5626;
  wire core__abc_21380_n5627;
  wire core__abc_21380_n5628;
  wire core__abc_21380_n5629;
  wire core__abc_21380_n5630;
  wire core__abc_21380_n5631;
  wire core__abc_21380_n5632;
  wire core__abc_21380_n5633;
  wire core__abc_21380_n5634;
  wire core__abc_21380_n5635;
  wire core__abc_21380_n5636;
  wire core__abc_21380_n5637;
  wire core__abc_21380_n5638;
  wire core__abc_21380_n5639;
  wire core__abc_21380_n5640;
  wire core__abc_21380_n5641;
  wire core__abc_21380_n5642;
  wire core__abc_21380_n5643;
  wire core__abc_21380_n5644;
  wire core__abc_21380_n5645;
  wire core__abc_21380_n5646;
  wire core__abc_21380_n5647;
  wire core__abc_21380_n5648;
  wire core__abc_21380_n5649;
  wire core__abc_21380_n5650;
  wire core__abc_21380_n5651;
  wire core__abc_21380_n5652;
  wire core__abc_21380_n5653;
  wire core__abc_21380_n5654;
  wire core__abc_21380_n5656;
  wire core__abc_21380_n5657;
  wire core__abc_21380_n5658;
  wire core__abc_21380_n5659;
  wire core__abc_21380_n5660;
  wire core__abc_21380_n5661;
  wire core__abc_21380_n5662;
  wire core__abc_21380_n5663;
  wire core__abc_21380_n5664;
  wire core__abc_21380_n5665;
  wire core__abc_21380_n5666;
  wire core__abc_21380_n5667;
  wire core__abc_21380_n5668;
  wire core__abc_21380_n5669;
  wire core__abc_21380_n5670;
  wire core__abc_21380_n5671;
  wire core__abc_21380_n5672;
  wire core__abc_21380_n5673;
  wire core__abc_21380_n5674;
  wire core__abc_21380_n5675;
  wire core__abc_21380_n5676;
  wire core__abc_21380_n5677;
  wire core__abc_21380_n5678;
  wire core__abc_21380_n5679;
  wire core__abc_21380_n5680;
  wire core__abc_21380_n5681;
  wire core__abc_21380_n5682;
  wire core__abc_21380_n5683;
  wire core__abc_21380_n5684;
  wire core__abc_21380_n5685;
  wire core__abc_21380_n5686;
  wire core__abc_21380_n5687;
  wire core__abc_21380_n5688;
  wire core__abc_21380_n5689;
  wire core__abc_21380_n5690;
  wire core__abc_21380_n5691;
  wire core__abc_21380_n5692;
  wire core__abc_21380_n5693;
  wire core__abc_21380_n5694;
  wire core__abc_21380_n5695;
  wire core__abc_21380_n5696;
  wire core__abc_21380_n5697;
  wire core__abc_21380_n5698;
  wire core__abc_21380_n5699;
  wire core__abc_21380_n5700;
  wire core__abc_21380_n5701;
  wire core__abc_21380_n5703;
  wire core__abc_21380_n5704;
  wire core__abc_21380_n5705;
  wire core__abc_21380_n5706;
  wire core__abc_21380_n5707;
  wire core__abc_21380_n5708;
  wire core__abc_21380_n5709;
  wire core__abc_21380_n5710;
  wire core__abc_21380_n5711;
  wire core__abc_21380_n5712;
  wire core__abc_21380_n5713;
  wire core__abc_21380_n5714;
  wire core__abc_21380_n5715;
  wire core__abc_21380_n5716;
  wire core__abc_21380_n5717;
  wire core__abc_21380_n5718;
  wire core__abc_21380_n5719;
  wire core__abc_21380_n5720;
  wire core__abc_21380_n5721;
  wire core__abc_21380_n5722;
  wire core__abc_21380_n5723;
  wire core__abc_21380_n5724;
  wire core__abc_21380_n5725;
  wire core__abc_21380_n5726;
  wire core__abc_21380_n5727;
  wire core__abc_21380_n5728;
  wire core__abc_21380_n5729;
  wire core__abc_21380_n5730;
  wire core__abc_21380_n5731;
  wire core__abc_21380_n5732;
  wire core__abc_21380_n5733;
  wire core__abc_21380_n5734;
  wire core__abc_21380_n5735;
  wire core__abc_21380_n5736;
  wire core__abc_21380_n5737;
  wire core__abc_21380_n5738;
  wire core__abc_21380_n5739;
  wire core__abc_21380_n5740;
  wire core__abc_21380_n5741;
  wire core__abc_21380_n5742;
  wire core__abc_21380_n5743;
  wire core__abc_21380_n5744;
  wire core__abc_21380_n5745;
  wire core__abc_21380_n5746;
  wire core__abc_21380_n5747;
  wire core__abc_21380_n5748;
  wire core__abc_21380_n5749;
  wire core__abc_21380_n5750;
  wire core__abc_21380_n5752;
  wire core__abc_21380_n5753;
  wire core__abc_21380_n5754;
  wire core__abc_21380_n5755;
  wire core__abc_21380_n5756;
  wire core__abc_21380_n5757;
  wire core__abc_21380_n5758;
  wire core__abc_21380_n5759;
  wire core__abc_21380_n5760;
  wire core__abc_21380_n5761;
  wire core__abc_21380_n5762;
  wire core__abc_21380_n5763;
  wire core__abc_21380_n5764;
  wire core__abc_21380_n5765;
  wire core__abc_21380_n5766;
  wire core__abc_21380_n5767;
  wire core__abc_21380_n5768;
  wire core__abc_21380_n5769;
  wire core__abc_21380_n5770;
  wire core__abc_21380_n5771;
  wire core__abc_21380_n5772;
  wire core__abc_21380_n5773;
  wire core__abc_21380_n5774;
  wire core__abc_21380_n5775;
  wire core__abc_21380_n5776;
  wire core__abc_21380_n5777;
  wire core__abc_21380_n5778;
  wire core__abc_21380_n5779;
  wire core__abc_21380_n5780;
  wire core__abc_21380_n5781;
  wire core__abc_21380_n5782;
  wire core__abc_21380_n5783;
  wire core__abc_21380_n5784;
  wire core__abc_21380_n5785;
  wire core__abc_21380_n5786;
  wire core__abc_21380_n5787;
  wire core__abc_21380_n5788;
  wire core__abc_21380_n5789;
  wire core__abc_21380_n5790;
  wire core__abc_21380_n5791;
  wire core__abc_21380_n5792;
  wire core__abc_21380_n5793;
  wire core__abc_21380_n5794;
  wire core__abc_21380_n5795;
  wire core__abc_21380_n5796;
  wire core__abc_21380_n5797;
  wire core__abc_21380_n5799;
  wire core__abc_21380_n5800;
  wire core__abc_21380_n5801;
  wire core__abc_21380_n5802;
  wire core__abc_21380_n5803;
  wire core__abc_21380_n5804;
  wire core__abc_21380_n5805;
  wire core__abc_21380_n5806;
  wire core__abc_21380_n5807;
  wire core__abc_21380_n5808;
  wire core__abc_21380_n5809;
  wire core__abc_21380_n5810;
  wire core__abc_21380_n5811;
  wire core__abc_21380_n5812;
  wire core__abc_21380_n5813;
  wire core__abc_21380_n5814;
  wire core__abc_21380_n5815;
  wire core__abc_21380_n5816;
  wire core__abc_21380_n5817;
  wire core__abc_21380_n5818;
  wire core__abc_21380_n5819;
  wire core__abc_21380_n5820;
  wire core__abc_21380_n5821;
  wire core__abc_21380_n5822;
  wire core__abc_21380_n5823;
  wire core__abc_21380_n5824;
  wire core__abc_21380_n5825;
  wire core__abc_21380_n5826;
  wire core__abc_21380_n5827;
  wire core__abc_21380_n5828;
  wire core__abc_21380_n5829;
  wire core__abc_21380_n5830;
  wire core__abc_21380_n5831;
  wire core__abc_21380_n5832;
  wire core__abc_21380_n5833;
  wire core__abc_21380_n5834;
  wire core__abc_21380_n5835;
  wire core__abc_21380_n5836;
  wire core__abc_21380_n5837;
  wire core__abc_21380_n5838;
  wire core__abc_21380_n5839;
  wire core__abc_21380_n5840;
  wire core__abc_21380_n5842;
  wire core__abc_21380_n5843;
  wire core__abc_21380_n5844;
  wire core__abc_21380_n5845;
  wire core__abc_21380_n5846;
  wire core__abc_21380_n5847;
  wire core__abc_21380_n5848;
  wire core__abc_21380_n5849;
  wire core__abc_21380_n5850;
  wire core__abc_21380_n5851;
  wire core__abc_21380_n5852;
  wire core__abc_21380_n5853;
  wire core__abc_21380_n5854;
  wire core__abc_21380_n5855;
  wire core__abc_21380_n5856;
  wire core__abc_21380_n5857;
  wire core__abc_21380_n5858;
  wire core__abc_21380_n5859;
  wire core__abc_21380_n5860;
  wire core__abc_21380_n5861;
  wire core__abc_21380_n5862;
  wire core__abc_21380_n5863;
  wire core__abc_21380_n5864;
  wire core__abc_21380_n5865;
  wire core__abc_21380_n5866;
  wire core__abc_21380_n5867;
  wire core__abc_21380_n5868;
  wire core__abc_21380_n5869;
  wire core__abc_21380_n5870;
  wire core__abc_21380_n5871;
  wire core__abc_21380_n5872;
  wire core__abc_21380_n5873;
  wire core__abc_21380_n5875;
  wire core__abc_21380_n5876;
  wire core__abc_21380_n5877;
  wire core__abc_21380_n5878;
  wire core__abc_21380_n5879;
  wire core__abc_21380_n5880;
  wire core__abc_21380_n5881;
  wire core__abc_21380_n5882;
  wire core__abc_21380_n5883;
  wire core__abc_21380_n5884;
  wire core__abc_21380_n5885;
  wire core__abc_21380_n5886;
  wire core__abc_21380_n5887;
  wire core__abc_21380_n5888;
  wire core__abc_21380_n5889;
  wire core__abc_21380_n5890;
  wire core__abc_21380_n5891;
  wire core__abc_21380_n5892;
  wire core__abc_21380_n5893;
  wire core__abc_21380_n5894;
  wire core__abc_21380_n5895;
  wire core__abc_21380_n5896;
  wire core__abc_21380_n5897;
  wire core__abc_21380_n5898;
  wire core__abc_21380_n5899;
  wire core__abc_21380_n5900;
  wire core__abc_21380_n5901;
  wire core__abc_21380_n5902;
  wire core__abc_21380_n5903;
  wire core__abc_21380_n5904;
  wire core__abc_21380_n5905;
  wire core__abc_21380_n5906;
  wire core__abc_21380_n5907;
  wire core__abc_21380_n5908;
  wire core__abc_21380_n5909;
  wire core__abc_21380_n5910;
  wire core__abc_21380_n5911;
  wire core__abc_21380_n5912;
  wire core__abc_21380_n5913;
  wire core__abc_21380_n5914;
  wire core__abc_21380_n5915;
  wire core__abc_21380_n5916;
  wire core__abc_21380_n5917;
  wire core__abc_21380_n5918;
  wire core__abc_21380_n5919;
  wire core__abc_21380_n5921;
  wire core__abc_21380_n5922;
  wire core__abc_21380_n5923;
  wire core__abc_21380_n5924;
  wire core__abc_21380_n5925;
  wire core__abc_21380_n5926;
  wire core__abc_21380_n5927;
  wire core__abc_21380_n5928;
  wire core__abc_21380_n5929;
  wire core__abc_21380_n5930;
  wire core__abc_21380_n5931;
  wire core__abc_21380_n5932;
  wire core__abc_21380_n5933;
  wire core__abc_21380_n5934;
  wire core__abc_21380_n5935;
  wire core__abc_21380_n5936;
  wire core__abc_21380_n5937;
  wire core__abc_21380_n5938;
  wire core__abc_21380_n5939;
  wire core__abc_21380_n5940;
  wire core__abc_21380_n5941;
  wire core__abc_21380_n5942;
  wire core__abc_21380_n5943;
  wire core__abc_21380_n5944;
  wire core__abc_21380_n5945;
  wire core__abc_21380_n5946;
  wire core__abc_21380_n5947;
  wire core__abc_21380_n5948;
  wire core__abc_21380_n5949;
  wire core__abc_21380_n5950;
  wire core__abc_21380_n5951;
  wire core__abc_21380_n5952;
  wire core__abc_21380_n5953;
  wire core__abc_21380_n5954;
  wire core__abc_21380_n5956;
  wire core__abc_21380_n5957;
  wire core__abc_21380_n5958;
  wire core__abc_21380_n5959;
  wire core__abc_21380_n5960;
  wire core__abc_21380_n5961;
  wire core__abc_21380_n5962;
  wire core__abc_21380_n5963;
  wire core__abc_21380_n5964;
  wire core__abc_21380_n5965;
  wire core__abc_21380_n5966;
  wire core__abc_21380_n5967;
  wire core__abc_21380_n5968;
  wire core__abc_21380_n5969;
  wire core__abc_21380_n5970;
  wire core__abc_21380_n5971;
  wire core__abc_21380_n5972;
  wire core__abc_21380_n5973;
  wire core__abc_21380_n5974;
  wire core__abc_21380_n5975;
  wire core__abc_21380_n5976;
  wire core__abc_21380_n5977;
  wire core__abc_21380_n5978;
  wire core__abc_21380_n5979;
  wire core__abc_21380_n5980;
  wire core__abc_21380_n5981;
  wire core__abc_21380_n5982;
  wire core__abc_21380_n5983;
  wire core__abc_21380_n5984;
  wire core__abc_21380_n5985;
  wire core__abc_21380_n5986;
  wire core__abc_21380_n5987;
  wire core__abc_21380_n5988;
  wire core__abc_21380_n5989;
  wire core__abc_21380_n5990;
  wire core__abc_21380_n5991;
  wire core__abc_21380_n5992;
  wire core__abc_21380_n5993;
  wire core__abc_21380_n5994;
  wire core__abc_21380_n5996;
  wire core__abc_21380_n5997;
  wire core__abc_21380_n5998;
  wire core__abc_21380_n5999;
  wire core__abc_21380_n6000;
  wire core__abc_21380_n6001;
  wire core__abc_21380_n6002;
  wire core__abc_21380_n6003;
  wire core__abc_21380_n6004;
  wire core__abc_21380_n6005;
  wire core__abc_21380_n6006;
  wire core__abc_21380_n6007;
  wire core__abc_21380_n6008;
  wire core__abc_21380_n6009;
  wire core__abc_21380_n6010;
  wire core__abc_21380_n6011;
  wire core__abc_21380_n6012;
  wire core__abc_21380_n6013;
  wire core__abc_21380_n6014;
  wire core__abc_21380_n6015;
  wire core__abc_21380_n6016;
  wire core__abc_21380_n6017;
  wire core__abc_21380_n6018;
  wire core__abc_21380_n6019;
  wire core__abc_21380_n6020;
  wire core__abc_21380_n6021;
  wire core__abc_21380_n6022;
  wire core__abc_21380_n6023;
  wire core__abc_21380_n6024;
  wire core__abc_21380_n6025;
  wire core__abc_21380_n6026;
  wire core__abc_21380_n6027;
  wire core__abc_21380_n6028;
  wire core__abc_21380_n6030;
  wire core__abc_21380_n6031;
  wire core__abc_21380_n6032;
  wire core__abc_21380_n6033;
  wire core__abc_21380_n6034;
  wire core__abc_21380_n6035;
  wire core__abc_21380_n6036;
  wire core__abc_21380_n6037;
  wire core__abc_21380_n6038;
  wire core__abc_21380_n6039;
  wire core__abc_21380_n6040;
  wire core__abc_21380_n6041;
  wire core__abc_21380_n6042;
  wire core__abc_21380_n6043;
  wire core__abc_21380_n6044;
  wire core__abc_21380_n6045;
  wire core__abc_21380_n6046;
  wire core__abc_21380_n6047;
  wire core__abc_21380_n6048;
  wire core__abc_21380_n6049;
  wire core__abc_21380_n6050;
  wire core__abc_21380_n6051;
  wire core__abc_21380_n6052;
  wire core__abc_21380_n6053;
  wire core__abc_21380_n6054;
  wire core__abc_21380_n6055;
  wire core__abc_21380_n6056;
  wire core__abc_21380_n6057;
  wire core__abc_21380_n6058;
  wire core__abc_21380_n6059;
  wire core__abc_21380_n6060;
  wire core__abc_21380_n6061;
  wire core__abc_21380_n6062;
  wire core__abc_21380_n6063;
  wire core__abc_21380_n6064;
  wire core__abc_21380_n6065;
  wire core__abc_21380_n6066;
  wire core__abc_21380_n6067;
  wire core__abc_21380_n6068;
  wire core__abc_21380_n6069;
  wire core__abc_21380_n6070;
  wire core__abc_21380_n6071;
  wire core__abc_21380_n6072;
  wire core__abc_21380_n6073;
  wire core__abc_21380_n6074;
  wire core__abc_21380_n6075;
  wire core__abc_21380_n6076;
  wire core__abc_21380_n6077;
  wire core__abc_21380_n6078;
  wire core__abc_21380_n6079;
  wire core__abc_21380_n6080;
  wire core__abc_21380_n6081;
  wire core__abc_21380_n6082;
  wire core__abc_21380_n6083;
  wire core__abc_21380_n6084;
  wire core__abc_21380_n6085;
  wire core__abc_21380_n6086;
  wire core__abc_21380_n6087;
  wire core__abc_21380_n6088;
  wire core__abc_21380_n6089;
  wire core__abc_21380_n6090;
  wire core__abc_21380_n6091;
  wire core__abc_21380_n6092;
  wire core__abc_21380_n6094;
  wire core__abc_21380_n6095;
  wire core__abc_21380_n6096;
  wire core__abc_21380_n6097;
  wire core__abc_21380_n6098;
  wire core__abc_21380_n6099;
  wire core__abc_21380_n6100;
  wire core__abc_21380_n6101;
  wire core__abc_21380_n6102;
  wire core__abc_21380_n6103;
  wire core__abc_21380_n6104;
  wire core__abc_21380_n6105;
  wire core__abc_21380_n6106;
  wire core__abc_21380_n6107;
  wire core__abc_21380_n6108;
  wire core__abc_21380_n6109;
  wire core__abc_21380_n6110;
  wire core__abc_21380_n6111;
  wire core__abc_21380_n6112;
  wire core__abc_21380_n6113;
  wire core__abc_21380_n6114;
  wire core__abc_21380_n6115;
  wire core__abc_21380_n6116;
  wire core__abc_21380_n6117;
  wire core__abc_21380_n6118;
  wire core__abc_21380_n6119;
  wire core__abc_21380_n6120;
  wire core__abc_21380_n6121;
  wire core__abc_21380_n6122;
  wire core__abc_21380_n6123;
  wire core__abc_21380_n6124;
  wire core__abc_21380_n6125;
  wire core__abc_21380_n6126;
  wire core__abc_21380_n6127;
  wire core__abc_21380_n6128;
  wire core__abc_21380_n6130;
  wire core__abc_21380_n6131;
  wire core__abc_21380_n6132;
  wire core__abc_21380_n6133;
  wire core__abc_21380_n6134;
  wire core__abc_21380_n6135;
  wire core__abc_21380_n6136;
  wire core__abc_21380_n6137;
  wire core__abc_21380_n6138;
  wire core__abc_21380_n6139;
  wire core__abc_21380_n6140;
  wire core__abc_21380_n6141;
  wire core__abc_21380_n6142;
  wire core__abc_21380_n6143;
  wire core__abc_21380_n6144;
  wire core__abc_21380_n6145;
  wire core__abc_21380_n6146;
  wire core__abc_21380_n6147;
  wire core__abc_21380_n6148;
  wire core__abc_21380_n6149;
  wire core__abc_21380_n6150;
  wire core__abc_21380_n6151;
  wire core__abc_21380_n6152;
  wire core__abc_21380_n6153;
  wire core__abc_21380_n6154;
  wire core__abc_21380_n6155;
  wire core__abc_21380_n6156;
  wire core__abc_21380_n6157;
  wire core__abc_21380_n6158;
  wire core__abc_21380_n6159;
  wire core__abc_21380_n6160;
  wire core__abc_21380_n6161;
  wire core__abc_21380_n6162;
  wire core__abc_21380_n6163;
  wire core__abc_21380_n6164;
  wire core__abc_21380_n6165;
  wire core__abc_21380_n6166;
  wire core__abc_21380_n6167;
  wire core__abc_21380_n6169;
  wire core__abc_21380_n6170;
  wire core__abc_21380_n6171;
  wire core__abc_21380_n6172;
  wire core__abc_21380_n6173;
  wire core__abc_21380_n6174;
  wire core__abc_21380_n6175;
  wire core__abc_21380_n6176;
  wire core__abc_21380_n6177;
  wire core__abc_21380_n6178;
  wire core__abc_21380_n6179;
  wire core__abc_21380_n6180;
  wire core__abc_21380_n6181;
  wire core__abc_21380_n6182;
  wire core__abc_21380_n6183;
  wire core__abc_21380_n6184;
  wire core__abc_21380_n6185;
  wire core__abc_21380_n6186;
  wire core__abc_21380_n6187;
  wire core__abc_21380_n6188;
  wire core__abc_21380_n6189;
  wire core__abc_21380_n6190;
  wire core__abc_21380_n6191;
  wire core__abc_21380_n6192;
  wire core__abc_21380_n6193;
  wire core__abc_21380_n6194;
  wire core__abc_21380_n6195;
  wire core__abc_21380_n6196;
  wire core__abc_21380_n6197;
  wire core__abc_21380_n6198;
  wire core__abc_21380_n6199;
  wire core__abc_21380_n6200;
  wire core__abc_21380_n6201;
  wire core__abc_21380_n6203;
  wire core__abc_21380_n6204;
  wire core__abc_21380_n6205;
  wire core__abc_21380_n6206;
  wire core__abc_21380_n6207;
  wire core__abc_21380_n6208;
  wire core__abc_21380_n6209;
  wire core__abc_21380_n6210;
  wire core__abc_21380_n6211;
  wire core__abc_21380_n6212;
  wire core__abc_21380_n6213;
  wire core__abc_21380_n6214;
  wire core__abc_21380_n6215;
  wire core__abc_21380_n6216;
  wire core__abc_21380_n6217;
  wire core__abc_21380_n6218;
  wire core__abc_21380_n6219;
  wire core__abc_21380_n6220;
  wire core__abc_21380_n6221;
  wire core__abc_21380_n6222;
  wire core__abc_21380_n6223;
  wire core__abc_21380_n6224;
  wire core__abc_21380_n6225;
  wire core__abc_21380_n6226;
  wire core__abc_21380_n6227;
  wire core__abc_21380_n6228;
  wire core__abc_21380_n6229;
  wire core__abc_21380_n6230;
  wire core__abc_21380_n6231;
  wire core__abc_21380_n6232;
  wire core__abc_21380_n6233;
  wire core__abc_21380_n6234;
  wire core__abc_21380_n6235;
  wire core__abc_21380_n6236;
  wire core__abc_21380_n6237;
  wire core__abc_21380_n6238;
  wire core__abc_21380_n6239;
  wire core__abc_21380_n6240;
  wire core__abc_21380_n6241;
  wire core__abc_21380_n6243;
  wire core__abc_21380_n6244;
  wire core__abc_21380_n6245;
  wire core__abc_21380_n6246;
  wire core__abc_21380_n6247;
  wire core__abc_21380_n6248;
  wire core__abc_21380_n6249;
  wire core__abc_21380_n6250;
  wire core__abc_21380_n6251;
  wire core__abc_21380_n6252;
  wire core__abc_21380_n6253;
  wire core__abc_21380_n6254;
  wire core__abc_21380_n6255;
  wire core__abc_21380_n6256;
  wire core__abc_21380_n6257;
  wire core__abc_21380_n6258;
  wire core__abc_21380_n6259;
  wire core__abc_21380_n6260;
  wire core__abc_21380_n6261;
  wire core__abc_21380_n6262;
  wire core__abc_21380_n6263;
  wire core__abc_21380_n6264;
  wire core__abc_21380_n6265;
  wire core__abc_21380_n6266;
  wire core__abc_21380_n6267;
  wire core__abc_21380_n6268;
  wire core__abc_21380_n6269;
  wire core__abc_21380_n6270;
  wire core__abc_21380_n6271;
  wire core__abc_21380_n6272;
  wire core__abc_21380_n6273;
  wire core__abc_21380_n6274;
  wire core__abc_21380_n6276;
  wire core__abc_21380_n6277;
  wire core__abc_21380_n6278;
  wire core__abc_21380_n6279;
  wire core__abc_21380_n6280;
  wire core__abc_21380_n6281;
  wire core__abc_21380_n6282;
  wire core__abc_21380_n6283;
  wire core__abc_21380_n6284;
  wire core__abc_21380_n6285;
  wire core__abc_21380_n6286;
  wire core__abc_21380_n6287;
  wire core__abc_21380_n6288;
  wire core__abc_21380_n6289;
  wire core__abc_21380_n6290;
  wire core__abc_21380_n6291;
  wire core__abc_21380_n6292;
  wire core__abc_21380_n6293;
  wire core__abc_21380_n6294;
  wire core__abc_21380_n6295;
  wire core__abc_21380_n6296;
  wire core__abc_21380_n6297;
  wire core__abc_21380_n6298;
  wire core__abc_21380_n6299;
  wire core__abc_21380_n6300;
  wire core__abc_21380_n6301;
  wire core__abc_21380_n6302;
  wire core__abc_21380_n6303;
  wire core__abc_21380_n6304;
  wire core__abc_21380_n6305;
  wire core__abc_21380_n6306;
  wire core__abc_21380_n6307;
  wire core__abc_21380_n6308;
  wire core__abc_21380_n6309;
  wire core__abc_21380_n6310;
  wire core__abc_21380_n6311;
  wire core__abc_21380_n6312;
  wire core__abc_21380_n6313;
  wire core__abc_21380_n6314;
  wire core__abc_21380_n6315;
  wire core__abc_21380_n6316;
  wire core__abc_21380_n6318;
  wire core__abc_21380_n6319;
  wire core__abc_21380_n6320;
  wire core__abc_21380_n6321;
  wire core__abc_21380_n6322;
  wire core__abc_21380_n6323;
  wire core__abc_21380_n6324;
  wire core__abc_21380_n6325;
  wire core__abc_21380_n6326;
  wire core__abc_21380_n6327;
  wire core__abc_21380_n6328;
  wire core__abc_21380_n6329;
  wire core__abc_21380_n6330;
  wire core__abc_21380_n6331;
  wire core__abc_21380_n6332;
  wire core__abc_21380_n6333;
  wire core__abc_21380_n6334;
  wire core__abc_21380_n6335;
  wire core__abc_21380_n6336;
  wire core__abc_21380_n6337;
  wire core__abc_21380_n6338;
  wire core__abc_21380_n6339;
  wire core__abc_21380_n6340;
  wire core__abc_21380_n6341;
  wire core__abc_21380_n6342;
  wire core__abc_21380_n6343;
  wire core__abc_21380_n6344;
  wire core__abc_21380_n6345;
  wire core__abc_21380_n6346;
  wire core__abc_21380_n6347;
  wire core__abc_21380_n6348;
  wire core__abc_21380_n6349;
  wire core__abc_21380_n6350;
  wire core__abc_21380_n6352;
  wire core__abc_21380_n6353;
  wire core__abc_21380_n6354;
  wire core__abc_21380_n6355;
  wire core__abc_21380_n6356;
  wire core__abc_21380_n6357;
  wire core__abc_21380_n6358;
  wire core__abc_21380_n6359;
  wire core__abc_21380_n6360;
  wire core__abc_21380_n6361;
  wire core__abc_21380_n6362;
  wire core__abc_21380_n6363;
  wire core__abc_21380_n6364;
  wire core__abc_21380_n6365;
  wire core__abc_21380_n6366;
  wire core__abc_21380_n6367;
  wire core__abc_21380_n6368;
  wire core__abc_21380_n6369;
  wire core__abc_21380_n6370;
  wire core__abc_21380_n6371;
  wire core__abc_21380_n6372;
  wire core__abc_21380_n6373;
  wire core__abc_21380_n6374;
  wire core__abc_21380_n6375;
  wire core__abc_21380_n6376;
  wire core__abc_21380_n6377;
  wire core__abc_21380_n6378;
  wire core__abc_21380_n6379;
  wire core__abc_21380_n6380;
  wire core__abc_21380_n6381;
  wire core__abc_21380_n6382;
  wire core__abc_21380_n6383;
  wire core__abc_21380_n6384;
  wire core__abc_21380_n6385;
  wire core__abc_21380_n6386;
  wire core__abc_21380_n6387;
  wire core__abc_21380_n6388;
  wire core__abc_21380_n6389;
  wire core__abc_21380_n6390;
  wire core__abc_21380_n6391;
  wire core__abc_21380_n6392;
  wire core__abc_21380_n6393;
  wire core__abc_21380_n6394;
  wire core__abc_21380_n6395;
  wire core__abc_21380_n6396;
  wire core__abc_21380_n6397;
  wire core__abc_21380_n6398;
  wire core__abc_21380_n6399;
  wire core__abc_21380_n6400;
  wire core__abc_21380_n6401;
  wire core__abc_21380_n6402;
  wire core__abc_21380_n6403;
  wire core__abc_21380_n6404;
  wire core__abc_21380_n6405;
  wire core__abc_21380_n6406;
  wire core__abc_21380_n6407;
  wire core__abc_21380_n6408;
  wire core__abc_21380_n6409;
  wire core__abc_21380_n6410;
  wire core__abc_21380_n6412;
  wire core__abc_21380_n6413;
  wire core__abc_21380_n6414;
  wire core__abc_21380_n6415;
  wire core__abc_21380_n6416;
  wire core__abc_21380_n6417;
  wire core__abc_21380_n6418;
  wire core__abc_21380_n6419;
  wire core__abc_21380_n6420;
  wire core__abc_21380_n6421;
  wire core__abc_21380_n6422;
  wire core__abc_21380_n6423;
  wire core__abc_21380_n6424;
  wire core__abc_21380_n6425;
  wire core__abc_21380_n6426;
  wire core__abc_21380_n6427;
  wire core__abc_21380_n6428;
  wire core__abc_21380_n6429;
  wire core__abc_21380_n6430;
  wire core__abc_21380_n6431;
  wire core__abc_21380_n6432;
  wire core__abc_21380_n6433;
  wire core__abc_21380_n6434;
  wire core__abc_21380_n6435;
  wire core__abc_21380_n6436;
  wire core__abc_21380_n6437;
  wire core__abc_21380_n6438;
  wire core__abc_21380_n6439;
  wire core__abc_21380_n6440;
  wire core__abc_21380_n6441;
  wire core__abc_21380_n6442;
  wire core__abc_21380_n6443;
  wire core__abc_21380_n6444;
  wire core__abc_21380_n6445;
  wire core__abc_21380_n6446;
  wire core__abc_21380_n6448;
  wire core__abc_21380_n6449;
  wire core__abc_21380_n6450;
  wire core__abc_21380_n6451;
  wire core__abc_21380_n6452;
  wire core__abc_21380_n6453;
  wire core__abc_21380_n6454;
  wire core__abc_21380_n6455;
  wire core__abc_21380_n6456;
  wire core__abc_21380_n6457;
  wire core__abc_21380_n6458;
  wire core__abc_21380_n6459;
  wire core__abc_21380_n6460;
  wire core__abc_21380_n6461;
  wire core__abc_21380_n6462;
  wire core__abc_21380_n6463;
  wire core__abc_21380_n6464;
  wire core__abc_21380_n6465;
  wire core__abc_21380_n6466;
  wire core__abc_21380_n6467;
  wire core__abc_21380_n6468;
  wire core__abc_21380_n6469;
  wire core__abc_21380_n6470;
  wire core__abc_21380_n6471;
  wire core__abc_21380_n6472;
  wire core__abc_21380_n6473;
  wire core__abc_21380_n6474;
  wire core__abc_21380_n6475;
  wire core__abc_21380_n6476;
  wire core__abc_21380_n6477;
  wire core__abc_21380_n6478;
  wire core__abc_21380_n6479;
  wire core__abc_21380_n6480;
  wire core__abc_21380_n6481;
  wire core__abc_21380_n6482;
  wire core__abc_21380_n6483;
  wire core__abc_21380_n6484;
  wire core__abc_21380_n6485;
  wire core__abc_21380_n6486;
  wire core__abc_21380_n6488;
  wire core__abc_21380_n6489;
  wire core__abc_21380_n6490;
  wire core__abc_21380_n6491;
  wire core__abc_21380_n6492;
  wire core__abc_21380_n6493;
  wire core__abc_21380_n6494;
  wire core__abc_21380_n6495;
  wire core__abc_21380_n6496;
  wire core__abc_21380_n6497;
  wire core__abc_21380_n6498;
  wire core__abc_21380_n6499;
  wire core__abc_21380_n6500;
  wire core__abc_21380_n6501;
  wire core__abc_21380_n6502;
  wire core__abc_21380_n6503;
  wire core__abc_21380_n6504;
  wire core__abc_21380_n6505;
  wire core__abc_21380_n6506;
  wire core__abc_21380_n6507;
  wire core__abc_21380_n6508;
  wire core__abc_21380_n6509;
  wire core__abc_21380_n6510;
  wire core__abc_21380_n6511;
  wire core__abc_21380_n6512;
  wire core__abc_21380_n6513;
  wire core__abc_21380_n6514;
  wire core__abc_21380_n6515;
  wire core__abc_21380_n6516;
  wire core__abc_21380_n6517;
  wire core__abc_21380_n6518;
  wire core__abc_21380_n6519;
  wire core__abc_21380_n6520;
  wire core__abc_21380_n6522;
  wire core__abc_21380_n6523;
  wire core__abc_21380_n6524;
  wire core__abc_21380_n6525;
  wire core__abc_21380_n6526;
  wire core__abc_21380_n6527;
  wire core__abc_21380_n6528;
  wire core__abc_21380_n6529;
  wire core__abc_21380_n6530;
  wire core__abc_21380_n6531;
  wire core__abc_21380_n6532;
  wire core__abc_21380_n6533;
  wire core__abc_21380_n6534;
  wire core__abc_21380_n6535;
  wire core__abc_21380_n6536;
  wire core__abc_21380_n6537;
  wire core__abc_21380_n6538;
  wire core__abc_21380_n6539;
  wire core__abc_21380_n6540;
  wire core__abc_21380_n6541;
  wire core__abc_21380_n6542;
  wire core__abc_21380_n6543;
  wire core__abc_21380_n6544;
  wire core__abc_21380_n6545;
  wire core__abc_21380_n6546;
  wire core__abc_21380_n6547;
  wire core__abc_21380_n6548;
  wire core__abc_21380_n6549;
  wire core__abc_21380_n6550;
  wire core__abc_21380_n6551;
  wire core__abc_21380_n6552;
  wire core__abc_21380_n6553;
  wire core__abc_21380_n6554;
  wire core__abc_21380_n6555;
  wire core__abc_21380_n6556;
  wire core__abc_21380_n6557;
  wire core__abc_21380_n6558;
  wire core__abc_21380_n6559;
  wire core__abc_21380_n6560;
  wire core__abc_21380_n6561;
  wire core__abc_21380_n6562;
  wire core__abc_21380_n6563;
  wire core__abc_21380_n6564;
  wire core__abc_21380_n6565;
  wire core__abc_21380_n6566;
  wire core__abc_21380_n6567;
  wire core__abc_21380_n6568;
  wire core__abc_21380_n6569;
  wire core__abc_21380_n6571;
  wire core__abc_21380_n6572;
  wire core__abc_21380_n6573;
  wire core__abc_21380_n6574;
  wire core__abc_21380_n6575;
  wire core__abc_21380_n6576;
  wire core__abc_21380_n6577;
  wire core__abc_21380_n6578;
  wire core__abc_21380_n6579;
  wire core__abc_21380_n6580;
  wire core__abc_21380_n6581;
  wire core__abc_21380_n6582;
  wire core__abc_21380_n6583;
  wire core__abc_21380_n6584;
  wire core__abc_21380_n6585;
  wire core__abc_21380_n6586;
  wire core__abc_21380_n6587;
  wire core__abc_21380_n6588;
  wire core__abc_21380_n6589;
  wire core__abc_21380_n6590;
  wire core__abc_21380_n6591;
  wire core__abc_21380_n6592;
  wire core__abc_21380_n6593;
  wire core__abc_21380_n6594;
  wire core__abc_21380_n6595;
  wire core__abc_21380_n6596;
  wire core__abc_21380_n6597;
  wire core__abc_21380_n6598;
  wire core__abc_21380_n6599;
  wire core__abc_21380_n6600;
  wire core__abc_21380_n6601;
  wire core__abc_21380_n6602;
  wire core__abc_21380_n6603;
  wire core__abc_21380_n6604;
  wire core__abc_21380_n6606;
  wire core__abc_21380_n6607;
  wire core__abc_21380_n6608;
  wire core__abc_21380_n6609;
  wire core__abc_21380_n6610;
  wire core__abc_21380_n6611;
  wire core__abc_21380_n6612;
  wire core__abc_21380_n6613;
  wire core__abc_21380_n6614;
  wire core__abc_21380_n6615;
  wire core__abc_21380_n6616;
  wire core__abc_21380_n6617;
  wire core__abc_21380_n6618;
  wire core__abc_21380_n6619;
  wire core__abc_21380_n6620;
  wire core__abc_21380_n6621;
  wire core__abc_21380_n6622;
  wire core__abc_21380_n6623;
  wire core__abc_21380_n6624;
  wire core__abc_21380_n6625;
  wire core__abc_21380_n6626;
  wire core__abc_21380_n6627;
  wire core__abc_21380_n6628;
  wire core__abc_21380_n6629;
  wire core__abc_21380_n6630;
  wire core__abc_21380_n6631;
  wire core__abc_21380_n6632;
  wire core__abc_21380_n6633;
  wire core__abc_21380_n6634;
  wire core__abc_21380_n6635;
  wire core__abc_21380_n6636;
  wire core__abc_21380_n6637;
  wire core__abc_21380_n6638;
  wire core__abc_21380_n6639;
  wire core__abc_21380_n6640;
  wire core__abc_21380_n6641;
  wire core__abc_21380_n6642;
  wire core__abc_21380_n6643;
  wire core__abc_21380_n6644;
  wire core__abc_21380_n6645;
  wire core__abc_21380_n6646;
  wire core__abc_21380_n6648;
  wire core__abc_21380_n6649;
  wire core__abc_21380_n6650;
  wire core__abc_21380_n6651;
  wire core__abc_21380_n6652;
  wire core__abc_21380_n6653;
  wire core__abc_21380_n6654;
  wire core__abc_21380_n6655;
  wire core__abc_21380_n6656;
  wire core__abc_21380_n6657;
  wire core__abc_21380_n6658;
  wire core__abc_21380_n6659;
  wire core__abc_21380_n6660;
  wire core__abc_21380_n6661;
  wire core__abc_21380_n6662;
  wire core__abc_21380_n6663;
  wire core__abc_21380_n6664;
  wire core__abc_21380_n6665;
  wire core__abc_21380_n6666;
  wire core__abc_21380_n6667;
  wire core__abc_21380_n6668;
  wire core__abc_21380_n6669;
  wire core__abc_21380_n6670;
  wire core__abc_21380_n6671;
  wire core__abc_21380_n6672;
  wire core__abc_21380_n6673;
  wire core__abc_21380_n6674;
  wire core__abc_21380_n6675;
  wire core__abc_21380_n6676;
  wire core__abc_21380_n6677;
  wire core__abc_21380_n6678;
  wire core__abc_21380_n6679;
  wire core__abc_21380_n6680;
  wire core__abc_21380_n6681;
  wire core__abc_21380_n6682;
  wire core__abc_21380_n6684;
  wire core__abc_21380_n6685;
  wire core__abc_21380_n6686;
  wire core__abc_21380_n6687;
  wire core__abc_21380_n6688;
  wire core__abc_21380_n6689;
  wire core__abc_21380_n6690;
  wire core__abc_21380_n6691;
  wire core__abc_21380_n6692;
  wire core__abc_21380_n6693;
  wire core__abc_21380_n6694;
  wire core__abc_21380_n6695;
  wire core__abc_21380_n6696;
  wire core__abc_21380_n6697;
  wire core__abc_21380_n6698;
  wire core__abc_21380_n6699;
  wire core__abc_21380_n6700;
  wire core__abc_21380_n6701;
  wire core__abc_21380_n6702;
  wire core__abc_21380_n6703;
  wire core__abc_21380_n6704;
  wire core__abc_21380_n6705;
  wire core__abc_21380_n6706;
  wire core__abc_21380_n6707;
  wire core__abc_21380_n6708;
  wire core__abc_21380_n6709;
  wire core__abc_21380_n6710;
  wire core__abc_21380_n6711;
  wire core__abc_21380_n6712;
  wire core__abc_21380_n6713;
  wire core__abc_21380_n6714;
  wire core__abc_21380_n6715;
  wire core__abc_21380_n6716;
  wire core__abc_21380_n6717;
  wire core__abc_21380_n6718;
  wire core__abc_21380_n6719;
  wire core__abc_21380_n6720;
  wire core__abc_21380_n6721;
  wire core__abc_21380_n6722;
  wire core__abc_21380_n6723;
  wire core__abc_21380_n6724;
  wire core__abc_21380_n6725;
  wire core__abc_21380_n6726;
  wire core__abc_21380_n6727;
  wire core__abc_21380_n6728;
  wire core__abc_21380_n6729;
  wire core__abc_21380_n6730;
  wire core__abc_21380_n6731;
  wire core__abc_21380_n6732;
  wire core__abc_21380_n6733;
  wire core__abc_21380_n6734;
  wire core__abc_21380_n6735;
  wire core__abc_21380_n6736;
  wire core__abc_21380_n6737;
  wire core__abc_21380_n6738;
  wire core__abc_21380_n6739;
  wire core__abc_21380_n6740;
  wire core__abc_21380_n6741;
  wire core__abc_21380_n6742;
  wire core__abc_21380_n6743;
  wire core__abc_21380_n6744;
  wire core__abc_21380_n6745;
  wire core__abc_21380_n6746;
  wire core__abc_21380_n6747;
  wire core__abc_21380_n6748;
  wire core__abc_21380_n6749;
  wire core__abc_21380_n6750;
  wire core__abc_21380_n6751;
  wire core__abc_21380_n6752;
  wire core__abc_21380_n6753;
  wire core__abc_21380_n6754;
  wire core__abc_21380_n6755;
  wire core__abc_21380_n6756;
  wire core__abc_21380_n6757;
  wire core__abc_21380_n6758;
  wire core__abc_21380_n6759;
  wire core__abc_21380_n6760;
  wire core__abc_21380_n6761;
  wire core__abc_21380_n6762;
  wire core__abc_21380_n6763;
  wire core__abc_21380_n6764;
  wire core__abc_21380_n6765;
  wire core__abc_21380_n6766;
  wire core__abc_21380_n6767;
  wire core__abc_21380_n6768;
  wire core__abc_21380_n6769;
  wire core__abc_21380_n6770;
  wire core__abc_21380_n6771;
  wire core__abc_21380_n6772;
  wire core__abc_21380_n6773;
  wire core__abc_21380_n6774;
  wire core__abc_21380_n6775;
  wire core__abc_21380_n6776;
  wire core__abc_21380_n6777;
  wire core__abc_21380_n6778;
  wire core__abc_21380_n6779;
  wire core__abc_21380_n6780;
  wire core__abc_21380_n6781;
  wire core__abc_21380_n6782;
  wire core__abc_21380_n6783;
  wire core__abc_21380_n6784;
  wire core__abc_21380_n6785;
  wire core__abc_21380_n6786;
  wire core__abc_21380_n6787;
  wire core__abc_21380_n6788;
  wire core__abc_21380_n6789;
  wire core__abc_21380_n6790;
  wire core__abc_21380_n6791;
  wire core__abc_21380_n6792;
  wire core__abc_21380_n6793;
  wire core__abc_21380_n6794;
  wire core__abc_21380_n6795;
  wire core__abc_21380_n6796;
  wire core__abc_21380_n6797;
  wire core__abc_21380_n6798;
  wire core__abc_21380_n6799;
  wire core__abc_21380_n6800;
  wire core__abc_21380_n6801;
  wire core__abc_21380_n6802;
  wire core__abc_21380_n6803;
  wire core__abc_21380_n6804;
  wire core__abc_21380_n6805;
  wire core__abc_21380_n6806;
  wire core__abc_21380_n6807;
  wire core__abc_21380_n6808;
  wire core__abc_21380_n6809;
  wire core__abc_21380_n6810;
  wire core__abc_21380_n6811;
  wire core__abc_21380_n6812;
  wire core__abc_21380_n6813;
  wire core__abc_21380_n6814;
  wire core__abc_21380_n6815;
  wire core__abc_21380_n6816;
  wire core__abc_21380_n6817;
  wire core__abc_21380_n6818;
  wire core__abc_21380_n6819;
  wire core__abc_21380_n6820;
  wire core__abc_21380_n6821;
  wire core__abc_21380_n6822;
  wire core__abc_21380_n6823;
  wire core__abc_21380_n6824;
  wire core__abc_21380_n6825;
  wire core__abc_21380_n6826;
  wire core__abc_21380_n6827;
  wire core__abc_21380_n6828;
  wire core__abc_21380_n6829;
  wire core__abc_21380_n6830;
  wire core__abc_21380_n6831;
  wire core__abc_21380_n6832;
  wire core__abc_21380_n6833;
  wire core__abc_21380_n6834;
  wire core__abc_21380_n6835;
  wire core__abc_21380_n6836;
  wire core__abc_21380_n6837;
  wire core__abc_21380_n6838;
  wire core__abc_21380_n6839;
  wire core__abc_21380_n6840;
  wire core__abc_21380_n6841;
  wire core__abc_21380_n6842;
  wire core__abc_21380_n6843;
  wire core__abc_21380_n6844;
  wire core__abc_21380_n6845;
  wire core__abc_21380_n6846;
  wire core__abc_21380_n6847;
  wire core__abc_21380_n6848;
  wire core__abc_21380_n6849;
  wire core__abc_21380_n6850;
  wire core__abc_21380_n6851;
  wire core__abc_21380_n6852;
  wire core__abc_21380_n6853;
  wire core__abc_21380_n6854;
  wire core__abc_21380_n6855;
  wire core__abc_21380_n6856;
  wire core__abc_21380_n6857;
  wire core__abc_21380_n6858;
  wire core__abc_21380_n6859;
  wire core__abc_21380_n6860;
  wire core__abc_21380_n6861;
  wire core__abc_21380_n6862;
  wire core__abc_21380_n6863;
  wire core__abc_21380_n6864;
  wire core__abc_21380_n6865;
  wire core__abc_21380_n6866;
  wire core__abc_21380_n6867;
  wire core__abc_21380_n6868;
  wire core__abc_21380_n6869;
  wire core__abc_21380_n6870;
  wire core__abc_21380_n6871;
  wire core__abc_21380_n6872;
  wire core__abc_21380_n6873;
  wire core__abc_21380_n6874;
  wire core__abc_21380_n6875;
  wire core__abc_21380_n6876;
  wire core__abc_21380_n6877;
  wire core__abc_21380_n6878;
  wire core__abc_21380_n6879;
  wire core__abc_21380_n6880;
  wire core__abc_21380_n6881;
  wire core__abc_21380_n6882;
  wire core__abc_21380_n6883;
  wire core__abc_21380_n6884;
  wire core__abc_21380_n6885;
  wire core__abc_21380_n6886;
  wire core__abc_21380_n6887;
  wire core__abc_21380_n6888;
  wire core__abc_21380_n6889;
  wire core__abc_21380_n6890;
  wire core__abc_21380_n6891;
  wire core__abc_21380_n6892;
  wire core__abc_21380_n6893;
  wire core__abc_21380_n6894;
  wire core__abc_21380_n6895;
  wire core__abc_21380_n6896;
  wire core__abc_21380_n6897;
  wire core__abc_21380_n6898;
  wire core__abc_21380_n6899;
  wire core__abc_21380_n6900;
  wire core__abc_21380_n6901;
  wire core__abc_21380_n6902;
  wire core__abc_21380_n6903;
  wire core__abc_21380_n6904;
  wire core__abc_21380_n6905;
  wire core__abc_21380_n6906;
  wire core__abc_21380_n6907;
  wire core__abc_21380_n6908;
  wire core__abc_21380_n6909;
  wire core__abc_21380_n6910;
  wire core__abc_21380_n6911;
  wire core__abc_21380_n6912;
  wire core__abc_21380_n6913;
  wire core__abc_21380_n6914;
  wire core__abc_21380_n6915;
  wire core__abc_21380_n6916;
  wire core__abc_21380_n6917;
  wire core__abc_21380_n6918;
  wire core__abc_21380_n6919;
  wire core__abc_21380_n6920;
  wire core__abc_21380_n6921;
  wire core__abc_21380_n6922;
  wire core__abc_21380_n6923;
  wire core__abc_21380_n6924;
  wire core__abc_21380_n6925;
  wire core__abc_21380_n6926;
  wire core__abc_21380_n6927;
  wire core__abc_21380_n6928;
  wire core__abc_21380_n6929;
  wire core__abc_21380_n6930;
  wire core__abc_21380_n6931;
  wire core__abc_21380_n6932;
  wire core__abc_21380_n6933;
  wire core__abc_21380_n6934;
  wire core__abc_21380_n6935;
  wire core__abc_21380_n6936;
  wire core__abc_21380_n6937;
  wire core__abc_21380_n6938;
  wire core__abc_21380_n6939;
  wire core__abc_21380_n6940;
  wire core__abc_21380_n6941;
  wire core__abc_21380_n6942;
  wire core__abc_21380_n6943;
  wire core__abc_21380_n6944;
  wire core__abc_21380_n6945;
  wire core__abc_21380_n6946;
  wire core__abc_21380_n6947;
  wire core__abc_21380_n6948;
  wire core__abc_21380_n6949;
  wire core__abc_21380_n6950;
  wire core__abc_21380_n6951;
  wire core__abc_21380_n6952;
  wire core__abc_21380_n6953;
  wire core__abc_21380_n6954;
  wire core__abc_21380_n6955;
  wire core__abc_21380_n6956;
  wire core__abc_21380_n6957;
  wire core__abc_21380_n6958;
  wire core__abc_21380_n6959;
  wire core__abc_21380_n6960;
  wire core__abc_21380_n6961;
  wire core__abc_21380_n6962;
  wire core__abc_21380_n6963;
  wire core__abc_21380_n6964;
  wire core__abc_21380_n6965;
  wire core__abc_21380_n6966;
  wire core__abc_21380_n6967;
  wire core__abc_21380_n6968;
  wire core__abc_21380_n6969;
  wire core__abc_21380_n6970;
  wire core__abc_21380_n6971;
  wire core__abc_21380_n6972;
  wire core__abc_21380_n6973;
  wire core__abc_21380_n6974;
  wire core__abc_21380_n6975;
  wire core__abc_21380_n6976;
  wire core__abc_21380_n6977;
  wire core__abc_21380_n6978;
  wire core__abc_21380_n6979;
  wire core__abc_21380_n6980;
  wire core__abc_21380_n6981;
  wire core__abc_21380_n6982;
  wire core__abc_21380_n6983;
  wire core__abc_21380_n6984;
  wire core__abc_21380_n6985;
  wire core__abc_21380_n6986;
  wire core__abc_21380_n6987;
  wire core__abc_21380_n6988;
  wire core__abc_21380_n6989;
  wire core__abc_21380_n6990;
  wire core__abc_21380_n6991;
  wire core__abc_21380_n6992;
  wire core__abc_21380_n6993;
  wire core__abc_21380_n6994;
  wire core__abc_21380_n6995;
  wire core__abc_21380_n6996;
  wire core__abc_21380_n6997;
  wire core__abc_21380_n6998;
  wire core__abc_21380_n6999;
  wire core__abc_21380_n7000;
  wire core__abc_21380_n7001;
  wire core__abc_21380_n7002;
  wire core__abc_21380_n7003;
  wire core__abc_21380_n7004;
  wire core__abc_21380_n7005;
  wire core__abc_21380_n7006;
  wire core__abc_21380_n7007;
  wire core__abc_21380_n7008;
  wire core__abc_21380_n7009;
  wire core__abc_21380_n7010;
  wire core__abc_21380_n7011;
  wire core__abc_21380_n7012;
  wire core__abc_21380_n7013;
  wire core__abc_21380_n7014;
  wire core__abc_21380_n7015;
  wire core__abc_21380_n7016;
  wire core__abc_21380_n7017;
  wire core__abc_21380_n7018;
  wire core__abc_21380_n7019;
  wire core__abc_21380_n7020;
  wire core__abc_21380_n7021;
  wire core__abc_21380_n7022;
  wire core__abc_21380_n7023;
  wire core__abc_21380_n7024;
  wire core__abc_21380_n7025;
  wire core__abc_21380_n7026;
  wire core__abc_21380_n7027;
  wire core__abc_21380_n7028;
  wire core__abc_21380_n7029;
  wire core__abc_21380_n7030;
  wire core__abc_21380_n7031;
  wire core__abc_21380_n7032;
  wire core__abc_21380_n7033;
  wire core__abc_21380_n7034;
  wire core__abc_21380_n7035;
  wire core__abc_21380_n7036;
  wire core__abc_21380_n7037;
  wire core__abc_21380_n7038;
  wire core__abc_21380_n7039;
  wire core__abc_21380_n7040;
  wire core__abc_21380_n7041;
  wire core__abc_21380_n7042;
  wire core__abc_21380_n7043;
  wire core__abc_21380_n7044;
  wire core__abc_21380_n7045;
  wire core__abc_21380_n7046;
  wire core__abc_21380_n7047;
  wire core__abc_21380_n7048;
  wire core__abc_21380_n7049;
  wire core__abc_21380_n7050;
  wire core__abc_21380_n7051;
  wire core__abc_21380_n7052;
  wire core__abc_21380_n7053;
  wire core__abc_21380_n7054;
  wire core__abc_21380_n7055;
  wire core__abc_21380_n7056;
  wire core__abc_21380_n7057;
  wire core__abc_21380_n7058;
  wire core__abc_21380_n7059;
  wire core__abc_21380_n7060;
  wire core__abc_21380_n7061;
  wire core__abc_21380_n7062;
  wire core__abc_21380_n7063;
  wire core__abc_21380_n7064;
  wire core__abc_21380_n7065;
  wire core__abc_21380_n7066;
  wire core__abc_21380_n7067;
  wire core__abc_21380_n7068;
  wire core__abc_21380_n7069;
  wire core__abc_21380_n7070;
  wire core__abc_21380_n7071;
  wire core__abc_21380_n7072;
  wire core__abc_21380_n7073;
  wire core__abc_21380_n7074;
  wire core__abc_21380_n7075;
  wire core__abc_21380_n7076;
  wire core__abc_21380_n7076_bF_buf0;
  wire core__abc_21380_n7076_bF_buf1;
  wire core__abc_21380_n7076_bF_buf2;
  wire core__abc_21380_n7076_bF_buf3;
  wire core__abc_21380_n7076_bF_buf4;
  wire core__abc_21380_n7076_bF_buf5;
  wire core__abc_21380_n7076_bF_buf6;
  wire core__abc_21380_n7077;
  wire core__abc_21380_n7078;
  wire core__abc_21380_n7079;
  wire core__abc_21380_n7080;
  wire core__abc_21380_n7081;
  wire core__abc_21380_n7082;
  wire core__abc_21380_n7083;
  wire core__abc_21380_n7084;
  wire core__abc_21380_n7085;
  wire core__abc_21380_n7086;
  wire core__abc_21380_n7087;
  wire core__abc_21380_n7087_bF_buf0;
  wire core__abc_21380_n7087_bF_buf1;
  wire core__abc_21380_n7087_bF_buf2;
  wire core__abc_21380_n7087_bF_buf3;
  wire core__abc_21380_n7087_bF_buf4;
  wire core__abc_21380_n7087_bF_buf5;
  wire core__abc_21380_n7087_bF_buf6;
  wire core__abc_21380_n7087_bF_buf7;
  wire core__abc_21380_n7088;
  wire core__abc_21380_n7089;
  wire core__abc_21380_n7091;
  wire core__abc_21380_n7092;
  wire core__abc_21380_n7093;
  wire core__abc_21380_n7094;
  wire core__abc_21380_n7095;
  wire core__abc_21380_n7096;
  wire core__abc_21380_n7097;
  wire core__abc_21380_n7098;
  wire core__abc_21380_n7099;
  wire core__abc_21380_n7100;
  wire core__abc_21380_n7101;
  wire core__abc_21380_n7102;
  wire core__abc_21380_n7103;
  wire core__abc_21380_n7104;
  wire core__abc_21380_n7105;
  wire core__abc_21380_n7106;
  wire core__abc_21380_n7107;
  wire core__abc_21380_n7108;
  wire core__abc_21380_n7109;
  wire core__abc_21380_n7110;
  wire core__abc_21380_n7111;
  wire core__abc_21380_n7112;
  wire core__abc_21380_n7113;
  wire core__abc_21380_n7115;
  wire core__abc_21380_n7116;
  wire core__abc_21380_n7117;
  wire core__abc_21380_n7118;
  wire core__abc_21380_n7119;
  wire core__abc_21380_n7120;
  wire core__abc_21380_n7121;
  wire core__abc_21380_n7122;
  wire core__abc_21380_n7123;
  wire core__abc_21380_n7124;
  wire core__abc_21380_n7125;
  wire core__abc_21380_n7126;
  wire core__abc_21380_n7127;
  wire core__abc_21380_n7128;
  wire core__abc_21380_n7129;
  wire core__abc_21380_n7130;
  wire core__abc_21380_n7131;
  wire core__abc_21380_n7132;
  wire core__abc_21380_n7133;
  wire core__abc_21380_n7134;
  wire core__abc_21380_n7135;
  wire core__abc_21380_n7136;
  wire core__abc_21380_n7137;
  wire core__abc_21380_n7138;
  wire core__abc_21380_n7139;
  wire core__abc_21380_n7140;
  wire core__abc_21380_n7141;
  wire core__abc_21380_n7143;
  wire core__abc_21380_n7144;
  wire core__abc_21380_n7145;
  wire core__abc_21380_n7146;
  wire core__abc_21380_n7147;
  wire core__abc_21380_n7148;
  wire core__abc_21380_n7149;
  wire core__abc_21380_n7150;
  wire core__abc_21380_n7151;
  wire core__abc_21380_n7152;
  wire core__abc_21380_n7153;
  wire core__abc_21380_n7154;
  wire core__abc_21380_n7155;
  wire core__abc_21380_n7156;
  wire core__abc_21380_n7157;
  wire core__abc_21380_n7158;
  wire core__abc_21380_n7159;
  wire core__abc_21380_n7160;
  wire core__abc_21380_n7161;
  wire core__abc_21380_n7162;
  wire core__abc_21380_n7163;
  wire core__abc_21380_n7164;
  wire core__abc_21380_n7165;
  wire core__abc_21380_n7166;
  wire core__abc_21380_n7168;
  wire core__abc_21380_n7169;
  wire core__abc_21380_n7170;
  wire core__abc_21380_n7171;
  wire core__abc_21380_n7172;
  wire core__abc_21380_n7173;
  wire core__abc_21380_n7174;
  wire core__abc_21380_n7175;
  wire core__abc_21380_n7176;
  wire core__abc_21380_n7177;
  wire core__abc_21380_n7178;
  wire core__abc_21380_n7179;
  wire core__abc_21380_n7180;
  wire core__abc_21380_n7181;
  wire core__abc_21380_n7182;
  wire core__abc_21380_n7183;
  wire core__abc_21380_n7184;
  wire core__abc_21380_n7185;
  wire core__abc_21380_n7186;
  wire core__abc_21380_n7187;
  wire core__abc_21380_n7188;
  wire core__abc_21380_n7189;
  wire core__abc_21380_n7190;
  wire core__abc_21380_n7191;
  wire core__abc_21380_n7192;
  wire core__abc_21380_n7193;
  wire core__abc_21380_n7194;
  wire core__abc_21380_n7195;
  wire core__abc_21380_n7196;
  wire core__abc_21380_n7197;
  wire core__abc_21380_n7198;
  wire core__abc_21380_n7200;
  wire core__abc_21380_n7201;
  wire core__abc_21380_n7202;
  wire core__abc_21380_n7203;
  wire core__abc_21380_n7204;
  wire core__abc_21380_n7205;
  wire core__abc_21380_n7206;
  wire core__abc_21380_n7207;
  wire core__abc_21380_n7208;
  wire core__abc_21380_n7209;
  wire core__abc_21380_n7210;
  wire core__abc_21380_n7211;
  wire core__abc_21380_n7212;
  wire core__abc_21380_n7213;
  wire core__abc_21380_n7214;
  wire core__abc_21380_n7215;
  wire core__abc_21380_n7216;
  wire core__abc_21380_n7217;
  wire core__abc_21380_n7218;
  wire core__abc_21380_n7219;
  wire core__abc_21380_n7220;
  wire core__abc_21380_n7221;
  wire core__abc_21380_n7222;
  wire core__abc_21380_n7223;
  wire core__abc_21380_n7224;
  wire core__abc_21380_n7225;
  wire core__abc_21380_n7227;
  wire core__abc_21380_n7228;
  wire core__abc_21380_n7229;
  wire core__abc_21380_n7230;
  wire core__abc_21380_n7231;
  wire core__abc_21380_n7232;
  wire core__abc_21380_n7233;
  wire core__abc_21380_n7234;
  wire core__abc_21380_n7235;
  wire core__abc_21380_n7236;
  wire core__abc_21380_n7237;
  wire core__abc_21380_n7238;
  wire core__abc_21380_n7239;
  wire core__abc_21380_n7240;
  wire core__abc_21380_n7241;
  wire core__abc_21380_n7242;
  wire core__abc_21380_n7243;
  wire core__abc_21380_n7244;
  wire core__abc_21380_n7245;
  wire core__abc_21380_n7246;
  wire core__abc_21380_n7247;
  wire core__abc_21380_n7248;
  wire core__abc_21380_n7249;
  wire core__abc_21380_n7250;
  wire core__abc_21380_n7251;
  wire core__abc_21380_n7253;
  wire core__abc_21380_n7254;
  wire core__abc_21380_n7255;
  wire core__abc_21380_n7256;
  wire core__abc_21380_n7257;
  wire core__abc_21380_n7258;
  wire core__abc_21380_n7259;
  wire core__abc_21380_n7260;
  wire core__abc_21380_n7261;
  wire core__abc_21380_n7262;
  wire core__abc_21380_n7263;
  wire core__abc_21380_n7264;
  wire core__abc_21380_n7265;
  wire core__abc_21380_n7266;
  wire core__abc_21380_n7267;
  wire core__abc_21380_n7268;
  wire core__abc_21380_n7269;
  wire core__abc_21380_n7270;
  wire core__abc_21380_n7271;
  wire core__abc_21380_n7272;
  wire core__abc_21380_n7273;
  wire core__abc_21380_n7274;
  wire core__abc_21380_n7275;
  wire core__abc_21380_n7277;
  wire core__abc_21380_n7278;
  wire core__abc_21380_n7279;
  wire core__abc_21380_n7280;
  wire core__abc_21380_n7281;
  wire core__abc_21380_n7282;
  wire core__abc_21380_n7283;
  wire core__abc_21380_n7284;
  wire core__abc_21380_n7285;
  wire core__abc_21380_n7286;
  wire core__abc_21380_n7287;
  wire core__abc_21380_n7288;
  wire core__abc_21380_n7289;
  wire core__abc_21380_n7290;
  wire core__abc_21380_n7291;
  wire core__abc_21380_n7292;
  wire core__abc_21380_n7293;
  wire core__abc_21380_n7294;
  wire core__abc_21380_n7295;
  wire core__abc_21380_n7296;
  wire core__abc_21380_n7297;
  wire core__abc_21380_n7298;
  wire core__abc_21380_n7299;
  wire core__abc_21380_n7300;
  wire core__abc_21380_n7301;
  wire core__abc_21380_n7302;
  wire core__abc_21380_n7303;
  wire core__abc_21380_n7304;
  wire core__abc_21380_n7305;
  wire core__abc_21380_n7306;
  wire core__abc_21380_n7307;
  wire core__abc_21380_n7308;
  wire core__abc_21380_n7309;
  wire core__abc_21380_n7310;
  wire core__abc_21380_n7311;
  wire core__abc_21380_n7312;
  wire core__abc_21380_n7313;
  wire core__abc_21380_n7314;
  wire core__abc_21380_n7315;
  wire core__abc_21380_n7317;
  wire core__abc_21380_n7318;
  wire core__abc_21380_n7319;
  wire core__abc_21380_n7320;
  wire core__abc_21380_n7321;
  wire core__abc_21380_n7322;
  wire core__abc_21380_n7323;
  wire core__abc_21380_n7324;
  wire core__abc_21380_n7325;
  wire core__abc_21380_n7326;
  wire core__abc_21380_n7327;
  wire core__abc_21380_n7328;
  wire core__abc_21380_n7329;
  wire core__abc_21380_n7330;
  wire core__abc_21380_n7331;
  wire core__abc_21380_n7332;
  wire core__abc_21380_n7333;
  wire core__abc_21380_n7334;
  wire core__abc_21380_n7335;
  wire core__abc_21380_n7336;
  wire core__abc_21380_n7337;
  wire core__abc_21380_n7338;
  wire core__abc_21380_n7339;
  wire core__abc_21380_n7340;
  wire core__abc_21380_n7341;
  wire core__abc_21380_n7342;
  wire core__abc_21380_n7343;
  wire core__abc_21380_n7345;
  wire core__abc_21380_n7346;
  wire core__abc_21380_n7347;
  wire core__abc_21380_n7348;
  wire core__abc_21380_n7349;
  wire core__abc_21380_n7350;
  wire core__abc_21380_n7351;
  wire core__abc_21380_n7352;
  wire core__abc_21380_n7353;
  wire core__abc_21380_n7354;
  wire core__abc_21380_n7355;
  wire core__abc_21380_n7356;
  wire core__abc_21380_n7357;
  wire core__abc_21380_n7358;
  wire core__abc_21380_n7359;
  wire core__abc_21380_n7360;
  wire core__abc_21380_n7361;
  wire core__abc_21380_n7362;
  wire core__abc_21380_n7363;
  wire core__abc_21380_n7364;
  wire core__abc_21380_n7365;
  wire core__abc_21380_n7366;
  wire core__abc_21380_n7367;
  wire core__abc_21380_n7368;
  wire core__abc_21380_n7369;
  wire core__abc_21380_n7370;
  wire core__abc_21380_n7371;
  wire core__abc_21380_n7373;
  wire core__abc_21380_n7374;
  wire core__abc_21380_n7375;
  wire core__abc_21380_n7376;
  wire core__abc_21380_n7377;
  wire core__abc_21380_n7378;
  wire core__abc_21380_n7379;
  wire core__abc_21380_n7380;
  wire core__abc_21380_n7381;
  wire core__abc_21380_n7382;
  wire core__abc_21380_n7383;
  wire core__abc_21380_n7384;
  wire core__abc_21380_n7385;
  wire core__abc_21380_n7386;
  wire core__abc_21380_n7387;
  wire core__abc_21380_n7388;
  wire core__abc_21380_n7389;
  wire core__abc_21380_n7390;
  wire core__abc_21380_n7391;
  wire core__abc_21380_n7392;
  wire core__abc_21380_n7393;
  wire core__abc_21380_n7394;
  wire core__abc_21380_n7396;
  wire core__abc_21380_n7397;
  wire core__abc_21380_n7398;
  wire core__abc_21380_n7399;
  wire core__abc_21380_n7400;
  wire core__abc_21380_n7401;
  wire core__abc_21380_n7402;
  wire core__abc_21380_n7403;
  wire core__abc_21380_n7404;
  wire core__abc_21380_n7405;
  wire core__abc_21380_n7406;
  wire core__abc_21380_n7407;
  wire core__abc_21380_n7408;
  wire core__abc_21380_n7409;
  wire core__abc_21380_n7410;
  wire core__abc_21380_n7411;
  wire core__abc_21380_n7412;
  wire core__abc_21380_n7413;
  wire core__abc_21380_n7414;
  wire core__abc_21380_n7415;
  wire core__abc_21380_n7416;
  wire core__abc_21380_n7417;
  wire core__abc_21380_n7418;
  wire core__abc_21380_n7419;
  wire core__abc_21380_n7420;
  wire core__abc_21380_n7421;
  wire core__abc_21380_n7422;
  wire core__abc_21380_n7423;
  wire core__abc_21380_n7424;
  wire core__abc_21380_n7425;
  wire core__abc_21380_n7427;
  wire core__abc_21380_n7428;
  wire core__abc_21380_n7429;
  wire core__abc_21380_n7430;
  wire core__abc_21380_n7431;
  wire core__abc_21380_n7432;
  wire core__abc_21380_n7433;
  wire core__abc_21380_n7434;
  wire core__abc_21380_n7435;
  wire core__abc_21380_n7436;
  wire core__abc_21380_n7437;
  wire core__abc_21380_n7438;
  wire core__abc_21380_n7439;
  wire core__abc_21380_n7440;
  wire core__abc_21380_n7441;
  wire core__abc_21380_n7442;
  wire core__abc_21380_n7443;
  wire core__abc_21380_n7444;
  wire core__abc_21380_n7445;
  wire core__abc_21380_n7446;
  wire core__abc_21380_n7447;
  wire core__abc_21380_n7448;
  wire core__abc_21380_n7449;
  wire core__abc_21380_n7450;
  wire core__abc_21380_n7451;
  wire core__abc_21380_n7453;
  wire core__abc_21380_n7454;
  wire core__abc_21380_n7455;
  wire core__abc_21380_n7456;
  wire core__abc_21380_n7457;
  wire core__abc_21380_n7458;
  wire core__abc_21380_n7459;
  wire core__abc_21380_n7460;
  wire core__abc_21380_n7461;
  wire core__abc_21380_n7462;
  wire core__abc_21380_n7463;
  wire core__abc_21380_n7464;
  wire core__abc_21380_n7465;
  wire core__abc_21380_n7466;
  wire core__abc_21380_n7467;
  wire core__abc_21380_n7468;
  wire core__abc_21380_n7469;
  wire core__abc_21380_n7470;
  wire core__abc_21380_n7471;
  wire core__abc_21380_n7472;
  wire core__abc_21380_n7473;
  wire core__abc_21380_n7474;
  wire core__abc_21380_n7475;
  wire core__abc_21380_n7476;
  wire core__abc_21380_n7477;
  wire core__abc_21380_n7478;
  wire core__abc_21380_n7479;
  wire core__abc_21380_n7480;
  wire core__abc_21380_n7482;
  wire core__abc_21380_n7483;
  wire core__abc_21380_n7484;
  wire core__abc_21380_n7485;
  wire core__abc_21380_n7486;
  wire core__abc_21380_n7487;
  wire core__abc_21380_n7488;
  wire core__abc_21380_n7489;
  wire core__abc_21380_n7490;
  wire core__abc_21380_n7491;
  wire core__abc_21380_n7492;
  wire core__abc_21380_n7493;
  wire core__abc_21380_n7494;
  wire core__abc_21380_n7495;
  wire core__abc_21380_n7496;
  wire core__abc_21380_n7497;
  wire core__abc_21380_n7498;
  wire core__abc_21380_n7499;
  wire core__abc_21380_n7500;
  wire core__abc_21380_n7501;
  wire core__abc_21380_n7502;
  wire core__abc_21380_n7503;
  wire core__abc_21380_n7505;
  wire core__abc_21380_n7506;
  wire core__abc_21380_n7507;
  wire core__abc_21380_n7508;
  wire core__abc_21380_n7509;
  wire core__abc_21380_n7510;
  wire core__abc_21380_n7511;
  wire core__abc_21380_n7512;
  wire core__abc_21380_n7513;
  wire core__abc_21380_n7514;
  wire core__abc_21380_n7515;
  wire core__abc_21380_n7516;
  wire core__abc_21380_n7517;
  wire core__abc_21380_n7518;
  wire core__abc_21380_n7519;
  wire core__abc_21380_n7520;
  wire core__abc_21380_n7521;
  wire core__abc_21380_n7522;
  wire core__abc_21380_n7523;
  wire core__abc_21380_n7524;
  wire core__abc_21380_n7525;
  wire core__abc_21380_n7526;
  wire core__abc_21380_n7527;
  wire core__abc_21380_n7528;
  wire core__abc_21380_n7529;
  wire core__abc_21380_n7530;
  wire core__abc_21380_n7531;
  wire core__abc_21380_n7532;
  wire core__abc_21380_n7533;
  wire core__abc_21380_n7534;
  wire core__abc_21380_n7535;
  wire core__abc_21380_n7536;
  wire core__abc_21380_n7537;
  wire core__abc_21380_n7538;
  wire core__abc_21380_n7539;
  wire core__abc_21380_n7540;
  wire core__abc_21380_n7541;
  wire core__abc_21380_n7542;
  wire core__abc_21380_n7543;
  wire core__abc_21380_n7544;
  wire core__abc_21380_n7545;
  wire core__abc_21380_n7547;
  wire core__abc_21380_n7548;
  wire core__abc_21380_n7549;
  wire core__abc_21380_n7550;
  wire core__abc_21380_n7551;
  wire core__abc_21380_n7552;
  wire core__abc_21380_n7553;
  wire core__abc_21380_n7554;
  wire core__abc_21380_n7555;
  wire core__abc_21380_n7556;
  wire core__abc_21380_n7557;
  wire core__abc_21380_n7558;
  wire core__abc_21380_n7559;
  wire core__abc_21380_n7560;
  wire core__abc_21380_n7561;
  wire core__abc_21380_n7562;
  wire core__abc_21380_n7563;
  wire core__abc_21380_n7564;
  wire core__abc_21380_n7565;
  wire core__abc_21380_n7566;
  wire core__abc_21380_n7567;
  wire core__abc_21380_n7568;
  wire core__abc_21380_n7569;
  wire core__abc_21380_n7570;
  wire core__abc_21380_n7571;
  wire core__abc_21380_n7573;
  wire core__abc_21380_n7574;
  wire core__abc_21380_n7575;
  wire core__abc_21380_n7576;
  wire core__abc_21380_n7577;
  wire core__abc_21380_n7578;
  wire core__abc_21380_n7579;
  wire core__abc_21380_n7580;
  wire core__abc_21380_n7581;
  wire core__abc_21380_n7582;
  wire core__abc_21380_n7583;
  wire core__abc_21380_n7584;
  wire core__abc_21380_n7585;
  wire core__abc_21380_n7586;
  wire core__abc_21380_n7587;
  wire core__abc_21380_n7588;
  wire core__abc_21380_n7589;
  wire core__abc_21380_n7590;
  wire core__abc_21380_n7591;
  wire core__abc_21380_n7592;
  wire core__abc_21380_n7593;
  wire core__abc_21380_n7594;
  wire core__abc_21380_n7595;
  wire core__abc_21380_n7596;
  wire core__abc_21380_n7597;
  wire core__abc_21380_n7598;
  wire core__abc_21380_n7599;
  wire core__abc_21380_n7601;
  wire core__abc_21380_n7602;
  wire core__abc_21380_n7603;
  wire core__abc_21380_n7604;
  wire core__abc_21380_n7605;
  wire core__abc_21380_n7606;
  wire core__abc_21380_n7607;
  wire core__abc_21380_n7608;
  wire core__abc_21380_n7609;
  wire core__abc_21380_n7610;
  wire core__abc_21380_n7611;
  wire core__abc_21380_n7612;
  wire core__abc_21380_n7613;
  wire core__abc_21380_n7614;
  wire core__abc_21380_n7615;
  wire core__abc_21380_n7616;
  wire core__abc_21380_n7617;
  wire core__abc_21380_n7618;
  wire core__abc_21380_n7619;
  wire core__abc_21380_n7620;
  wire core__abc_21380_n7621;
  wire core__abc_21380_n7622;
  wire core__abc_21380_n7624;
  wire core__abc_21380_n7625;
  wire core__abc_21380_n7626;
  wire core__abc_21380_n7627;
  wire core__abc_21380_n7628;
  wire core__abc_21380_n7629;
  wire core__abc_21380_n7630;
  wire core__abc_21380_n7631;
  wire core__abc_21380_n7632;
  wire core__abc_21380_n7633;
  wire core__abc_21380_n7634;
  wire core__abc_21380_n7635;
  wire core__abc_21380_n7636;
  wire core__abc_21380_n7637;
  wire core__abc_21380_n7638;
  wire core__abc_21380_n7639;
  wire core__abc_21380_n7640;
  wire core__abc_21380_n7641;
  wire core__abc_21380_n7642;
  wire core__abc_21380_n7643;
  wire core__abc_21380_n7644;
  wire core__abc_21380_n7645;
  wire core__abc_21380_n7646;
  wire core__abc_21380_n7647;
  wire core__abc_21380_n7648;
  wire core__abc_21380_n7649;
  wire core__abc_21380_n7650;
  wire core__abc_21380_n7651;
  wire core__abc_21380_n7652;
  wire core__abc_21380_n7653;
  wire core__abc_21380_n7655;
  wire core__abc_21380_n7656;
  wire core__abc_21380_n7657;
  wire core__abc_21380_n7658;
  wire core__abc_21380_n7659;
  wire core__abc_21380_n7660;
  wire core__abc_21380_n7661;
  wire core__abc_21380_n7662;
  wire core__abc_21380_n7663;
  wire core__abc_21380_n7664;
  wire core__abc_21380_n7665;
  wire core__abc_21380_n7666;
  wire core__abc_21380_n7667;
  wire core__abc_21380_n7668;
  wire core__abc_21380_n7669;
  wire core__abc_21380_n7670;
  wire core__abc_21380_n7671;
  wire core__abc_21380_n7672;
  wire core__abc_21380_n7673;
  wire core__abc_21380_n7674;
  wire core__abc_21380_n7675;
  wire core__abc_21380_n7676;
  wire core__abc_21380_n7678;
  wire core__abc_21380_n7679;
  wire core__abc_21380_n7680;
  wire core__abc_21380_n7681;
  wire core__abc_21380_n7682;
  wire core__abc_21380_n7683;
  wire core__abc_21380_n7684;
  wire core__abc_21380_n7685;
  wire core__abc_21380_n7686;
  wire core__abc_21380_n7687;
  wire core__abc_21380_n7688;
  wire core__abc_21380_n7689;
  wire core__abc_21380_n7690;
  wire core__abc_21380_n7691;
  wire core__abc_21380_n7692;
  wire core__abc_21380_n7693;
  wire core__abc_21380_n7694;
  wire core__abc_21380_n7695;
  wire core__abc_21380_n7696;
  wire core__abc_21380_n7697;
  wire core__abc_21380_n7698;
  wire core__abc_21380_n7699;
  wire core__abc_21380_n7700;
  wire core__abc_21380_n7701;
  wire core__abc_21380_n7702;
  wire core__abc_21380_n7703;
  wire core__abc_21380_n7704;
  wire core__abc_21380_n7706;
  wire core__abc_21380_n7707;
  wire core__abc_21380_n7708;
  wire core__abc_21380_n7709;
  wire core__abc_21380_n7710;
  wire core__abc_21380_n7711;
  wire core__abc_21380_n7712;
  wire core__abc_21380_n7713;
  wire core__abc_21380_n7714;
  wire core__abc_21380_n7715;
  wire core__abc_21380_n7716;
  wire core__abc_21380_n7717;
  wire core__abc_21380_n7718;
  wire core__abc_21380_n7719;
  wire core__abc_21380_n7720;
  wire core__abc_21380_n7721;
  wire core__abc_21380_n7722;
  wire core__abc_21380_n7723;
  wire core__abc_21380_n7724;
  wire core__abc_21380_n7725;
  wire core__abc_21380_n7726;
  wire core__abc_21380_n7727;
  wire core__abc_21380_n7728;
  wire core__abc_21380_n7729;
  wire core__abc_21380_n7731;
  wire core__abc_21380_n7732;
  wire core__abc_21380_n7733;
  wire core__abc_21380_n7734;
  wire core__abc_21380_n7735;
  wire core__abc_21380_n7736;
  wire core__abc_21380_n7737;
  wire core__abc_21380_n7738;
  wire core__abc_21380_n7739;
  wire core__abc_21380_n7740;
  wire core__abc_21380_n7741;
  wire core__abc_21380_n7742;
  wire core__abc_21380_n7743;
  wire core__abc_21380_n7744;
  wire core__abc_21380_n7745;
  wire core__abc_21380_n7746;
  wire core__abc_21380_n7747;
  wire core__abc_21380_n7748;
  wire core__abc_21380_n7749;
  wire core__abc_21380_n7750;
  wire core__abc_21380_n7751;
  wire core__abc_21380_n7752;
  wire core__abc_21380_n7753;
  wire core__abc_21380_n7754;
  wire core__abc_21380_n7755;
  wire core__abc_21380_n7756;
  wire core__abc_21380_n7757;
  wire core__abc_21380_n7758;
  wire core__abc_21380_n7759;
  wire core__abc_21380_n7760;
  wire core__abc_21380_n7761;
  wire core__abc_21380_n7762;
  wire core__abc_21380_n7763;
  wire core__abc_21380_n7764;
  wire core__abc_21380_n7765;
  wire core__abc_21380_n7766;
  wire core__abc_21380_n7768;
  wire core__abc_21380_n7769;
  wire core__abc_21380_n7770;
  wire core__abc_21380_n7771;
  wire core__abc_21380_n7772;
  wire core__abc_21380_n7773;
  wire core__abc_21380_n7774;
  wire core__abc_21380_n7775;
  wire core__abc_21380_n7776;
  wire core__abc_21380_n7777;
  wire core__abc_21380_n7778;
  wire core__abc_21380_n7779;
  wire core__abc_21380_n7780;
  wire core__abc_21380_n7781;
  wire core__abc_21380_n7782;
  wire core__abc_21380_n7783;
  wire core__abc_21380_n7784;
  wire core__abc_21380_n7785;
  wire core__abc_21380_n7786;
  wire core__abc_21380_n7787;
  wire core__abc_21380_n7788;
  wire core__abc_21380_n7789;
  wire core__abc_21380_n7790;
  wire core__abc_21380_n7791;
  wire core__abc_21380_n7792;
  wire core__abc_21380_n7793;
  wire core__abc_21380_n7794;
  wire core__abc_21380_n7796;
  wire core__abc_21380_n7797;
  wire core__abc_21380_n7798;
  wire core__abc_21380_n7799;
  wire core__abc_21380_n7800;
  wire core__abc_21380_n7801;
  wire core__abc_21380_n7802;
  wire core__abc_21380_n7803;
  wire core__abc_21380_n7804;
  wire core__abc_21380_n7805;
  wire core__abc_21380_n7806;
  wire core__abc_21380_n7807;
  wire core__abc_21380_n7808;
  wire core__abc_21380_n7809;
  wire core__abc_21380_n7810;
  wire core__abc_21380_n7811;
  wire core__abc_21380_n7812;
  wire core__abc_21380_n7813;
  wire core__abc_21380_n7814;
  wire core__abc_21380_n7815;
  wire core__abc_21380_n7816;
  wire core__abc_21380_n7817;
  wire core__abc_21380_n7818;
  wire core__abc_21380_n7819;
  wire core__abc_21380_n7820;
  wire core__abc_21380_n7821;
  wire core__abc_21380_n7823;
  wire core__abc_21380_n7824;
  wire core__abc_21380_n7825;
  wire core__abc_21380_n7826;
  wire core__abc_21380_n7827;
  wire core__abc_21380_n7828;
  wire core__abc_21380_n7829;
  wire core__abc_21380_n7830;
  wire core__abc_21380_n7831;
  wire core__abc_21380_n7832;
  wire core__abc_21380_n7833;
  wire core__abc_21380_n7834;
  wire core__abc_21380_n7835;
  wire core__abc_21380_n7836;
  wire core__abc_21380_n7837;
  wire core__abc_21380_n7838;
  wire core__abc_21380_n7839;
  wire core__abc_21380_n7840;
  wire core__abc_21380_n7841;
  wire core__abc_21380_n7842;
  wire core__abc_21380_n7843;
  wire core__abc_21380_n7844;
  wire core__abc_21380_n7845;
  wire core__abc_21380_n7846;
  wire core__abc_21380_n7847;
  wire core__abc_21380_n7848;
  wire core__abc_21380_n7849;
  wire core__abc_21380_n7851;
  wire core__abc_21380_n7852;
  wire core__abc_21380_n7853;
  wire core__abc_21380_n7854;
  wire core__abc_21380_n7855;
  wire core__abc_21380_n7856;
  wire core__abc_21380_n7857;
  wire core__abc_21380_n7858;
  wire core__abc_21380_n7859;
  wire core__abc_21380_n7860;
  wire core__abc_21380_n7861;
  wire core__abc_21380_n7862;
  wire core__abc_21380_n7863;
  wire core__abc_21380_n7864;
  wire core__abc_21380_n7865;
  wire core__abc_21380_n7866;
  wire core__abc_21380_n7867;
  wire core__abc_21380_n7868;
  wire core__abc_21380_n7869;
  wire core__abc_21380_n7870;
  wire core__abc_21380_n7871;
  wire core__abc_21380_n7872;
  wire core__abc_21380_n7873;
  wire core__abc_21380_n7874;
  wire core__abc_21380_n7875;
  wire core__abc_21380_n7876;
  wire core__abc_21380_n7877;
  wire core__abc_21380_n7878;
  wire core__abc_21380_n7879;
  wire core__abc_21380_n7880;
  wire core__abc_21380_n7881;
  wire core__abc_21380_n7882;
  wire core__abc_21380_n7883;
  wire core__abc_21380_n7884;
  wire core__abc_21380_n7885;
  wire core__abc_21380_n7887;
  wire core__abc_21380_n7888;
  wire core__abc_21380_n7889;
  wire core__abc_21380_n7890;
  wire core__abc_21380_n7891;
  wire core__abc_21380_n7892;
  wire core__abc_21380_n7893;
  wire core__abc_21380_n7894;
  wire core__abc_21380_n7895;
  wire core__abc_21380_n7896;
  wire core__abc_21380_n7897;
  wire core__abc_21380_n7898;
  wire core__abc_21380_n7899;
  wire core__abc_21380_n7900;
  wire core__abc_21380_n7901;
  wire core__abc_21380_n7902;
  wire core__abc_21380_n7903;
  wire core__abc_21380_n7904;
  wire core__abc_21380_n7905;
  wire core__abc_21380_n7906;
  wire core__abc_21380_n7907;
  wire core__abc_21380_n7908;
  wire core__abc_21380_n7909;
  wire core__abc_21380_n7910;
  wire core__abc_21380_n7912;
  wire core__abc_21380_n7913;
  wire core__abc_21380_n7914;
  wire core__abc_21380_n7915;
  wire core__abc_21380_n7916;
  wire core__abc_21380_n7917;
  wire core__abc_21380_n7918;
  wire core__abc_21380_n7919;
  wire core__abc_21380_n7920;
  wire core__abc_21380_n7921;
  wire core__abc_21380_n7922;
  wire core__abc_21380_n7923;
  wire core__abc_21380_n7924;
  wire core__abc_21380_n7925;
  wire core__abc_21380_n7926;
  wire core__abc_21380_n7927;
  wire core__abc_21380_n7928;
  wire core__abc_21380_n7929;
  wire core__abc_21380_n7930;
  wire core__abc_21380_n7931;
  wire core__abc_21380_n7932;
  wire core__abc_21380_n7933;
  wire core__abc_21380_n7934;
  wire core__abc_21380_n7935;
  wire core__abc_21380_n7936;
  wire core__abc_21380_n7937;
  wire core__abc_21380_n7938;
  wire core__abc_21380_n7939;
  wire core__abc_21380_n7940;
  wire core__abc_21380_n7941;
  wire core__abc_21380_n7943;
  wire core__abc_21380_n7944;
  wire core__abc_21380_n7945;
  wire core__abc_21380_n7946;
  wire core__abc_21380_n7947;
  wire core__abc_21380_n7948;
  wire core__abc_21380_n7949;
  wire core__abc_21380_n7950;
  wire core__abc_21380_n7951;
  wire core__abc_21380_n7952;
  wire core__abc_21380_n7953;
  wire core__abc_21380_n7954;
  wire core__abc_21380_n7955;
  wire core__abc_21380_n7956;
  wire core__abc_21380_n7957;
  wire core__abc_21380_n7958;
  wire core__abc_21380_n7959;
  wire core__abc_21380_n7960;
  wire core__abc_21380_n7961;
  wire core__abc_21380_n7962;
  wire core__abc_21380_n7963;
  wire core__abc_21380_n7964;
  wire core__abc_21380_n7965;
  wire core__abc_21380_n7967;
  wire core__abc_21380_n7968;
  wire core__abc_21380_n7969;
  wire core__abc_21380_n7970;
  wire core__abc_21380_n7971;
  wire core__abc_21380_n7972;
  wire core__abc_21380_n7973;
  wire core__abc_21380_n7974;
  wire core__abc_21380_n7975;
  wire core__abc_21380_n7976;
  wire core__abc_21380_n7977;
  wire core__abc_21380_n7978;
  wire core__abc_21380_n7980;
  wire core__abc_21380_n7981;
  wire core__abc_21380_n7982;
  wire core__abc_21380_n7983;
  wire core__abc_21380_n7984;
  wire core__abc_21380_n7985;
  wire core__abc_21380_n7986;
  wire core__abc_21380_n7987;
  wire core__abc_21380_n7988;
  wire core__abc_21380_n7990;
  wire core__abc_21380_n7991;
  wire core__abc_21380_n7992;
  wire core__abc_21380_n7993;
  wire core__abc_21380_n7994;
  wire core__abc_21380_n7995;
  wire core__abc_21380_n7996;
  wire core__abc_21380_n7997;
  wire core__abc_21380_n7998;
  wire core__abc_21380_n7999;
  wire core__abc_21380_n8001;
  wire core__abc_21380_n8002;
  wire core__abc_21380_n8003;
  wire core__abc_21380_n8004;
  wire core__abc_21380_n8005;
  wire core__abc_21380_n8006;
  wire core__abc_21380_n8007;
  wire core__abc_21380_n8008;
  wire core__abc_21380_n8009;
  wire core__abc_21380_n8010;
  wire core__abc_21380_n8011;
  wire core__abc_21380_n8013;
  wire core__abc_21380_n8014;
  wire core__abc_21380_n8015;
  wire core__abc_21380_n8016;
  wire core__abc_21380_n8017;
  wire core__abc_21380_n8018;
  wire core__abc_21380_n8019;
  wire core__abc_21380_n8020;
  wire core__abc_21380_n8021;
  wire core__abc_21380_n8022;
  wire core__abc_21380_n8023;
  wire core__abc_21380_n8025;
  wire core__abc_21380_n8026;
  wire core__abc_21380_n8027;
  wire core__abc_21380_n8028;
  wire core__abc_21380_n8029;
  wire core__abc_21380_n8030;
  wire core__abc_21380_n8031;
  wire core__abc_21380_n8032;
  wire core__abc_21380_n8033;
  wire core__abc_21380_n8034;
  wire core__abc_21380_n8035;
  wire core__abc_21380_n8036;
  wire core__abc_21380_n8038;
  wire core__abc_21380_n8039;
  wire core__abc_21380_n8040;
  wire core__abc_21380_n8041;
  wire core__abc_21380_n8042;
  wire core__abc_21380_n8043;
  wire core__abc_21380_n8044;
  wire core__abc_21380_n8045;
  wire core__abc_21380_n8046;
  wire core__abc_21380_n8047;
  wire core__abc_21380_n8048;
  wire core__abc_21380_n8049;
  wire core__abc_21380_n8050;
  wire core__abc_21380_n8052;
  wire core__abc_21380_n8053;
  wire core__abc_21380_n8054;
  wire core__abc_21380_n8055;
  wire core__abc_21380_n8056;
  wire core__abc_21380_n8057;
  wire core__abc_21380_n8058;
  wire core__abc_21380_n8059;
  wire core__abc_21380_n8060;
  wire core__abc_21380_n8061;
  wire core__abc_21380_n8062;
  wire core__abc_21380_n8063;
  wire core__abc_21380_n8064;
  wire core__abc_21380_n8065;
  wire core__abc_21380_n8067;
  wire core__abc_21380_n8068;
  wire core__abc_21380_n8069;
  wire core__abc_21380_n8070;
  wire core__abc_21380_n8071;
  wire core__abc_21380_n8072;
  wire core__abc_21380_n8073;
  wire core__abc_21380_n8074;
  wire core__abc_21380_n8075;
  wire core__abc_21380_n8076;
  wire core__abc_21380_n8077;
  wire core__abc_21380_n8078;
  wire core__abc_21380_n8079;
  wire core__abc_21380_n8080;
  wire core__abc_21380_n8082;
  wire core__abc_21380_n8083;
  wire core__abc_21380_n8084;
  wire core__abc_21380_n8085;
  wire core__abc_21380_n8086;
  wire core__abc_21380_n8087;
  wire core__abc_21380_n8088;
  wire core__abc_21380_n8089;
  wire core__abc_21380_n8090;
  wire core__abc_21380_n8091;
  wire core__abc_21380_n8092;
  wire core__abc_21380_n8093;
  wire core__abc_21380_n8094;
  wire core__abc_21380_n8095;
  wire core__abc_21380_n8096;
  wire core__abc_21380_n8097;
  wire core__abc_21380_n8099;
  wire core__abc_21380_n8100;
  wire core__abc_21380_n8101;
  wire core__abc_21380_n8102;
  wire core__abc_21380_n8103;
  wire core__abc_21380_n8104;
  wire core__abc_21380_n8105;
  wire core__abc_21380_n8106;
  wire core__abc_21380_n8107;
  wire core__abc_21380_n8108;
  wire core__abc_21380_n8109;
  wire core__abc_21380_n8110;
  wire core__abc_21380_n8111;
  wire core__abc_21380_n8112;
  wire core__abc_21380_n8113;
  wire core__abc_21380_n8115;
  wire core__abc_21380_n8116;
  wire core__abc_21380_n8117;
  wire core__abc_21380_n8118;
  wire core__abc_21380_n8119;
  wire core__abc_21380_n8120;
  wire core__abc_21380_n8121;
  wire core__abc_21380_n8122;
  wire core__abc_21380_n8123;
  wire core__abc_21380_n8124;
  wire core__abc_21380_n8125;
  wire core__abc_21380_n8126;
  wire core__abc_21380_n8127;
  wire core__abc_21380_n8128;
  wire core__abc_21380_n8130;
  wire core__abc_21380_n8131;
  wire core__abc_21380_n8132;
  wire core__abc_21380_n8133;
  wire core__abc_21380_n8134;
  wire core__abc_21380_n8135;
  wire core__abc_21380_n8136;
  wire core__abc_21380_n8137;
  wire core__abc_21380_n8138;
  wire core__abc_21380_n8139;
  wire core__abc_21380_n8140;
  wire core__abc_21380_n8141;
  wire core__abc_21380_n8142;
  wire core__abc_21380_n8144;
  wire core__abc_21380_n8145;
  wire core__abc_21380_n8146;
  wire core__abc_21380_n8147;
  wire core__abc_21380_n8148;
  wire core__abc_21380_n8149;
  wire core__abc_21380_n8150;
  wire core__abc_21380_n8151;
  wire core__abc_21380_n8152;
  wire core__abc_21380_n8153;
  wire core__abc_21380_n8154;
  wire core__abc_21380_n8155;
  wire core__abc_21380_n8156;
  wire core__abc_21380_n8157;
  wire core__abc_21380_n8158;
  wire core__abc_21380_n8159;
  wire core__abc_21380_n8161;
  wire core__abc_21380_n8162;
  wire core__abc_21380_n8163;
  wire core__abc_21380_n8164;
  wire core__abc_21380_n8165;
  wire core__abc_21380_n8166;
  wire core__abc_21380_n8167;
  wire core__abc_21380_n8168;
  wire core__abc_21380_n8169;
  wire core__abc_21380_n8170;
  wire core__abc_21380_n8171;
  wire core__abc_21380_n8172;
  wire core__abc_21380_n8173;
  wire core__abc_21380_n8174;
  wire core__abc_21380_n8175;
  wire core__abc_21380_n8177;
  wire core__abc_21380_n8178;
  wire core__abc_21380_n8179;
  wire core__abc_21380_n8180;
  wire core__abc_21380_n8181;
  wire core__abc_21380_n8182;
  wire core__abc_21380_n8183;
  wire core__abc_21380_n8184;
  wire core__abc_21380_n8185;
  wire core__abc_21380_n8186;
  wire core__abc_21380_n8187;
  wire core__abc_21380_n8188;
  wire core__abc_21380_n8189;
  wire core__abc_21380_n8190;
  wire core__abc_21380_n8191;
  wire core__abc_21380_n8193;
  wire core__abc_21380_n8194;
  wire core__abc_21380_n8195;
  wire core__abc_21380_n8196;
  wire core__abc_21380_n8197;
  wire core__abc_21380_n8198;
  wire core__abc_21380_n8199;
  wire core__abc_21380_n8200;
  wire core__abc_21380_n8201;
  wire core__abc_21380_n8202;
  wire core__abc_21380_n8203;
  wire core__abc_21380_n8204;
  wire core__abc_21380_n8205;
  wire core__abc_21380_n8206;
  wire core__abc_21380_n8208;
  wire core__abc_21380_n8209;
  wire core__abc_21380_n8210;
  wire core__abc_21380_n8211;
  wire core__abc_21380_n8212;
  wire core__abc_21380_n8213;
  wire core__abc_21380_n8214;
  wire core__abc_21380_n8215;
  wire core__abc_21380_n8216;
  wire core__abc_21380_n8217;
  wire core__abc_21380_n8218;
  wire core__abc_21380_n8219;
  wire core__abc_21380_n8220;
  wire core__abc_21380_n8221;
  wire core__abc_21380_n8223;
  wire core__abc_21380_n8224;
  wire core__abc_21380_n8225;
  wire core__abc_21380_n8226;
  wire core__abc_21380_n8227;
  wire core__abc_21380_n8228;
  wire core__abc_21380_n8229;
  wire core__abc_21380_n8230;
  wire core__abc_21380_n8231;
  wire core__abc_21380_n8232;
  wire core__abc_21380_n8233;
  wire core__abc_21380_n8234;
  wire core__abc_21380_n8235;
  wire core__abc_21380_n8236;
  wire core__abc_21380_n8237;
  wire core__abc_21380_n8239;
  wire core__abc_21380_n8240;
  wire core__abc_21380_n8241;
  wire core__abc_21380_n8242;
  wire core__abc_21380_n8243;
  wire core__abc_21380_n8244;
  wire core__abc_21380_n8245;
  wire core__abc_21380_n8246;
  wire core__abc_21380_n8247;
  wire core__abc_21380_n8248;
  wire core__abc_21380_n8249;
  wire core__abc_21380_n8250;
  wire core__abc_21380_n8251;
  wire core__abc_21380_n8252;
  wire core__abc_21380_n8253;
  wire core__abc_21380_n8254;
  wire core__abc_21380_n8256;
  wire core__abc_21380_n8257;
  wire core__abc_21380_n8258;
  wire core__abc_21380_n8259;
  wire core__abc_21380_n8260;
  wire core__abc_21380_n8261;
  wire core__abc_21380_n8262;
  wire core__abc_21380_n8263;
  wire core__abc_21380_n8264;
  wire core__abc_21380_n8265;
  wire core__abc_21380_n8266;
  wire core__abc_21380_n8267;
  wire core__abc_21380_n8268;
  wire core__abc_21380_n8269;
  wire core__abc_21380_n8270;
  wire core__abc_21380_n8272;
  wire core__abc_21380_n8273;
  wire core__abc_21380_n8274;
  wire core__abc_21380_n8275;
  wire core__abc_21380_n8276;
  wire core__abc_21380_n8277;
  wire core__abc_21380_n8278;
  wire core__abc_21380_n8279;
  wire core__abc_21380_n8280;
  wire core__abc_21380_n8281;
  wire core__abc_21380_n8282;
  wire core__abc_21380_n8283;
  wire core__abc_21380_n8284;
  wire core__abc_21380_n8285;
  wire core__abc_21380_n8286;
  wire core__abc_21380_n8288;
  wire core__abc_21380_n8289;
  wire core__abc_21380_n8290;
  wire core__abc_21380_n8291;
  wire core__abc_21380_n8292;
  wire core__abc_21380_n8293;
  wire core__abc_21380_n8294;
  wire core__abc_21380_n8295;
  wire core__abc_21380_n8296;
  wire core__abc_21380_n8297;
  wire core__abc_21380_n8298;
  wire core__abc_21380_n8299;
  wire core__abc_21380_n8300;
  wire core__abc_21380_n8301;
  wire core__abc_21380_n8302;
  wire core__abc_21380_n8303;
  wire core__abc_21380_n8305;
  wire core__abc_21380_n8306;
  wire core__abc_21380_n8307;
  wire core__abc_21380_n8308;
  wire core__abc_21380_n8309;
  wire core__abc_21380_n8310;
  wire core__abc_21380_n8311;
  wire core__abc_21380_n8312;
  wire core__abc_21380_n8313;
  wire core__abc_21380_n8314;
  wire core__abc_21380_n8315;
  wire core__abc_21380_n8316;
  wire core__abc_21380_n8317;
  wire core__abc_21380_n8318;
  wire core__abc_21380_n8320;
  wire core__abc_21380_n8321;
  wire core__abc_21380_n8322;
  wire core__abc_21380_n8323;
  wire core__abc_21380_n8324;
  wire core__abc_21380_n8325;
  wire core__abc_21380_n8326;
  wire core__abc_21380_n8327;
  wire core__abc_21380_n8328;
  wire core__abc_21380_n8329;
  wire core__abc_21380_n8330;
  wire core__abc_21380_n8331;
  wire core__abc_21380_n8332;
  wire core__abc_21380_n8334;
  wire core__abc_21380_n8335;
  wire core__abc_21380_n8336;
  wire core__abc_21380_n8337;
  wire core__abc_21380_n8338;
  wire core__abc_21380_n8339;
  wire core__abc_21380_n8340;
  wire core__abc_21380_n8341;
  wire core__abc_21380_n8342;
  wire core__abc_21380_n8343;
  wire core__abc_21380_n8344;
  wire core__abc_21380_n8345;
  wire core__abc_21380_n8346;
  wire core__abc_21380_n8347;
  wire core__abc_21380_n8348;
  wire core__abc_21380_n8350;
  wire core__abc_21380_n8351;
  wire core__abc_21380_n8352;
  wire core__abc_21380_n8353;
  wire core__abc_21380_n8354;
  wire core__abc_21380_n8355;
  wire core__abc_21380_n8356;
  wire core__abc_21380_n8357;
  wire core__abc_21380_n8358;
  wire core__abc_21380_n8359;
  wire core__abc_21380_n8360;
  wire core__abc_21380_n8361;
  wire core__abc_21380_n8362;
  wire core__abc_21380_n8363;
  wire core__abc_21380_n8364;
  wire core__abc_21380_n8365;
  wire core__abc_21380_n8367;
  wire core__abc_21380_n8368;
  wire core__abc_21380_n8369;
  wire core__abc_21380_n8370;
  wire core__abc_21380_n8371;
  wire core__abc_21380_n8372;
  wire core__abc_21380_n8373;
  wire core__abc_21380_n8374;
  wire core__abc_21380_n8375;
  wire core__abc_21380_n8376;
  wire core__abc_21380_n8377;
  wire core__abc_21380_n8378;
  wire core__abc_21380_n8379;
  wire core__abc_21380_n8380;
  wire core__abc_21380_n8381;
  wire core__abc_21380_n8383;
  wire core__abc_21380_n8384;
  wire core__abc_21380_n8385;
  wire core__abc_21380_n8386;
  wire core__abc_21380_n8387;
  wire core__abc_21380_n8388;
  wire core__abc_21380_n8389;
  wire core__abc_21380_n8390;
  wire core__abc_21380_n8391;
  wire core__abc_21380_n8392;
  wire core__abc_21380_n8393;
  wire core__abc_21380_n8394;
  wire core__abc_21380_n8395;
  wire core__abc_21380_n8396;
  wire core__abc_21380_n8397;
  wire core__abc_21380_n8399;
  wire core__abc_21380_n8400;
  wire core__abc_21380_n8401;
  wire core__abc_21380_n8402;
  wire core__abc_21380_n8403;
  wire core__abc_21380_n8404;
  wire core__abc_21380_n8405;
  wire core__abc_21380_n8406;
  wire core__abc_21380_n8407;
  wire core__abc_21380_n8408;
  wire core__abc_21380_n8409;
  wire core__abc_21380_n8410;
  wire core__abc_21380_n8411;
  wire core__abc_21380_n8412;
  wire core__abc_21380_n8413;
  wire core__abc_21380_n8414;
  wire core__abc_21380_n8416;
  wire core__abc_21380_n8417;
  wire core__abc_21380_n8418;
  wire core__abc_21380_n8419;
  wire core__abc_21380_n8420;
  wire core__abc_21380_n8421;
  wire core__abc_21380_n8422;
  wire core__abc_21380_n8423;
  wire core__abc_21380_n8424;
  wire core__abc_21380_n8425;
  wire core__abc_21380_n8426;
  wire core__abc_21380_n8427;
  wire core__abc_21380_n8428;
  wire core__abc_21380_n8429;
  wire core__abc_21380_n8430;
  wire core__abc_21380_n8431;
  wire core__abc_21380_n8433;
  wire core__abc_21380_n8434;
  wire core__abc_21380_n8435;
  wire core__abc_21380_n8436;
  wire core__abc_21380_n8437;
  wire core__abc_21380_n8438;
  wire core__abc_21380_n8439;
  wire core__abc_21380_n8440;
  wire core__abc_21380_n8441;
  wire core__abc_21380_n8442;
  wire core__abc_21380_n8443;
  wire core__abc_21380_n8444;
  wire core__abc_21380_n8445;
  wire core__abc_21380_n8446;
  wire core__abc_21380_n8448;
  wire core__abc_21380_n8449;
  wire core__abc_21380_n8450;
  wire core__abc_21380_n8451;
  wire core__abc_21380_n8452;
  wire core__abc_21380_n8453;
  wire core__abc_21380_n8454;
  wire core__abc_21380_n8454_bF_buf0;
  wire core__abc_21380_n8454_bF_buf1;
  wire core__abc_21380_n8454_bF_buf2;
  wire core__abc_21380_n8454_bF_buf3;
  wire core__abc_21380_n8454_bF_buf4;
  wire core__abc_21380_n8454_bF_buf5;
  wire core__abc_21380_n8454_bF_buf6;
  wire core__abc_21380_n8454_bF_buf7;
  wire core__abc_21380_n8455;
  wire core__abc_21380_n8455_bF_buf0;
  wire core__abc_21380_n8455_bF_buf1;
  wire core__abc_21380_n8455_bF_buf2;
  wire core__abc_21380_n8455_bF_buf3;
  wire core__abc_21380_n8455_bF_buf4;
  wire core__abc_21380_n8455_bF_buf5;
  wire core__abc_21380_n8455_bF_buf6;
  wire core__abc_21380_n8455_bF_buf7;
  wire core__abc_21380_n8456;
  wire core__abc_21380_n8456_bF_buf0;
  wire core__abc_21380_n8456_bF_buf1;
  wire core__abc_21380_n8456_bF_buf2;
  wire core__abc_21380_n8456_bF_buf3;
  wire core__abc_21380_n8456_bF_buf4;
  wire core__abc_21380_n8456_bF_buf5;
  wire core__abc_21380_n8456_bF_buf6;
  wire core__abc_21380_n8456_bF_buf7;
  wire core__abc_21380_n8457;
  wire core__abc_21380_n8458;
  wire core__abc_21380_n8459;
  wire core__abc_21380_n8460;
  wire core__abc_21380_n8461;
  wire core__abc_21380_n8462;
  wire core__abc_21380_n8464;
  wire core__abc_21380_n8465;
  wire core__abc_21380_n8466;
  wire core__abc_21380_n8467;
  wire core__abc_21380_n8468;
  wire core__abc_21380_n8469;
  wire core__abc_21380_n8470;
  wire core__abc_21380_n8471;
  wire core__abc_21380_n8472;
  wire core__abc_21380_n8473;
  wire core__abc_21380_n8474;
  wire core__abc_21380_n8475;
  wire core__abc_21380_n8476;
  wire core__abc_21380_n8477;
  wire core__abc_21380_n8478;
  wire core__abc_21380_n8480;
  wire core__abc_21380_n8481;
  wire core__abc_21380_n8482;
  wire core__abc_21380_n8483;
  wire core__abc_21380_n8484;
  wire core__abc_21380_n8485;
  wire core__abc_21380_n8486;
  wire core__abc_21380_n8487;
  wire core__abc_21380_n8488;
  wire core__abc_21380_n8489;
  wire core__abc_21380_n8490;
  wire core__abc_21380_n8491;
  wire core__abc_21380_n8492;
  wire core__abc_21380_n8493;
  wire core__abc_21380_n8494;
  wire core__abc_21380_n8495;
  wire core__abc_21380_n8497;
  wire core__abc_21380_n8498;
  wire core__abc_21380_n8499;
  wire core__abc_21380_n8500;
  wire core__abc_21380_n8501;
  wire core__abc_21380_n8502;
  wire core__abc_21380_n8503;
  wire core__abc_21380_n8504;
  wire core__abc_21380_n8505;
  wire core__abc_21380_n8506;
  wire core__abc_21380_n8507;
  wire core__abc_21380_n8508;
  wire core__abc_21380_n8509;
  wire core__abc_21380_n8510;
  wire core__abc_21380_n8511;
  wire core__abc_21380_n8512;
  wire core__abc_21380_n8514;
  wire core__abc_21380_n8515;
  wire core__abc_21380_n8516;
  wire core__abc_21380_n8517;
  wire core__abc_21380_n8518;
  wire core__abc_21380_n8519;
  wire core__abc_21380_n8520;
  wire core__abc_21380_n8521;
  wire core__abc_21380_n8522;
  wire core__abc_21380_n8523;
  wire core__abc_21380_n8524;
  wire core__abc_21380_n8525;
  wire core__abc_21380_n8527;
  wire core__abc_21380_n8528;
  wire core__abc_21380_n8529;
  wire core__abc_21380_n8530;
  wire core__abc_21380_n8531;
  wire core__abc_21380_n8532;
  wire core__abc_21380_n8533;
  wire core__abc_21380_n8534;
  wire core__abc_21380_n8535;
  wire core__abc_21380_n8536;
  wire core__abc_21380_n8537;
  wire core__abc_21380_n8538;
  wire core__abc_21380_n8539;
  wire core__abc_21380_n8540;
  wire core__abc_21380_n8541;
  wire core__abc_21380_n8543;
  wire core__abc_21380_n8544;
  wire core__abc_21380_n8545;
  wire core__abc_21380_n8546;
  wire core__abc_21380_n8547;
  wire core__abc_21380_n8548;
  wire core__abc_21380_n8549;
  wire core__abc_21380_n8550;
  wire core__abc_21380_n8551;
  wire core__abc_21380_n8552;
  wire core__abc_21380_n8553;
  wire core__abc_21380_n8554;
  wire core__abc_21380_n8555;
  wire core__abc_21380_n8556;
  wire core__abc_21380_n8557;
  wire core__abc_21380_n8559;
  wire core__abc_21380_n8560;
  wire core__abc_21380_n8561;
  wire core__abc_21380_n8562;
  wire core__abc_21380_n8563;
  wire core__abc_21380_n8564;
  wire core__abc_21380_n8565;
  wire core__abc_21380_n8566;
  wire core__abc_21380_n8567;
  wire core__abc_21380_n8568;
  wire core__abc_21380_n8569;
  wire core__abc_21380_n8570;
  wire core__abc_21380_n8571;
  wire core__abc_21380_n8572;
  wire core__abc_21380_n8573;
  wire core__abc_21380_n8574;
  wire core__abc_21380_n8576;
  wire core__abc_21380_n8577;
  wire core__abc_21380_n8578;
  wire core__abc_21380_n8579;
  wire core__abc_21380_n8580;
  wire core__abc_21380_n8581;
  wire core__abc_21380_n8582;
  wire core__abc_21380_n8583;
  wire core__abc_21380_n8584;
  wire core__abc_21380_n8585;
  wire core__abc_21380_n8587;
  wire core__abc_21380_n8588;
  wire core__abc_21380_n8589;
  wire core__abc_21380_n8590;
  wire core__abc_21380_n8591;
  wire core__abc_21380_n8592;
  wire core__abc_21380_n8593;
  wire core__abc_21380_n8594;
  wire core__abc_21380_n8595;
  wire core__abc_21380_n8596;
  wire core__abc_21380_n8597;
  wire core__abc_21380_n8598;
  wire core__abc_21380_n8600;
  wire core__abc_21380_n8601;
  wire core__abc_21380_n8602;
  wire core__abc_21380_n8603;
  wire core__abc_21380_n8604;
  wire core__abc_21380_n8605;
  wire core__abc_21380_n8606;
  wire core__abc_21380_n8607;
  wire core__abc_21380_n8608;
  wire core__abc_21380_n8609;
  wire core__abc_21380_n8610;
  wire core__abc_21380_n8612;
  wire core__abc_21380_n8613;
  wire core__abc_21380_n8614;
  wire core__abc_21380_n8615;
  wire core__abc_21380_n8616;
  wire core__abc_21380_n8617;
  wire core__abc_21380_n8618;
  wire core__abc_21380_n8619;
  wire core__abc_21380_n8620;
  wire core__abc_21380_n8621;
  wire core__abc_21380_n8622;
  wire core__abc_21380_n8623;
  wire core__abc_21380_n8624;
  wire core__abc_21380_n8626;
  wire core__abc_21380_n8627;
  wire core__abc_21380_n8628;
  wire core__abc_21380_n8629;
  wire core__abc_21380_n8630;
  wire core__abc_21380_n8631;
  wire core__abc_21380_n8632;
  wire core__abc_21380_n8633;
  wire core__abc_21380_n8634;
  wire core__abc_21380_n8635;
  wire core__abc_21380_n8637;
  wire core__abc_21380_n8638;
  wire core__abc_21380_n8639;
  wire core__abc_21380_n8640;
  wire core__abc_21380_n8641;
  wire core__abc_21380_n8642;
  wire core__abc_21380_n8643;
  wire core__abc_21380_n8644;
  wire core__abc_21380_n8645;
  wire core__abc_21380_n8646;
  wire core__abc_21380_n8648;
  wire core__abc_21380_n8649;
  wire core__abc_21380_n8650;
  wire core__abc_21380_n8651;
  wire core__abc_21380_n8652;
  wire core__abc_21380_n8653;
  wire core__abc_21380_n8654;
  wire core__abc_21380_n8655;
  wire core__abc_21380_n8656;
  wire core__abc_21380_n8657;
  wire core__abc_21380_n8658;
  wire core__abc_21380_n8660;
  wire core__abc_21380_n8661;
  wire core__abc_21380_n8662;
  wire core__abc_21380_n8663;
  wire core__abc_21380_n8664;
  wire core__abc_21380_n8665;
  wire core__abc_21380_n8666;
  wire core__abc_21380_n8667;
  wire core__abc_21380_n8668;
  wire core__abc_21380_n8669;
  wire core__abc_21380_n8671;
  wire core__abc_21380_n8672;
  wire core__abc_21380_n8673;
  wire core__abc_21380_n8674;
  wire core__abc_21380_n8675;
  wire core__abc_21380_n8676;
  wire core__abc_21380_n8677;
  wire core__abc_21380_n8678;
  wire core__abc_21380_n8679;
  wire core__abc_21380_n8680;
  wire core__abc_21380_n8682;
  wire core__abc_21380_n8683;
  wire core__abc_21380_n8684;
  wire core__abc_21380_n8685;
  wire core__abc_21380_n8686;
  wire core__abc_21380_n8687;
  wire core__abc_21380_n8688;
  wire core__abc_21380_n8689;
  wire core__abc_21380_n8690;
  wire core__abc_21380_n8691;
  wire core__abc_21380_n8692;
  wire core__abc_21380_n8694;
  wire core__abc_21380_n8695;
  wire core__abc_21380_n8696;
  wire core__abc_21380_n8697;
  wire core__abc_21380_n8698;
  wire core__abc_21380_n8699;
  wire core__abc_21380_n8700;
  wire core__abc_21380_n8701;
  wire core__abc_21380_n8702;
  wire core__abc_21380_n8703;
  wire core__abc_21380_n8705;
  wire core__abc_21380_n8706;
  wire core__abc_21380_n8707;
  wire core__abc_21380_n8708;
  wire core__abc_21380_n8709;
  wire core__abc_21380_n8710;
  wire core__abc_21380_n8711;
  wire core__abc_21380_n8712;
  wire core__abc_21380_n8713;
  wire core__abc_21380_n8714;
  wire core__abc_21380_n8716;
  wire core__abc_21380_n8717;
  wire core__abc_21380_n8718;
  wire core__abc_21380_n8719;
  wire core__abc_21380_n8720;
  wire core__abc_21380_n8721;
  wire core__abc_21380_n8722;
  wire core__abc_21380_n8723;
  wire core__abc_21380_n8724;
  wire core__abc_21380_n8725;
  wire core__abc_21380_n8726;
  wire core__abc_21380_n8727;
  wire core__abc_21380_n8728;
  wire core__abc_21380_n8730;
  wire core__abc_21380_n8731;
  wire core__abc_21380_n8732;
  wire core__abc_21380_n8733;
  wire core__abc_21380_n8734;
  wire core__abc_21380_n8735;
  wire core__abc_21380_n8736;
  wire core__abc_21380_n8737;
  wire core__abc_21380_n8738;
  wire core__abc_21380_n8739;
  wire core__abc_21380_n8740;
  wire core__abc_21380_n8742;
  wire core__abc_21380_n8743;
  wire core__abc_21380_n8744;
  wire core__abc_21380_n8745;
  wire core__abc_21380_n8746;
  wire core__abc_21380_n8747;
  wire core__abc_21380_n8748;
  wire core__abc_21380_n8749;
  wire core__abc_21380_n8750;
  wire core__abc_21380_n8751;
  wire core__abc_21380_n8753;
  wire core__abc_21380_n8754;
  wire core__abc_21380_n8755;
  wire core__abc_21380_n8756;
  wire core__abc_21380_n8757;
  wire core__abc_21380_n8758;
  wire core__abc_21380_n8759;
  wire core__abc_21380_n8760;
  wire core__abc_21380_n8761;
  wire core__abc_21380_n8762;
  wire core__abc_21380_n8763;
  wire core__abc_21380_n8765;
  wire core__abc_21380_n8766;
  wire core__abc_21380_n8767;
  wire core__abc_21380_n8768;
  wire core__abc_21380_n8769;
  wire core__abc_21380_n8770;
  wire core__abc_21380_n8771;
  wire core__abc_21380_n8772;
  wire core__abc_21380_n8773;
  wire core__abc_21380_n8774;
  wire core__abc_21380_n8775;
  wire core__abc_21380_n8777;
  wire core__abc_21380_n8778;
  wire core__abc_21380_n8779;
  wire core__abc_21380_n8780;
  wire core__abc_21380_n8781;
  wire core__abc_21380_n8782;
  wire core__abc_21380_n8783;
  wire core__abc_21380_n8784;
  wire core__abc_21380_n8785;
  wire core__abc_21380_n8786;
  wire core__abc_21380_n8787;
  wire core__abc_21380_n8788;
  wire core__abc_21380_n8789;
  wire core__abc_21380_n8791;
  wire core__abc_21380_n8792;
  wire core__abc_21380_n8793;
  wire core__abc_21380_n8794;
  wire core__abc_21380_n8795;
  wire core__abc_21380_n8796;
  wire core__abc_21380_n8797;
  wire core__abc_21380_n8798;
  wire core__abc_21380_n8799;
  wire core__abc_21380_n8800;
  wire core__abc_21380_n8801;
  wire core__abc_21380_n8802;
  wire core__abc_21380_n8804;
  wire core__abc_21380_n8805;
  wire core__abc_21380_n8806;
  wire core__abc_21380_n8807;
  wire core__abc_21380_n8808;
  wire core__abc_21380_n8809;
  wire core__abc_21380_n8810;
  wire core__abc_21380_n8811;
  wire core__abc_21380_n8812;
  wire core__abc_21380_n8813;
  wire core__abc_21380_n8814;
  wire core__abc_21380_n8816;
  wire core__abc_21380_n8817;
  wire core__abc_21380_n8818;
  wire core__abc_21380_n8819;
  wire core__abc_21380_n8820;
  wire core__abc_21380_n8821;
  wire core__abc_21380_n8822;
  wire core__abc_21380_n8823;
  wire core__abc_21380_n8824;
  wire core__abc_21380_n8825;
  wire core__abc_21380_n8826;
  wire core__abc_21380_n8827;
  wire core__abc_21380_n8829;
  wire core__abc_21380_n8830;
  wire core__abc_21380_n8831;
  wire core__abc_21380_n8832;
  wire core__abc_21380_n8833;
  wire core__abc_21380_n8834;
  wire core__abc_21380_n8835;
  wire core__abc_21380_n8836;
  wire core__abc_21380_n8837;
  wire core__abc_21380_n8838;
  wire core__abc_21380_n8839;
  wire core__abc_21380_n8841;
  wire core__abc_21380_n8842;
  wire core__abc_21380_n8843;
  wire core__abc_21380_n8844;
  wire core__abc_21380_n8845;
  wire core__abc_21380_n8846;
  wire core__abc_21380_n8847;
  wire core__abc_21380_n8848;
  wire core__abc_21380_n8849;
  wire core__abc_21380_n8850;
  wire core__abc_21380_n8852;
  wire core__abc_21380_n8853;
  wire core__abc_21380_n8854;
  wire core__abc_21380_n8855;
  wire core__abc_21380_n8856;
  wire core__abc_21380_n8857;
  wire core__abc_21380_n8858;
  wire core__abc_21380_n8859;
  wire core__abc_21380_n8860;
  wire core__abc_21380_n8861;
  wire core__abc_21380_n8862;
  wire core__abc_21380_n8864;
  wire core__abc_21380_n8865;
  wire core__abc_21380_n8866;
  wire core__abc_21380_n8867;
  wire core__abc_21380_n8868;
  wire core__abc_21380_n8869;
  wire core__abc_21380_n8870;
  wire core__abc_21380_n8871;
  wire core__abc_21380_n8872;
  wire core__abc_21380_n8873;
  wire core__abc_21380_n8874;
  wire core__abc_21380_n8875;
  wire core__abc_21380_n8876;
  wire core__abc_21380_n8878;
  wire core__abc_21380_n8879;
  wire core__abc_21380_n8880;
  wire core__abc_21380_n8881;
  wire core__abc_21380_n8882;
  wire core__abc_21380_n8883;
  wire core__abc_21380_n8884;
  wire core__abc_21380_n8885;
  wire core__abc_21380_n8886;
  wire core__abc_21380_n8887;
  wire core__abc_21380_n8888;
  wire core__abc_21380_n8890;
  wire core__abc_21380_n8891;
  wire core__abc_21380_n8892;
  wire core__abc_21380_n8893;
  wire core__abc_21380_n8894;
  wire core__abc_21380_n8895;
  wire core__abc_21380_n8896;
  wire core__abc_21380_n8897;
  wire core__abc_21380_n8898;
  wire core__abc_21380_n8899;
  wire core__abc_21380_n8901;
  wire core__abc_21380_n8902;
  wire core__abc_21380_n8903;
  wire core__abc_21380_n8904;
  wire core__abc_21380_n8905;
  wire core__abc_21380_n8906;
  wire core__abc_21380_n8907;
  wire core__abc_21380_n8908;
  wire core__abc_21380_n8909;
  wire core__abc_21380_n8910;
  wire core__abc_21380_n8912;
  wire core__abc_21380_n8913;
  wire core__abc_21380_n8914;
  wire core__abc_21380_n8915;
  wire core__abc_21380_n8916;
  wire core__abc_21380_n8917;
  wire core__abc_21380_n8918;
  wire core__abc_21380_n8919;
  wire core__abc_21380_n8920;
  wire core__abc_21380_n8921;
  wire core__abc_21380_n8922;
  wire core__abc_21380_n8923;
  wire core__abc_21380_n8925;
  wire core__abc_21380_n8926;
  wire core__abc_21380_n8927;
  wire core__abc_21380_n8928;
  wire core__abc_21380_n8929;
  wire core__abc_21380_n8930;
  wire core__abc_21380_n8931;
  wire core__abc_21380_n8932;
  wire core__abc_21380_n8933;
  wire core__abc_21380_n8934;
  wire core__abc_21380_n8935;
  wire core__abc_21380_n8937;
  wire core__abc_21380_n8938;
  wire core__abc_21380_n8939;
  wire core__abc_21380_n8940;
  wire core__abc_21380_n8941;
  wire core__abc_21380_n8942;
  wire core__abc_21380_n8943;
  wire core__abc_21380_n8944;
  wire core__abc_21380_n8945;
  wire core__abc_21380_n8946;
  wire core__abc_21380_n8948;
  wire core__abc_21380_n8949;
  wire core__abc_21380_n8950;
  wire core__abc_21380_n8951;
  wire core__abc_21380_n8952;
  wire core__abc_21380_n8953;
  wire core__abc_21380_n8954;
  wire core__abc_21380_n8955;
  wire core__abc_21380_n8956;
  wire core__abc_21380_n8957;
  wire core__abc_21380_n8958;
  wire core__abc_21380_n8960;
  wire core__abc_21380_n8961;
  wire core__abc_21380_n8962;
  wire core__abc_21380_n8963;
  wire core__abc_21380_n8964;
  wire core__abc_21380_n8965;
  wire core__abc_21380_n8966;
  wire core__abc_21380_n8967;
  wire core__abc_21380_n8968;
  wire core__abc_21380_n8969;
  wire core__abc_21380_n8971;
  wire core__abc_21380_n8972;
  wire core__abc_21380_n8973;
  wire core__abc_21380_n8974;
  wire core__abc_21380_n8975;
  wire core__abc_21380_n8976;
  wire core__abc_21380_n8977;
  wire core__abc_21380_n8978;
  wire core__abc_21380_n8979;
  wire core__abc_21380_n8980;
  wire core__abc_21380_n8981;
  wire core__abc_21380_n8982;
  wire core__abc_21380_n8983;
  wire core__abc_21380_n8985;
  wire core__abc_21380_n8986;
  wire core__abc_21380_n8987;
  wire core__abc_21380_n8988;
  wire core__abc_21380_n8989;
  wire core__abc_21380_n8990;
  wire core__abc_21380_n8991;
  wire core__abc_21380_n8992;
  wire core__abc_21380_n8993;
  wire core__abc_21380_n8994;
  wire core__abc_21380_n8995;
  wire core__abc_21380_n8997;
  wire core__abc_21380_n8998;
  wire core__abc_21380_n8999;
  wire core__abc_21380_n9000;
  wire core__abc_21380_n9001;
  wire core__abc_21380_n9002;
  wire core__abc_21380_n9003;
  wire core__abc_21380_n9004;
  wire core__abc_21380_n9005;
  wire core__abc_21380_n9006;
  wire core__abc_21380_n9008;
  wire core__abc_21380_n9009;
  wire core__abc_21380_n9010;
  wire core__abc_21380_n9011;
  wire core__abc_21380_n9012;
  wire core__abc_21380_n9013;
  wire core__abc_21380_n9014;
  wire core__abc_21380_n9015;
  wire core__abc_21380_n9016;
  wire core__abc_21380_n9017;
  wire core__abc_21380_n9018;
  wire core__abc_21380_n9019;
  wire core__abc_21380_n9020;
  wire core__abc_21380_n9021;
  wire core__abc_21380_n9023;
  wire core__abc_21380_n9024;
  wire core__abc_21380_n9025;
  wire core__abc_21380_n9026;
  wire core__abc_21380_n9027;
  wire core__abc_21380_n9028;
  wire core__abc_21380_n9029;
  wire core__abc_21380_n9030;
  wire core__abc_21380_n9031;
  wire core__abc_21380_n9032;
  wire core__abc_21380_n9034;
  wire core__abc_21380_n9035;
  wire core__abc_21380_n9036;
  wire core__abc_21380_n9037;
  wire core__abc_21380_n9038;
  wire core__abc_21380_n9039;
  wire core__abc_21380_n9040;
  wire core__abc_21380_n9041;
  wire core__abc_21380_n9042;
  wire core__abc_21380_n9043;
  wire core__abc_21380_n9045;
  wire core__abc_21380_n9046;
  wire core__abc_21380_n9047;
  wire core__abc_21380_n9048;
  wire core__abc_21380_n9049;
  wire core__abc_21380_n9050;
  wire core__abc_21380_n9051;
  wire core__abc_21380_n9052;
  wire core__abc_21380_n9053;
  wire core__abc_21380_n9054;
  wire core__abc_21380_n9056;
  wire core__abc_21380_n9057;
  wire core__abc_21380_n9058;
  wire core__abc_21380_n9059;
  wire core__abc_21380_n9060;
  wire core__abc_21380_n9061;
  wire core__abc_21380_n9062;
  wire core__abc_21380_n9063;
  wire core__abc_21380_n9064;
  wire core__abc_21380_n9065;
  wire core__abc_21380_n9067;
  wire core__abc_21380_n9068;
  wire core__abc_21380_n9069;
  wire core__abc_21380_n9070;
  wire core__abc_21380_n9071;
  wire core__abc_21380_n9072;
  wire core__abc_21380_n9073;
  wire core__abc_21380_n9074;
  wire core__abc_21380_n9075;
  wire core__abc_21380_n9076;
  wire core__abc_21380_n9077;
  wire core__abc_21380_n9078;
  wire core__abc_21380_n9079;
  wire core__abc_21380_n9081;
  wire core__abc_21380_n9082;
  wire core__abc_21380_n9083;
  wire core__abc_21380_n9084;
  wire core__abc_21380_n9085;
  wire core__abc_21380_n9086;
  wire core__abc_21380_n9087;
  wire core__abc_21380_n9088;
  wire core__abc_21380_n9089;
  wire core__abc_21380_n9090;
  wire core__abc_21380_n9092;
  wire core__abc_21380_n9093;
  wire core__abc_21380_n9094;
  wire core__abc_21380_n9095;
  wire core__abc_21380_n9096;
  wire core__abc_21380_n9097;
  wire core__abc_21380_n9098;
  wire core__abc_21380_n9099;
  wire core__abc_21380_n9100;
  wire core__abc_21380_n9101;
  wire core__abc_21380_n9102;
  wire core__abc_21380_n9103;
  wire core__abc_21380_n9104;
  wire core__abc_21380_n9106;
  wire core__abc_21380_n9107;
  wire core__abc_21380_n9108;
  wire core__abc_21380_n9109;
  wire core__abc_21380_n9110;
  wire core__abc_21380_n9111;
  wire core__abc_21380_n9112;
  wire core__abc_21380_n9113;
  wire core__abc_21380_n9114;
  wire core__abc_21380_n9115;
  wire core__abc_21380_n9117;
  wire core__abc_21380_n9118;
  wire core__abc_21380_n9119;
  wire core__abc_21380_n9120;
  wire core__abc_21380_n9121;
  wire core__abc_21380_n9122;
  wire core__abc_21380_n9123;
  wire core__abc_21380_n9124;
  wire core__abc_21380_n9125;
  wire core__abc_21380_n9126;
  wire core__abc_21380_n9127;
  wire core__abc_21380_n9129;
  wire core__abc_21380_n9130;
  wire core__abc_21380_n9131;
  wire core__abc_21380_n9132;
  wire core__abc_21380_n9133;
  wire core__abc_21380_n9134;
  wire core__abc_21380_n9135;
  wire core__abc_21380_n9136;
  wire core__abc_21380_n9137;
  wire core__abc_21380_n9138;
  wire core__abc_21380_n9140;
  wire core__abc_21380_n9141;
  wire core__abc_21380_n9142;
  wire core__abc_21380_n9143;
  wire core__abc_21380_n9144;
  wire core__abc_21380_n9145;
  wire core__abc_21380_n9146;
  wire core__abc_21380_n9147;
  wire core__abc_21380_n9148;
  wire core__abc_21380_n9149;
  wire core__abc_21380_n9151;
  wire core__abc_21380_n9152;
  wire core__abc_21380_n9153;
  wire core__abc_21380_n9154;
  wire core__abc_21380_n9155;
  wire core__abc_21380_n9156;
  wire core__abc_21380_n9157;
  wire core__abc_21380_n9158;
  wire core__abc_21380_n9159;
  wire core__abc_21380_n9160;
  wire core__abc_21380_n9162;
  wire core__abc_21380_n9163;
  wire core__abc_21380_n9164;
  wire core__abc_21380_n9165;
  wire core__abc_21380_n9166;
  wire core__abc_21380_n9167;
  wire core__abc_21380_n9168;
  wire core__abc_21380_n9169;
  wire core__abc_21380_n9170;
  wire core__abc_21380_n9171;
  wire core__abc_21380_n9173;
  wire core__abc_21380_n9174;
  wire core__abc_21380_n9175;
  wire core__abc_21380_n9176;
  wire core__abc_21380_n9177;
  wire core__abc_21380_n9178;
  wire core__abc_21380_n9179;
  wire core__abc_21380_n9180;
  wire core__abc_21380_n9181;
  wire core__abc_21380_n9182;
  wire core__abc_21380_n9184;
  wire core__abc_21380_n9185;
  wire core__abc_21380_n9186;
  wire core__abc_21380_n9187;
  wire core__abc_21380_n9188;
  wire core__abc_21380_n9189;
  wire core__abc_21380_n9190;
  wire core__abc_21380_n9191;
  wire core__abc_21380_n9192;
  wire core__abc_21380_n9193;
  wire core__abc_21380_n9195;
  wire core__abc_21380_n9196;
  wire core__abc_21380_n9197;
  wire core__abc_21380_n9198;
  wire core__abc_21380_n9199;
  wire core__abc_21380_n9200;
  wire core__abc_21380_n9201;
  wire core__abc_21380_n9202;
  wire core__abc_21380_n9203;
  wire core__abc_21380_n9204;
  wire core__abc_21380_n9205;
  wire core__abc_21380_n9207;
  wire core__abc_21380_n9208;
  wire core__abc_21380_n9209;
  wire core__abc_21380_n9210;
  wire core__abc_21380_n9211;
  wire core__abc_21380_n9212;
  wire core__abc_21380_n9213;
  wire core__abc_21380_n9214;
  wire core__abc_21380_n9215;
  wire core__abc_21380_n9216;
  wire core__abc_21380_n9218;
  wire core__abc_21380_n9219;
  wire core__abc_21380_n9220;
  wire core__abc_21380_n9221;
  wire core__abc_21380_n9222;
  wire core__abc_21380_n9223;
  wire core__abc_21380_n9224;
  wire core__abc_21380_n9225;
  wire core__abc_21380_n9226;
  wire core__abc_21380_n9227;
  wire core__abc_21380_n9228;
  wire core__abc_21380_n9230;
  wire core__abc_21380_n9231;
  wire core__abc_21380_n9232;
  wire core__abc_21380_n9233;
  wire core__abc_21380_n9234;
  wire core__abc_21380_n9235;
  wire core__abc_21380_n9236;
  wire core__abc_21380_n9237;
  wire core__abc_21380_n9238;
  wire core__abc_21380_n9239;
  wire core__abc_21380_n9240;
  wire core__abc_21380_n9241;
  wire core__abc_21380_n9242;
  wire core__abc_21380_n9244;
  wire core__abc_21380_n9245;
  wire core__abc_21380_n9245_bF_buf0;
  wire core__abc_21380_n9245_bF_buf1;
  wire core__abc_21380_n9245_bF_buf2;
  wire core__abc_21380_n9245_bF_buf3;
  wire core__abc_21380_n9245_bF_buf4;
  wire core__abc_21380_n9245_bF_buf5;
  wire core__abc_21380_n9245_bF_buf6;
  wire core__abc_21380_n9245_bF_buf7;
  wire core__abc_21380_n9246;
  wire core__abc_21380_n9246_bF_buf0;
  wire core__abc_21380_n9246_bF_buf1;
  wire core__abc_21380_n9246_bF_buf2;
  wire core__abc_21380_n9246_bF_buf3;
  wire core__abc_21380_n9246_bF_buf4;
  wire core__abc_21380_n9246_bF_buf5;
  wire core__abc_21380_n9246_bF_buf6;
  wire core__abc_21380_n9246_bF_buf7;
  wire core__abc_21380_n9247;
  wire core__abc_21380_n9248;
  wire core__abc_21380_n9248_bF_buf0;
  wire core__abc_21380_n9248_bF_buf1;
  wire core__abc_21380_n9248_bF_buf2;
  wire core__abc_21380_n9248_bF_buf3;
  wire core__abc_21380_n9248_bF_buf4;
  wire core__abc_21380_n9248_bF_buf5;
  wire core__abc_21380_n9248_bF_buf6;
  wire core__abc_21380_n9248_bF_buf7;
  wire core__abc_21380_n9249;
  wire core__abc_21380_n9250;
  wire core__abc_21380_n9251;
  wire core__abc_21380_n9252;
  wire core__abc_21380_n9253;
  wire core__abc_21380_n9254;
  wire core__abc_21380_n9255;
  wire core__abc_21380_n9256;
  wire core__abc_21380_n9257;
  wire core__abc_21380_n9258;
  wire core__abc_21380_n9260;
  wire core__abc_21380_n9261;
  wire core__abc_21380_n9262;
  wire core__abc_21380_n9263;
  wire core__abc_21380_n9264;
  wire core__abc_21380_n9265;
  wire core__abc_21380_n9266;
  wire core__abc_21380_n9267;
  wire core__abc_21380_n9268;
  wire core__abc_21380_n9269;
  wire core__abc_21380_n9270;
  wire core__abc_21380_n9272;
  wire core__abc_21380_n9273;
  wire core__abc_21380_n9274;
  wire core__abc_21380_n9275;
  wire core__abc_21380_n9276;
  wire core__abc_21380_n9277;
  wire core__abc_21380_n9278;
  wire core__abc_21380_n9279;
  wire core__abc_21380_n9280;
  wire core__abc_21380_n9281;
  wire core__abc_21380_n9282;
  wire core__abc_21380_n9283;
  wire core__abc_21380_n9284;
  wire core__abc_21380_n9286;
  wire core__abc_21380_n9287;
  wire core__abc_21380_n9288;
  wire core__abc_21380_n9289;
  wire core__abc_21380_n9290;
  wire core__abc_21380_n9291;
  wire core__abc_21380_n9292;
  wire core__abc_21380_n9293;
  wire core__abc_21380_n9294;
  wire core__abc_21380_n9295;
  wire core__abc_21380_n9296;
  wire core__abc_21380_n9298;
  wire core__abc_21380_n9299;
  wire core__abc_21380_n9300;
  wire core__abc_21380_n9301;
  wire core__abc_21380_n9302;
  wire core__abc_21380_n9303;
  wire core__abc_21380_n9304;
  wire core__abc_21380_n9305;
  wire core__abc_21380_n9306;
  wire core__abc_21380_n9307;
  wire core__abc_21380_n9308;
  wire core__abc_21380_n9309;
  wire core__abc_21380_n9310;
  wire core__abc_21380_n9312;
  wire core__abc_21380_n9313;
  wire core__abc_21380_n9314;
  wire core__abc_21380_n9315;
  wire core__abc_21380_n9316;
  wire core__abc_21380_n9317;
  wire core__abc_21380_n9318;
  wire core__abc_21380_n9319;
  wire core__abc_21380_n9320;
  wire core__abc_21380_n9321;
  wire core__abc_21380_n9322;
  wire core__abc_21380_n9324;
  wire core__abc_21380_n9325;
  wire core__abc_21380_n9326;
  wire core__abc_21380_n9327;
  wire core__abc_21380_n9328;
  wire core__abc_21380_n9329;
  wire core__abc_21380_n9330;
  wire core__abc_21380_n9331;
  wire core__abc_21380_n9332;
  wire core__abc_21380_n9333;
  wire core__abc_21380_n9334;
  wire core__abc_21380_n9336;
  wire core__abc_21380_n9337;
  wire core__abc_21380_n9338;
  wire core__abc_21380_n9339;
  wire core__abc_21380_n9340;
  wire core__abc_21380_n9341;
  wire core__abc_21380_n9342;
  wire core__abc_21380_n9343;
  wire core__abc_21380_n9344;
  wire core__abc_21380_n9345;
  wire core__abc_21380_n9346;
  wire core__abc_21380_n9348;
  wire core__abc_21380_n9349;
  wire core__abc_21380_n9350;
  wire core__abc_21380_n9351;
  wire core__abc_21380_n9352;
  wire core__abc_21380_n9353;
  wire core__abc_21380_n9354;
  wire core__abc_21380_n9355;
  wire core__abc_21380_n9356;
  wire core__abc_21380_n9357;
  wire core__abc_21380_n9358;
  wire core__abc_21380_n9359;
  wire core__abc_21380_n9360;
  wire core__abc_21380_n9362;
  wire core__abc_21380_n9363;
  wire core__abc_21380_n9364;
  wire core__abc_21380_n9365;
  wire core__abc_21380_n9366;
  wire core__abc_21380_n9367;
  wire core__abc_21380_n9368;
  wire core__abc_21380_n9369;
  wire core__abc_21380_n9370;
  wire core__abc_21380_n9371;
  wire core__abc_21380_n9372;
  wire core__abc_21380_n9373;
  wire core__abc_21380_n9375;
  wire core__abc_21380_n9376;
  wire core__abc_21380_n9377;
  wire core__abc_21380_n9378;
  wire core__abc_21380_n9379;
  wire core__abc_21380_n9380;
  wire core__abc_21380_n9381;
  wire core__abc_21380_n9382;
  wire core__abc_21380_n9383;
  wire core__abc_21380_n9384;
  wire core__abc_21380_n9385;
  wire core__abc_21380_n9386;
  wire core__abc_21380_n9387;
  wire core__abc_21380_n9389;
  wire core__abc_21380_n9390;
  wire core__abc_21380_n9391;
  wire core__abc_21380_n9392;
  wire core__abc_21380_n9393;
  wire core__abc_21380_n9394;
  wire core__abc_21380_n9395;
  wire core__abc_21380_n9396;
  wire core__abc_21380_n9397;
  wire core__abc_21380_n9398;
  wire core__abc_21380_n9399;
  wire core__abc_21380_n9400;
  wire core__abc_21380_n9402;
  wire core__abc_21380_n9403;
  wire core__abc_21380_n9404;
  wire core__abc_21380_n9405;
  wire core__abc_21380_n9406;
  wire core__abc_21380_n9407;
  wire core__abc_21380_n9408;
  wire core__abc_21380_n9409;
  wire core__abc_21380_n9410;
  wire core__abc_21380_n9411;
  wire core__abc_21380_n9412;
  wire core__abc_21380_n9413;
  wire core__abc_21380_n9415;
  wire core__abc_21380_n9416;
  wire core__abc_21380_n9417;
  wire core__abc_21380_n9418;
  wire core__abc_21380_n9419;
  wire core__abc_21380_n9420;
  wire core__abc_21380_n9421;
  wire core__abc_21380_n9422;
  wire core__abc_21380_n9423;
  wire core__abc_21380_n9424;
  wire core__abc_21380_n9425;
  wire core__abc_21380_n9427;
  wire core__abc_21380_n9428;
  wire core__abc_21380_n9429;
  wire core__abc_21380_n9430;
  wire core__abc_21380_n9431;
  wire core__abc_21380_n9432;
  wire core__abc_21380_n9433;
  wire core__abc_21380_n9434;
  wire core__abc_21380_n9435;
  wire core__abc_21380_n9436;
  wire core__abc_21380_n9437;
  wire core__abc_21380_n9439;
  wire core__abc_21380_n9440;
  wire core__abc_21380_n9441;
  wire core__abc_21380_n9442;
  wire core__abc_21380_n9443;
  wire core__abc_21380_n9444;
  wire core__abc_21380_n9445;
  wire core__abc_21380_n9446;
  wire core__abc_21380_n9447;
  wire core__abc_21380_n9448;
  wire core__abc_21380_n9449;
  wire core__abc_21380_n9451;
  wire core__abc_21380_n9452;
  wire core__abc_21380_n9453;
  wire core__abc_21380_n9454;
  wire core__abc_21380_n9455;
  wire core__abc_21380_n9456;
  wire core__abc_21380_n9457;
  wire core__abc_21380_n9458;
  wire core__abc_21380_n9459;
  wire core__abc_21380_n9460;
  wire core__abc_21380_n9461;
  wire core__abc_21380_n9463;
  wire core__abc_21380_n9464;
  wire core__abc_21380_n9465;
  wire core__abc_21380_n9466;
  wire core__abc_21380_n9467;
  wire core__abc_21380_n9468;
  wire core__abc_21380_n9469;
  wire core__abc_21380_n9470;
  wire core__abc_21380_n9471;
  wire core__abc_21380_n9472;
  wire core__abc_21380_n9473;
  wire core__abc_21380_n9474;
  wire core__abc_21380_n9475;
  wire core__abc_21380_n9477;
  wire core__abc_21380_n9478;
  wire core__abc_21380_n9479;
  wire core__abc_21380_n9480;
  wire core__abc_21380_n9481;
  wire core__abc_21380_n9482;
  wire core__abc_21380_n9483;
  wire core__abc_21380_n9484;
  wire core__abc_21380_n9485;
  wire core__abc_21380_n9486;
  wire core__abc_21380_n9487;
  wire core__abc_21380_n9488;
  wire core__abc_21380_n9489;
  wire core__abc_21380_n9491;
  wire core__abc_21380_n9492;
  wire core__abc_21380_n9493;
  wire core__abc_21380_n9494;
  wire core__abc_21380_n9495;
  wire core__abc_21380_n9496;
  wire core__abc_21380_n9497;
  wire core__abc_21380_n9498;
  wire core__abc_21380_n9499;
  wire core__abc_21380_n9500;
  wire core__abc_21380_n9501;
  wire core__abc_21380_n9503;
  wire core__abc_21380_n9504;
  wire core__abc_21380_n9505;
  wire core__abc_21380_n9506;
  wire core__abc_21380_n9507;
  wire core__abc_21380_n9508;
  wire core__abc_21380_n9509;
  wire core__abc_21380_n9510;
  wire core__abc_21380_n9511;
  wire core__abc_21380_n9512;
  wire core__abc_21380_n9513;
  wire core__abc_21380_n9514;
  wire core__abc_21380_n9515;
  wire core__abc_21380_n9517;
  wire core__abc_21380_n9518;
  wire core__abc_21380_n9519;
  wire core__abc_21380_n9520;
  wire core__abc_21380_n9521;
  wire core__abc_21380_n9522;
  wire core__abc_21380_n9523;
  wire core__abc_21380_n9524;
  wire core__abc_21380_n9525;
  wire core__abc_21380_n9526;
  wire core__abc_21380_n9527;
  wire core__abc_21380_n9529;
  wire core__abc_21380_n9530;
  wire core__abc_21380_n9531;
  wire core__abc_21380_n9532;
  wire core__abc_21380_n9533;
  wire core__abc_21380_n9534;
  wire core__abc_21380_n9535;
  wire core__abc_21380_n9536;
  wire core__abc_21380_n9537;
  wire core__abc_21380_n9538;
  wire core__abc_21380_n9539;
  wire core__abc_21380_n9541;
  wire core__abc_21380_n9542;
  wire core__abc_21380_n9543;
  wire core__abc_21380_n9544;
  wire core__abc_21380_n9545;
  wire core__abc_21380_n9546;
  wire core__abc_21380_n9547;
  wire core__abc_21380_n9548;
  wire core__abc_21380_n9549;
  wire core__abc_21380_n9550;
  wire core__abc_21380_n9551;
  wire core__abc_21380_n9553;
  wire core__abc_21380_n9554;
  wire core__abc_21380_n9555;
  wire core__abc_21380_n9556;
  wire core__abc_21380_n9557;
  wire core__abc_21380_n9558;
  wire core__abc_21380_n9559;
  wire core__abc_21380_n9560;
  wire core__abc_21380_n9561;
  wire core__abc_21380_n9562;
  wire core__abc_21380_n9563;
  wire core__abc_21380_n9565;
  wire core__abc_21380_n9566;
  wire core__abc_21380_n9567;
  wire core__abc_21380_n9568;
  wire core__abc_21380_n9569;
  wire core__abc_21380_n9570;
  wire core__abc_21380_n9571;
  wire core__abc_21380_n9572;
  wire core__abc_21380_n9573;
  wire core__abc_21380_n9574;
  wire core__abc_21380_n9575;
  wire core__abc_21380_n9576;
  wire core__abc_21380_n9578;
  wire core__abc_21380_n9579;
  wire core__abc_21380_n9580;
  wire core__abc_21380_n9581;
  wire core__abc_21380_n9582;
  wire core__abc_21380_n9583;
  wire core__abc_21380_n9584;
  wire core__abc_21380_n9585;
  wire core__abc_21380_n9586;
  wire core__abc_21380_n9587;
  wire core__abc_21380_n9588;
  wire core__abc_21380_n9589;
  wire core__abc_21380_n9591;
  wire core__abc_21380_n9592;
  wire core__abc_21380_n9593;
  wire core__abc_21380_n9594;
  wire core__abc_21380_n9595;
  wire core__abc_21380_n9596;
  wire core__abc_21380_n9597;
  wire core__abc_21380_n9598;
  wire core__abc_21380_n9599;
  wire core__abc_21380_n9600;
  wire core__abc_21380_n9601;
  wire core__abc_21380_n9602;
  wire core__abc_21380_n9604;
  wire core__abc_21380_n9605;
  wire core__abc_21380_n9606;
  wire core__abc_21380_n9607;
  wire core__abc_21380_n9608;
  wire core__abc_21380_n9609;
  wire core__abc_21380_n9610;
  wire core__abc_21380_n9611;
  wire core__abc_21380_n9612;
  wire core__abc_21380_n9613;
  wire core__abc_21380_n9614;
  wire core__abc_21380_n9615;
  wire core__abc_21380_n9616;
  wire core__abc_21380_n9618;
  wire core__abc_21380_n9619;
  wire core__abc_21380_n9620;
  wire core__abc_21380_n9621;
  wire core__abc_21380_n9622;
  wire core__abc_21380_n9623;
  wire core__abc_21380_n9624;
  wire core__abc_21380_n9625;
  wire core__abc_21380_n9626;
  wire core__abc_21380_n9627;
  wire core__abc_21380_n9628;
  wire core__abc_21380_n9630;
  wire core__abc_21380_n9631;
  wire core__abc_21380_n9632;
  wire core__abc_21380_n9633;
  wire core__abc_21380_n9634;
  wire core__abc_21380_n9635;
  wire core__abc_21380_n9636;
  wire core__abc_21380_n9637;
  wire core__abc_21380_n9638;
  wire core__abc_21380_n9639;
  wire core__abc_21380_n9640;
  wire core__abc_21380_n9642;
  wire core__abc_21380_n9643;
  wire core__abc_21380_n9644;
  wire core__abc_21380_n9645;
  wire core__abc_21380_n9646;
  wire core__abc_21380_n9647;
  wire core__abc_21380_n9648;
  wire core__abc_21380_n9649;
  wire core__abc_21380_n9650;
  wire core__abc_21380_n9651;
  wire core__abc_21380_n9652;
  wire core__abc_21380_n9654;
  wire core__abc_21380_n9655;
  wire core__abc_21380_n9656;
  wire core__abc_21380_n9657;
  wire core__abc_21380_n9658;
  wire core__abc_21380_n9659;
  wire core__abc_21380_n9660;
  wire core__abc_21380_n9661;
  wire core__abc_21380_n9662;
  wire core__abc_21380_n9663;
  wire core__abc_21380_n9664;
  wire core__abc_21380_n9666;
  wire core__abc_21380_n9667;
  wire core__abc_21380_n9668;
  wire core__abc_21380_n9669;
  wire core__abc_21380_n9670;
  wire core__abc_21380_n9671;
  wire core__abc_21380_n9672;
  wire core__abc_21380_n9673;
  wire core__abc_21380_n9674;
  wire core__abc_21380_n9675;
  wire core__abc_21380_n9676;
  wire core__abc_21380_n9678;
  wire core__abc_21380_n9679;
  wire core__abc_21380_n9680;
  wire core__abc_21380_n9681;
  wire core__abc_21380_n9682;
  wire core__abc_21380_n9683;
  wire core__abc_21380_n9684;
  wire core__abc_21380_n9685;
  wire core__abc_21380_n9686;
  wire core__abc_21380_n9687;
  wire core__abc_21380_n9688;
  wire core__abc_21380_n9690;
  wire core__abc_21380_n9691;
  wire core__abc_21380_n9692;
  wire core__abc_21380_n9693;
  wire core__abc_21380_n9694;
  wire core__abc_21380_n9695;
  wire core__abc_21380_n9696;
  wire core__abc_21380_n9697;
  wire core__abc_21380_n9698;
  wire core__abc_21380_n9699;
  wire core__abc_21380_n9700;
  wire core__abc_21380_n9702;
  wire core__abc_21380_n9703;
  wire core__abc_21380_n9704;
  wire core__abc_21380_n9705;
  wire core__abc_21380_n9706;
  wire core__abc_21380_n9707;
  wire core__abc_21380_n9708;
  wire core__abc_21380_n9709;
  wire core__abc_21380_n9710;
  wire core__abc_21380_n9711;
  wire core__abc_21380_n9712;
  wire core__abc_21380_n9714;
  wire core__abc_21380_n9715;
  wire core__abc_21380_n9716;
  wire core__abc_21380_n9717;
  wire core__abc_21380_n9718;
  wire core__abc_21380_n9719;
  wire core__abc_21380_n9720;
  wire core__abc_21380_n9721;
  wire core__abc_21380_n9722;
  wire core__abc_21380_n9723;
  wire core__abc_21380_n9724;
  wire core__abc_21380_n9726;
  wire core__abc_21380_n9727;
  wire core__abc_21380_n9728;
  wire core__abc_21380_n9729;
  wire core__abc_21380_n9730;
  wire core__abc_21380_n9731;
  wire core__abc_21380_n9732;
  wire core__abc_21380_n9733;
  wire core__abc_21380_n9734;
  wire core__abc_21380_n9735;
  wire core__abc_21380_n9736;
  wire core__abc_21380_n9738;
  wire core__abc_21380_n9739;
  wire core__abc_21380_n9740;
  wire core__abc_21380_n9741;
  wire core__abc_21380_n9742;
  wire core__abc_21380_n9743;
  wire core__abc_21380_n9744;
  wire core__abc_21380_n9745;
  wire core__abc_21380_n9746;
  wire core__abc_21380_n9747;
  wire core__abc_21380_n9748;
  wire core__abc_21380_n9750;
  wire core__abc_21380_n9751;
  wire core__abc_21380_n9752;
  wire core__abc_21380_n9753;
  wire core__abc_21380_n9754;
  wire core__abc_21380_n9755;
  wire core__abc_21380_n9756;
  wire core__abc_21380_n9757;
  wire core__abc_21380_n9758;
  wire core__abc_21380_n9759;
  wire core__abc_21380_n9760;
  wire core__abc_21380_n9762;
  wire core__abc_21380_n9763;
  wire core__abc_21380_n9764;
  wire core__abc_21380_n9765;
  wire core__abc_21380_n9766;
  wire core__abc_21380_n9767;
  wire core__abc_21380_n9768;
  wire core__abc_21380_n9769;
  wire core__abc_21380_n9770;
  wire core__abc_21380_n9771;
  wire core__abc_21380_n9772;
  wire core__abc_21380_n9773;
  wire core__abc_21380_n9775;
  wire core__abc_21380_n9776;
  wire core__abc_21380_n9777;
  wire core__abc_21380_n9778;
  wire core__abc_21380_n9779;
  wire core__abc_21380_n9780;
  wire core__abc_21380_n9781;
  wire core__abc_21380_n9782;
  wire core__abc_21380_n9783;
  wire core__abc_21380_n9784;
  wire core__abc_21380_n9785;
  wire core__abc_21380_n9787;
  wire core__abc_21380_n9788;
  wire core__abc_21380_n9789;
  wire core__abc_21380_n9790;
  wire core__abc_21380_n9791;
  wire core__abc_21380_n9792;
  wire core__abc_21380_n9793;
  wire core__abc_21380_n9794;
  wire core__abc_21380_n9795;
  wire core__abc_21380_n9796;
  wire core__abc_21380_n9797;
  wire core__abc_21380_n9798;
  wire core__abc_21380_n9799;
  wire core__abc_21380_n9801;
  wire core__abc_21380_n9802;
  wire core__abc_21380_n9803;
  wire core__abc_21380_n9804;
  wire core__abc_21380_n9805;
  wire core__abc_21380_n9806;
  wire core__abc_21380_n9807;
  wire core__abc_21380_n9808;
  wire core__abc_21380_n9809;
  wire core__abc_21380_n9810;
  wire core__abc_21380_n9811;
  wire core__abc_21380_n9813;
  wire core__abc_21380_n9814;
  wire core__abc_21380_n9815;
  wire core__abc_21380_n9816;
  wire core__abc_21380_n9817;
  wire core__abc_21380_n9818;
  wire core__abc_21380_n9819;
  wire core__abc_21380_n9820;
  wire core__abc_21380_n9821;
  wire core__abc_21380_n9822;
  wire core__abc_21380_n9823;
  wire core__abc_21380_n9825;
  wire core__abc_21380_n9826;
  wire core__abc_21380_n9827;
  wire core__abc_21380_n9828;
  wire core__abc_21380_n9829;
  wire core__abc_21380_n9830;
  wire core__abc_21380_n9831;
  wire core__abc_21380_n9832;
  wire core__abc_21380_n9833;
  wire core__abc_21380_n9834;
  wire core__abc_21380_n9835;
  wire core__abc_21380_n9837;
  wire core__abc_21380_n9838;
  wire core__abc_21380_n9839;
  wire core__abc_21380_n9840;
  wire core__abc_21380_n9841;
  wire core__abc_21380_n9842;
  wire core__abc_21380_n9843;
  wire core__abc_21380_n9844;
  wire core__abc_21380_n9845;
  wire core__abc_21380_n9846;
  wire core__abc_21380_n9847;
  wire core__abc_21380_n9849;
  wire core__abc_21380_n9850;
  wire core__abc_21380_n9851;
  wire core__abc_21380_n9852;
  wire core__abc_21380_n9853;
  wire core__abc_21380_n9854;
  wire core__abc_21380_n9855;
  wire core__abc_21380_n9856;
  wire core__abc_21380_n9857;
  wire core__abc_21380_n9858;
  wire core__abc_21380_n9859;
  wire core__abc_21380_n9861;
  wire core__abc_21380_n9862;
  wire core__abc_21380_n9863;
  wire core__abc_21380_n9864;
  wire core__abc_21380_n9865;
  wire core__abc_21380_n9866;
  wire core__abc_21380_n9867;
  wire core__abc_21380_n9868;
  wire core__abc_21380_n9869;
  wire core__abc_21380_n9870;
  wire core__abc_21380_n9871;
  wire core__abc_21380_n9872;
  wire core__abc_21380_n9873;
  wire core__abc_21380_n9875;
  wire core__abc_21380_n9876;
  wire core__abc_21380_n9877;
  wire core__abc_21380_n9878;
  wire core__abc_21380_n9879;
  wire core__abc_21380_n9880;
  wire core__abc_21380_n9881;
  wire core__abc_21380_n9882;
  wire core__abc_21380_n9883;
  wire core__abc_21380_n9884;
  wire core__abc_21380_n9885;
  wire core__abc_21380_n9886;
  wire core__abc_21380_n9887;
  wire core__abc_21380_n9889;
  wire core__abc_21380_n9890;
  wire core__abc_21380_n9891;
  wire core__abc_21380_n9892;
  wire core__abc_21380_n9893;
  wire core__abc_21380_n9894;
  wire core__abc_21380_n9895;
  wire core__abc_21380_n9896;
  wire core__abc_21380_n9897;
  wire core__abc_21380_n9898;
  wire core__abc_21380_n9899;
  wire core__abc_21380_n9901;
  wire core__abc_21380_n9902;
  wire core__abc_21380_n9903;
  wire core__abc_21380_n9904;
  wire core__abc_21380_n9905;
  wire core__abc_21380_n9906;
  wire core__abc_21380_n9907;
  wire core__abc_21380_n9908;
  wire core__abc_21380_n9909;
  wire core__abc_21380_n9910;
  wire core__abc_21380_n9911;
  wire core__abc_21380_n9912;
  wire core__abc_21380_n9914;
  wire core__abc_21380_n9915;
  wire core__abc_21380_n9916;
  wire core__abc_21380_n9917;
  wire core__abc_21380_n9918;
  wire core__abc_21380_n9919;
  wire core__abc_21380_n9920;
  wire core__abc_21380_n9921;
  wire core__abc_21380_n9922;
  wire core__abc_21380_n9923;
  wire core__abc_21380_n9924;
  wire core__abc_21380_n9926;
  wire core__abc_21380_n9927;
  wire core__abc_21380_n9928;
  wire core__abc_21380_n9929;
  wire core__abc_21380_n9930;
  wire core__abc_21380_n9931;
  wire core__abc_21380_n9932;
  wire core__abc_21380_n9933;
  wire core__abc_21380_n9934;
  wire core__abc_21380_n9935;
  wire core__abc_21380_n9936;
  wire core__abc_21380_n9938;
  wire core__abc_21380_n9939;
  wire core__abc_21380_n9940;
  wire core__abc_21380_n9941;
  wire core__abc_21380_n9942;
  wire core__abc_21380_n9943;
  wire core__abc_21380_n9944;
  wire core__abc_21380_n9945;
  wire core__abc_21380_n9946;
  wire core__abc_21380_n9947;
  wire core__abc_21380_n9948;
  wire core__abc_21380_n9950;
  wire core__abc_21380_n9951;
  wire core__abc_21380_n9952;
  wire core__abc_21380_n9953;
  wire core__abc_21380_n9954;
  wire core__abc_21380_n9955;
  wire core__abc_21380_n9956;
  wire core__abc_21380_n9957;
  wire core__abc_21380_n9958;
  wire core__abc_21380_n9959;
  wire core__abc_21380_n9960;
  wire core__abc_21380_n9961;
  wire core__abc_21380_n9962;
  wire core__abc_21380_n9964;
  wire core__abc_21380_n9965;
  wire core__abc_21380_n9966;
  wire core__abc_21380_n9967;
  wire core__abc_21380_n9968;
  wire core__abc_21380_n9969;
  wire core__abc_21380_n9970;
  wire core__abc_21380_n9971;
  wire core__abc_21380_n9972;
  wire core__abc_21380_n9973;
  wire core__abc_21380_n9974;
  wire core__abc_21380_n9975;
  wire core__abc_21380_n9976;
  wire core__abc_21380_n9978;
  wire core__abc_21380_n9979;
  wire core__abc_21380_n9980;
  wire core__abc_21380_n9981;
  wire core__abc_21380_n9982;
  wire core__abc_21380_n9983;
  wire core__abc_21380_n9984;
  wire core__abc_21380_n9985;
  wire core__abc_21380_n9986;
  wire core__abc_21380_n9987;
  wire core__abc_21380_n9988;
  wire core__abc_21380_n9989;
  wire core__abc_21380_n9991;
  wire core__abc_21380_n9992;
  wire core__abc_21380_n9993;
  wire core__abc_21380_n9994;
  wire core__abc_21380_n9995;
  wire core__abc_21380_n9996;
  wire core__abc_21380_n9997;
  wire core__abc_21380_n9998;
  wire core__abc_21380_n9999;
  wire core_compress;
  wire core_compression_rounds_0_;
  wire core_compression_rounds_1_;
  wire core_compression_rounds_2_;
  wire core_compression_rounds_3_;
  wire core_final_rounds_0_;
  wire core_final_rounds_1_;
  wire core_final_rounds_2_;
  wire core_final_rounds_3_;
  wire core_finalize;
  wire core_initalize;
  wire core_key_0_;
  wire core_key_100_;
  wire core_key_101_;
  wire core_key_102_;
  wire core_key_103_;
  wire core_key_104_;
  wire core_key_105_;
  wire core_key_106_;
  wire core_key_107_;
  wire core_key_108_;
  wire core_key_109_;
  wire core_key_10_;
  wire core_key_110_;
  wire core_key_111_;
  wire core_key_112_;
  wire core_key_113_;
  wire core_key_114_;
  wire core_key_115_;
  wire core_key_116_;
  wire core_key_117_;
  wire core_key_118_;
  wire core_key_119_;
  wire core_key_11_;
  wire core_key_120_;
  wire core_key_121_;
  wire core_key_122_;
  wire core_key_123_;
  wire core_key_124_;
  wire core_key_125_;
  wire core_key_126_;
  wire core_key_127_;
  wire core_key_12_;
  wire core_key_13_;
  wire core_key_14_;
  wire core_key_15_;
  wire core_key_16_;
  wire core_key_17_;
  wire core_key_18_;
  wire core_key_19_;
  wire core_key_1_;
  wire core_key_20_;
  wire core_key_21_;
  wire core_key_22_;
  wire core_key_23_;
  wire core_key_24_;
  wire core_key_25_;
  wire core_key_26_;
  wire core_key_27_;
  wire core_key_28_;
  wire core_key_29_;
  wire core_key_2_;
  wire core_key_30_;
  wire core_key_31_;
  wire core_key_32_;
  wire core_key_33_;
  wire core_key_34_;
  wire core_key_35_;
  wire core_key_36_;
  wire core_key_37_;
  wire core_key_38_;
  wire core_key_39_;
  wire core_key_3_;
  wire core_key_40_;
  wire core_key_41_;
  wire core_key_42_;
  wire core_key_43_;
  wire core_key_44_;
  wire core_key_45_;
  wire core_key_46_;
  wire core_key_47_;
  wire core_key_48_;
  wire core_key_49_;
  wire core_key_4_;
  wire core_key_50_;
  wire core_key_51_;
  wire core_key_52_;
  wire core_key_53_;
  wire core_key_54_;
  wire core_key_55_;
  wire core_key_56_;
  wire core_key_57_;
  wire core_key_58_;
  wire core_key_59_;
  wire core_key_5_;
  wire core_key_60_;
  wire core_key_61_;
  wire core_key_62_;
  wire core_key_63_;
  wire core_key_64_;
  wire core_key_65_;
  wire core_key_66_;
  wire core_key_67_;
  wire core_key_68_;
  wire core_key_69_;
  wire core_key_6_;
  wire core_key_70_;
  wire core_key_71_;
  wire core_key_72_;
  wire core_key_73_;
  wire core_key_74_;
  wire core_key_75_;
  wire core_key_76_;
  wire core_key_77_;
  wire core_key_78_;
  wire core_key_79_;
  wire core_key_7_;
  wire core_key_80_;
  wire core_key_81_;
  wire core_key_82_;
  wire core_key_83_;
  wire core_key_84_;
  wire core_key_85_;
  wire core_key_86_;
  wire core_key_87_;
  wire core_key_88_;
  wire core_key_89_;
  wire core_key_8_;
  wire core_key_90_;
  wire core_key_91_;
  wire core_key_92_;
  wire core_key_93_;
  wire core_key_94_;
  wire core_key_95_;
  wire core_key_96_;
  wire core_key_97_;
  wire core_key_98_;
  wire core_key_99_;
  wire core_key_9_;
  wire core_long;
  wire core_loop_ctr_reg_0_;
  wire core_loop_ctr_reg_0__FF_INPUT;
  wire core_loop_ctr_reg_1_;
  wire core_loop_ctr_reg_1__FF_INPUT;
  wire core_loop_ctr_reg_2_;
  wire core_loop_ctr_reg_2__FF_INPUT;
  wire core_loop_ctr_reg_3_;
  wire core_loop_ctr_reg_3__FF_INPUT;
  wire core_mi_0_;
  wire core_mi_10_;
  wire core_mi_11_;
  wire core_mi_12_;
  wire core_mi_13_;
  wire core_mi_14_;
  wire core_mi_15_;
  wire core_mi_16_;
  wire core_mi_17_;
  wire core_mi_18_;
  wire core_mi_19_;
  wire core_mi_1_;
  wire core_mi_20_;
  wire core_mi_21_;
  wire core_mi_22_;
  wire core_mi_23_;
  wire core_mi_24_;
  wire core_mi_25_;
  wire core_mi_26_;
  wire core_mi_27_;
  wire core_mi_28_;
  wire core_mi_29_;
  wire core_mi_2_;
  wire core_mi_30_;
  wire core_mi_31_;
  wire core_mi_32_;
  wire core_mi_33_;
  wire core_mi_34_;
  wire core_mi_35_;
  wire core_mi_36_;
  wire core_mi_37_;
  wire core_mi_38_;
  wire core_mi_39_;
  wire core_mi_3_;
  wire core_mi_40_;
  wire core_mi_41_;
  wire core_mi_42_;
  wire core_mi_43_;
  wire core_mi_44_;
  wire core_mi_45_;
  wire core_mi_46_;
  wire core_mi_47_;
  wire core_mi_48_;
  wire core_mi_49_;
  wire core_mi_4_;
  wire core_mi_50_;
  wire core_mi_51_;
  wire core_mi_52_;
  wire core_mi_53_;
  wire core_mi_54_;
  wire core_mi_55_;
  wire core_mi_56_;
  wire core_mi_57_;
  wire core_mi_58_;
  wire core_mi_59_;
  wire core_mi_5_;
  wire core_mi_60_;
  wire core_mi_61_;
  wire core_mi_62_;
  wire core_mi_63_;
  wire core_mi_6_;
  wire core_mi_7_;
  wire core_mi_8_;
  wire core_mi_9_;
  wire core_mi_reg_0_;
  wire core_mi_reg_0__FF_INPUT;
  wire core_mi_reg_10_;
  wire core_mi_reg_10__FF_INPUT;
  wire core_mi_reg_11_;
  wire core_mi_reg_11__FF_INPUT;
  wire core_mi_reg_12_;
  wire core_mi_reg_12__FF_INPUT;
  wire core_mi_reg_13_;
  wire core_mi_reg_13__FF_INPUT;
  wire core_mi_reg_14_;
  wire core_mi_reg_14__FF_INPUT;
  wire core_mi_reg_15_;
  wire core_mi_reg_15__FF_INPUT;
  wire core_mi_reg_16_;
  wire core_mi_reg_16__FF_INPUT;
  wire core_mi_reg_17_;
  wire core_mi_reg_17__FF_INPUT;
  wire core_mi_reg_18_;
  wire core_mi_reg_18__FF_INPUT;
  wire core_mi_reg_19_;
  wire core_mi_reg_19__FF_INPUT;
  wire core_mi_reg_1_;
  wire core_mi_reg_1__FF_INPUT;
  wire core_mi_reg_20_;
  wire core_mi_reg_20__FF_INPUT;
  wire core_mi_reg_21_;
  wire core_mi_reg_21__FF_INPUT;
  wire core_mi_reg_22_;
  wire core_mi_reg_22__FF_INPUT;
  wire core_mi_reg_23_;
  wire core_mi_reg_23__FF_INPUT;
  wire core_mi_reg_24_;
  wire core_mi_reg_24__FF_INPUT;
  wire core_mi_reg_25_;
  wire core_mi_reg_25__FF_INPUT;
  wire core_mi_reg_26_;
  wire core_mi_reg_26__FF_INPUT;
  wire core_mi_reg_27_;
  wire core_mi_reg_27__FF_INPUT;
  wire core_mi_reg_28_;
  wire core_mi_reg_28__FF_INPUT;
  wire core_mi_reg_29_;
  wire core_mi_reg_29__FF_INPUT;
  wire core_mi_reg_2_;
  wire core_mi_reg_2__FF_INPUT;
  wire core_mi_reg_30_;
  wire core_mi_reg_30__FF_INPUT;
  wire core_mi_reg_31_;
  wire core_mi_reg_31__FF_INPUT;
  wire core_mi_reg_32_;
  wire core_mi_reg_32__FF_INPUT;
  wire core_mi_reg_33_;
  wire core_mi_reg_33__FF_INPUT;
  wire core_mi_reg_34_;
  wire core_mi_reg_34__FF_INPUT;
  wire core_mi_reg_35_;
  wire core_mi_reg_35__FF_INPUT;
  wire core_mi_reg_36_;
  wire core_mi_reg_36__FF_INPUT;
  wire core_mi_reg_37_;
  wire core_mi_reg_37__FF_INPUT;
  wire core_mi_reg_38_;
  wire core_mi_reg_38__FF_INPUT;
  wire core_mi_reg_39_;
  wire core_mi_reg_39__FF_INPUT;
  wire core_mi_reg_3_;
  wire core_mi_reg_3__FF_INPUT;
  wire core_mi_reg_40_;
  wire core_mi_reg_40__FF_INPUT;
  wire core_mi_reg_41_;
  wire core_mi_reg_41__FF_INPUT;
  wire core_mi_reg_42_;
  wire core_mi_reg_42__FF_INPUT;
  wire core_mi_reg_43_;
  wire core_mi_reg_43__FF_INPUT;
  wire core_mi_reg_44_;
  wire core_mi_reg_44__FF_INPUT;
  wire core_mi_reg_45_;
  wire core_mi_reg_45__FF_INPUT;
  wire core_mi_reg_46_;
  wire core_mi_reg_46__FF_INPUT;
  wire core_mi_reg_47_;
  wire core_mi_reg_47__FF_INPUT;
  wire core_mi_reg_48_;
  wire core_mi_reg_48__FF_INPUT;
  wire core_mi_reg_49_;
  wire core_mi_reg_49__FF_INPUT;
  wire core_mi_reg_4_;
  wire core_mi_reg_4__FF_INPUT;
  wire core_mi_reg_50_;
  wire core_mi_reg_50__FF_INPUT;
  wire core_mi_reg_51_;
  wire core_mi_reg_51__FF_INPUT;
  wire core_mi_reg_52_;
  wire core_mi_reg_52__FF_INPUT;
  wire core_mi_reg_53_;
  wire core_mi_reg_53__FF_INPUT;
  wire core_mi_reg_54_;
  wire core_mi_reg_54__FF_INPUT;
  wire core_mi_reg_55_;
  wire core_mi_reg_55__FF_INPUT;
  wire core_mi_reg_56_;
  wire core_mi_reg_56__FF_INPUT;
  wire core_mi_reg_57_;
  wire core_mi_reg_57__FF_INPUT;
  wire core_mi_reg_58_;
  wire core_mi_reg_58__FF_INPUT;
  wire core_mi_reg_59_;
  wire core_mi_reg_59__FF_INPUT;
  wire core_mi_reg_5_;
  wire core_mi_reg_5__FF_INPUT;
  wire core_mi_reg_60_;
  wire core_mi_reg_60__FF_INPUT;
  wire core_mi_reg_61_;
  wire core_mi_reg_61__FF_INPUT;
  wire core_mi_reg_62_;
  wire core_mi_reg_62__FF_INPUT;
  wire core_mi_reg_63_;
  wire core_mi_reg_63__FF_INPUT;
  wire core_mi_reg_6_;
  wire core_mi_reg_6__FF_INPUT;
  wire core_mi_reg_7_;
  wire core_mi_reg_7__FF_INPUT;
  wire core_mi_reg_8_;
  wire core_mi_reg_8__FF_INPUT;
  wire core_mi_reg_9_;
  wire core_mi_reg_9__FF_INPUT;
  wire core_ready;
  wire core_ready_reg_FF_INPUT;
  wire core_siphash_ctrl_reg_0_;
  wire core_siphash_ctrl_reg_1_;
  wire core_siphash_ctrl_reg_2_;
  wire core_siphash_ctrl_reg_3_;
  wire core_siphash_ctrl_reg_4_;
  wire core_siphash_ctrl_reg_5_;
  wire core_siphash_ctrl_reg_6_;
  wire core_siphash_valid_reg;
  wire core_siphash_valid_reg_FF_INPUT;
  wire core_siphash_valid_reg_bF_buf0;
  wire core_siphash_valid_reg_bF_buf1;
  wire core_siphash_valid_reg_bF_buf10;
  wire core_siphash_valid_reg_bF_buf2;
  wire core_siphash_valid_reg_bF_buf3;
  wire core_siphash_valid_reg_bF_buf4;
  wire core_siphash_valid_reg_bF_buf5;
  wire core_siphash_valid_reg_bF_buf6;
  wire core_siphash_valid_reg_bF_buf7;
  wire core_siphash_valid_reg_bF_buf8;
  wire core_siphash_valid_reg_bF_buf9;
  wire core_siphash_word0_reg_0__FF_INPUT;
  wire core_siphash_word0_reg_10__FF_INPUT;
  wire core_siphash_word0_reg_11__FF_INPUT;
  wire core_siphash_word0_reg_12__FF_INPUT;
  wire core_siphash_word0_reg_13__FF_INPUT;
  wire core_siphash_word0_reg_14__FF_INPUT;
  wire core_siphash_word0_reg_15__FF_INPUT;
  wire core_siphash_word0_reg_16__FF_INPUT;
  wire core_siphash_word0_reg_17__FF_INPUT;
  wire core_siphash_word0_reg_18__FF_INPUT;
  wire core_siphash_word0_reg_19__FF_INPUT;
  wire core_siphash_word0_reg_1__FF_INPUT;
  wire core_siphash_word0_reg_20__FF_INPUT;
  wire core_siphash_word0_reg_21__FF_INPUT;
  wire core_siphash_word0_reg_22__FF_INPUT;
  wire core_siphash_word0_reg_23__FF_INPUT;
  wire core_siphash_word0_reg_24__FF_INPUT;
  wire core_siphash_word0_reg_25__FF_INPUT;
  wire core_siphash_word0_reg_26__FF_INPUT;
  wire core_siphash_word0_reg_27__FF_INPUT;
  wire core_siphash_word0_reg_28__FF_INPUT;
  wire core_siphash_word0_reg_29__FF_INPUT;
  wire core_siphash_word0_reg_2__FF_INPUT;
  wire core_siphash_word0_reg_30__FF_INPUT;
  wire core_siphash_word0_reg_31__FF_INPUT;
  wire core_siphash_word0_reg_32__FF_INPUT;
  wire core_siphash_word0_reg_33__FF_INPUT;
  wire core_siphash_word0_reg_34__FF_INPUT;
  wire core_siphash_word0_reg_35__FF_INPUT;
  wire core_siphash_word0_reg_36__FF_INPUT;
  wire core_siphash_word0_reg_37__FF_INPUT;
  wire core_siphash_word0_reg_38__FF_INPUT;
  wire core_siphash_word0_reg_39__FF_INPUT;
  wire core_siphash_word0_reg_3__FF_INPUT;
  wire core_siphash_word0_reg_40__FF_INPUT;
  wire core_siphash_word0_reg_41__FF_INPUT;
  wire core_siphash_word0_reg_42__FF_INPUT;
  wire core_siphash_word0_reg_43__FF_INPUT;
  wire core_siphash_word0_reg_44__FF_INPUT;
  wire core_siphash_word0_reg_45__FF_INPUT;
  wire core_siphash_word0_reg_46__FF_INPUT;
  wire core_siphash_word0_reg_47__FF_INPUT;
  wire core_siphash_word0_reg_48__FF_INPUT;
  wire core_siphash_word0_reg_49__FF_INPUT;
  wire core_siphash_word0_reg_4__FF_INPUT;
  wire core_siphash_word0_reg_50__FF_INPUT;
  wire core_siphash_word0_reg_51__FF_INPUT;
  wire core_siphash_word0_reg_52__FF_INPUT;
  wire core_siphash_word0_reg_53__FF_INPUT;
  wire core_siphash_word0_reg_54__FF_INPUT;
  wire core_siphash_word0_reg_55__FF_INPUT;
  wire core_siphash_word0_reg_56__FF_INPUT;
  wire core_siphash_word0_reg_57__FF_INPUT;
  wire core_siphash_word0_reg_58__FF_INPUT;
  wire core_siphash_word0_reg_59__FF_INPUT;
  wire core_siphash_word0_reg_5__FF_INPUT;
  wire core_siphash_word0_reg_60__FF_INPUT;
  wire core_siphash_word0_reg_61__FF_INPUT;
  wire core_siphash_word0_reg_62__FF_INPUT;
  wire core_siphash_word0_reg_63__FF_INPUT;
  wire core_siphash_word0_reg_6__FF_INPUT;
  wire core_siphash_word0_reg_7__FF_INPUT;
  wire core_siphash_word0_reg_8__FF_INPUT;
  wire core_siphash_word0_reg_9__FF_INPUT;
  wire core_siphash_word1_reg_0__FF_INPUT;
  wire core_siphash_word1_reg_10__FF_INPUT;
  wire core_siphash_word1_reg_11__FF_INPUT;
  wire core_siphash_word1_reg_12__FF_INPUT;
  wire core_siphash_word1_reg_13__FF_INPUT;
  wire core_siphash_word1_reg_14__FF_INPUT;
  wire core_siphash_word1_reg_15__FF_INPUT;
  wire core_siphash_word1_reg_16__FF_INPUT;
  wire core_siphash_word1_reg_17__FF_INPUT;
  wire core_siphash_word1_reg_18__FF_INPUT;
  wire core_siphash_word1_reg_19__FF_INPUT;
  wire core_siphash_word1_reg_1__FF_INPUT;
  wire core_siphash_word1_reg_20__FF_INPUT;
  wire core_siphash_word1_reg_21__FF_INPUT;
  wire core_siphash_word1_reg_22__FF_INPUT;
  wire core_siphash_word1_reg_23__FF_INPUT;
  wire core_siphash_word1_reg_24__FF_INPUT;
  wire core_siphash_word1_reg_25__FF_INPUT;
  wire core_siphash_word1_reg_26__FF_INPUT;
  wire core_siphash_word1_reg_27__FF_INPUT;
  wire core_siphash_word1_reg_28__FF_INPUT;
  wire core_siphash_word1_reg_29__FF_INPUT;
  wire core_siphash_word1_reg_2__FF_INPUT;
  wire core_siphash_word1_reg_30__FF_INPUT;
  wire core_siphash_word1_reg_31__FF_INPUT;
  wire core_siphash_word1_reg_32__FF_INPUT;
  wire core_siphash_word1_reg_33__FF_INPUT;
  wire core_siphash_word1_reg_34__FF_INPUT;
  wire core_siphash_word1_reg_35__FF_INPUT;
  wire core_siphash_word1_reg_36__FF_INPUT;
  wire core_siphash_word1_reg_37__FF_INPUT;
  wire core_siphash_word1_reg_38__FF_INPUT;
  wire core_siphash_word1_reg_39__FF_INPUT;
  wire core_siphash_word1_reg_3__FF_INPUT;
  wire core_siphash_word1_reg_40__FF_INPUT;
  wire core_siphash_word1_reg_41__FF_INPUT;
  wire core_siphash_word1_reg_42__FF_INPUT;
  wire core_siphash_word1_reg_43__FF_INPUT;
  wire core_siphash_word1_reg_44__FF_INPUT;
  wire core_siphash_word1_reg_45__FF_INPUT;
  wire core_siphash_word1_reg_46__FF_INPUT;
  wire core_siphash_word1_reg_47__FF_INPUT;
  wire core_siphash_word1_reg_48__FF_INPUT;
  wire core_siphash_word1_reg_49__FF_INPUT;
  wire core_siphash_word1_reg_4__FF_INPUT;
  wire core_siphash_word1_reg_50__FF_INPUT;
  wire core_siphash_word1_reg_51__FF_INPUT;
  wire core_siphash_word1_reg_52__FF_INPUT;
  wire core_siphash_word1_reg_53__FF_INPUT;
  wire core_siphash_word1_reg_54__FF_INPUT;
  wire core_siphash_word1_reg_55__FF_INPUT;
  wire core_siphash_word1_reg_56__FF_INPUT;
  wire core_siphash_word1_reg_57__FF_INPUT;
  wire core_siphash_word1_reg_58__FF_INPUT;
  wire core_siphash_word1_reg_59__FF_INPUT;
  wire core_siphash_word1_reg_5__FF_INPUT;
  wire core_siphash_word1_reg_60__FF_INPUT;
  wire core_siphash_word1_reg_61__FF_INPUT;
  wire core_siphash_word1_reg_62__FF_INPUT;
  wire core_siphash_word1_reg_63__FF_INPUT;
  wire core_siphash_word1_reg_6__FF_INPUT;
  wire core_siphash_word1_reg_7__FF_INPUT;
  wire core_siphash_word1_reg_8__FF_INPUT;
  wire core_siphash_word1_reg_9__FF_INPUT;
  wire core_siphash_word1_we;
  wire core_siphash_word1_we_bF_buf0;
  wire core_siphash_word1_we_bF_buf1;
  wire core_siphash_word1_we_bF_buf2;
  wire core_siphash_word1_we_bF_buf3;
  wire core_siphash_word1_we_bF_buf4;
  wire core_siphash_word1_we_bF_buf5;
  wire core_siphash_word1_we_bF_buf6;
  wire core_siphash_word1_we_bF_buf7;
  wire core_siphash_word_0_;
  wire core_siphash_word_100_;
  wire core_siphash_word_101_;
  wire core_siphash_word_102_;
  wire core_siphash_word_103_;
  wire core_siphash_word_104_;
  wire core_siphash_word_105_;
  wire core_siphash_word_106_;
  wire core_siphash_word_107_;
  wire core_siphash_word_108_;
  wire core_siphash_word_109_;
  wire core_siphash_word_10_;
  wire core_siphash_word_110_;
  wire core_siphash_word_111_;
  wire core_siphash_word_112_;
  wire core_siphash_word_113_;
  wire core_siphash_word_114_;
  wire core_siphash_word_115_;
  wire core_siphash_word_116_;
  wire core_siphash_word_117_;
  wire core_siphash_word_118_;
  wire core_siphash_word_119_;
  wire core_siphash_word_11_;
  wire core_siphash_word_120_;
  wire core_siphash_word_121_;
  wire core_siphash_word_122_;
  wire core_siphash_word_123_;
  wire core_siphash_word_124_;
  wire core_siphash_word_125_;
  wire core_siphash_word_126_;
  wire core_siphash_word_127_;
  wire core_siphash_word_12_;
  wire core_siphash_word_13_;
  wire core_siphash_word_14_;
  wire core_siphash_word_15_;
  wire core_siphash_word_16_;
  wire core_siphash_word_17_;
  wire core_siphash_word_18_;
  wire core_siphash_word_19_;
  wire core_siphash_word_1_;
  wire core_siphash_word_20_;
  wire core_siphash_word_21_;
  wire core_siphash_word_22_;
  wire core_siphash_word_23_;
  wire core_siphash_word_24_;
  wire core_siphash_word_25_;
  wire core_siphash_word_26_;
  wire core_siphash_word_27_;
  wire core_siphash_word_28_;
  wire core_siphash_word_29_;
  wire core_siphash_word_2_;
  wire core_siphash_word_30_;
  wire core_siphash_word_31_;
  wire core_siphash_word_32_;
  wire core_siphash_word_33_;
  wire core_siphash_word_34_;
  wire core_siphash_word_35_;
  wire core_siphash_word_36_;
  wire core_siphash_word_37_;
  wire core_siphash_word_38_;
  wire core_siphash_word_39_;
  wire core_siphash_word_3_;
  wire core_siphash_word_40_;
  wire core_siphash_word_41_;
  wire core_siphash_word_42_;
  wire core_siphash_word_43_;
  wire core_siphash_word_44_;
  wire core_siphash_word_45_;
  wire core_siphash_word_46_;
  wire core_siphash_word_47_;
  wire core_siphash_word_48_;
  wire core_siphash_word_49_;
  wire core_siphash_word_4_;
  wire core_siphash_word_50_;
  wire core_siphash_word_51_;
  wire core_siphash_word_52_;
  wire core_siphash_word_53_;
  wire core_siphash_word_54_;
  wire core_siphash_word_55_;
  wire core_siphash_word_56_;
  wire core_siphash_word_57_;
  wire core_siphash_word_58_;
  wire core_siphash_word_59_;
  wire core_siphash_word_5_;
  wire core_siphash_word_60_;
  wire core_siphash_word_61_;
  wire core_siphash_word_62_;
  wire core_siphash_word_63_;
  wire core_siphash_word_64_;
  wire core_siphash_word_65_;
  wire core_siphash_word_66_;
  wire core_siphash_word_67_;
  wire core_siphash_word_68_;
  wire core_siphash_word_69_;
  wire core_siphash_word_6_;
  wire core_siphash_word_70_;
  wire core_siphash_word_71_;
  wire core_siphash_word_72_;
  wire core_siphash_word_73_;
  wire core_siphash_word_74_;
  wire core_siphash_word_75_;
  wire core_siphash_word_76_;
  wire core_siphash_word_77_;
  wire core_siphash_word_78_;
  wire core_siphash_word_79_;
  wire core_siphash_word_7_;
  wire core_siphash_word_80_;
  wire core_siphash_word_81_;
  wire core_siphash_word_82_;
  wire core_siphash_word_83_;
  wire core_siphash_word_84_;
  wire core_siphash_word_85_;
  wire core_siphash_word_86_;
  wire core_siphash_word_87_;
  wire core_siphash_word_88_;
  wire core_siphash_word_89_;
  wire core_siphash_word_8_;
  wire core_siphash_word_90_;
  wire core_siphash_word_91_;
  wire core_siphash_word_92_;
  wire core_siphash_word_93_;
  wire core_siphash_word_94_;
  wire core_siphash_word_95_;
  wire core_siphash_word_96_;
  wire core_siphash_word_97_;
  wire core_siphash_word_98_;
  wire core_siphash_word_99_;
  wire core_siphash_word_9_;
  wire core_v0_reg_0_;
  wire core_v0_reg_0__FF_INPUT;
  wire core_v0_reg_10_;
  wire core_v0_reg_10__FF_INPUT;
  wire core_v0_reg_11_;
  wire core_v0_reg_11__FF_INPUT;
  wire core_v0_reg_12_;
  wire core_v0_reg_12__FF_INPUT;
  wire core_v0_reg_13_;
  wire core_v0_reg_13__FF_INPUT;
  wire core_v0_reg_14_;
  wire core_v0_reg_14__FF_INPUT;
  wire core_v0_reg_15_;
  wire core_v0_reg_15__FF_INPUT;
  wire core_v0_reg_16_;
  wire core_v0_reg_16__FF_INPUT;
  wire core_v0_reg_17_;
  wire core_v0_reg_17__FF_INPUT;
  wire core_v0_reg_18_;
  wire core_v0_reg_18__FF_INPUT;
  wire core_v0_reg_19_;
  wire core_v0_reg_19__FF_INPUT;
  wire core_v0_reg_1_;
  wire core_v0_reg_1__FF_INPUT;
  wire core_v0_reg_20_;
  wire core_v0_reg_20__FF_INPUT;
  wire core_v0_reg_21_;
  wire core_v0_reg_21__FF_INPUT;
  wire core_v0_reg_22_;
  wire core_v0_reg_22__FF_INPUT;
  wire core_v0_reg_23_;
  wire core_v0_reg_23__FF_INPUT;
  wire core_v0_reg_24_;
  wire core_v0_reg_24__FF_INPUT;
  wire core_v0_reg_25_;
  wire core_v0_reg_25__FF_INPUT;
  wire core_v0_reg_26_;
  wire core_v0_reg_26__FF_INPUT;
  wire core_v0_reg_27_;
  wire core_v0_reg_27__FF_INPUT;
  wire core_v0_reg_28_;
  wire core_v0_reg_28__FF_INPUT;
  wire core_v0_reg_29_;
  wire core_v0_reg_29__FF_INPUT;
  wire core_v0_reg_2_;
  wire core_v0_reg_2__FF_INPUT;
  wire core_v0_reg_30_;
  wire core_v0_reg_30__FF_INPUT;
  wire core_v0_reg_31_;
  wire core_v0_reg_31__FF_INPUT;
  wire core_v0_reg_32_;
  wire core_v0_reg_32__FF_INPUT;
  wire core_v0_reg_33_;
  wire core_v0_reg_33__FF_INPUT;
  wire core_v0_reg_34_;
  wire core_v0_reg_34__FF_INPUT;
  wire core_v0_reg_35_;
  wire core_v0_reg_35__FF_INPUT;
  wire core_v0_reg_36_;
  wire core_v0_reg_36__FF_INPUT;
  wire core_v0_reg_37_;
  wire core_v0_reg_37__FF_INPUT;
  wire core_v0_reg_38_;
  wire core_v0_reg_38__FF_INPUT;
  wire core_v0_reg_39_;
  wire core_v0_reg_39__FF_INPUT;
  wire core_v0_reg_3_;
  wire core_v0_reg_3__FF_INPUT;
  wire core_v0_reg_40_;
  wire core_v0_reg_40__FF_INPUT;
  wire core_v0_reg_41_;
  wire core_v0_reg_41__FF_INPUT;
  wire core_v0_reg_42_;
  wire core_v0_reg_42__FF_INPUT;
  wire core_v0_reg_43_;
  wire core_v0_reg_43__FF_INPUT;
  wire core_v0_reg_44_;
  wire core_v0_reg_44__FF_INPUT;
  wire core_v0_reg_45_;
  wire core_v0_reg_45__FF_INPUT;
  wire core_v0_reg_46_;
  wire core_v0_reg_46__FF_INPUT;
  wire core_v0_reg_47_;
  wire core_v0_reg_47__FF_INPUT;
  wire core_v0_reg_48_;
  wire core_v0_reg_48__FF_INPUT;
  wire core_v0_reg_49_;
  wire core_v0_reg_49__FF_INPUT;
  wire core_v0_reg_4_;
  wire core_v0_reg_4__FF_INPUT;
  wire core_v0_reg_50_;
  wire core_v0_reg_50__FF_INPUT;
  wire core_v0_reg_51_;
  wire core_v0_reg_51__FF_INPUT;
  wire core_v0_reg_52_;
  wire core_v0_reg_52__FF_INPUT;
  wire core_v0_reg_53_;
  wire core_v0_reg_53__FF_INPUT;
  wire core_v0_reg_54_;
  wire core_v0_reg_54__FF_INPUT;
  wire core_v0_reg_55_;
  wire core_v0_reg_55__FF_INPUT;
  wire core_v0_reg_56_;
  wire core_v0_reg_56__FF_INPUT;
  wire core_v0_reg_57_;
  wire core_v0_reg_57__FF_INPUT;
  wire core_v0_reg_58_;
  wire core_v0_reg_58__FF_INPUT;
  wire core_v0_reg_59_;
  wire core_v0_reg_59__FF_INPUT;
  wire core_v0_reg_5_;
  wire core_v0_reg_5__FF_INPUT;
  wire core_v0_reg_60_;
  wire core_v0_reg_60__FF_INPUT;
  wire core_v0_reg_61_;
  wire core_v0_reg_61__FF_INPUT;
  wire core_v0_reg_62_;
  wire core_v0_reg_62__FF_INPUT;
  wire core_v0_reg_63_;
  wire core_v0_reg_63__FF_INPUT;
  wire core_v0_reg_6_;
  wire core_v0_reg_6__FF_INPUT;
  wire core_v0_reg_7_;
  wire core_v0_reg_7__FF_INPUT;
  wire core_v0_reg_8_;
  wire core_v0_reg_8__FF_INPUT;
  wire core_v0_reg_9_;
  wire core_v0_reg_9__FF_INPUT;
  wire core_v1_reg_0_;
  wire core_v1_reg_0__FF_INPUT;
  wire core_v1_reg_10_;
  wire core_v1_reg_10__FF_INPUT;
  wire core_v1_reg_11_;
  wire core_v1_reg_11__FF_INPUT;
  wire core_v1_reg_12_;
  wire core_v1_reg_12__FF_INPUT;
  wire core_v1_reg_13_;
  wire core_v1_reg_13__FF_INPUT;
  wire core_v1_reg_14_;
  wire core_v1_reg_14__FF_INPUT;
  wire core_v1_reg_15_;
  wire core_v1_reg_15__FF_INPUT;
  wire core_v1_reg_16_;
  wire core_v1_reg_16__FF_INPUT;
  wire core_v1_reg_17_;
  wire core_v1_reg_17__FF_INPUT;
  wire core_v1_reg_18_;
  wire core_v1_reg_18__FF_INPUT;
  wire core_v1_reg_19_;
  wire core_v1_reg_19__FF_INPUT;
  wire core_v1_reg_1_;
  wire core_v1_reg_1__FF_INPUT;
  wire core_v1_reg_20_;
  wire core_v1_reg_20__FF_INPUT;
  wire core_v1_reg_21_;
  wire core_v1_reg_21__FF_INPUT;
  wire core_v1_reg_22_;
  wire core_v1_reg_22__FF_INPUT;
  wire core_v1_reg_23_;
  wire core_v1_reg_23__FF_INPUT;
  wire core_v1_reg_24_;
  wire core_v1_reg_24__FF_INPUT;
  wire core_v1_reg_25_;
  wire core_v1_reg_25__FF_INPUT;
  wire core_v1_reg_26_;
  wire core_v1_reg_26__FF_INPUT;
  wire core_v1_reg_27_;
  wire core_v1_reg_27__FF_INPUT;
  wire core_v1_reg_28_;
  wire core_v1_reg_28__FF_INPUT;
  wire core_v1_reg_29_;
  wire core_v1_reg_29__FF_INPUT;
  wire core_v1_reg_2_;
  wire core_v1_reg_2__FF_INPUT;
  wire core_v1_reg_30_;
  wire core_v1_reg_30__FF_INPUT;
  wire core_v1_reg_31_;
  wire core_v1_reg_31__FF_INPUT;
  wire core_v1_reg_32_;
  wire core_v1_reg_32__FF_INPUT;
  wire core_v1_reg_33_;
  wire core_v1_reg_33__FF_INPUT;
  wire core_v1_reg_34_;
  wire core_v1_reg_34__FF_INPUT;
  wire core_v1_reg_35_;
  wire core_v1_reg_35__FF_INPUT;
  wire core_v1_reg_36_;
  wire core_v1_reg_36__FF_INPUT;
  wire core_v1_reg_37_;
  wire core_v1_reg_37__FF_INPUT;
  wire core_v1_reg_38_;
  wire core_v1_reg_38__FF_INPUT;
  wire core_v1_reg_39_;
  wire core_v1_reg_39__FF_INPUT;
  wire core_v1_reg_3_;
  wire core_v1_reg_3__FF_INPUT;
  wire core_v1_reg_40_;
  wire core_v1_reg_40__FF_INPUT;
  wire core_v1_reg_41_;
  wire core_v1_reg_41__FF_INPUT;
  wire core_v1_reg_42_;
  wire core_v1_reg_42__FF_INPUT;
  wire core_v1_reg_43_;
  wire core_v1_reg_43__FF_INPUT;
  wire core_v1_reg_44_;
  wire core_v1_reg_44__FF_INPUT;
  wire core_v1_reg_45_;
  wire core_v1_reg_45__FF_INPUT;
  wire core_v1_reg_46_;
  wire core_v1_reg_46__FF_INPUT;
  wire core_v1_reg_47_;
  wire core_v1_reg_47__FF_INPUT;
  wire core_v1_reg_48_;
  wire core_v1_reg_48__FF_INPUT;
  wire core_v1_reg_49_;
  wire core_v1_reg_49__FF_INPUT;
  wire core_v1_reg_4_;
  wire core_v1_reg_4__FF_INPUT;
  wire core_v1_reg_50_;
  wire core_v1_reg_50__FF_INPUT;
  wire core_v1_reg_51_;
  wire core_v1_reg_51__FF_INPUT;
  wire core_v1_reg_52_;
  wire core_v1_reg_52__FF_INPUT;
  wire core_v1_reg_53_;
  wire core_v1_reg_53__FF_INPUT;
  wire core_v1_reg_54_;
  wire core_v1_reg_54__FF_INPUT;
  wire core_v1_reg_55_;
  wire core_v1_reg_55__FF_INPUT;
  wire core_v1_reg_56_;
  wire core_v1_reg_56__FF_INPUT;
  wire core_v1_reg_57_;
  wire core_v1_reg_57__FF_INPUT;
  wire core_v1_reg_58_;
  wire core_v1_reg_58__FF_INPUT;
  wire core_v1_reg_59_;
  wire core_v1_reg_59__FF_INPUT;
  wire core_v1_reg_5_;
  wire core_v1_reg_5__FF_INPUT;
  wire core_v1_reg_60_;
  wire core_v1_reg_60__FF_INPUT;
  wire core_v1_reg_61_;
  wire core_v1_reg_61__FF_INPUT;
  wire core_v1_reg_62_;
  wire core_v1_reg_62__FF_INPUT;
  wire core_v1_reg_63_;
  wire core_v1_reg_63__FF_INPUT;
  wire core_v1_reg_6_;
  wire core_v1_reg_6__FF_INPUT;
  wire core_v1_reg_7_;
  wire core_v1_reg_7__FF_INPUT;
  wire core_v1_reg_8_;
  wire core_v1_reg_8__FF_INPUT;
  wire core_v1_reg_9_;
  wire core_v1_reg_9__FF_INPUT;
  wire core_v2_reg_0_;
  wire core_v2_reg_0__FF_INPUT;
  wire core_v2_reg_10_;
  wire core_v2_reg_10__FF_INPUT;
  wire core_v2_reg_11_;
  wire core_v2_reg_11__FF_INPUT;
  wire core_v2_reg_12_;
  wire core_v2_reg_12__FF_INPUT;
  wire core_v2_reg_13_;
  wire core_v2_reg_13__FF_INPUT;
  wire core_v2_reg_14_;
  wire core_v2_reg_14__FF_INPUT;
  wire core_v2_reg_15_;
  wire core_v2_reg_15__FF_INPUT;
  wire core_v2_reg_16_;
  wire core_v2_reg_16__FF_INPUT;
  wire core_v2_reg_17_;
  wire core_v2_reg_17__FF_INPUT;
  wire core_v2_reg_18_;
  wire core_v2_reg_18__FF_INPUT;
  wire core_v2_reg_19_;
  wire core_v2_reg_19__FF_INPUT;
  wire core_v2_reg_1_;
  wire core_v2_reg_1__FF_INPUT;
  wire core_v2_reg_20_;
  wire core_v2_reg_20__FF_INPUT;
  wire core_v2_reg_21_;
  wire core_v2_reg_21__FF_INPUT;
  wire core_v2_reg_22_;
  wire core_v2_reg_22__FF_INPUT;
  wire core_v2_reg_23_;
  wire core_v2_reg_23__FF_INPUT;
  wire core_v2_reg_24_;
  wire core_v2_reg_24__FF_INPUT;
  wire core_v2_reg_25_;
  wire core_v2_reg_25__FF_INPUT;
  wire core_v2_reg_26_;
  wire core_v2_reg_26__FF_INPUT;
  wire core_v2_reg_27_;
  wire core_v2_reg_27__FF_INPUT;
  wire core_v2_reg_28_;
  wire core_v2_reg_28__FF_INPUT;
  wire core_v2_reg_29_;
  wire core_v2_reg_29__FF_INPUT;
  wire core_v2_reg_2_;
  wire core_v2_reg_2__FF_INPUT;
  wire core_v2_reg_30_;
  wire core_v2_reg_30__FF_INPUT;
  wire core_v2_reg_31_;
  wire core_v2_reg_31__FF_INPUT;
  wire core_v2_reg_32_;
  wire core_v2_reg_32__FF_INPUT;
  wire core_v2_reg_33_;
  wire core_v2_reg_33__FF_INPUT;
  wire core_v2_reg_34_;
  wire core_v2_reg_34__FF_INPUT;
  wire core_v2_reg_35_;
  wire core_v2_reg_35__FF_INPUT;
  wire core_v2_reg_36_;
  wire core_v2_reg_36__FF_INPUT;
  wire core_v2_reg_37_;
  wire core_v2_reg_37__FF_INPUT;
  wire core_v2_reg_38_;
  wire core_v2_reg_38__FF_INPUT;
  wire core_v2_reg_39_;
  wire core_v2_reg_39__FF_INPUT;
  wire core_v2_reg_3_;
  wire core_v2_reg_3__FF_INPUT;
  wire core_v2_reg_40_;
  wire core_v2_reg_40__FF_INPUT;
  wire core_v2_reg_41_;
  wire core_v2_reg_41__FF_INPUT;
  wire core_v2_reg_42_;
  wire core_v2_reg_42__FF_INPUT;
  wire core_v2_reg_43_;
  wire core_v2_reg_43__FF_INPUT;
  wire core_v2_reg_44_;
  wire core_v2_reg_44__FF_INPUT;
  wire core_v2_reg_45_;
  wire core_v2_reg_45__FF_INPUT;
  wire core_v2_reg_46_;
  wire core_v2_reg_46__FF_INPUT;
  wire core_v2_reg_47_;
  wire core_v2_reg_47__FF_INPUT;
  wire core_v2_reg_48_;
  wire core_v2_reg_48__FF_INPUT;
  wire core_v2_reg_49_;
  wire core_v2_reg_49__FF_INPUT;
  wire core_v2_reg_4_;
  wire core_v2_reg_4__FF_INPUT;
  wire core_v2_reg_50_;
  wire core_v2_reg_50__FF_INPUT;
  wire core_v2_reg_51_;
  wire core_v2_reg_51__FF_INPUT;
  wire core_v2_reg_52_;
  wire core_v2_reg_52__FF_INPUT;
  wire core_v2_reg_53_;
  wire core_v2_reg_53__FF_INPUT;
  wire core_v2_reg_54_;
  wire core_v2_reg_54__FF_INPUT;
  wire core_v2_reg_55_;
  wire core_v2_reg_55__FF_INPUT;
  wire core_v2_reg_56_;
  wire core_v2_reg_56__FF_INPUT;
  wire core_v2_reg_57_;
  wire core_v2_reg_57__FF_INPUT;
  wire core_v2_reg_58_;
  wire core_v2_reg_58__FF_INPUT;
  wire core_v2_reg_59_;
  wire core_v2_reg_59__FF_INPUT;
  wire core_v2_reg_5_;
  wire core_v2_reg_5__FF_INPUT;
  wire core_v2_reg_60_;
  wire core_v2_reg_60__FF_INPUT;
  wire core_v2_reg_61_;
  wire core_v2_reg_61__FF_INPUT;
  wire core_v2_reg_62_;
  wire core_v2_reg_62__FF_INPUT;
  wire core_v2_reg_63_;
  wire core_v2_reg_63__FF_INPUT;
  wire core_v2_reg_6_;
  wire core_v2_reg_6__FF_INPUT;
  wire core_v2_reg_7_;
  wire core_v2_reg_7__FF_INPUT;
  wire core_v2_reg_8_;
  wire core_v2_reg_8__FF_INPUT;
  wire core_v2_reg_9_;
  wire core_v2_reg_9__FF_INPUT;
  wire core_v3_reg_0_;
  wire core_v3_reg_0__FF_INPUT;
  wire core_v3_reg_10_;
  wire core_v3_reg_10__FF_INPUT;
  wire core_v3_reg_11_;
  wire core_v3_reg_11__FF_INPUT;
  wire core_v3_reg_12_;
  wire core_v3_reg_12__FF_INPUT;
  wire core_v3_reg_13_;
  wire core_v3_reg_13__FF_INPUT;
  wire core_v3_reg_14_;
  wire core_v3_reg_14__FF_INPUT;
  wire core_v3_reg_15_;
  wire core_v3_reg_15__FF_INPUT;
  wire core_v3_reg_16_;
  wire core_v3_reg_16__FF_INPUT;
  wire core_v3_reg_17_;
  wire core_v3_reg_17__FF_INPUT;
  wire core_v3_reg_18_;
  wire core_v3_reg_18__FF_INPUT;
  wire core_v3_reg_19_;
  wire core_v3_reg_19__FF_INPUT;
  wire core_v3_reg_1_;
  wire core_v3_reg_1__FF_INPUT;
  wire core_v3_reg_20_;
  wire core_v3_reg_20__FF_INPUT;
  wire core_v3_reg_21_;
  wire core_v3_reg_21__FF_INPUT;
  wire core_v3_reg_22_;
  wire core_v3_reg_22__FF_INPUT;
  wire core_v3_reg_23_;
  wire core_v3_reg_23__FF_INPUT;
  wire core_v3_reg_24_;
  wire core_v3_reg_24__FF_INPUT;
  wire core_v3_reg_25_;
  wire core_v3_reg_25__FF_INPUT;
  wire core_v3_reg_26_;
  wire core_v3_reg_26__FF_INPUT;
  wire core_v3_reg_27_;
  wire core_v3_reg_27__FF_INPUT;
  wire core_v3_reg_28_;
  wire core_v3_reg_28__FF_INPUT;
  wire core_v3_reg_29_;
  wire core_v3_reg_29__FF_INPUT;
  wire core_v3_reg_2_;
  wire core_v3_reg_2__FF_INPUT;
  wire core_v3_reg_30_;
  wire core_v3_reg_30__FF_INPUT;
  wire core_v3_reg_31_;
  wire core_v3_reg_31__FF_INPUT;
  wire core_v3_reg_32_;
  wire core_v3_reg_32__FF_INPUT;
  wire core_v3_reg_33_;
  wire core_v3_reg_33__FF_INPUT;
  wire core_v3_reg_34_;
  wire core_v3_reg_34__FF_INPUT;
  wire core_v3_reg_35_;
  wire core_v3_reg_35__FF_INPUT;
  wire core_v3_reg_36_;
  wire core_v3_reg_36__FF_INPUT;
  wire core_v3_reg_37_;
  wire core_v3_reg_37__FF_INPUT;
  wire core_v3_reg_38_;
  wire core_v3_reg_38__FF_INPUT;
  wire core_v3_reg_39_;
  wire core_v3_reg_39__FF_INPUT;
  wire core_v3_reg_3_;
  wire core_v3_reg_3__FF_INPUT;
  wire core_v3_reg_40_;
  wire core_v3_reg_40__FF_INPUT;
  wire core_v3_reg_41_;
  wire core_v3_reg_41__FF_INPUT;
  wire core_v3_reg_42_;
  wire core_v3_reg_42__FF_INPUT;
  wire core_v3_reg_43_;
  wire core_v3_reg_43__FF_INPUT;
  wire core_v3_reg_44_;
  wire core_v3_reg_44__FF_INPUT;
  wire core_v3_reg_45_;
  wire core_v3_reg_45__FF_INPUT;
  wire core_v3_reg_46_;
  wire core_v3_reg_46__FF_INPUT;
  wire core_v3_reg_47_;
  wire core_v3_reg_47__FF_INPUT;
  wire core_v3_reg_48_;
  wire core_v3_reg_48__FF_INPUT;
  wire core_v3_reg_49_;
  wire core_v3_reg_49__FF_INPUT;
  wire core_v3_reg_4_;
  wire core_v3_reg_4__FF_INPUT;
  wire core_v3_reg_50_;
  wire core_v3_reg_50__FF_INPUT;
  wire core_v3_reg_51_;
  wire core_v3_reg_51__FF_INPUT;
  wire core_v3_reg_52_;
  wire core_v3_reg_52__FF_INPUT;
  wire core_v3_reg_53_;
  wire core_v3_reg_53__FF_INPUT;
  wire core_v3_reg_54_;
  wire core_v3_reg_54__FF_INPUT;
  wire core_v3_reg_55_;
  wire core_v3_reg_55__FF_INPUT;
  wire core_v3_reg_56_;
  wire core_v3_reg_56__FF_INPUT;
  wire core_v3_reg_57_;
  wire core_v3_reg_57__FF_INPUT;
  wire core_v3_reg_58_;
  wire core_v3_reg_58__FF_INPUT;
  wire core_v3_reg_59_;
  wire core_v3_reg_59__FF_INPUT;
  wire core_v3_reg_5_;
  wire core_v3_reg_5__FF_INPUT;
  wire core_v3_reg_60_;
  wire core_v3_reg_60__FF_INPUT;
  wire core_v3_reg_61_;
  wire core_v3_reg_61__FF_INPUT;
  wire core_v3_reg_62_;
  wire core_v3_reg_62__FF_INPUT;
  wire core_v3_reg_63_;
  wire core_v3_reg_63__FF_INPUT;
  wire core_v3_reg_6_;
  wire core_v3_reg_6__FF_INPUT;
  wire core_v3_reg_7_;
  wire core_v3_reg_7__FF_INPUT;
  wire core_v3_reg_8_;
  wire core_v3_reg_8__FF_INPUT;
  wire core_v3_reg_9_;
  wire core_v3_reg_9__FF_INPUT;
  input cs;
  wire ctrl_reg_0__FF_INPUT;
  wire ctrl_reg_1__FF_INPUT;
  wire ctrl_reg_2__FF_INPUT;
  wire key0_reg_0__FF_INPUT;
  wire key0_reg_10__FF_INPUT;
  wire key0_reg_11__FF_INPUT;
  wire key0_reg_12__FF_INPUT;
  wire key0_reg_13__FF_INPUT;
  wire key0_reg_14__FF_INPUT;
  wire key0_reg_15__FF_INPUT;
  wire key0_reg_16__FF_INPUT;
  wire key0_reg_17__FF_INPUT;
  wire key0_reg_18__FF_INPUT;
  wire key0_reg_19__FF_INPUT;
  wire key0_reg_1__FF_INPUT;
  wire key0_reg_20__FF_INPUT;
  wire key0_reg_21__FF_INPUT;
  wire key0_reg_22__FF_INPUT;
  wire key0_reg_23__FF_INPUT;
  wire key0_reg_24__FF_INPUT;
  wire key0_reg_25__FF_INPUT;
  wire key0_reg_26__FF_INPUT;
  wire key0_reg_27__FF_INPUT;
  wire key0_reg_28__FF_INPUT;
  wire key0_reg_29__FF_INPUT;
  wire key0_reg_2__FF_INPUT;
  wire key0_reg_30__FF_INPUT;
  wire key0_reg_31__FF_INPUT;
  wire key0_reg_3__FF_INPUT;
  wire key0_reg_4__FF_INPUT;
  wire key0_reg_5__FF_INPUT;
  wire key0_reg_6__FF_INPUT;
  wire key0_reg_7__FF_INPUT;
  wire key0_reg_8__FF_INPUT;
  wire key0_reg_9__FF_INPUT;
  wire key1_reg_0__FF_INPUT;
  wire key1_reg_10__FF_INPUT;
  wire key1_reg_11__FF_INPUT;
  wire key1_reg_12__FF_INPUT;
  wire key1_reg_13__FF_INPUT;
  wire key1_reg_14__FF_INPUT;
  wire key1_reg_15__FF_INPUT;
  wire key1_reg_16__FF_INPUT;
  wire key1_reg_17__FF_INPUT;
  wire key1_reg_18__FF_INPUT;
  wire key1_reg_19__FF_INPUT;
  wire key1_reg_1__FF_INPUT;
  wire key1_reg_20__FF_INPUT;
  wire key1_reg_21__FF_INPUT;
  wire key1_reg_22__FF_INPUT;
  wire key1_reg_23__FF_INPUT;
  wire key1_reg_24__FF_INPUT;
  wire key1_reg_25__FF_INPUT;
  wire key1_reg_26__FF_INPUT;
  wire key1_reg_27__FF_INPUT;
  wire key1_reg_28__FF_INPUT;
  wire key1_reg_29__FF_INPUT;
  wire key1_reg_2__FF_INPUT;
  wire key1_reg_30__FF_INPUT;
  wire key1_reg_31__FF_INPUT;
  wire key1_reg_3__FF_INPUT;
  wire key1_reg_4__FF_INPUT;
  wire key1_reg_5__FF_INPUT;
  wire key1_reg_6__FF_INPUT;
  wire key1_reg_7__FF_INPUT;
  wire key1_reg_8__FF_INPUT;
  wire key1_reg_9__FF_INPUT;
  wire key2_reg_0__FF_INPUT;
  wire key2_reg_10__FF_INPUT;
  wire key2_reg_11__FF_INPUT;
  wire key2_reg_12__FF_INPUT;
  wire key2_reg_13__FF_INPUT;
  wire key2_reg_14__FF_INPUT;
  wire key2_reg_15__FF_INPUT;
  wire key2_reg_16__FF_INPUT;
  wire key2_reg_17__FF_INPUT;
  wire key2_reg_18__FF_INPUT;
  wire key2_reg_19__FF_INPUT;
  wire key2_reg_1__FF_INPUT;
  wire key2_reg_20__FF_INPUT;
  wire key2_reg_21__FF_INPUT;
  wire key2_reg_22__FF_INPUT;
  wire key2_reg_23__FF_INPUT;
  wire key2_reg_24__FF_INPUT;
  wire key2_reg_25__FF_INPUT;
  wire key2_reg_26__FF_INPUT;
  wire key2_reg_27__FF_INPUT;
  wire key2_reg_28__FF_INPUT;
  wire key2_reg_29__FF_INPUT;
  wire key2_reg_2__FF_INPUT;
  wire key2_reg_30__FF_INPUT;
  wire key2_reg_31__FF_INPUT;
  wire key2_reg_3__FF_INPUT;
  wire key2_reg_4__FF_INPUT;
  wire key2_reg_5__FF_INPUT;
  wire key2_reg_6__FF_INPUT;
  wire key2_reg_7__FF_INPUT;
  wire key2_reg_8__FF_INPUT;
  wire key2_reg_9__FF_INPUT;
  wire key3_reg_0__FF_INPUT;
  wire key3_reg_10__FF_INPUT;
  wire key3_reg_11__FF_INPUT;
  wire key3_reg_12__FF_INPUT;
  wire key3_reg_13__FF_INPUT;
  wire key3_reg_14__FF_INPUT;
  wire key3_reg_15__FF_INPUT;
  wire key3_reg_16__FF_INPUT;
  wire key3_reg_17__FF_INPUT;
  wire key3_reg_18__FF_INPUT;
  wire key3_reg_19__FF_INPUT;
  wire key3_reg_1__FF_INPUT;
  wire key3_reg_20__FF_INPUT;
  wire key3_reg_21__FF_INPUT;
  wire key3_reg_22__FF_INPUT;
  wire key3_reg_23__FF_INPUT;
  wire key3_reg_24__FF_INPUT;
  wire key3_reg_25__FF_INPUT;
  wire key3_reg_26__FF_INPUT;
  wire key3_reg_27__FF_INPUT;
  wire key3_reg_28__FF_INPUT;
  wire key3_reg_29__FF_INPUT;
  wire key3_reg_2__FF_INPUT;
  wire key3_reg_30__FF_INPUT;
  wire key3_reg_31__FF_INPUT;
  wire key3_reg_3__FF_INPUT;
  wire key3_reg_4__FF_INPUT;
  wire key3_reg_5__FF_INPUT;
  wire key3_reg_6__FF_INPUT;
  wire key3_reg_7__FF_INPUT;
  wire key3_reg_8__FF_INPUT;
  wire key3_reg_9__FF_INPUT;
  wire long_reg_FF_INPUT;
  wire mi0_reg_0__FF_INPUT;
  wire mi0_reg_10__FF_INPUT;
  wire mi0_reg_11__FF_INPUT;
  wire mi0_reg_12__FF_INPUT;
  wire mi0_reg_13__FF_INPUT;
  wire mi0_reg_14__FF_INPUT;
  wire mi0_reg_15__FF_INPUT;
  wire mi0_reg_16__FF_INPUT;
  wire mi0_reg_17__FF_INPUT;
  wire mi0_reg_18__FF_INPUT;
  wire mi0_reg_19__FF_INPUT;
  wire mi0_reg_1__FF_INPUT;
  wire mi0_reg_20__FF_INPUT;
  wire mi0_reg_21__FF_INPUT;
  wire mi0_reg_22__FF_INPUT;
  wire mi0_reg_23__FF_INPUT;
  wire mi0_reg_24__FF_INPUT;
  wire mi0_reg_25__FF_INPUT;
  wire mi0_reg_26__FF_INPUT;
  wire mi0_reg_27__FF_INPUT;
  wire mi0_reg_28__FF_INPUT;
  wire mi0_reg_29__FF_INPUT;
  wire mi0_reg_2__FF_INPUT;
  wire mi0_reg_30__FF_INPUT;
  wire mi0_reg_31__FF_INPUT;
  wire mi0_reg_3__FF_INPUT;
  wire mi0_reg_4__FF_INPUT;
  wire mi0_reg_5__FF_INPUT;
  wire mi0_reg_6__FF_INPUT;
  wire mi0_reg_7__FF_INPUT;
  wire mi0_reg_8__FF_INPUT;
  wire mi0_reg_9__FF_INPUT;
  wire mi1_reg_0__FF_INPUT;
  wire mi1_reg_10__FF_INPUT;
  wire mi1_reg_11__FF_INPUT;
  wire mi1_reg_12__FF_INPUT;
  wire mi1_reg_13__FF_INPUT;
  wire mi1_reg_14__FF_INPUT;
  wire mi1_reg_15__FF_INPUT;
  wire mi1_reg_16__FF_INPUT;
  wire mi1_reg_17__FF_INPUT;
  wire mi1_reg_18__FF_INPUT;
  wire mi1_reg_19__FF_INPUT;
  wire mi1_reg_1__FF_INPUT;
  wire mi1_reg_20__FF_INPUT;
  wire mi1_reg_21__FF_INPUT;
  wire mi1_reg_22__FF_INPUT;
  wire mi1_reg_23__FF_INPUT;
  wire mi1_reg_24__FF_INPUT;
  wire mi1_reg_25__FF_INPUT;
  wire mi1_reg_26__FF_INPUT;
  wire mi1_reg_27__FF_INPUT;
  wire mi1_reg_28__FF_INPUT;
  wire mi1_reg_29__FF_INPUT;
  wire mi1_reg_2__FF_INPUT;
  wire mi1_reg_30__FF_INPUT;
  wire mi1_reg_31__FF_INPUT;
  wire mi1_reg_3__FF_INPUT;
  wire mi1_reg_4__FF_INPUT;
  wire mi1_reg_5__FF_INPUT;
  wire mi1_reg_6__FF_INPUT;
  wire mi1_reg_7__FF_INPUT;
  wire mi1_reg_8__FF_INPUT;
  wire mi1_reg_9__FF_INPUT;
  wire param_reg_0__FF_INPUT;
  wire param_reg_1__FF_INPUT;
  wire param_reg_2__FF_INPUT;
  wire param_reg_3__FF_INPUT;
  wire param_reg_4__FF_INPUT;
  wire param_reg_5__FF_INPUT;
  wire param_reg_6__FF_INPUT;
  wire param_reg_7__FF_INPUT;
  output \read_data[0] ;
  output \read_data[10] ;
  output \read_data[11] ;
  output \read_data[12] ;
  output \read_data[13] ;
  output \read_data[14] ;
  output \read_data[15] ;
  output \read_data[16] ;
  output \read_data[17] ;
  output \read_data[18] ;
  output \read_data[19] ;
  output \read_data[1] ;
  output \read_data[20] ;
  output \read_data[21] ;
  output \read_data[22] ;
  output \read_data[23] ;
  output \read_data[24] ;
  output \read_data[25] ;
  output \read_data[26] ;
  output \read_data[27] ;
  output \read_data[28] ;
  output \read_data[29] ;
  output \read_data[2] ;
  output \read_data[30] ;
  output \read_data[31] ;
  output \read_data[3] ;
  output \read_data[4] ;
  output \read_data[5] ;
  output \read_data[6] ;
  output \read_data[7] ;
  output \read_data[8] ;
  output \read_data[9] ;
  input reset_n;
  wire reset_n_bF_buf0;
  wire reset_n_bF_buf1;
  wire reset_n_bF_buf10;
  wire reset_n_bF_buf11;
  wire reset_n_bF_buf12;
  wire reset_n_bF_buf13;
  wire reset_n_bF_buf14;
  wire reset_n_bF_buf15;
  wire reset_n_bF_buf16;
  wire reset_n_bF_buf17;
  wire reset_n_bF_buf18;
  wire reset_n_bF_buf19;
  wire reset_n_bF_buf2;
  wire reset_n_bF_buf20;
  wire reset_n_bF_buf21;
  wire reset_n_bF_buf22;
  wire reset_n_bF_buf23;
  wire reset_n_bF_buf24;
  wire reset_n_bF_buf25;
  wire reset_n_bF_buf26;
  wire reset_n_bF_buf27;
  wire reset_n_bF_buf28;
  wire reset_n_bF_buf29;
  wire reset_n_bF_buf3;
  wire reset_n_bF_buf30;
  wire reset_n_bF_buf31;
  wire reset_n_bF_buf32;
  wire reset_n_bF_buf33;
  wire reset_n_bF_buf34;
  wire reset_n_bF_buf35;
  wire reset_n_bF_buf36;
  wire reset_n_bF_buf37;
  wire reset_n_bF_buf38;
  wire reset_n_bF_buf39;
  wire reset_n_bF_buf4;
  wire reset_n_bF_buf40;
  wire reset_n_bF_buf41;
  wire reset_n_bF_buf42;
  wire reset_n_bF_buf43;
  wire reset_n_bF_buf44;
  wire reset_n_bF_buf45;
  wire reset_n_bF_buf46;
  wire reset_n_bF_buf47;
  wire reset_n_bF_buf48;
  wire reset_n_bF_buf49;
  wire reset_n_bF_buf5;
  wire reset_n_bF_buf50;
  wire reset_n_bF_buf51;
  wire reset_n_bF_buf52;
  wire reset_n_bF_buf53;
  wire reset_n_bF_buf54;
  wire reset_n_bF_buf55;
  wire reset_n_bF_buf56;
  wire reset_n_bF_buf57;
  wire reset_n_bF_buf58;
  wire reset_n_bF_buf59;
  wire reset_n_bF_buf6;
  wire reset_n_bF_buf60;
  wire reset_n_bF_buf61;
  wire reset_n_bF_buf62;
  wire reset_n_bF_buf63;
  wire reset_n_bF_buf64;
  wire reset_n_bF_buf65;
  wire reset_n_bF_buf66;
  wire reset_n_bF_buf67;
  wire reset_n_bF_buf68;
  wire reset_n_bF_buf69;
  wire reset_n_bF_buf7;
  wire reset_n_bF_buf70;
  wire reset_n_bF_buf71;
  wire reset_n_bF_buf72;
  wire reset_n_bF_buf73;
  wire reset_n_bF_buf74;
  wire reset_n_bF_buf75;
  wire reset_n_bF_buf76;
  wire reset_n_bF_buf77;
  wire reset_n_bF_buf78;
  wire reset_n_bF_buf79;
  wire reset_n_bF_buf8;
  wire reset_n_bF_buf80;
  wire reset_n_bF_buf81;
  wire reset_n_bF_buf82;
  wire reset_n_bF_buf83;
  wire reset_n_bF_buf84;
  wire reset_n_bF_buf9;
  wire reset_n_hier0_bF_buf0;
  wire reset_n_hier0_bF_buf1;
  wire reset_n_hier0_bF_buf2;
  wire reset_n_hier0_bF_buf3;
  wire reset_n_hier0_bF_buf4;
  wire reset_n_hier0_bF_buf5;
  wire reset_n_hier0_bF_buf6;
  wire reset_n_hier0_bF_buf7;
  wire reset_n_hier0_bF_buf8;
  input we;
  wire word0_reg_0_;
  wire word0_reg_0__FF_INPUT;
  wire word0_reg_10_;
  wire word0_reg_10__FF_INPUT;
  wire word0_reg_11_;
  wire word0_reg_11__FF_INPUT;
  wire word0_reg_12_;
  wire word0_reg_12__FF_INPUT;
  wire word0_reg_13_;
  wire word0_reg_13__FF_INPUT;
  wire word0_reg_14_;
  wire word0_reg_14__FF_INPUT;
  wire word0_reg_15_;
  wire word0_reg_15__FF_INPUT;
  wire word0_reg_16_;
  wire word0_reg_16__FF_INPUT;
  wire word0_reg_17_;
  wire word0_reg_17__FF_INPUT;
  wire word0_reg_18_;
  wire word0_reg_18__FF_INPUT;
  wire word0_reg_19_;
  wire word0_reg_19__FF_INPUT;
  wire word0_reg_1_;
  wire word0_reg_1__FF_INPUT;
  wire word0_reg_20_;
  wire word0_reg_20__FF_INPUT;
  wire word0_reg_21_;
  wire word0_reg_21__FF_INPUT;
  wire word0_reg_22_;
  wire word0_reg_22__FF_INPUT;
  wire word0_reg_23_;
  wire word0_reg_23__FF_INPUT;
  wire word0_reg_24_;
  wire word0_reg_24__FF_INPUT;
  wire word0_reg_25_;
  wire word0_reg_25__FF_INPUT;
  wire word0_reg_26_;
  wire word0_reg_26__FF_INPUT;
  wire word0_reg_27_;
  wire word0_reg_27__FF_INPUT;
  wire word0_reg_28_;
  wire word0_reg_28__FF_INPUT;
  wire word0_reg_29_;
  wire word0_reg_29__FF_INPUT;
  wire word0_reg_2_;
  wire word0_reg_2__FF_INPUT;
  wire word0_reg_30_;
  wire word0_reg_30__FF_INPUT;
  wire word0_reg_31_;
  wire word0_reg_31__FF_INPUT;
  wire word0_reg_3_;
  wire word0_reg_3__FF_INPUT;
  wire word0_reg_4_;
  wire word0_reg_4__FF_INPUT;
  wire word0_reg_5_;
  wire word0_reg_5__FF_INPUT;
  wire word0_reg_6_;
  wire word0_reg_6__FF_INPUT;
  wire word0_reg_7_;
  wire word0_reg_7__FF_INPUT;
  wire word0_reg_8_;
  wire word0_reg_8__FF_INPUT;
  wire word0_reg_9_;
  wire word0_reg_9__FF_INPUT;
  wire word1_reg_0_;
  wire word1_reg_0__FF_INPUT;
  wire word1_reg_10_;
  wire word1_reg_10__FF_INPUT;
  wire word1_reg_11_;
  wire word1_reg_11__FF_INPUT;
  wire word1_reg_12_;
  wire word1_reg_12__FF_INPUT;
  wire word1_reg_13_;
  wire word1_reg_13__FF_INPUT;
  wire word1_reg_14_;
  wire word1_reg_14__FF_INPUT;
  wire word1_reg_15_;
  wire word1_reg_15__FF_INPUT;
  wire word1_reg_16_;
  wire word1_reg_16__FF_INPUT;
  wire word1_reg_17_;
  wire word1_reg_17__FF_INPUT;
  wire word1_reg_18_;
  wire word1_reg_18__FF_INPUT;
  wire word1_reg_19_;
  wire word1_reg_19__FF_INPUT;
  wire word1_reg_1_;
  wire word1_reg_1__FF_INPUT;
  wire word1_reg_20_;
  wire word1_reg_20__FF_INPUT;
  wire word1_reg_21_;
  wire word1_reg_21__FF_INPUT;
  wire word1_reg_22_;
  wire word1_reg_22__FF_INPUT;
  wire word1_reg_23_;
  wire word1_reg_23__FF_INPUT;
  wire word1_reg_24_;
  wire word1_reg_24__FF_INPUT;
  wire word1_reg_25_;
  wire word1_reg_25__FF_INPUT;
  wire word1_reg_26_;
  wire word1_reg_26__FF_INPUT;
  wire word1_reg_27_;
  wire word1_reg_27__FF_INPUT;
  wire word1_reg_28_;
  wire word1_reg_28__FF_INPUT;
  wire word1_reg_29_;
  wire word1_reg_29__FF_INPUT;
  wire word1_reg_2_;
  wire word1_reg_2__FF_INPUT;
  wire word1_reg_30_;
  wire word1_reg_30__FF_INPUT;
  wire word1_reg_31_;
  wire word1_reg_31__FF_INPUT;
  wire word1_reg_3_;
  wire word1_reg_3__FF_INPUT;
  wire word1_reg_4_;
  wire word1_reg_4__FF_INPUT;
  wire word1_reg_5_;
  wire word1_reg_5__FF_INPUT;
  wire word1_reg_6_;
  wire word1_reg_6__FF_INPUT;
  wire word1_reg_7_;
  wire word1_reg_7__FF_INPUT;
  wire word1_reg_8_;
  wire word1_reg_8__FF_INPUT;
  wire word1_reg_9_;
  wire word1_reg_9__FF_INPUT;
  wire word2_reg_0_;
  wire word2_reg_0__FF_INPUT;
  wire word2_reg_10_;
  wire word2_reg_10__FF_INPUT;
  wire word2_reg_11_;
  wire word2_reg_11__FF_INPUT;
  wire word2_reg_12_;
  wire word2_reg_12__FF_INPUT;
  wire word2_reg_13_;
  wire word2_reg_13__FF_INPUT;
  wire word2_reg_14_;
  wire word2_reg_14__FF_INPUT;
  wire word2_reg_15_;
  wire word2_reg_15__FF_INPUT;
  wire word2_reg_16_;
  wire word2_reg_16__FF_INPUT;
  wire word2_reg_17_;
  wire word2_reg_17__FF_INPUT;
  wire word2_reg_18_;
  wire word2_reg_18__FF_INPUT;
  wire word2_reg_19_;
  wire word2_reg_19__FF_INPUT;
  wire word2_reg_1_;
  wire word2_reg_1__FF_INPUT;
  wire word2_reg_20_;
  wire word2_reg_20__FF_INPUT;
  wire word2_reg_21_;
  wire word2_reg_21__FF_INPUT;
  wire word2_reg_22_;
  wire word2_reg_22__FF_INPUT;
  wire word2_reg_23_;
  wire word2_reg_23__FF_INPUT;
  wire word2_reg_24_;
  wire word2_reg_24__FF_INPUT;
  wire word2_reg_25_;
  wire word2_reg_25__FF_INPUT;
  wire word2_reg_26_;
  wire word2_reg_26__FF_INPUT;
  wire word2_reg_27_;
  wire word2_reg_27__FF_INPUT;
  wire word2_reg_28_;
  wire word2_reg_28__FF_INPUT;
  wire word2_reg_29_;
  wire word2_reg_29__FF_INPUT;
  wire word2_reg_2_;
  wire word2_reg_2__FF_INPUT;
  wire word2_reg_30_;
  wire word2_reg_30__FF_INPUT;
  wire word2_reg_31_;
  wire word2_reg_31__FF_INPUT;
  wire word2_reg_3_;
  wire word2_reg_3__FF_INPUT;
  wire word2_reg_4_;
  wire word2_reg_4__FF_INPUT;
  wire word2_reg_5_;
  wire word2_reg_5__FF_INPUT;
  wire word2_reg_6_;
  wire word2_reg_6__FF_INPUT;
  wire word2_reg_7_;
  wire word2_reg_7__FF_INPUT;
  wire word2_reg_8_;
  wire word2_reg_8__FF_INPUT;
  wire word2_reg_9_;
  wire word2_reg_9__FF_INPUT;
  wire word3_reg_0_;
  wire word3_reg_0__FF_INPUT;
  wire word3_reg_10_;
  wire word3_reg_10__FF_INPUT;
  wire word3_reg_11_;
  wire word3_reg_11__FF_INPUT;
  wire word3_reg_12_;
  wire word3_reg_12__FF_INPUT;
  wire word3_reg_13_;
  wire word3_reg_13__FF_INPUT;
  wire word3_reg_14_;
  wire word3_reg_14__FF_INPUT;
  wire word3_reg_15_;
  wire word3_reg_15__FF_INPUT;
  wire word3_reg_16_;
  wire word3_reg_16__FF_INPUT;
  wire word3_reg_17_;
  wire word3_reg_17__FF_INPUT;
  wire word3_reg_18_;
  wire word3_reg_18__FF_INPUT;
  wire word3_reg_19_;
  wire word3_reg_19__FF_INPUT;
  wire word3_reg_1_;
  wire word3_reg_1__FF_INPUT;
  wire word3_reg_20_;
  wire word3_reg_20__FF_INPUT;
  wire word3_reg_21_;
  wire word3_reg_21__FF_INPUT;
  wire word3_reg_22_;
  wire word3_reg_22__FF_INPUT;
  wire word3_reg_23_;
  wire word3_reg_23__FF_INPUT;
  wire word3_reg_24_;
  wire word3_reg_24__FF_INPUT;
  wire word3_reg_25_;
  wire word3_reg_25__FF_INPUT;
  wire word3_reg_26_;
  wire word3_reg_26__FF_INPUT;
  wire word3_reg_27_;
  wire word3_reg_27__FF_INPUT;
  wire word3_reg_28_;
  wire word3_reg_28__FF_INPUT;
  wire word3_reg_29_;
  wire word3_reg_29__FF_INPUT;
  wire word3_reg_2_;
  wire word3_reg_2__FF_INPUT;
  wire word3_reg_30_;
  wire word3_reg_30__FF_INPUT;
  wire word3_reg_31_;
  wire word3_reg_31__FF_INPUT;
  wire word3_reg_3_;
  wire word3_reg_3__FF_INPUT;
  wire word3_reg_4_;
  wire word3_reg_4__FF_INPUT;
  wire word3_reg_5_;
  wire word3_reg_5__FF_INPUT;
  wire word3_reg_6_;
  wire word3_reg_6__FF_INPUT;
  wire word3_reg_7_;
  wire word3_reg_7__FF_INPUT;
  wire word3_reg_8_;
  wire word3_reg_8__FF_INPUT;
  wire word3_reg_9_;
  wire word3_reg_9__FF_INPUT;
  input \write_data[0] ;
  input \write_data[10] ;
  input \write_data[11] ;
  input \write_data[12] ;
  input \write_data[13] ;
  input \write_data[14] ;
  input \write_data[15] ;
  input \write_data[16] ;
  input \write_data[17] ;
  input \write_data[18] ;
  input \write_data[19] ;
  input \write_data[1] ;
  input \write_data[20] ;
  input \write_data[21] ;
  input \write_data[22] ;
  input \write_data[23] ;
  input \write_data[24] ;
  input \write_data[25] ;
  input \write_data[26] ;
  input \write_data[27] ;
  input \write_data[28] ;
  input \write_data[29] ;
  input \write_data[2] ;
  input \write_data[30] ;
  input \write_data[31] ;
  input \write_data[3] ;
  input \write_data[4] ;
  input \write_data[5] ;
  input \write_data[6] ;
  input \write_data[7] ;
  input \write_data[8] ;
  input \write_data[9] ;
  AND2X2 AND2X2_1 ( .A(_abc_19068_n870_1), .B(\addr[3] ), .Y(_abc_19068_n871_1) );
  AND2X2 AND2X2_10 ( .A(_abc_19068_n881), .B(_abc_19068_n884), .Y(_abc_19068_n885_1) );
  AND2X2 AND2X2_100 ( .A(_abc_19068_n885_1), .B(core_final_rounds_0_), .Y(_abc_19068_n1043) );
  AND2X2 AND2X2_1000 ( .A(_abc_19068_n2511), .B(_abc_19068_n2508), .Y(key3_reg_4__FF_INPUT) );
  AND2X2 AND2X2_1001 ( .A(_abc_19068_n2487_bF_buf4), .B(_abc_19068_n2165), .Y(_abc_19068_n2514) );
  AND2X2 AND2X2_1002 ( .A(_abc_19068_n2515), .B(reset_n_bF_buf57), .Y(_abc_19068_n2516) );
  AND2X2 AND2X2_1003 ( .A(_abc_19068_n2516), .B(_abc_19068_n2513), .Y(key3_reg_5__FF_INPUT) );
  AND2X2 AND2X2_1004 ( .A(_abc_19068_n2487_bF_buf2), .B(_abc_19068_n2171), .Y(_abc_19068_n2519) );
  AND2X2 AND2X2_1005 ( .A(_abc_19068_n2520), .B(reset_n_bF_buf56), .Y(_abc_19068_n2521) );
  AND2X2 AND2X2_1006 ( .A(_abc_19068_n2521), .B(_abc_19068_n2518), .Y(key3_reg_6__FF_INPUT) );
  AND2X2 AND2X2_1007 ( .A(_abc_19068_n2487_bF_buf0), .B(_abc_19068_n2177), .Y(_abc_19068_n2524) );
  AND2X2 AND2X2_1008 ( .A(_abc_19068_n2525), .B(reset_n_bF_buf55), .Y(_abc_19068_n2526) );
  AND2X2 AND2X2_1009 ( .A(_abc_19068_n2526), .B(_abc_19068_n2523), .Y(key3_reg_7__FF_INPUT) );
  AND2X2 AND2X2_101 ( .A(_abc_19068_n926_bF_buf0), .B(core_key_4_), .Y(_abc_19068_n1044_1) );
  AND2X2 AND2X2_1010 ( .A(_abc_19068_n2487_bF_buf6), .B(_abc_19068_n2183), .Y(_abc_19068_n2529) );
  AND2X2 AND2X2_1011 ( .A(_abc_19068_n2530), .B(reset_n_bF_buf54), .Y(_abc_19068_n2531) );
  AND2X2 AND2X2_1012 ( .A(_abc_19068_n2531), .B(_abc_19068_n2528), .Y(key3_reg_8__FF_INPUT) );
  AND2X2 AND2X2_1013 ( .A(_abc_19068_n2487_bF_buf4), .B(_abc_19068_n2189), .Y(_abc_19068_n2534) );
  AND2X2 AND2X2_1014 ( .A(_abc_19068_n2535), .B(reset_n_bF_buf53), .Y(_abc_19068_n2536) );
  AND2X2 AND2X2_1015 ( .A(_abc_19068_n2536), .B(_abc_19068_n2533), .Y(key3_reg_9__FF_INPUT) );
  AND2X2 AND2X2_1016 ( .A(_abc_19068_n2487_bF_buf2), .B(_abc_19068_n2195), .Y(_abc_19068_n2539) );
  AND2X2 AND2X2_1017 ( .A(_abc_19068_n2540), .B(reset_n_bF_buf52), .Y(_abc_19068_n2541) );
  AND2X2 AND2X2_1018 ( .A(_abc_19068_n2541), .B(_abc_19068_n2538), .Y(key3_reg_10__FF_INPUT) );
  AND2X2 AND2X2_1019 ( .A(_abc_19068_n2487_bF_buf0), .B(_abc_19068_n2201), .Y(_abc_19068_n2544) );
  AND2X2 AND2X2_102 ( .A(_abc_19068_n924_1_bF_buf0), .B(core_key_36_), .Y(_abc_19068_n1046) );
  AND2X2 AND2X2_1020 ( .A(_abc_19068_n2545), .B(reset_n_bF_buf51), .Y(_abc_19068_n2546) );
  AND2X2 AND2X2_1021 ( .A(_abc_19068_n2546), .B(_abc_19068_n2543), .Y(key3_reg_11__FF_INPUT) );
  AND2X2 AND2X2_1022 ( .A(_abc_19068_n2487_bF_buf6), .B(_abc_19068_n2207), .Y(_abc_19068_n2549) );
  AND2X2 AND2X2_1023 ( .A(_abc_19068_n2550), .B(reset_n_bF_buf50), .Y(_abc_19068_n2551) );
  AND2X2 AND2X2_1024 ( .A(_abc_19068_n2551), .B(_abc_19068_n2548), .Y(key3_reg_12__FF_INPUT) );
  AND2X2 AND2X2_1025 ( .A(_abc_19068_n2487_bF_buf4), .B(_abc_19068_n2213), .Y(_abc_19068_n2554) );
  AND2X2 AND2X2_1026 ( .A(_abc_19068_n2555), .B(reset_n_bF_buf49), .Y(_abc_19068_n2556) );
  AND2X2 AND2X2_1027 ( .A(_abc_19068_n2556), .B(_abc_19068_n2553), .Y(key3_reg_13__FF_INPUT) );
  AND2X2 AND2X2_1028 ( .A(_abc_19068_n2487_bF_buf2), .B(_abc_19068_n2219), .Y(_abc_19068_n2559) );
  AND2X2 AND2X2_1029 ( .A(_abc_19068_n2560), .B(reset_n_bF_buf48), .Y(_abc_19068_n2561) );
  AND2X2 AND2X2_103 ( .A(_abc_19068_n939_1_bF_buf0), .B(core_key_68_), .Y(_abc_19068_n1047_1) );
  AND2X2 AND2X2_1030 ( .A(_abc_19068_n2561), .B(_abc_19068_n2558), .Y(key3_reg_14__FF_INPUT) );
  AND2X2 AND2X2_1031 ( .A(_abc_19068_n2487_bF_buf0), .B(_abc_19068_n2225), .Y(_abc_19068_n2564) );
  AND2X2 AND2X2_1032 ( .A(_abc_19068_n2565), .B(reset_n_bF_buf47), .Y(_abc_19068_n2566) );
  AND2X2 AND2X2_1033 ( .A(_abc_19068_n2566), .B(_abc_19068_n2563), .Y(key3_reg_15__FF_INPUT) );
  AND2X2 AND2X2_1034 ( .A(_abc_19068_n2487_bF_buf6), .B(_abc_19068_n2231), .Y(_abc_19068_n2569) );
  AND2X2 AND2X2_1035 ( .A(_abc_19068_n2570), .B(reset_n_bF_buf46), .Y(_abc_19068_n2571) );
  AND2X2 AND2X2_1036 ( .A(_abc_19068_n2571), .B(_abc_19068_n2568), .Y(key3_reg_16__FF_INPUT) );
  AND2X2 AND2X2_1037 ( .A(_abc_19068_n2487_bF_buf4), .B(_abc_19068_n2237), .Y(_abc_19068_n2574) );
  AND2X2 AND2X2_1038 ( .A(_abc_19068_n2575), .B(reset_n_bF_buf45), .Y(_abc_19068_n2576) );
  AND2X2 AND2X2_1039 ( .A(_abc_19068_n2576), .B(_abc_19068_n2573), .Y(key3_reg_17__FF_INPUT) );
  AND2X2 AND2X2_104 ( .A(_abc_19068_n923_bF_buf0), .B(_abc_19068_n1050_1), .Y(_auto_iopadmap_cc_313_execute_30317_4_) );
  AND2X2 AND2X2_1040 ( .A(_abc_19068_n2487_bF_buf2), .B(_abc_19068_n2243), .Y(_abc_19068_n2579) );
  AND2X2 AND2X2_1041 ( .A(_abc_19068_n2580), .B(reset_n_bF_buf44), .Y(_abc_19068_n2581) );
  AND2X2 AND2X2_1042 ( .A(_abc_19068_n2581), .B(_abc_19068_n2578), .Y(key3_reg_18__FF_INPUT) );
  AND2X2 AND2X2_1043 ( .A(_abc_19068_n2487_bF_buf0), .B(_abc_19068_n2249), .Y(_abc_19068_n2584) );
  AND2X2 AND2X2_1044 ( .A(_abc_19068_n2585), .B(reset_n_bF_buf43), .Y(_abc_19068_n2586) );
  AND2X2 AND2X2_1045 ( .A(_abc_19068_n2586), .B(_abc_19068_n2583), .Y(key3_reg_19__FF_INPUT) );
  AND2X2 AND2X2_1046 ( .A(_abc_19068_n2487_bF_buf6), .B(_abc_19068_n2255), .Y(_abc_19068_n2589) );
  AND2X2 AND2X2_1047 ( .A(_abc_19068_n2590), .B(reset_n_bF_buf42), .Y(_abc_19068_n2591) );
  AND2X2 AND2X2_1048 ( .A(_abc_19068_n2591), .B(_abc_19068_n2588), .Y(key3_reg_20__FF_INPUT) );
  AND2X2 AND2X2_1049 ( .A(_abc_19068_n2487_bF_buf4), .B(_abc_19068_n2261), .Y(_abc_19068_n2594) );
  AND2X2 AND2X2_105 ( .A(_abc_19068_n945_1_bF_buf4), .B(core_mi_5_), .Y(_abc_19068_n1052) );
  AND2X2 AND2X2_1050 ( .A(_abc_19068_n2595), .B(reset_n_bF_buf41), .Y(_abc_19068_n2596) );
  AND2X2 AND2X2_1051 ( .A(_abc_19068_n2596), .B(_abc_19068_n2593), .Y(key3_reg_21__FF_INPUT) );
  AND2X2 AND2X2_1052 ( .A(_abc_19068_n2487_bF_buf2), .B(_abc_19068_n2267), .Y(_abc_19068_n2599) );
  AND2X2 AND2X2_1053 ( .A(_abc_19068_n2600), .B(reset_n_bF_buf40), .Y(_abc_19068_n2601) );
  AND2X2 AND2X2_1054 ( .A(_abc_19068_n2601), .B(_abc_19068_n2598), .Y(key3_reg_22__FF_INPUT) );
  AND2X2 AND2X2_1055 ( .A(_abc_19068_n2487_bF_buf0), .B(_abc_19068_n2273), .Y(_abc_19068_n2604) );
  AND2X2 AND2X2_1056 ( .A(_abc_19068_n2605), .B(reset_n_bF_buf39), .Y(_abc_19068_n2606) );
  AND2X2 AND2X2_1057 ( .A(_abc_19068_n2606), .B(_abc_19068_n2603), .Y(key3_reg_23__FF_INPUT) );
  AND2X2 AND2X2_1058 ( .A(_abc_19068_n2487_bF_buf6), .B(_abc_19068_n2279), .Y(_abc_19068_n2609) );
  AND2X2 AND2X2_1059 ( .A(_abc_19068_n2610), .B(reset_n_bF_buf38), .Y(_abc_19068_n2611) );
  AND2X2 AND2X2_106 ( .A(_abc_19068_n915_1_bF_buf3), .B(core_mi_37_), .Y(_abc_19068_n1053_1) );
  AND2X2 AND2X2_1060 ( .A(_abc_19068_n2611), .B(_abc_19068_n2608), .Y(key3_reg_24__FF_INPUT) );
  AND2X2 AND2X2_1061 ( .A(_abc_19068_n2487_bF_buf4), .B(_abc_19068_n2285), .Y(_abc_19068_n2614) );
  AND2X2 AND2X2_1062 ( .A(_abc_19068_n2615), .B(reset_n_bF_buf37), .Y(_abc_19068_n2616) );
  AND2X2 AND2X2_1063 ( .A(_abc_19068_n2616), .B(_abc_19068_n2613), .Y(key3_reg_25__FF_INPUT) );
  AND2X2 AND2X2_1064 ( .A(_abc_19068_n2487_bF_buf2), .B(_abc_19068_n2291), .Y(_abc_19068_n2619) );
  AND2X2 AND2X2_1065 ( .A(_abc_19068_n2620), .B(reset_n_bF_buf36), .Y(_abc_19068_n2621) );
  AND2X2 AND2X2_1066 ( .A(_abc_19068_n2621), .B(_abc_19068_n2618), .Y(key3_reg_26__FF_INPUT) );
  AND2X2 AND2X2_1067 ( .A(_abc_19068_n2487_bF_buf0), .B(_abc_19068_n2297), .Y(_abc_19068_n2624) );
  AND2X2 AND2X2_1068 ( .A(_abc_19068_n2625), .B(reset_n_bF_buf35), .Y(_abc_19068_n2626) );
  AND2X2 AND2X2_1069 ( .A(_abc_19068_n2626), .B(_abc_19068_n2623), .Y(key3_reg_27__FF_INPUT) );
  AND2X2 AND2X2_107 ( .A(_abc_19068_n902_bF_buf3), .B(word2_reg_5_), .Y(_abc_19068_n1056_1) );
  AND2X2 AND2X2_1070 ( .A(_abc_19068_n2487_bF_buf6), .B(_abc_19068_n2303), .Y(_abc_19068_n2629) );
  AND2X2 AND2X2_1071 ( .A(_abc_19068_n2630), .B(reset_n_bF_buf34), .Y(_abc_19068_n2631) );
  AND2X2 AND2X2_1072 ( .A(_abc_19068_n2631), .B(_abc_19068_n2628), .Y(key3_reg_28__FF_INPUT) );
  AND2X2 AND2X2_1073 ( .A(_abc_19068_n2487_bF_buf4), .B(_abc_19068_n2309), .Y(_abc_19068_n2634) );
  AND2X2 AND2X2_1074 ( .A(_abc_19068_n2635), .B(reset_n_bF_buf33), .Y(_abc_19068_n2636) );
  AND2X2 AND2X2_1075 ( .A(_abc_19068_n2636), .B(_abc_19068_n2633), .Y(key3_reg_29__FF_INPUT) );
  AND2X2 AND2X2_1076 ( .A(_abc_19068_n2487_bF_buf2), .B(_abc_19068_n2315), .Y(_abc_19068_n2639) );
  AND2X2 AND2X2_1077 ( .A(_abc_19068_n2640), .B(reset_n_bF_buf32), .Y(_abc_19068_n2641) );
  AND2X2 AND2X2_1078 ( .A(_abc_19068_n2641), .B(_abc_19068_n2638), .Y(key3_reg_30__FF_INPUT) );
  AND2X2 AND2X2_1079 ( .A(_abc_19068_n2487_bF_buf0), .B(_abc_19068_n2321), .Y(_abc_19068_n2644) );
  AND2X2 AND2X2_108 ( .A(_abc_19068_n885_1), .B(core_final_rounds_1_), .Y(_abc_19068_n1057_1) );
  AND2X2 AND2X2_1080 ( .A(_abc_19068_n2645), .B(reset_n_bF_buf31), .Y(_abc_19068_n2646) );
  AND2X2 AND2X2_1081 ( .A(_abc_19068_n2646), .B(_abc_19068_n2643), .Y(key3_reg_31__FF_INPUT) );
  AND2X2 AND2X2_1082 ( .A(_abc_19068_n939_1_bF_buf2), .B(_abc_19068_n2132), .Y(_abc_19068_n2648) );
  AND2X2 AND2X2_1083 ( .A(_abc_19068_n2648_bF_buf6), .B(_abc_19068_n2135), .Y(_abc_19068_n2650) );
  AND2X2 AND2X2_1084 ( .A(_abc_19068_n2651), .B(reset_n_bF_buf30), .Y(_abc_19068_n2652) );
  AND2X2 AND2X2_1085 ( .A(_abc_19068_n2652), .B(_abc_19068_n2649), .Y(key2_reg_0__FF_INPUT) );
  AND2X2 AND2X2_1086 ( .A(_abc_19068_n2648_bF_buf4), .B(_abc_19068_n2141), .Y(_abc_19068_n2655) );
  AND2X2 AND2X2_1087 ( .A(_abc_19068_n2656), .B(reset_n_bF_buf29), .Y(_abc_19068_n2657) );
  AND2X2 AND2X2_1088 ( .A(_abc_19068_n2657), .B(_abc_19068_n2654), .Y(key2_reg_1__FF_INPUT) );
  AND2X2 AND2X2_1089 ( .A(_abc_19068_n2648_bF_buf2), .B(_abc_19068_n2147), .Y(_abc_19068_n2660) );
  AND2X2 AND2X2_109 ( .A(_abc_19068_n897_1_bF_buf3), .B(word0_reg_5_), .Y(_abc_19068_n1058) );
  AND2X2 AND2X2_1090 ( .A(_abc_19068_n2661), .B(reset_n_bF_buf28), .Y(_abc_19068_n2662) );
  AND2X2 AND2X2_1091 ( .A(_abc_19068_n2662), .B(_abc_19068_n2659), .Y(key2_reg_2__FF_INPUT) );
  AND2X2 AND2X2_1092 ( .A(_abc_19068_n2648_bF_buf0), .B(_abc_19068_n2153), .Y(_abc_19068_n2665) );
  AND2X2 AND2X2_1093 ( .A(_abc_19068_n2666), .B(reset_n_bF_buf27), .Y(_abc_19068_n2667) );
  AND2X2 AND2X2_1094 ( .A(_abc_19068_n2667), .B(_abc_19068_n2664), .Y(key2_reg_3__FF_INPUT) );
  AND2X2 AND2X2_1095 ( .A(_abc_19068_n2648_bF_buf6), .B(_abc_19068_n2159), .Y(_abc_19068_n2670) );
  AND2X2 AND2X2_1096 ( .A(_abc_19068_n2671), .B(reset_n_bF_buf26), .Y(_abc_19068_n2672) );
  AND2X2 AND2X2_1097 ( .A(_abc_19068_n2672), .B(_abc_19068_n2669), .Y(key2_reg_4__FF_INPUT) );
  AND2X2 AND2X2_1098 ( .A(_abc_19068_n2648_bF_buf4), .B(_abc_19068_n2165), .Y(_abc_19068_n2675) );
  AND2X2 AND2X2_1099 ( .A(_abc_19068_n2676), .B(reset_n_bF_buf25), .Y(_abc_19068_n2677) );
  AND2X2 AND2X2_11 ( .A(_abc_19068_n886_1), .B(_abc_19068_n872), .Y(_abc_19068_n887) );
  AND2X2 AND2X2_110 ( .A(_abc_19068_n941_bF_buf4), .B(core_key_101_), .Y(_abc_19068_n1062_1) );
  AND2X2 AND2X2_1100 ( .A(_abc_19068_n2677), .B(_abc_19068_n2674), .Y(key2_reg_5__FF_INPUT) );
  AND2X2 AND2X2_1101 ( .A(_abc_19068_n2648_bF_buf2), .B(_abc_19068_n2171), .Y(_abc_19068_n2680) );
  AND2X2 AND2X2_1102 ( .A(_abc_19068_n2681), .B(reset_n_bF_buf24), .Y(_abc_19068_n2682) );
  AND2X2 AND2X2_1103 ( .A(_abc_19068_n2682), .B(_abc_19068_n2679), .Y(key2_reg_6__FF_INPUT) );
  AND2X2 AND2X2_1104 ( .A(_abc_19068_n2648_bF_buf0), .B(_abc_19068_n2177), .Y(_abc_19068_n2685) );
  AND2X2 AND2X2_1105 ( .A(_abc_19068_n2686), .B(reset_n_bF_buf23), .Y(_abc_19068_n2687) );
  AND2X2 AND2X2_1106 ( .A(_abc_19068_n2687), .B(_abc_19068_n2684), .Y(key2_reg_7__FF_INPUT) );
  AND2X2 AND2X2_1107 ( .A(_abc_19068_n2648_bF_buf6), .B(_abc_19068_n2183), .Y(_abc_19068_n2690) );
  AND2X2 AND2X2_1108 ( .A(_abc_19068_n2691), .B(reset_n_bF_buf22), .Y(_abc_19068_n2692) );
  AND2X2 AND2X2_1109 ( .A(_abc_19068_n2692), .B(_abc_19068_n2689), .Y(key2_reg_8__FF_INPUT) );
  AND2X2 AND2X2_111 ( .A(_abc_19068_n939_1_bF_buf4), .B(core_key_69_), .Y(_abc_19068_n1063_1) );
  AND2X2 AND2X2_1110 ( .A(_abc_19068_n2648_bF_buf4), .B(_abc_19068_n2189), .Y(_abc_19068_n2695) );
  AND2X2 AND2X2_1111 ( .A(_abc_19068_n2696), .B(reset_n_bF_buf21), .Y(_abc_19068_n2697) );
  AND2X2 AND2X2_1112 ( .A(_abc_19068_n2697), .B(_abc_19068_n2694), .Y(key2_reg_9__FF_INPUT) );
  AND2X2 AND2X2_1113 ( .A(_abc_19068_n2648_bF_buf2), .B(_abc_19068_n2195), .Y(_abc_19068_n2700) );
  AND2X2 AND2X2_1114 ( .A(_abc_19068_n2701), .B(reset_n_bF_buf20), .Y(_abc_19068_n2702) );
  AND2X2 AND2X2_1115 ( .A(_abc_19068_n2702), .B(_abc_19068_n2699), .Y(key2_reg_10__FF_INPUT) );
  AND2X2 AND2X2_1116 ( .A(_abc_19068_n2648_bF_buf0), .B(_abc_19068_n2201), .Y(_abc_19068_n2705) );
  AND2X2 AND2X2_1117 ( .A(_abc_19068_n2706), .B(reset_n_bF_buf19), .Y(_abc_19068_n2707) );
  AND2X2 AND2X2_1118 ( .A(_abc_19068_n2707), .B(_abc_19068_n2704), .Y(key2_reg_11__FF_INPUT) );
  AND2X2 AND2X2_1119 ( .A(_abc_19068_n2648_bF_buf6), .B(_abc_19068_n2207), .Y(_abc_19068_n2710) );
  AND2X2 AND2X2_112 ( .A(_abc_19068_n926_bF_buf4), .B(core_key_5_), .Y(_abc_19068_n1065_1) );
  AND2X2 AND2X2_1120 ( .A(_abc_19068_n2711), .B(reset_n_bF_buf18), .Y(_abc_19068_n2712) );
  AND2X2 AND2X2_1121 ( .A(_abc_19068_n2712), .B(_abc_19068_n2709), .Y(key2_reg_12__FF_INPUT) );
  AND2X2 AND2X2_1122 ( .A(_abc_19068_n2648_bF_buf4), .B(_abc_19068_n2213), .Y(_abc_19068_n2715) );
  AND2X2 AND2X2_1123 ( .A(_abc_19068_n2716), .B(reset_n_bF_buf17), .Y(_abc_19068_n2717) );
  AND2X2 AND2X2_1124 ( .A(_abc_19068_n2717), .B(_abc_19068_n2714), .Y(key2_reg_13__FF_INPUT) );
  AND2X2 AND2X2_1125 ( .A(_abc_19068_n2648_bF_buf2), .B(_abc_19068_n2219), .Y(_abc_19068_n2720) );
  AND2X2 AND2X2_1126 ( .A(_abc_19068_n2721), .B(reset_n_bF_buf16), .Y(_abc_19068_n2722) );
  AND2X2 AND2X2_1127 ( .A(_abc_19068_n2722), .B(_abc_19068_n2719), .Y(key2_reg_14__FF_INPUT) );
  AND2X2 AND2X2_1128 ( .A(_abc_19068_n2648_bF_buf0), .B(_abc_19068_n2225), .Y(_abc_19068_n2725) );
  AND2X2 AND2X2_1129 ( .A(_abc_19068_n2726), .B(reset_n_bF_buf15), .Y(_abc_19068_n2727) );
  AND2X2 AND2X2_113 ( .A(_abc_19068_n924_1_bF_buf4), .B(core_key_37_), .Y(_abc_19068_n1066_1) );
  AND2X2 AND2X2_1130 ( .A(_abc_19068_n2727), .B(_abc_19068_n2724), .Y(key2_reg_15__FF_INPUT) );
  AND2X2 AND2X2_1131 ( .A(_abc_19068_n2648_bF_buf6), .B(_abc_19068_n2231), .Y(_abc_19068_n2730) );
  AND2X2 AND2X2_1132 ( .A(_abc_19068_n2731), .B(reset_n_bF_buf14), .Y(_abc_19068_n2732) );
  AND2X2 AND2X2_1133 ( .A(_abc_19068_n2732), .B(_abc_19068_n2729), .Y(key2_reg_16__FF_INPUT) );
  AND2X2 AND2X2_1134 ( .A(_abc_19068_n2648_bF_buf4), .B(_abc_19068_n2237), .Y(_abc_19068_n2735) );
  AND2X2 AND2X2_1135 ( .A(_abc_19068_n2736), .B(reset_n_bF_buf13), .Y(_abc_19068_n2737) );
  AND2X2 AND2X2_1136 ( .A(_abc_19068_n2737), .B(_abc_19068_n2734), .Y(key2_reg_17__FF_INPUT) );
  AND2X2 AND2X2_1137 ( .A(_abc_19068_n2648_bF_buf2), .B(_abc_19068_n2243), .Y(_abc_19068_n2740) );
  AND2X2 AND2X2_1138 ( .A(_abc_19068_n2741), .B(reset_n_bF_buf12), .Y(_abc_19068_n2742) );
  AND2X2 AND2X2_1139 ( .A(_abc_19068_n2742), .B(_abc_19068_n2739), .Y(key2_reg_18__FF_INPUT) );
  AND2X2 AND2X2_114 ( .A(_abc_19068_n916_1_bF_buf3), .B(word1_reg_5_), .Y(_abc_19068_n1068_1) );
  AND2X2 AND2X2_1140 ( .A(_abc_19068_n2648_bF_buf0), .B(_abc_19068_n2249), .Y(_abc_19068_n2745) );
  AND2X2 AND2X2_1141 ( .A(_abc_19068_n2746), .B(reset_n_bF_buf11), .Y(_abc_19068_n2747) );
  AND2X2 AND2X2_1142 ( .A(_abc_19068_n2747), .B(_abc_19068_n2744), .Y(key2_reg_19__FF_INPUT) );
  AND2X2 AND2X2_1143 ( .A(_abc_19068_n2648_bF_buf6), .B(_abc_19068_n2255), .Y(_abc_19068_n2750) );
  AND2X2 AND2X2_1144 ( .A(_abc_19068_n2751), .B(reset_n_bF_buf10), .Y(_abc_19068_n2752) );
  AND2X2 AND2X2_1145 ( .A(_abc_19068_n2752), .B(_abc_19068_n2749), .Y(key2_reg_20__FF_INPUT) );
  AND2X2 AND2X2_1146 ( .A(_abc_19068_n2648_bF_buf4), .B(_abc_19068_n2261), .Y(_abc_19068_n2755) );
  AND2X2 AND2X2_1147 ( .A(_abc_19068_n2756), .B(reset_n_bF_buf9), .Y(_abc_19068_n2757) );
  AND2X2 AND2X2_1148 ( .A(_abc_19068_n2757), .B(_abc_19068_n2754), .Y(key2_reg_21__FF_INPUT) );
  AND2X2 AND2X2_1149 ( .A(_abc_19068_n2648_bF_buf2), .B(_abc_19068_n2267), .Y(_abc_19068_n2760) );
  AND2X2 AND2X2_115 ( .A(_abc_19068_n899_bF_buf3), .B(word3_reg_5_), .Y(_abc_19068_n1069_1) );
  AND2X2 AND2X2_1150 ( .A(_abc_19068_n2761), .B(reset_n_bF_buf8), .Y(_abc_19068_n2762) );
  AND2X2 AND2X2_1151 ( .A(_abc_19068_n2762), .B(_abc_19068_n2759), .Y(key2_reg_22__FF_INPUT) );
  AND2X2 AND2X2_1152 ( .A(_abc_19068_n2648_bF_buf0), .B(_abc_19068_n2273), .Y(_abc_19068_n2765) );
  AND2X2 AND2X2_1153 ( .A(_abc_19068_n2766), .B(reset_n_bF_buf7), .Y(_abc_19068_n2767) );
  AND2X2 AND2X2_1154 ( .A(_abc_19068_n2767), .B(_abc_19068_n2764), .Y(key2_reg_23__FF_INPUT) );
  AND2X2 AND2X2_1155 ( .A(_abc_19068_n2648_bF_buf6), .B(_abc_19068_n2279), .Y(_abc_19068_n2770) );
  AND2X2 AND2X2_1156 ( .A(_abc_19068_n2771), .B(reset_n_bF_buf6), .Y(_abc_19068_n2772) );
  AND2X2 AND2X2_1157 ( .A(_abc_19068_n2772), .B(_abc_19068_n2769), .Y(key2_reg_24__FF_INPUT) );
  AND2X2 AND2X2_1158 ( .A(_abc_19068_n2648_bF_buf4), .B(_abc_19068_n2285), .Y(_abc_19068_n2775) );
  AND2X2 AND2X2_1159 ( .A(_abc_19068_n2776), .B(reset_n_bF_buf5), .Y(_abc_19068_n2777) );
  AND2X2 AND2X2_116 ( .A(_abc_19068_n1073), .B(_abc_19068_n923_bF_buf4), .Y(_auto_iopadmap_cc_313_execute_30317_5_) );
  AND2X2 AND2X2_1160 ( .A(_abc_19068_n2777), .B(_abc_19068_n2774), .Y(key2_reg_25__FF_INPUT) );
  AND2X2 AND2X2_1161 ( .A(_abc_19068_n2648_bF_buf2), .B(_abc_19068_n2291), .Y(_abc_19068_n2780) );
  AND2X2 AND2X2_1162 ( .A(_abc_19068_n2781), .B(reset_n_bF_buf4), .Y(_abc_19068_n2782) );
  AND2X2 AND2X2_1163 ( .A(_abc_19068_n2782), .B(_abc_19068_n2779), .Y(key2_reg_26__FF_INPUT) );
  AND2X2 AND2X2_1164 ( .A(_abc_19068_n2648_bF_buf0), .B(_abc_19068_n2297), .Y(_abc_19068_n2785) );
  AND2X2 AND2X2_1165 ( .A(_abc_19068_n2786), .B(reset_n_bF_buf3), .Y(_abc_19068_n2787) );
  AND2X2 AND2X2_1166 ( .A(_abc_19068_n2787), .B(_abc_19068_n2784), .Y(key2_reg_27__FF_INPUT) );
  AND2X2 AND2X2_1167 ( .A(_abc_19068_n2648_bF_buf6), .B(_abc_19068_n2303), .Y(_abc_19068_n2790) );
  AND2X2 AND2X2_1168 ( .A(_abc_19068_n2791), .B(reset_n_bF_buf2), .Y(_abc_19068_n2792) );
  AND2X2 AND2X2_1169 ( .A(_abc_19068_n2792), .B(_abc_19068_n2789), .Y(key2_reg_28__FF_INPUT) );
  AND2X2 AND2X2_117 ( .A(_abc_19068_n897_1_bF_buf2), .B(word0_reg_6_), .Y(_abc_19068_n1075_1) );
  AND2X2 AND2X2_1170 ( .A(_abc_19068_n2648_bF_buf4), .B(_abc_19068_n2309), .Y(_abc_19068_n2795) );
  AND2X2 AND2X2_1171 ( .A(_abc_19068_n2796), .B(reset_n_bF_buf1), .Y(_abc_19068_n2797) );
  AND2X2 AND2X2_1172 ( .A(_abc_19068_n2797), .B(_abc_19068_n2794), .Y(key2_reg_29__FF_INPUT) );
  AND2X2 AND2X2_1173 ( .A(_abc_19068_n2648_bF_buf2), .B(_abc_19068_n2315), .Y(_abc_19068_n2800) );
  AND2X2 AND2X2_1174 ( .A(_abc_19068_n2801), .B(reset_n_bF_buf0), .Y(_abc_19068_n2802) );
  AND2X2 AND2X2_1175 ( .A(_abc_19068_n2802), .B(_abc_19068_n2799), .Y(key2_reg_30__FF_INPUT) );
  AND2X2 AND2X2_1176 ( .A(_abc_19068_n2648_bF_buf0), .B(_abc_19068_n2321), .Y(_abc_19068_n2805) );
  AND2X2 AND2X2_1177 ( .A(_abc_19068_n2806), .B(reset_n_bF_buf84), .Y(_abc_19068_n2807) );
  AND2X2 AND2X2_1178 ( .A(_abc_19068_n2807), .B(_abc_19068_n2804), .Y(key2_reg_31__FF_INPUT) );
  AND2X2 AND2X2_1179 ( .A(_abc_19068_n924_1_bF_buf2), .B(_abc_19068_n2132), .Y(_abc_19068_n2809) );
  AND2X2 AND2X2_118 ( .A(_abc_19068_n915_1_bF_buf2), .B(core_mi_38_), .Y(_abc_19068_n1076) );
  AND2X2 AND2X2_1180 ( .A(_abc_19068_n2809_bF_buf6), .B(_abc_19068_n2135), .Y(_abc_19068_n2811) );
  AND2X2 AND2X2_1181 ( .A(_abc_19068_n2812), .B(reset_n_bF_buf83), .Y(_abc_19068_n2813) );
  AND2X2 AND2X2_1182 ( .A(_abc_19068_n2813), .B(_abc_19068_n2810), .Y(key1_reg_0__FF_INPUT) );
  AND2X2 AND2X2_1183 ( .A(_abc_19068_n2809_bF_buf4), .B(_abc_19068_n2141), .Y(_abc_19068_n2816) );
  AND2X2 AND2X2_1184 ( .A(_abc_19068_n2817), .B(reset_n_bF_buf82), .Y(_abc_19068_n2818) );
  AND2X2 AND2X2_1185 ( .A(_abc_19068_n2818), .B(_abc_19068_n2815), .Y(key1_reg_1__FF_INPUT) );
  AND2X2 AND2X2_1186 ( .A(_abc_19068_n2809_bF_buf2), .B(_abc_19068_n2147), .Y(_abc_19068_n2821) );
  AND2X2 AND2X2_1187 ( .A(_abc_19068_n2822), .B(reset_n_bF_buf81), .Y(_abc_19068_n2823) );
  AND2X2 AND2X2_1188 ( .A(_abc_19068_n2823), .B(_abc_19068_n2820), .Y(key1_reg_2__FF_INPUT) );
  AND2X2 AND2X2_1189 ( .A(_abc_19068_n2809_bF_buf0), .B(_abc_19068_n2153), .Y(_abc_19068_n2826) );
  AND2X2 AND2X2_119 ( .A(_abc_19068_n945_1_bF_buf3), .B(core_mi_6_), .Y(_abc_19068_n1078_1) );
  AND2X2 AND2X2_1190 ( .A(_abc_19068_n2827), .B(reset_n_bF_buf80), .Y(_abc_19068_n2828) );
  AND2X2 AND2X2_1191 ( .A(_abc_19068_n2828), .B(_abc_19068_n2825), .Y(key1_reg_3__FF_INPUT) );
  AND2X2 AND2X2_1192 ( .A(_abc_19068_n2809_bF_buf6), .B(_abc_19068_n2159), .Y(_abc_19068_n2831) );
  AND2X2 AND2X2_1193 ( .A(_abc_19068_n2832), .B(reset_n_bF_buf79), .Y(_abc_19068_n2833) );
  AND2X2 AND2X2_1194 ( .A(_abc_19068_n2833), .B(_abc_19068_n2830), .Y(key1_reg_4__FF_INPUT) );
  AND2X2 AND2X2_1195 ( .A(_abc_19068_n2809_bF_buf4), .B(_abc_19068_n2165), .Y(_abc_19068_n2836) );
  AND2X2 AND2X2_1196 ( .A(_abc_19068_n2837), .B(reset_n_bF_buf78), .Y(_abc_19068_n2838) );
  AND2X2 AND2X2_1197 ( .A(_abc_19068_n2838), .B(_abc_19068_n2835), .Y(key1_reg_5__FF_INPUT) );
  AND2X2 AND2X2_1198 ( .A(_abc_19068_n2809_bF_buf2), .B(_abc_19068_n2171), .Y(_abc_19068_n2841) );
  AND2X2 AND2X2_1199 ( .A(_abc_19068_n2842), .B(reset_n_bF_buf77), .Y(_abc_19068_n2843) );
  AND2X2 AND2X2_12 ( .A(_abc_19068_n887), .B(_abc_19068_n871_1), .Y(_abc_19068_n888_1) );
  AND2X2 AND2X2_120 ( .A(_abc_19068_n941_bF_buf3), .B(core_key_102_), .Y(_abc_19068_n1079) );
  AND2X2 AND2X2_1200 ( .A(_abc_19068_n2843), .B(_abc_19068_n2840), .Y(key1_reg_6__FF_INPUT) );
  AND2X2 AND2X2_1201 ( .A(_abc_19068_n2809_bF_buf0), .B(_abc_19068_n2177), .Y(_abc_19068_n2846) );
  AND2X2 AND2X2_1202 ( .A(_abc_19068_n2847), .B(reset_n_bF_buf76), .Y(_abc_19068_n2848) );
  AND2X2 AND2X2_1203 ( .A(_abc_19068_n2848), .B(_abc_19068_n2845), .Y(key1_reg_7__FF_INPUT) );
  AND2X2 AND2X2_1204 ( .A(_abc_19068_n2809_bF_buf6), .B(_abc_19068_n2183), .Y(_abc_19068_n2851) );
  AND2X2 AND2X2_1205 ( .A(_abc_19068_n2852), .B(reset_n_bF_buf75), .Y(_abc_19068_n2853) );
  AND2X2 AND2X2_1206 ( .A(_abc_19068_n2853), .B(_abc_19068_n2850), .Y(key1_reg_8__FF_INPUT) );
  AND2X2 AND2X2_1207 ( .A(_abc_19068_n2809_bF_buf4), .B(_abc_19068_n2189), .Y(_abc_19068_n2856) );
  AND2X2 AND2X2_1208 ( .A(_abc_19068_n2857), .B(reset_n_bF_buf74), .Y(_abc_19068_n2858) );
  AND2X2 AND2X2_1209 ( .A(_abc_19068_n2858), .B(_abc_19068_n2855), .Y(key1_reg_9__FF_INPUT) );
  AND2X2 AND2X2_121 ( .A(_abc_19068_n916_1_bF_buf2), .B(word1_reg_6_), .Y(_abc_19068_n1082) );
  AND2X2 AND2X2_1210 ( .A(_abc_19068_n2809_bF_buf2), .B(_abc_19068_n2195), .Y(_abc_19068_n2861) );
  AND2X2 AND2X2_1211 ( .A(_abc_19068_n2862), .B(reset_n_bF_buf73), .Y(_abc_19068_n2863) );
  AND2X2 AND2X2_1212 ( .A(_abc_19068_n2863), .B(_abc_19068_n2860), .Y(key1_reg_10__FF_INPUT) );
  AND2X2 AND2X2_1213 ( .A(_abc_19068_n2809_bF_buf0), .B(_abc_19068_n2201), .Y(_abc_19068_n2866) );
  AND2X2 AND2X2_1214 ( .A(_abc_19068_n2867), .B(reset_n_bF_buf72), .Y(_abc_19068_n2868) );
  AND2X2 AND2X2_1215 ( .A(_abc_19068_n2868), .B(_abc_19068_n2865), .Y(key1_reg_11__FF_INPUT) );
  AND2X2 AND2X2_1216 ( .A(_abc_19068_n2809_bF_buf6), .B(_abc_19068_n2207), .Y(_abc_19068_n2871) );
  AND2X2 AND2X2_1217 ( .A(_abc_19068_n2872), .B(reset_n_bF_buf71), .Y(_abc_19068_n2873) );
  AND2X2 AND2X2_1218 ( .A(_abc_19068_n2873), .B(_abc_19068_n2870), .Y(key1_reg_12__FF_INPUT) );
  AND2X2 AND2X2_1219 ( .A(_abc_19068_n2809_bF_buf4), .B(_abc_19068_n2213), .Y(_abc_19068_n2876) );
  AND2X2 AND2X2_122 ( .A(_abc_19068_n902_bF_buf2), .B(word2_reg_6_), .Y(_abc_19068_n1083_1) );
  AND2X2 AND2X2_1220 ( .A(_abc_19068_n2877), .B(reset_n_bF_buf70), .Y(_abc_19068_n2878) );
  AND2X2 AND2X2_1221 ( .A(_abc_19068_n2878), .B(_abc_19068_n2875), .Y(key1_reg_13__FF_INPUT) );
  AND2X2 AND2X2_1222 ( .A(_abc_19068_n2809_bF_buf2), .B(_abc_19068_n2219), .Y(_abc_19068_n2881) );
  AND2X2 AND2X2_1223 ( .A(_abc_19068_n2882), .B(reset_n_bF_buf69), .Y(_abc_19068_n2883) );
  AND2X2 AND2X2_1224 ( .A(_abc_19068_n2883), .B(_abc_19068_n2880), .Y(key1_reg_14__FF_INPUT) );
  AND2X2 AND2X2_1225 ( .A(_abc_19068_n2809_bF_buf0), .B(_abc_19068_n2225), .Y(_abc_19068_n2886) );
  AND2X2 AND2X2_1226 ( .A(_abc_19068_n2887), .B(reset_n_bF_buf68), .Y(_abc_19068_n2888) );
  AND2X2 AND2X2_1227 ( .A(_abc_19068_n2888), .B(_abc_19068_n2885), .Y(key1_reg_15__FF_INPUT) );
  AND2X2 AND2X2_1228 ( .A(_abc_19068_n2809_bF_buf6), .B(_abc_19068_n2231), .Y(_abc_19068_n2891) );
  AND2X2 AND2X2_1229 ( .A(_abc_19068_n2892), .B(reset_n_bF_buf67), .Y(_abc_19068_n2893) );
  AND2X2 AND2X2_123 ( .A(_abc_19068_n899_bF_buf2), .B(word3_reg_6_), .Y(_abc_19068_n1085) );
  AND2X2 AND2X2_1230 ( .A(_abc_19068_n2893), .B(_abc_19068_n2890), .Y(key1_reg_16__FF_INPUT) );
  AND2X2 AND2X2_1231 ( .A(_abc_19068_n2809_bF_buf4), .B(_abc_19068_n2237), .Y(_abc_19068_n2896) );
  AND2X2 AND2X2_1232 ( .A(_abc_19068_n2897), .B(reset_n_bF_buf66), .Y(_abc_19068_n2898) );
  AND2X2 AND2X2_1233 ( .A(_abc_19068_n2898), .B(_abc_19068_n2895), .Y(key1_reg_17__FF_INPUT) );
  AND2X2 AND2X2_1234 ( .A(_abc_19068_n2809_bF_buf2), .B(_abc_19068_n2243), .Y(_abc_19068_n2901) );
  AND2X2 AND2X2_1235 ( .A(_abc_19068_n2902), .B(reset_n_bF_buf65), .Y(_abc_19068_n2903) );
  AND2X2 AND2X2_1236 ( .A(_abc_19068_n2903), .B(_abc_19068_n2900), .Y(key1_reg_18__FF_INPUT) );
  AND2X2 AND2X2_1237 ( .A(_abc_19068_n2809_bF_buf0), .B(_abc_19068_n2249), .Y(_abc_19068_n2906) );
  AND2X2 AND2X2_1238 ( .A(_abc_19068_n2907), .B(reset_n_bF_buf64), .Y(_abc_19068_n2908) );
  AND2X2 AND2X2_1239 ( .A(_abc_19068_n2908), .B(_abc_19068_n2905), .Y(key1_reg_19__FF_INPUT) );
  AND2X2 AND2X2_124 ( .A(_abc_19068_n885_1), .B(core_final_rounds_2_), .Y(_abc_19068_n1089_1) );
  AND2X2 AND2X2_1240 ( .A(_abc_19068_n2809_bF_buf6), .B(_abc_19068_n2255), .Y(_abc_19068_n2911) );
  AND2X2 AND2X2_1241 ( .A(_abc_19068_n2912), .B(reset_n_bF_buf63), .Y(_abc_19068_n2913) );
  AND2X2 AND2X2_1242 ( .A(_abc_19068_n2913), .B(_abc_19068_n2910), .Y(key1_reg_20__FF_INPUT) );
  AND2X2 AND2X2_1243 ( .A(_abc_19068_n2809_bF_buf4), .B(_abc_19068_n2261), .Y(_abc_19068_n2916) );
  AND2X2 AND2X2_1244 ( .A(_abc_19068_n2917), .B(reset_n_bF_buf62), .Y(_abc_19068_n2918) );
  AND2X2 AND2X2_1245 ( .A(_abc_19068_n2918), .B(_abc_19068_n2915), .Y(key1_reg_21__FF_INPUT) );
  AND2X2 AND2X2_1246 ( .A(_abc_19068_n2809_bF_buf2), .B(_abc_19068_n2267), .Y(_abc_19068_n2921) );
  AND2X2 AND2X2_1247 ( .A(_abc_19068_n2922), .B(reset_n_bF_buf61), .Y(_abc_19068_n2923) );
  AND2X2 AND2X2_1248 ( .A(_abc_19068_n2923), .B(_abc_19068_n2920), .Y(key1_reg_22__FF_INPUT) );
  AND2X2 AND2X2_1249 ( .A(_abc_19068_n2809_bF_buf0), .B(_abc_19068_n2273), .Y(_abc_19068_n2926) );
  AND2X2 AND2X2_125 ( .A(_abc_19068_n926_bF_buf3), .B(core_key_6_), .Y(_abc_19068_n1090_1) );
  AND2X2 AND2X2_1250 ( .A(_abc_19068_n2927), .B(reset_n_bF_buf60), .Y(_abc_19068_n2928) );
  AND2X2 AND2X2_1251 ( .A(_abc_19068_n2928), .B(_abc_19068_n2925), .Y(key1_reg_23__FF_INPUT) );
  AND2X2 AND2X2_1252 ( .A(_abc_19068_n2809_bF_buf6), .B(_abc_19068_n2279), .Y(_abc_19068_n2931) );
  AND2X2 AND2X2_1253 ( .A(_abc_19068_n2932), .B(reset_n_bF_buf59), .Y(_abc_19068_n2933) );
  AND2X2 AND2X2_1254 ( .A(_abc_19068_n2933), .B(_abc_19068_n2930), .Y(key1_reg_24__FF_INPUT) );
  AND2X2 AND2X2_1255 ( .A(_abc_19068_n2809_bF_buf4), .B(_abc_19068_n2285), .Y(_abc_19068_n2936) );
  AND2X2 AND2X2_1256 ( .A(_abc_19068_n2937), .B(reset_n_bF_buf58), .Y(_abc_19068_n2938) );
  AND2X2 AND2X2_1257 ( .A(_abc_19068_n2938), .B(_abc_19068_n2935), .Y(key1_reg_25__FF_INPUT) );
  AND2X2 AND2X2_1258 ( .A(_abc_19068_n2809_bF_buf2), .B(_abc_19068_n2291), .Y(_abc_19068_n2941) );
  AND2X2 AND2X2_1259 ( .A(_abc_19068_n2942), .B(reset_n_bF_buf57), .Y(_abc_19068_n2943) );
  AND2X2 AND2X2_126 ( .A(_abc_19068_n924_1_bF_buf3), .B(core_key_38_), .Y(_abc_19068_n1092_1) );
  AND2X2 AND2X2_1260 ( .A(_abc_19068_n2943), .B(_abc_19068_n2940), .Y(key1_reg_26__FF_INPUT) );
  AND2X2 AND2X2_1261 ( .A(_abc_19068_n2809_bF_buf0), .B(_abc_19068_n2297), .Y(_abc_19068_n2946) );
  AND2X2 AND2X2_1262 ( .A(_abc_19068_n2947), .B(reset_n_bF_buf56), .Y(_abc_19068_n2948) );
  AND2X2 AND2X2_1263 ( .A(_abc_19068_n2948), .B(_abc_19068_n2945), .Y(key1_reg_27__FF_INPUT) );
  AND2X2 AND2X2_1264 ( .A(_abc_19068_n2809_bF_buf6), .B(_abc_19068_n2303), .Y(_abc_19068_n2951) );
  AND2X2 AND2X2_1265 ( .A(_abc_19068_n2952), .B(reset_n_bF_buf55), .Y(_abc_19068_n2953) );
  AND2X2 AND2X2_1266 ( .A(_abc_19068_n2953), .B(_abc_19068_n2950), .Y(key1_reg_28__FF_INPUT) );
  AND2X2 AND2X2_1267 ( .A(_abc_19068_n2809_bF_buf4), .B(_abc_19068_n2309), .Y(_abc_19068_n2956) );
  AND2X2 AND2X2_1268 ( .A(_abc_19068_n2957), .B(reset_n_bF_buf54), .Y(_abc_19068_n2958) );
  AND2X2 AND2X2_1269 ( .A(_abc_19068_n2958), .B(_abc_19068_n2955), .Y(key1_reg_29__FF_INPUT) );
  AND2X2 AND2X2_127 ( .A(_abc_19068_n939_1_bF_buf3), .B(core_key_70_), .Y(_abc_19068_n1093_1) );
  AND2X2 AND2X2_1270 ( .A(_abc_19068_n2809_bF_buf2), .B(_abc_19068_n2315), .Y(_abc_19068_n2961) );
  AND2X2 AND2X2_1271 ( .A(_abc_19068_n2962), .B(reset_n_bF_buf53), .Y(_abc_19068_n2963) );
  AND2X2 AND2X2_1272 ( .A(_abc_19068_n2963), .B(_abc_19068_n2960), .Y(key1_reg_30__FF_INPUT) );
  AND2X2 AND2X2_1273 ( .A(_abc_19068_n2809_bF_buf0), .B(_abc_19068_n2321), .Y(_abc_19068_n2966) );
  AND2X2 AND2X2_1274 ( .A(_abc_19068_n2967), .B(reset_n_bF_buf52), .Y(_abc_19068_n2968) );
  AND2X2 AND2X2_1275 ( .A(_abc_19068_n2968), .B(_abc_19068_n2965), .Y(key1_reg_31__FF_INPUT) );
  AND2X2 AND2X2_1276 ( .A(_abc_19068_n926_bF_buf2), .B(_abc_19068_n2132), .Y(_abc_19068_n2970) );
  AND2X2 AND2X2_1277 ( .A(_abc_19068_n2970_bF_buf6), .B(_abc_19068_n2135), .Y(_abc_19068_n2972) );
  AND2X2 AND2X2_1278 ( .A(_abc_19068_n2973), .B(reset_n_bF_buf51), .Y(_abc_19068_n2974) );
  AND2X2 AND2X2_1279 ( .A(_abc_19068_n2974), .B(_abc_19068_n2971), .Y(key0_reg_0__FF_INPUT) );
  AND2X2 AND2X2_128 ( .A(_abc_19068_n923_bF_buf3), .B(_abc_19068_n1096_1), .Y(_auto_iopadmap_cc_313_execute_30317_6_) );
  AND2X2 AND2X2_1280 ( .A(_abc_19068_n2970_bF_buf4), .B(_abc_19068_n2141), .Y(_abc_19068_n2977) );
  AND2X2 AND2X2_1281 ( .A(_abc_19068_n2978), .B(reset_n_bF_buf50), .Y(_abc_19068_n2979) );
  AND2X2 AND2X2_1282 ( .A(_abc_19068_n2979), .B(_abc_19068_n2976), .Y(key0_reg_1__FF_INPUT) );
  AND2X2 AND2X2_1283 ( .A(_abc_19068_n2970_bF_buf2), .B(_abc_19068_n2147), .Y(_abc_19068_n2982) );
  AND2X2 AND2X2_1284 ( .A(_abc_19068_n2983), .B(reset_n_bF_buf49), .Y(_abc_19068_n2984) );
  AND2X2 AND2X2_1285 ( .A(_abc_19068_n2984), .B(_abc_19068_n2981), .Y(key0_reg_2__FF_INPUT) );
  AND2X2 AND2X2_1286 ( .A(_abc_19068_n2970_bF_buf0), .B(_abc_19068_n2153), .Y(_abc_19068_n2987) );
  AND2X2 AND2X2_1287 ( .A(_abc_19068_n2988), .B(reset_n_bF_buf48), .Y(_abc_19068_n2989) );
  AND2X2 AND2X2_1288 ( .A(_abc_19068_n2989), .B(_abc_19068_n2986), .Y(key0_reg_3__FF_INPUT) );
  AND2X2 AND2X2_1289 ( .A(_abc_19068_n2970_bF_buf6), .B(_abc_19068_n2159), .Y(_abc_19068_n2992) );
  AND2X2 AND2X2_129 ( .A(_abc_19068_n897_1_bF_buf1), .B(word0_reg_7_), .Y(_abc_19068_n1098_1) );
  AND2X2 AND2X2_1290 ( .A(_abc_19068_n2993), .B(reset_n_bF_buf47), .Y(_abc_19068_n2994) );
  AND2X2 AND2X2_1291 ( .A(_abc_19068_n2994), .B(_abc_19068_n2991), .Y(key0_reg_4__FF_INPUT) );
  AND2X2 AND2X2_1292 ( .A(_abc_19068_n2970_bF_buf4), .B(_abc_19068_n2165), .Y(_abc_19068_n2997) );
  AND2X2 AND2X2_1293 ( .A(_abc_19068_n2998), .B(reset_n_bF_buf46), .Y(_abc_19068_n2999) );
  AND2X2 AND2X2_1294 ( .A(_abc_19068_n2999), .B(_abc_19068_n2996), .Y(key0_reg_5__FF_INPUT) );
  AND2X2 AND2X2_1295 ( .A(_abc_19068_n2970_bF_buf2), .B(_abc_19068_n2171), .Y(_abc_19068_n3002) );
  AND2X2 AND2X2_1296 ( .A(_abc_19068_n3003), .B(reset_n_bF_buf45), .Y(_abc_19068_n3004) );
  AND2X2 AND2X2_1297 ( .A(_abc_19068_n3004), .B(_abc_19068_n3001), .Y(key0_reg_6__FF_INPUT) );
  AND2X2 AND2X2_1298 ( .A(_abc_19068_n2970_bF_buf0), .B(_abc_19068_n2177), .Y(_abc_19068_n3007) );
  AND2X2 AND2X2_1299 ( .A(_abc_19068_n3008), .B(reset_n_bF_buf44), .Y(_abc_19068_n3009) );
  AND2X2 AND2X2_13 ( .A(_abc_19068_n881), .B(_abc_19068_n888_1), .Y(_abc_19068_n889_1) );
  AND2X2 AND2X2_130 ( .A(_abc_19068_n916_1_bF_buf1), .B(word1_reg_7_), .Y(_abc_19068_n1099_1) );
  AND2X2 AND2X2_1300 ( .A(_abc_19068_n3009), .B(_abc_19068_n3006), .Y(key0_reg_7__FF_INPUT) );
  AND2X2 AND2X2_1301 ( .A(_abc_19068_n2970_bF_buf6), .B(_abc_19068_n2183), .Y(_abc_19068_n3012) );
  AND2X2 AND2X2_1302 ( .A(_abc_19068_n3013), .B(reset_n_bF_buf43), .Y(_abc_19068_n3014) );
  AND2X2 AND2X2_1303 ( .A(_abc_19068_n3014), .B(_abc_19068_n3011), .Y(key0_reg_8__FF_INPUT) );
  AND2X2 AND2X2_1304 ( .A(_abc_19068_n2970_bF_buf4), .B(_abc_19068_n2189), .Y(_abc_19068_n3017) );
  AND2X2 AND2X2_1305 ( .A(_abc_19068_n3018), .B(reset_n_bF_buf42), .Y(_abc_19068_n3019) );
  AND2X2 AND2X2_1306 ( .A(_abc_19068_n3019), .B(_abc_19068_n3016), .Y(key0_reg_9__FF_INPUT) );
  AND2X2 AND2X2_1307 ( .A(_abc_19068_n2970_bF_buf2), .B(_abc_19068_n2195), .Y(_abc_19068_n3022) );
  AND2X2 AND2X2_1308 ( .A(_abc_19068_n3023), .B(reset_n_bF_buf41), .Y(_abc_19068_n3024) );
  AND2X2 AND2X2_1309 ( .A(_abc_19068_n3024), .B(_abc_19068_n3021), .Y(key0_reg_10__FF_INPUT) );
  AND2X2 AND2X2_131 ( .A(_abc_19068_n915_1_bF_buf1), .B(core_mi_39_), .Y(_abc_19068_n1101_1) );
  AND2X2 AND2X2_1310 ( .A(_abc_19068_n2970_bF_buf0), .B(_abc_19068_n2201), .Y(_abc_19068_n3027) );
  AND2X2 AND2X2_1311 ( .A(_abc_19068_n3028), .B(reset_n_bF_buf40), .Y(_abc_19068_n3029) );
  AND2X2 AND2X2_1312 ( .A(_abc_19068_n3029), .B(_abc_19068_n3026), .Y(key0_reg_11__FF_INPUT) );
  AND2X2 AND2X2_1313 ( .A(_abc_19068_n2970_bF_buf6), .B(_abc_19068_n2207), .Y(_abc_19068_n3032) );
  AND2X2 AND2X2_1314 ( .A(_abc_19068_n3033), .B(reset_n_bF_buf39), .Y(_abc_19068_n3034) );
  AND2X2 AND2X2_1315 ( .A(_abc_19068_n3034), .B(_abc_19068_n3031), .Y(key0_reg_12__FF_INPUT) );
  AND2X2 AND2X2_1316 ( .A(_abc_19068_n2970_bF_buf4), .B(_abc_19068_n2213), .Y(_abc_19068_n3037) );
  AND2X2 AND2X2_1317 ( .A(_abc_19068_n3038), .B(reset_n_bF_buf38), .Y(_abc_19068_n3039) );
  AND2X2 AND2X2_1318 ( .A(_abc_19068_n3039), .B(_abc_19068_n3036), .Y(key0_reg_13__FF_INPUT) );
  AND2X2 AND2X2_1319 ( .A(_abc_19068_n2970_bF_buf2), .B(_abc_19068_n2219), .Y(_abc_19068_n3042) );
  AND2X2 AND2X2_132 ( .A(_abc_19068_n945_1_bF_buf2), .B(core_mi_7_), .Y(_abc_19068_n1102_1) );
  AND2X2 AND2X2_1320 ( .A(_abc_19068_n3043), .B(reset_n_bF_buf37), .Y(_abc_19068_n3044) );
  AND2X2 AND2X2_1321 ( .A(_abc_19068_n3044), .B(_abc_19068_n3041), .Y(key0_reg_14__FF_INPUT) );
  AND2X2 AND2X2_1322 ( .A(_abc_19068_n2970_bF_buf0), .B(_abc_19068_n2225), .Y(_abc_19068_n3047) );
  AND2X2 AND2X2_1323 ( .A(_abc_19068_n3048), .B(reset_n_bF_buf36), .Y(_abc_19068_n3049) );
  AND2X2 AND2X2_1324 ( .A(_abc_19068_n3049), .B(_abc_19068_n3046), .Y(key0_reg_15__FF_INPUT) );
  AND2X2 AND2X2_1325 ( .A(_abc_19068_n2970_bF_buf6), .B(_abc_19068_n2231), .Y(_abc_19068_n3052) );
  AND2X2 AND2X2_1326 ( .A(_abc_19068_n3053), .B(reset_n_bF_buf35), .Y(_abc_19068_n3054) );
  AND2X2 AND2X2_1327 ( .A(_abc_19068_n3054), .B(_abc_19068_n3051), .Y(key0_reg_16__FF_INPUT) );
  AND2X2 AND2X2_1328 ( .A(_abc_19068_n2970_bF_buf4), .B(_abc_19068_n2237), .Y(_abc_19068_n3057) );
  AND2X2 AND2X2_1329 ( .A(_abc_19068_n3058), .B(reset_n_bF_buf34), .Y(_abc_19068_n3059) );
  AND2X2 AND2X2_133 ( .A(_abc_19068_n924_1_bF_buf2), .B(core_key_39_), .Y(_abc_19068_n1105_1) );
  AND2X2 AND2X2_1330 ( .A(_abc_19068_n3059), .B(_abc_19068_n3056), .Y(key0_reg_17__FF_INPUT) );
  AND2X2 AND2X2_1331 ( .A(_abc_19068_n2970_bF_buf2), .B(_abc_19068_n2243), .Y(_abc_19068_n3062) );
  AND2X2 AND2X2_1332 ( .A(_abc_19068_n3063), .B(reset_n_bF_buf33), .Y(_abc_19068_n3064) );
  AND2X2 AND2X2_1333 ( .A(_abc_19068_n3064), .B(_abc_19068_n3061), .Y(key0_reg_18__FF_INPUT) );
  AND2X2 AND2X2_1334 ( .A(_abc_19068_n2970_bF_buf0), .B(_abc_19068_n2249), .Y(_abc_19068_n3067) );
  AND2X2 AND2X2_1335 ( .A(_abc_19068_n3068), .B(reset_n_bF_buf32), .Y(_abc_19068_n3069) );
  AND2X2 AND2X2_1336 ( .A(_abc_19068_n3069), .B(_abc_19068_n3066), .Y(key0_reg_19__FF_INPUT) );
  AND2X2 AND2X2_1337 ( .A(_abc_19068_n2970_bF_buf6), .B(_abc_19068_n2255), .Y(_abc_19068_n3072) );
  AND2X2 AND2X2_1338 ( .A(_abc_19068_n3073), .B(reset_n_bF_buf31), .Y(_abc_19068_n3074) );
  AND2X2 AND2X2_1339 ( .A(_abc_19068_n3074), .B(_abc_19068_n3071), .Y(key0_reg_20__FF_INPUT) );
  AND2X2 AND2X2_134 ( .A(_abc_19068_n885_1), .B(core_final_rounds_3_), .Y(_abc_19068_n1106) );
  AND2X2 AND2X2_1340 ( .A(_abc_19068_n2970_bF_buf4), .B(_abc_19068_n2261), .Y(_abc_19068_n3077) );
  AND2X2 AND2X2_1341 ( .A(_abc_19068_n3078), .B(reset_n_bF_buf30), .Y(_abc_19068_n3079) );
  AND2X2 AND2X2_1342 ( .A(_abc_19068_n3079), .B(_abc_19068_n3076), .Y(key0_reg_21__FF_INPUT) );
  AND2X2 AND2X2_1343 ( .A(_abc_19068_n2970_bF_buf2), .B(_abc_19068_n2267), .Y(_abc_19068_n3082) );
  AND2X2 AND2X2_1344 ( .A(_abc_19068_n3083), .B(reset_n_bF_buf29), .Y(_abc_19068_n3084) );
  AND2X2 AND2X2_1345 ( .A(_abc_19068_n3084), .B(_abc_19068_n3081), .Y(key0_reg_22__FF_INPUT) );
  AND2X2 AND2X2_1346 ( .A(_abc_19068_n2970_bF_buf0), .B(_abc_19068_n2273), .Y(_abc_19068_n3087) );
  AND2X2 AND2X2_1347 ( .A(_abc_19068_n3088), .B(reset_n_bF_buf28), .Y(_abc_19068_n3089) );
  AND2X2 AND2X2_1348 ( .A(_abc_19068_n3089), .B(_abc_19068_n3086), .Y(key0_reg_23__FF_INPUT) );
  AND2X2 AND2X2_1349 ( .A(_abc_19068_n2970_bF_buf6), .B(_abc_19068_n2279), .Y(_abc_19068_n3092) );
  AND2X2 AND2X2_135 ( .A(_abc_19068_n926_bF_buf2), .B(core_key_7_), .Y(_abc_19068_n1107_1) );
  AND2X2 AND2X2_1350 ( .A(_abc_19068_n3093), .B(reset_n_bF_buf27), .Y(_abc_19068_n3094) );
  AND2X2 AND2X2_1351 ( .A(_abc_19068_n3094), .B(_abc_19068_n3091), .Y(key0_reg_24__FF_INPUT) );
  AND2X2 AND2X2_1352 ( .A(_abc_19068_n2970_bF_buf4), .B(_abc_19068_n2285), .Y(_abc_19068_n3097) );
  AND2X2 AND2X2_1353 ( .A(_abc_19068_n3098), .B(reset_n_bF_buf26), .Y(_abc_19068_n3099) );
  AND2X2 AND2X2_1354 ( .A(_abc_19068_n3099), .B(_abc_19068_n3096), .Y(key0_reg_25__FF_INPUT) );
  AND2X2 AND2X2_1355 ( .A(_abc_19068_n2970_bF_buf2), .B(_abc_19068_n2291), .Y(_abc_19068_n3102) );
  AND2X2 AND2X2_1356 ( .A(_abc_19068_n3103), .B(reset_n_bF_buf25), .Y(_abc_19068_n3104) );
  AND2X2 AND2X2_1357 ( .A(_abc_19068_n3104), .B(_abc_19068_n3101), .Y(key0_reg_26__FF_INPUT) );
  AND2X2 AND2X2_1358 ( .A(_abc_19068_n2970_bF_buf0), .B(_abc_19068_n2297), .Y(_abc_19068_n3107) );
  AND2X2 AND2X2_1359 ( .A(_abc_19068_n3108), .B(reset_n_bF_buf24), .Y(_abc_19068_n3109) );
  AND2X2 AND2X2_136 ( .A(_abc_19068_n899_bF_buf1), .B(word3_reg_7_), .Y(_abc_19068_n1110_1) );
  AND2X2 AND2X2_1360 ( .A(_abc_19068_n3109), .B(_abc_19068_n3106), .Y(key0_reg_27__FF_INPUT) );
  AND2X2 AND2X2_1361 ( .A(_abc_19068_n2970_bF_buf6), .B(_abc_19068_n2303), .Y(_abc_19068_n3112) );
  AND2X2 AND2X2_1362 ( .A(_abc_19068_n3113), .B(reset_n_bF_buf23), .Y(_abc_19068_n3114) );
  AND2X2 AND2X2_1363 ( .A(_abc_19068_n3114), .B(_abc_19068_n3111), .Y(key0_reg_28__FF_INPUT) );
  AND2X2 AND2X2_1364 ( .A(_abc_19068_n2970_bF_buf4), .B(_abc_19068_n2309), .Y(_abc_19068_n3117) );
  AND2X2 AND2X2_1365 ( .A(_abc_19068_n3118), .B(reset_n_bF_buf22), .Y(_abc_19068_n3119) );
  AND2X2 AND2X2_1366 ( .A(_abc_19068_n3119), .B(_abc_19068_n3116), .Y(key0_reg_29__FF_INPUT) );
  AND2X2 AND2X2_1367 ( .A(_abc_19068_n2970_bF_buf2), .B(_abc_19068_n2315), .Y(_abc_19068_n3122) );
  AND2X2 AND2X2_1368 ( .A(_abc_19068_n3123), .B(reset_n_bF_buf21), .Y(_abc_19068_n3124) );
  AND2X2 AND2X2_1369 ( .A(_abc_19068_n3124), .B(_abc_19068_n3121), .Y(key0_reg_30__FF_INPUT) );
  AND2X2 AND2X2_137 ( .A(_abc_19068_n902_bF_buf1), .B(word2_reg_7_), .Y(_abc_19068_n1111_1) );
  AND2X2 AND2X2_1370 ( .A(_abc_19068_n2970_bF_buf0), .B(_abc_19068_n2321), .Y(_abc_19068_n3127) );
  AND2X2 AND2X2_1371 ( .A(_abc_19068_n3128), .B(reset_n_bF_buf20), .Y(_abc_19068_n3129) );
  AND2X2 AND2X2_1372 ( .A(_abc_19068_n3129), .B(_abc_19068_n3126), .Y(key0_reg_31__FF_INPUT) );
  AND2X2 AND2X2_1373 ( .A(_abc_19068_n885_1), .B(_abc_19068_n2132), .Y(_abc_19068_n3131) );
  AND2X2 AND2X2_1374 ( .A(_abc_19068_n3131), .B(\write_data[0] ), .Y(_abc_19068_n3132) );
  AND2X2 AND2X2_1375 ( .A(_abc_19068_n3133), .B(core_compression_rounds_0_), .Y(_abc_19068_n3134) );
  AND2X2 AND2X2_1376 ( .A(_abc_19068_n3135), .B(reset_n_bF_buf19), .Y(param_reg_0__FF_INPUT) );
  AND2X2 AND2X2_1377 ( .A(_abc_19068_n3133), .B(core_compression_rounds_1_), .Y(_abc_19068_n3137) );
  AND2X2 AND2X2_1378 ( .A(_abc_19068_n3131), .B(\write_data[1] ), .Y(_abc_19068_n3139) );
  AND2X2 AND2X2_1379 ( .A(_abc_19068_n3131), .B(\write_data[2] ), .Y(_abc_19068_n3142) );
  AND2X2 AND2X2_138 ( .A(_abc_19068_n941_bF_buf2), .B(core_key_103_), .Y(_abc_19068_n1113_1) );
  AND2X2 AND2X2_1380 ( .A(_abc_19068_n3133), .B(core_compression_rounds_2_), .Y(_abc_19068_n3143) );
  AND2X2 AND2X2_1381 ( .A(_abc_19068_n3144), .B(reset_n_bF_buf17), .Y(param_reg_2__FF_INPUT) );
  AND2X2 AND2X2_1382 ( .A(_abc_19068_n3131), .B(\write_data[3] ), .Y(_abc_19068_n3146) );
  AND2X2 AND2X2_1383 ( .A(_abc_19068_n3133), .B(core_compression_rounds_3_), .Y(_abc_19068_n3147) );
  AND2X2 AND2X2_1384 ( .A(_abc_19068_n3148), .B(reset_n_bF_buf16), .Y(param_reg_3__FF_INPUT) );
  AND2X2 AND2X2_1385 ( .A(_abc_19068_n3131), .B(\write_data[4] ), .Y(_abc_19068_n3150) );
  AND2X2 AND2X2_1386 ( .A(_abc_19068_n3133), .B(core_final_rounds_0_), .Y(_abc_19068_n3151) );
  AND2X2 AND2X2_1387 ( .A(_abc_19068_n3152), .B(reset_n_bF_buf15), .Y(param_reg_4__FF_INPUT) );
  AND2X2 AND2X2_1388 ( .A(_abc_19068_n3131), .B(\write_data[5] ), .Y(_abc_19068_n3154) );
  AND2X2 AND2X2_1389 ( .A(_abc_19068_n3133), .B(core_final_rounds_1_), .Y(_abc_19068_n3155) );
  AND2X2 AND2X2_139 ( .A(_abc_19068_n939_1_bF_buf2), .B(core_key_71_), .Y(_abc_19068_n1114_1) );
  AND2X2 AND2X2_1390 ( .A(_abc_19068_n3156), .B(reset_n_bF_buf14), .Y(param_reg_5__FF_INPUT) );
  AND2X2 AND2X2_1391 ( .A(_abc_19068_n3133), .B(core_final_rounds_2_), .Y(_abc_19068_n3158) );
  AND2X2 AND2X2_1392 ( .A(_abc_19068_n3131), .B(\write_data[6] ), .Y(_abc_19068_n3159) );
  AND2X2 AND2X2_1393 ( .A(_abc_19068_n3131), .B(\write_data[7] ), .Y(_abc_19068_n3162) );
  AND2X2 AND2X2_1394 ( .A(_abc_19068_n3133), .B(core_final_rounds_3_), .Y(_abc_19068_n3163) );
  AND2X2 AND2X2_1395 ( .A(_abc_19068_n3164), .B(reset_n_bF_buf13), .Y(param_reg_7__FF_INPUT) );
  AND2X2 AND2X2_1396 ( .A(_abc_19068_n2132), .B(reset_n_bF_buf12), .Y(_abc_19068_n3166) );
  AND2X2 AND2X2_1397 ( .A(_abc_19068_n3166), .B(\write_data[0] ), .Y(_abc_19068_n3167) );
  AND2X2 AND2X2_1398 ( .A(_abc_19068_n889_1), .B(_abc_19068_n3167), .Y(ctrl_reg_0__FF_INPUT) );
  AND2X2 AND2X2_1399 ( .A(_abc_19068_n3166), .B(\write_data[1] ), .Y(_abc_19068_n3169) );
  AND2X2 AND2X2_14 ( .A(_abc_19068_n892_1), .B(_abc_19068_n870_1), .Y(_abc_19068_n893) );
  AND2X2 AND2X2_140 ( .A(_abc_19068_n923_bF_buf2), .B(_abc_19068_n1118), .Y(_auto_iopadmap_cc_313_execute_30317_7_) );
  AND2X2 AND2X2_1400 ( .A(_abc_19068_n889_1), .B(_abc_19068_n3169), .Y(ctrl_reg_1__FF_INPUT) );
  AND2X2 AND2X2_1401 ( .A(_abc_19068_n3166), .B(\write_data[2] ), .Y(_abc_19068_n3171) );
  AND2X2 AND2X2_1402 ( .A(_abc_19068_n889_1), .B(_abc_19068_n3171), .Y(ctrl_reg_2__FF_INPUT) );
  AND2X2 AND2X2_1403 ( .A(_abc_19068_n900_1), .B(_abc_19068_n2132), .Y(_abc_19068_n3173) );
  AND2X2 AND2X2_1404 ( .A(_abc_19068_n3173), .B(_abc_19068_n871_1), .Y(_abc_19068_n3174) );
  AND2X2 AND2X2_1405 ( .A(_abc_19068_n3174), .B(_abc_19068_n881), .Y(_abc_19068_n3175) );
  AND2X2 AND2X2_1406 ( .A(_abc_19068_n3175), .B(_abc_19068_n2135), .Y(_abc_19068_n3176) );
  AND2X2 AND2X2_1407 ( .A(_abc_19068_n3178), .B(reset_n_bF_buf11), .Y(_abc_19068_n3179) );
  AND2X2 AND2X2_1408 ( .A(_abc_19068_n3179), .B(_abc_19068_n3177), .Y(long_reg_FF_INPUT) );
  AND2X2 AND2X2_1409 ( .A(core__abc_21380_n1130_1), .B(core__abc_21380_n1131), .Y(core__abc_21380_n1132_1) );
  AND2X2 AND2X2_141 ( .A(_abc_19068_n916_1_bF_buf0), .B(word1_reg_8_), .Y(_abc_19068_n1120_1) );
  AND2X2 AND2X2_1410 ( .A(core__abc_21380_n1133_1), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n1135) );
  AND2X2 AND2X2_1411 ( .A(core__abc_21380_n1136_1), .B(core__abc_21380_n1137_1), .Y(core__abc_21380_n1138_1) );
  AND2X2 AND2X2_1412 ( .A(core__abc_21380_n1135), .B(core__abc_21380_n1138_1), .Y(core__abc_21380_n1139) );
  AND2X2 AND2X2_1413 ( .A(core__abc_21380_n1142_1), .B(core__abc_21380_n1139), .Y(core__abc_21380_n1143) );
  AND2X2 AND2X2_1414 ( .A(core__abc_21380_n1145_1), .B(core__abc_21380_n1144_1), .Y(core__abc_21380_n1146_1) );
  AND2X2 AND2X2_1415 ( .A(core__abc_21380_n1143), .B(core__abc_21380_n1146_1), .Y(core__abc_21380_n1147) );
  AND2X2 AND2X2_1416 ( .A(core__abc_21380_n1150_1), .B(core__abc_21380_n1151), .Y(core__abc_21380_n1152_1) );
  AND2X2 AND2X2_1417 ( .A(core__abc_21380_n1152_1), .B(core__abc_21380_n1149_1), .Y(core__abc_21380_n1153_1) );
  AND2X2 AND2X2_1418 ( .A(core__abc_21380_n1153_1), .B(core__abc_21380_n1148_1), .Y(core__abc_21380_n1154_1) );
  AND2X2 AND2X2_1419 ( .A(core__abc_21380_n1156_1), .B(core__abc_21380_n1158_1), .Y(core__abc_21380_n1159) );
  AND2X2 AND2X2_142 ( .A(_abc_19068_n897_1_bF_buf0), .B(word0_reg_8_), .Y(_abc_19068_n1121) );
  AND2X2 AND2X2_1420 ( .A(core__abc_21380_n1160_1), .B(core__abc_21380_n1155), .Y(core__abc_21380_n1161_1) );
  AND2X2 AND2X2_1421 ( .A(core_compression_rounds_0_), .B(core_loop_ctr_reg_0_), .Y(core__abc_21380_n1163) );
  AND2X2 AND2X2_1422 ( .A(core__abc_21380_n1159), .B(core__abc_21380_n1151), .Y(core__abc_21380_n1164_1) );
  AND2X2 AND2X2_1423 ( .A(core__abc_21380_n1168_1), .B(core__abc_21380_n1169_1), .Y(core__abc_21380_n1170_1) );
  AND2X2 AND2X2_1424 ( .A(core__abc_21380_n1170_1), .B(core_loop_ctr_reg_2_), .Y(core__abc_21380_n1171) );
  AND2X2 AND2X2_1425 ( .A(core__abc_21380_n1172_1), .B(core__abc_21380_n1173_1), .Y(core__abc_21380_n1174_1) );
  AND2X2 AND2X2_1426 ( .A(core__abc_21380_n1167), .B(core__abc_21380_n1174_1), .Y(core__abc_21380_n1175) );
  AND2X2 AND2X2_1427 ( .A(core__abc_21380_n1168_1), .B(core_compression_rounds_3_), .Y(core__abc_21380_n1176_1) );
  AND2X2 AND2X2_1428 ( .A(core__abc_21380_n1178_1), .B(core_loop_ctr_reg_3_), .Y(core__abc_21380_n1179) );
  AND2X2 AND2X2_1429 ( .A(core__abc_21380_n1177_1), .B(core__abc_21380_n1180_1), .Y(core__abc_21380_n1181_1) );
  AND2X2 AND2X2_143 ( .A(_abc_19068_n939_1_bF_buf1), .B(core_key_72_), .Y(_abc_19068_n1123_1) );
  AND2X2 AND2X2_1430 ( .A(core__abc_21380_n1183), .B(core__abc_21380_n1175), .Y(core__abc_21380_n1184_1) );
  AND2X2 AND2X2_1431 ( .A(core__abc_21380_n1184_1), .B(core_siphash_ctrl_reg_4_), .Y(core__abc_21380_n1185_1) );
  AND2X2 AND2X2_1432 ( .A(core__abc_21380_n1188_1), .B(core__abc_21380_n1189_1), .Y(core__abc_21380_n1190_1) );
  AND2X2 AND2X2_1433 ( .A(core__abc_21380_n1190_1), .B(core__abc_21380_n1187), .Y(core__abc_21380_n1191) );
  AND2X2 AND2X2_1434 ( .A(core__abc_21380_n1191), .B(core__abc_21380_n1186_1), .Y(core__abc_21380_n1192_1) );
  AND2X2 AND2X2_1435 ( .A(core_loop_ctr_reg_0_), .B(core_final_rounds_0_), .Y(core__abc_21380_n1193_1) );
  AND2X2 AND2X2_1436 ( .A(core__abc_21380_n1195), .B(core__abc_21380_n1196_1), .Y(core__abc_21380_n1197_1) );
  AND2X2 AND2X2_1437 ( .A(core__abc_21380_n1198_1), .B(core__abc_21380_n1155), .Y(core__abc_21380_n1199) );
  AND2X2 AND2X2_1438 ( .A(core__abc_21380_n1197_1), .B(core__abc_21380_n1189_1), .Y(core__abc_21380_n1200_1) );
  AND2X2 AND2X2_1439 ( .A(core__abc_21380_n1205_1), .B(core__abc_21380_n1206_1), .Y(core__abc_21380_n1207) );
  AND2X2 AND2X2_144 ( .A(_abc_19068_n924_1_bF_buf1), .B(core_key_40_), .Y(_abc_19068_n1124) );
  AND2X2 AND2X2_1440 ( .A(core__abc_21380_n1209_1), .B(core__abc_21380_n1210_1), .Y(core__abc_21380_n1211) );
  AND2X2 AND2X2_1441 ( .A(core__abc_21380_n1203), .B(core__abc_21380_n1211), .Y(core__abc_21380_n1212_1) );
  AND2X2 AND2X2_1442 ( .A(core__abc_21380_n1205_1), .B(core_final_rounds_3_), .Y(core__abc_21380_n1213_1) );
  AND2X2 AND2X2_1443 ( .A(core__abc_21380_n1215), .B(core_loop_ctr_reg_3_), .Y(core__abc_21380_n1216_1) );
  AND2X2 AND2X2_1444 ( .A(core__abc_21380_n1214_1), .B(core__abc_21380_n1180_1), .Y(core__abc_21380_n1217_1) );
  AND2X2 AND2X2_1445 ( .A(core__abc_21380_n1219), .B(core__abc_21380_n1212_1), .Y(core__abc_21380_n1220_1) );
  AND2X2 AND2X2_1446 ( .A(core__abc_21380_n1220_1), .B(core__abc_21380_n1140_1), .Y(core__abc_21380_n1221_1) );
  AND2X2 AND2X2_1447 ( .A(core__abc_21380_n1225_1), .B(reset_n_bF_buf10), .Y(core__abc_21380_n1226_1) );
  AND2X2 AND2X2_1448 ( .A(core__abc_21380_n1144_1), .B(core_siphash_ctrl_reg_0_), .Y(core__abc_21380_n1227) );
  AND2X2 AND2X2_1449 ( .A(core__abc_21380_n1226_1), .B(core__abc_21380_n1227), .Y(core__abc_21380_n1228_1) );
  AND2X2 AND2X2_145 ( .A(_abc_19068_n926_bF_buf1), .B(core_key_8_), .Y(_abc_19068_n1125_1) );
  AND2X2 AND2X2_1450 ( .A(core__abc_21380_n1228_1), .B(core__abc_21380_n1132_1), .Y(core__abc_21380_n1229_1) );
  AND2X2 AND2X2_1451 ( .A(core__abc_21380_n1230_1), .B(core__abc_21380_n1140_1), .Y(core__abc_21380_n1231) );
  AND2X2 AND2X2_1452 ( .A(core__abc_21380_n1232_1), .B(core_siphash_ctrl_reg_4_), .Y(core__abc_21380_n1233_1) );
  AND2X2 AND2X2_1453 ( .A(core_initalize), .B(core_siphash_ctrl_reg_0_), .Y(core__abc_21380_n1234_1) );
  AND2X2 AND2X2_1454 ( .A(core__abc_21380_n1226_1), .B(core__abc_21380_n1236_1), .Y(core__abc_21380_n1237_1) );
  AND2X2 AND2X2_1455 ( .A(core__abc_21380_n1238_1), .B(reset_n_bF_buf9), .Y(core__abc_21380_n1239) );
  AND2X2 AND2X2_1456 ( .A(core__abc_21380_n1239), .B(core_siphash_ctrl_reg_0_), .Y(core__abc_21380_n1240_1) );
  AND2X2 AND2X2_1457 ( .A(core_siphash_ctrl_reg_5_), .B(reset_n_bF_buf7), .Y(core__abc_21380_n1248_1) );
  AND2X2 AND2X2_1458 ( .A(core_siphash_ctrl_reg_3_), .B(reset_n_bF_buf6), .Y(core__abc_21380_n1249_1) );
  AND2X2 AND2X2_1459 ( .A(core__abc_21380_n1238_1), .B(core__abc_21380_n1249_1), .Y(core__abc_21380_n1250_1) );
  AND2X2 AND2X2_146 ( .A(_abc_19068_n941_bF_buf1), .B(core_key_104_), .Y(_abc_19068_n1129_1) );
  AND2X2 AND2X2_1460 ( .A(core__abc_21380_n1239), .B(core_siphash_ctrl_reg_4_), .Y(core__abc_21380_n1252_1) );
  AND2X2 AND2X2_1461 ( .A(core__abc_21380_n1228_1), .B(core_compress), .Y(core__abc_21380_n1253_1) );
  AND2X2 AND2X2_1462 ( .A(core__abc_21380_n1131), .B(core_finalize), .Y(core__abc_21380_n1255) );
  AND2X2 AND2X2_1463 ( .A(core__abc_21380_n1228_1), .B(core__abc_21380_n1255), .Y(core__abc_21380_n1256_1) );
  AND2X2 AND2X2_1464 ( .A(core__abc_21380_n1239), .B(core_siphash_ctrl_reg_6_), .Y(core__abc_21380_n1257_1) );
  AND2X2 AND2X2_1465 ( .A(core_v0_reg_0_), .B(core_v1_reg_0_), .Y(core__abc_21380_n1260_1) );
  AND2X2 AND2X2_1466 ( .A(core__abc_21380_n1261_1), .B(core__abc_21380_n1259), .Y(core__abc_21380_n1262_1) );
  AND2X2 AND2X2_1467 ( .A(core__abc_21380_n1263), .B(core__abc_21380_n1264_1), .Y(core__abc_21380_n1265_1) );
  AND2X2 AND2X2_1468 ( .A(core_v3_reg_0_), .B(core_v2_reg_0_), .Y(core__abc_21380_n1266_1) );
  AND2X2 AND2X2_1469 ( .A(core__abc_21380_n1269_1), .B(core__abc_21380_n1271), .Y(core__abc_21380_n1272_1) );
  AND2X2 AND2X2_147 ( .A(_abc_19068_n902_bF_buf0), .B(word2_reg_8_), .Y(_abc_19068_n1130) );
  AND2X2 AND2X2_1470 ( .A(core__abc_21380_n1274_1), .B(reset_n_bF_buf5), .Y(core__abc_21380_n1275) );
  AND2X2 AND2X2_1471 ( .A(core__abc_21380_n1273_1), .B(core__abc_21380_n1275), .Y(core_siphash_word1_reg_0__FF_INPUT) );
  AND2X2 AND2X2_1472 ( .A(core_v0_reg_1_), .B(core_v1_reg_1_), .Y(core__abc_21380_n1278_1) );
  AND2X2 AND2X2_1473 ( .A(core__abc_21380_n1279), .B(core__abc_21380_n1277_1), .Y(core__abc_21380_n1280_1) );
  AND2X2 AND2X2_1474 ( .A(core_v3_reg_1_), .B(core_v2_reg_1_), .Y(core__abc_21380_n1281_1) );
  AND2X2 AND2X2_1475 ( .A(core__abc_21380_n1282_1), .B(core__abc_21380_n1283), .Y(core__abc_21380_n1284_1) );
  AND2X2 AND2X2_1476 ( .A(core__abc_21380_n1288_1), .B(core__abc_21380_n1289), .Y(core__abc_21380_n1290) );
  AND2X2 AND2X2_1477 ( .A(core__abc_21380_n1287), .B(core__abc_21380_n1292), .Y(core__abc_21380_n1293) );
  AND2X2 AND2X2_1478 ( .A(core__abc_21380_n1295), .B(reset_n_bF_buf4), .Y(core__abc_21380_n1296) );
  AND2X2 AND2X2_1479 ( .A(core__abc_21380_n1294), .B(core__abc_21380_n1296), .Y(core_siphash_word1_reg_1__FF_INPUT) );
  AND2X2 AND2X2_148 ( .A(_abc_19068_n899_bF_buf0), .B(word3_reg_8_), .Y(_abc_19068_n1131_1) );
  AND2X2 AND2X2_1480 ( .A(core__abc_21380_n1298), .B(core__abc_21380_n1299), .Y(core__abc_21380_n1300) );
  AND2X2 AND2X2_1481 ( .A(core_v0_reg_2_), .B(core_v1_reg_2_), .Y(core__abc_21380_n1301) );
  AND2X2 AND2X2_1482 ( .A(core_v3_reg_2_), .B(core_v2_reg_2_), .Y(core__abc_21380_n1304) );
  AND2X2 AND2X2_1483 ( .A(core__abc_21380_n1305), .B(core__abc_21380_n1306), .Y(core__abc_21380_n1307) );
  AND2X2 AND2X2_1484 ( .A(core__abc_21380_n1310), .B(core__abc_21380_n1311), .Y(core__abc_21380_n1312) );
  AND2X2 AND2X2_1485 ( .A(core__abc_21380_n1314), .B(reset_n_bF_buf3), .Y(core__abc_21380_n1315) );
  AND2X2 AND2X2_1486 ( .A(core__abc_21380_n1313), .B(core__abc_21380_n1315), .Y(core_siphash_word1_reg_2__FF_INPUT) );
  AND2X2 AND2X2_1487 ( .A(core_v0_reg_3_), .B(core_v1_reg_3_), .Y(core__abc_21380_n1317) );
  AND2X2 AND2X2_1488 ( .A(core__abc_21380_n1318), .B(core__abc_21380_n1319), .Y(core__abc_21380_n1320) );
  AND2X2 AND2X2_1489 ( .A(core_v2_reg_3_), .B(core_v3_reg_3_), .Y(core__abc_21380_n1323) );
  AND2X2 AND2X2_149 ( .A(_abc_19068_n945_1_bF_buf1), .B(core_mi_8_), .Y(_abc_19068_n1133) );
  AND2X2 AND2X2_1490 ( .A(core__abc_21380_n1324), .B(core__abc_21380_n1325), .Y(core__abc_21380_n1326) );
  AND2X2 AND2X2_1491 ( .A(core__abc_21380_n1322), .B(core__abc_21380_n1327), .Y(core__abc_21380_n1328) );
  AND2X2 AND2X2_1492 ( .A(core__abc_21380_n1329), .B(core__abc_21380_n1321), .Y(core__abc_21380_n1330) );
  AND2X2 AND2X2_1493 ( .A(core__abc_21380_n1333), .B(reset_n_bF_buf2), .Y(core__abc_21380_n1334) );
  AND2X2 AND2X2_1494 ( .A(core__abc_21380_n1332), .B(core__abc_21380_n1334), .Y(core_siphash_word1_reg_3__FF_INPUT) );
  AND2X2 AND2X2_1495 ( .A(core_v0_reg_4_), .B(core_v1_reg_4_), .Y(core__abc_21380_n1337) );
  AND2X2 AND2X2_1496 ( .A(core__abc_21380_n1338), .B(core__abc_21380_n1336), .Y(core__abc_21380_n1339) );
  AND2X2 AND2X2_1497 ( .A(core_v3_reg_4_), .B(core_v2_reg_4_), .Y(core__abc_21380_n1340) );
  AND2X2 AND2X2_1498 ( .A(core__abc_21380_n1341), .B(core__abc_21380_n1342), .Y(core__abc_21380_n1343) );
  AND2X2 AND2X2_1499 ( .A(core__abc_21380_n1346), .B(core__abc_21380_n1348), .Y(core__abc_21380_n1349) );
  AND2X2 AND2X2_15 ( .A(_abc_19068_n893), .B(_abc_19068_n887), .Y(_abc_19068_n894_1) );
  AND2X2 AND2X2_150 ( .A(_abc_19068_n915_1_bF_buf0), .B(core_mi_40_), .Y(_abc_19068_n1134_1) );
  AND2X2 AND2X2_1500 ( .A(core__abc_21380_n1351), .B(reset_n_bF_buf1), .Y(core__abc_21380_n1352) );
  AND2X2 AND2X2_1501 ( .A(core__abc_21380_n1350), .B(core__abc_21380_n1352), .Y(core_siphash_word1_reg_4__FF_INPUT) );
  AND2X2 AND2X2_1502 ( .A(core_v0_reg_5_), .B(core_v1_reg_5_), .Y(core__abc_21380_n1354) );
  AND2X2 AND2X2_1503 ( .A(core__abc_21380_n1355), .B(core__abc_21380_n1356), .Y(core__abc_21380_n1357) );
  AND2X2 AND2X2_1504 ( .A(core_v2_reg_5_), .B(core_v3_reg_5_), .Y(core__abc_21380_n1360) );
  AND2X2 AND2X2_1505 ( .A(core__abc_21380_n1361), .B(core__abc_21380_n1362), .Y(core__abc_21380_n1363) );
  AND2X2 AND2X2_1506 ( .A(core__abc_21380_n1359), .B(core__abc_21380_n1364), .Y(core__abc_21380_n1365) );
  AND2X2 AND2X2_1507 ( .A(core__abc_21380_n1366), .B(core__abc_21380_n1358), .Y(core__abc_21380_n1367) );
  AND2X2 AND2X2_1508 ( .A(core__abc_21380_n1370), .B(reset_n_bF_buf0), .Y(core__abc_21380_n1371) );
  AND2X2 AND2X2_1509 ( .A(core__abc_21380_n1369), .B(core__abc_21380_n1371), .Y(core_siphash_word1_reg_5__FF_INPUT) );
  AND2X2 AND2X2_151 ( .A(_abc_19068_n923_bF_buf1), .B(_abc_19068_n1138), .Y(_auto_iopadmap_cc_313_execute_30317_8_) );
  AND2X2 AND2X2_1510 ( .A(core__abc_21380_n1373), .B(core__abc_21380_n1374), .Y(core__abc_21380_n1375) );
  AND2X2 AND2X2_1511 ( .A(core_v0_reg_6_), .B(core_v1_reg_6_), .Y(core__abc_21380_n1376) );
  AND2X2 AND2X2_1512 ( .A(core_v3_reg_6_), .B(core_v2_reg_6_), .Y(core__abc_21380_n1379) );
  AND2X2 AND2X2_1513 ( .A(core__abc_21380_n1380), .B(core__abc_21380_n1381), .Y(core__abc_21380_n1382) );
  AND2X2 AND2X2_1514 ( .A(core__abc_21380_n1385), .B(core__abc_21380_n1386), .Y(core__abc_21380_n1387) );
  AND2X2 AND2X2_1515 ( .A(core__abc_21380_n1389), .B(reset_n_bF_buf84), .Y(core__abc_21380_n1390) );
  AND2X2 AND2X2_1516 ( .A(core__abc_21380_n1388), .B(core__abc_21380_n1390), .Y(core_siphash_word1_reg_6__FF_INPUT) );
  AND2X2 AND2X2_1517 ( .A(core__abc_21380_n1392), .B(core__abc_21380_n1393), .Y(core__abc_21380_n1394) );
  AND2X2 AND2X2_1518 ( .A(core_v0_reg_7_), .B(core_v1_reg_7_), .Y(core__abc_21380_n1395) );
  AND2X2 AND2X2_1519 ( .A(core_v3_reg_7_), .B(core_v2_reg_7_), .Y(core__abc_21380_n1398) );
  AND2X2 AND2X2_152 ( .A(_abc_19068_n916_1_bF_buf4), .B(word1_reg_9_), .Y(_abc_19068_n1140_1) );
  AND2X2 AND2X2_1520 ( .A(core__abc_21380_n1399), .B(core__abc_21380_n1400), .Y(core__abc_21380_n1401) );
  AND2X2 AND2X2_1521 ( .A(core__abc_21380_n1404), .B(core__abc_21380_n1405), .Y(core__abc_21380_n1406) );
  AND2X2 AND2X2_1522 ( .A(core__abc_21380_n1408), .B(reset_n_bF_buf83), .Y(core__abc_21380_n1409) );
  AND2X2 AND2X2_1523 ( .A(core__abc_21380_n1407), .B(core__abc_21380_n1409), .Y(core_siphash_word1_reg_7__FF_INPUT) );
  AND2X2 AND2X2_1524 ( .A(core_v0_reg_8_), .B(core_v1_reg_8_), .Y(core__abc_21380_n1411) );
  AND2X2 AND2X2_1525 ( .A(core__abc_21380_n1412), .B(core__abc_21380_n1413), .Y(core__abc_21380_n1414) );
  AND2X2 AND2X2_1526 ( .A(core_v2_reg_8_), .B(core_v3_reg_8_), .Y(core__abc_21380_n1415) );
  AND2X2 AND2X2_1527 ( .A(core__abc_21380_n1416), .B(core__abc_21380_n1417), .Y(core__abc_21380_n1418) );
  AND2X2 AND2X2_1528 ( .A(core__abc_21380_n1419), .B(core__abc_21380_n1414), .Y(core__abc_21380_n1420) );
  AND2X2 AND2X2_1529 ( .A(core__abc_21380_n1421), .B(core__abc_21380_n1418), .Y(core__abc_21380_n1422) );
  AND2X2 AND2X2_153 ( .A(_abc_19068_n897_1_bF_buf4), .B(word0_reg_9_), .Y(_abc_19068_n1141) );
  AND2X2 AND2X2_1530 ( .A(core__abc_21380_n1425), .B(reset_n_bF_buf82), .Y(core__abc_21380_n1426) );
  AND2X2 AND2X2_1531 ( .A(core__abc_21380_n1424), .B(core__abc_21380_n1426), .Y(core_siphash_word1_reg_8__FF_INPUT) );
  AND2X2 AND2X2_1532 ( .A(core_v0_reg_9_), .B(core_v1_reg_9_), .Y(core__abc_21380_n1428) );
  AND2X2 AND2X2_1533 ( .A(core__abc_21380_n1430), .B(core__abc_21380_n1431), .Y(core__abc_21380_n1432) );
  AND2X2 AND2X2_1534 ( .A(core__abc_21380_n1433), .B(core__abc_21380_n1429), .Y(core__abc_21380_n1434) );
  AND2X2 AND2X2_1535 ( .A(core_v2_reg_9_), .B(core_v3_reg_9_), .Y(core__abc_21380_n1435) );
  AND2X2 AND2X2_1536 ( .A(core__abc_21380_n1436), .B(core__abc_21380_n1437), .Y(core__abc_21380_n1438) );
  AND2X2 AND2X2_1537 ( .A(core__abc_21380_n1439), .B(core__abc_21380_n1434), .Y(core__abc_21380_n1440) );
  AND2X2 AND2X2_1538 ( .A(core__abc_21380_n1441), .B(core__abc_21380_n1438), .Y(core__abc_21380_n1442) );
  AND2X2 AND2X2_1539 ( .A(core__abc_21380_n1445), .B(reset_n_bF_buf81), .Y(core__abc_21380_n1446) );
  AND2X2 AND2X2_154 ( .A(_abc_19068_n941_bF_buf0), .B(core_key_105_), .Y(_abc_19068_n1143) );
  AND2X2 AND2X2_1540 ( .A(core__abc_21380_n1444), .B(core__abc_21380_n1446), .Y(core_siphash_word1_reg_9__FF_INPUT) );
  AND2X2 AND2X2_1541 ( .A(core_v0_reg_10_), .B(core_v1_reg_10_), .Y(core__abc_21380_n1449) );
  AND2X2 AND2X2_1542 ( .A(core__abc_21380_n1450), .B(core__abc_21380_n1448), .Y(core__abc_21380_n1451) );
  AND2X2 AND2X2_1543 ( .A(core_v3_reg_10_), .B(core_v2_reg_10_), .Y(core__abc_21380_n1452) );
  AND2X2 AND2X2_1544 ( .A(core__abc_21380_n1453), .B(core__abc_21380_n1454), .Y(core__abc_21380_n1455) );
  AND2X2 AND2X2_1545 ( .A(core__abc_21380_n1459), .B(core__abc_21380_n1456), .Y(core__abc_21380_n1460) );
  AND2X2 AND2X2_1546 ( .A(core__abc_21380_n1462), .B(reset_n_bF_buf80), .Y(core__abc_21380_n1463) );
  AND2X2 AND2X2_1547 ( .A(core__abc_21380_n1461), .B(core__abc_21380_n1463), .Y(core_siphash_word1_reg_10__FF_INPUT) );
  AND2X2 AND2X2_1548 ( .A(core_v0_reg_11_), .B(core_v1_reg_11_), .Y(core__abc_21380_n1466) );
  AND2X2 AND2X2_1549 ( .A(core__abc_21380_n1467), .B(core__abc_21380_n1465), .Y(core__abc_21380_n1468) );
  AND2X2 AND2X2_155 ( .A(_abc_19068_n924_1_bF_buf0), .B(core_key_41_), .Y(_abc_19068_n1144_1) );
  AND2X2 AND2X2_1550 ( .A(core_v3_reg_11_), .B(core_v2_reg_11_), .Y(core__abc_21380_n1469) );
  AND2X2 AND2X2_1551 ( .A(core__abc_21380_n1470), .B(core__abc_21380_n1471), .Y(core__abc_21380_n1472) );
  AND2X2 AND2X2_1552 ( .A(core__abc_21380_n1476), .B(core__abc_21380_n1473), .Y(core__abc_21380_n1477) );
  AND2X2 AND2X2_1553 ( .A(core__abc_21380_n1479), .B(reset_n_bF_buf79), .Y(core__abc_21380_n1480) );
  AND2X2 AND2X2_1554 ( .A(core__abc_21380_n1478), .B(core__abc_21380_n1480), .Y(core_siphash_word1_reg_11__FF_INPUT) );
  AND2X2 AND2X2_1555 ( .A(core_v0_reg_12_), .B(core_v1_reg_12_), .Y(core__abc_21380_n1482) );
  AND2X2 AND2X2_1556 ( .A(core__abc_21380_n1483), .B(core__abc_21380_n1484), .Y(core__abc_21380_n1485) );
  AND2X2 AND2X2_1557 ( .A(core_v2_reg_12_), .B(core_v3_reg_12_), .Y(core__abc_21380_n1488) );
  AND2X2 AND2X2_1558 ( .A(core__abc_21380_n1489), .B(core__abc_21380_n1490), .Y(core__abc_21380_n1491) );
  AND2X2 AND2X2_1559 ( .A(core__abc_21380_n1487), .B(core__abc_21380_n1492), .Y(core__abc_21380_n1493) );
  AND2X2 AND2X2_156 ( .A(_abc_19068_n926_bF_buf0), .B(core_key_9_), .Y(_abc_19068_n1145) );
  AND2X2 AND2X2_1560 ( .A(core__abc_21380_n1486), .B(core__abc_21380_n1491), .Y(core__abc_21380_n1494) );
  AND2X2 AND2X2_1561 ( .A(core__abc_21380_n1497), .B(reset_n_bF_buf78), .Y(core__abc_21380_n1498) );
  AND2X2 AND2X2_1562 ( .A(core__abc_21380_n1496), .B(core__abc_21380_n1498), .Y(core_siphash_word1_reg_12__FF_INPUT) );
  AND2X2 AND2X2_1563 ( .A(core__abc_21380_n1500), .B(core__abc_21380_n1501), .Y(core__abc_21380_n1502) );
  AND2X2 AND2X2_1564 ( .A(core_v0_reg_13_), .B(core_v1_reg_13_), .Y(core__abc_21380_n1503) );
  AND2X2 AND2X2_1565 ( .A(core_v3_reg_13_), .B(core_v2_reg_13_), .Y(core__abc_21380_n1506) );
  AND2X2 AND2X2_1566 ( .A(core__abc_21380_n1507), .B(core__abc_21380_n1508), .Y(core__abc_21380_n1509) );
  AND2X2 AND2X2_1567 ( .A(core__abc_21380_n1510), .B(core__abc_21380_n1512), .Y(core__abc_21380_n1513) );
  AND2X2 AND2X2_1568 ( .A(core__abc_21380_n1515), .B(reset_n_bF_buf77), .Y(core__abc_21380_n1516) );
  AND2X2 AND2X2_1569 ( .A(core__abc_21380_n1514), .B(core__abc_21380_n1516), .Y(core_siphash_word1_reg_13__FF_INPUT) );
  AND2X2 AND2X2_157 ( .A(_abc_19068_n939_1_bF_buf0), .B(core_key_73_), .Y(_abc_19068_n1149_1) );
  AND2X2 AND2X2_1570 ( .A(core__abc_21380_n1518), .B(core__abc_21380_n1519), .Y(core__abc_21380_n1520) );
  AND2X2 AND2X2_1571 ( .A(core_v0_reg_14_), .B(core_v1_reg_14_), .Y(core__abc_21380_n1521) );
  AND2X2 AND2X2_1572 ( .A(core_v3_reg_14_), .B(core_v2_reg_14_), .Y(core__abc_21380_n1524) );
  AND2X2 AND2X2_1573 ( .A(core__abc_21380_n1525), .B(core__abc_21380_n1526), .Y(core__abc_21380_n1527) );
  AND2X2 AND2X2_1574 ( .A(core__abc_21380_n1528), .B(core__abc_21380_n1530), .Y(core__abc_21380_n1531) );
  AND2X2 AND2X2_1575 ( .A(core__abc_21380_n1533), .B(reset_n_bF_buf76), .Y(core__abc_21380_n1534) );
  AND2X2 AND2X2_1576 ( .A(core__abc_21380_n1532), .B(core__abc_21380_n1534), .Y(core_siphash_word1_reg_14__FF_INPUT) );
  AND2X2 AND2X2_1577 ( .A(core__abc_21380_n1536), .B(core__abc_21380_n1537), .Y(core__abc_21380_n1538) );
  AND2X2 AND2X2_1578 ( .A(core_v0_reg_15_), .B(core_v1_reg_15_), .Y(core__abc_21380_n1540) );
  AND2X2 AND2X2_1579 ( .A(core__abc_21380_n1539), .B(core__abc_21380_n1541), .Y(core__abc_21380_n1542) );
  AND2X2 AND2X2_158 ( .A(_abc_19068_n899_bF_buf4), .B(word3_reg_9_), .Y(_abc_19068_n1150_1) );
  AND2X2 AND2X2_1580 ( .A(core_v3_reg_15_), .B(core_v2_reg_15_), .Y(core__abc_21380_n1543) );
  AND2X2 AND2X2_1581 ( .A(core__abc_21380_n1544), .B(core__abc_21380_n1545), .Y(core__abc_21380_n1546) );
  AND2X2 AND2X2_1582 ( .A(core__abc_21380_n1550), .B(core__abc_21380_n1547), .Y(core__abc_21380_n1551) );
  AND2X2 AND2X2_1583 ( .A(core__abc_21380_n1553), .B(reset_n_bF_buf75), .Y(core__abc_21380_n1554) );
  AND2X2 AND2X2_1584 ( .A(core__abc_21380_n1552), .B(core__abc_21380_n1554), .Y(core_siphash_word1_reg_15__FF_INPUT) );
  AND2X2 AND2X2_1585 ( .A(core_v0_reg_16_), .B(core_v1_reg_16_), .Y(core__abc_21380_n1556) );
  AND2X2 AND2X2_1586 ( .A(core__abc_21380_n1557), .B(core__abc_21380_n1558), .Y(core__abc_21380_n1559) );
  AND2X2 AND2X2_1587 ( .A(core_v2_reg_16_), .B(core_v3_reg_16_), .Y(core__abc_21380_n1562) );
  AND2X2 AND2X2_1588 ( .A(core__abc_21380_n1563), .B(core__abc_21380_n1564), .Y(core__abc_21380_n1565) );
  AND2X2 AND2X2_1589 ( .A(core__abc_21380_n1561), .B(core__abc_21380_n1566), .Y(core__abc_21380_n1567) );
  AND2X2 AND2X2_159 ( .A(_abc_19068_n902_bF_buf4), .B(word2_reg_9_), .Y(_abc_19068_n1151) );
  AND2X2 AND2X2_1590 ( .A(core__abc_21380_n1560), .B(core__abc_21380_n1565), .Y(core__abc_21380_n1568) );
  AND2X2 AND2X2_1591 ( .A(core__abc_21380_n1571), .B(reset_n_bF_buf74), .Y(core__abc_21380_n1572) );
  AND2X2 AND2X2_1592 ( .A(core__abc_21380_n1570), .B(core__abc_21380_n1572), .Y(core_siphash_word1_reg_16__FF_INPUT) );
  AND2X2 AND2X2_1593 ( .A(core_v0_reg_17_), .B(core_v1_reg_17_), .Y(core__abc_21380_n1574) );
  AND2X2 AND2X2_1594 ( .A(core__abc_21380_n1576), .B(core__abc_21380_n1577), .Y(core__abc_21380_n1578) );
  AND2X2 AND2X2_1595 ( .A(core__abc_21380_n1579), .B(core__abc_21380_n1575), .Y(core__abc_21380_n1580) );
  AND2X2 AND2X2_1596 ( .A(core_v2_reg_17_), .B(core_v3_reg_17_), .Y(core__abc_21380_n1581) );
  AND2X2 AND2X2_1597 ( .A(core__abc_21380_n1582), .B(core__abc_21380_n1583), .Y(core__abc_21380_n1584) );
  AND2X2 AND2X2_1598 ( .A(core__abc_21380_n1585), .B(core__abc_21380_n1580), .Y(core__abc_21380_n1586) );
  AND2X2 AND2X2_1599 ( .A(core__abc_21380_n1587), .B(core__abc_21380_n1584), .Y(core__abc_21380_n1588) );
  AND2X2 AND2X2_16 ( .A(_abc_19068_n878), .B(\addr[5] ), .Y(_abc_19068_n895_1) );
  AND2X2 AND2X2_160 ( .A(_abc_19068_n945_1_bF_buf0), .B(core_mi_9_), .Y(_abc_19068_n1153_1) );
  AND2X2 AND2X2_1600 ( .A(core__abc_21380_n1591), .B(reset_n_bF_buf73), .Y(core__abc_21380_n1592) );
  AND2X2 AND2X2_1601 ( .A(core__abc_21380_n1590), .B(core__abc_21380_n1592), .Y(core_siphash_word1_reg_17__FF_INPUT) );
  AND2X2 AND2X2_1602 ( .A(core_v0_reg_18_), .B(core_v1_reg_18_), .Y(core__abc_21380_n1595) );
  AND2X2 AND2X2_1603 ( .A(core__abc_21380_n1596), .B(core__abc_21380_n1594), .Y(core__abc_21380_n1597) );
  AND2X2 AND2X2_1604 ( .A(core_v3_reg_18_), .B(core_v2_reg_18_), .Y(core__abc_21380_n1598) );
  AND2X2 AND2X2_1605 ( .A(core__abc_21380_n1599), .B(core__abc_21380_n1600), .Y(core__abc_21380_n1601) );
  AND2X2 AND2X2_1606 ( .A(core__abc_21380_n1605), .B(core__abc_21380_n1602), .Y(core__abc_21380_n1606) );
  AND2X2 AND2X2_1607 ( .A(core__abc_21380_n1608), .B(reset_n_bF_buf72), .Y(core__abc_21380_n1609) );
  AND2X2 AND2X2_1608 ( .A(core__abc_21380_n1607), .B(core__abc_21380_n1609), .Y(core_siphash_word1_reg_18__FF_INPUT) );
  AND2X2 AND2X2_1609 ( .A(core_v0_reg_19_), .B(core_v1_reg_19_), .Y(core__abc_21380_n1611) );
  AND2X2 AND2X2_161 ( .A(_abc_19068_n915_1_bF_buf4), .B(core_mi_41_), .Y(_abc_19068_n1154) );
  AND2X2 AND2X2_1610 ( .A(core__abc_21380_n1612), .B(core__abc_21380_n1613), .Y(core__abc_21380_n1614) );
  AND2X2 AND2X2_1611 ( .A(core_v2_reg_19_), .B(core_v3_reg_19_), .Y(core__abc_21380_n1615) );
  AND2X2 AND2X2_1612 ( .A(core__abc_21380_n1616), .B(core__abc_21380_n1617), .Y(core__abc_21380_n1618) );
  AND2X2 AND2X2_1613 ( .A(core__abc_21380_n1619), .B(core__abc_21380_n1614), .Y(core__abc_21380_n1620) );
  AND2X2 AND2X2_1614 ( .A(core__abc_21380_n1621), .B(core__abc_21380_n1618), .Y(core__abc_21380_n1622) );
  AND2X2 AND2X2_1615 ( .A(core__abc_21380_n1625), .B(reset_n_bF_buf71), .Y(core__abc_21380_n1626) );
  AND2X2 AND2X2_1616 ( .A(core__abc_21380_n1624), .B(core__abc_21380_n1626), .Y(core_siphash_word1_reg_19__FF_INPUT) );
  AND2X2 AND2X2_1617 ( .A(core__abc_21380_n1628), .B(core__abc_21380_n1629), .Y(core__abc_21380_n1630) );
  AND2X2 AND2X2_1618 ( .A(core_v0_reg_20_), .B(core_v1_reg_20_), .Y(core__abc_21380_n1631) );
  AND2X2 AND2X2_1619 ( .A(core_v3_reg_20_), .B(core_v2_reg_20_), .Y(core__abc_21380_n1634) );
  AND2X2 AND2X2_162 ( .A(_abc_19068_n923_bF_buf0), .B(_abc_19068_n1158_1), .Y(_auto_iopadmap_cc_313_execute_30317_9_) );
  AND2X2 AND2X2_1620 ( .A(core__abc_21380_n1635), .B(core__abc_21380_n1636), .Y(core__abc_21380_n1637) );
  AND2X2 AND2X2_1621 ( .A(core__abc_21380_n1638), .B(core__abc_21380_n1640), .Y(core__abc_21380_n1641) );
  AND2X2 AND2X2_1622 ( .A(core__abc_21380_n1643), .B(reset_n_bF_buf70), .Y(core__abc_21380_n1644) );
  AND2X2 AND2X2_1623 ( .A(core__abc_21380_n1642), .B(core__abc_21380_n1644), .Y(core_siphash_word1_reg_20__FF_INPUT) );
  AND2X2 AND2X2_1624 ( .A(core__abc_21380_n1646), .B(core__abc_21380_n1647), .Y(core__abc_21380_n1648) );
  AND2X2 AND2X2_1625 ( .A(core_v0_reg_21_), .B(core_v1_reg_21_), .Y(core__abc_21380_n1649_1) );
  AND2X2 AND2X2_1626 ( .A(core_v3_reg_21_), .B(core_v2_reg_21_), .Y(core__abc_21380_n1652) );
  AND2X2 AND2X2_1627 ( .A(core__abc_21380_n1653), .B(core__abc_21380_n1654), .Y(core__abc_21380_n1655_1) );
  AND2X2 AND2X2_1628 ( .A(core__abc_21380_n1656), .B(core__abc_21380_n1658), .Y(core__abc_21380_n1659) );
  AND2X2 AND2X2_1629 ( .A(core__abc_21380_n1661), .B(reset_n_bF_buf69), .Y(core__abc_21380_n1662) );
  AND2X2 AND2X2_163 ( .A(_abc_19068_n916_1_bF_buf3), .B(word1_reg_10_), .Y(_abc_19068_n1160) );
  AND2X2 AND2X2_1630 ( .A(core__abc_21380_n1660), .B(core__abc_21380_n1662), .Y(core_siphash_word1_reg_21__FF_INPUT) );
  AND2X2 AND2X2_1631 ( .A(core__abc_21380_n1664), .B(core__abc_21380_n1665), .Y(core__abc_21380_n1666) );
  AND2X2 AND2X2_1632 ( .A(core_v0_reg_22_), .B(core_v1_reg_22_), .Y(core__abc_21380_n1667) );
  AND2X2 AND2X2_1633 ( .A(core_v3_reg_22_), .B(core_v2_reg_22_), .Y(core__abc_21380_n1670) );
  AND2X2 AND2X2_1634 ( .A(core__abc_21380_n1671), .B(core__abc_21380_n1672), .Y(core__abc_21380_n1673) );
  AND2X2 AND2X2_1635 ( .A(core__abc_21380_n1674), .B(core__abc_21380_n1676), .Y(core__abc_21380_n1677) );
  AND2X2 AND2X2_1636 ( .A(core__abc_21380_n1679), .B(reset_n_bF_buf68), .Y(core__abc_21380_n1680) );
  AND2X2 AND2X2_1637 ( .A(core__abc_21380_n1678), .B(core__abc_21380_n1680), .Y(core_siphash_word1_reg_22__FF_INPUT) );
  AND2X2 AND2X2_1638 ( .A(core__abc_21380_n1682), .B(core__abc_21380_n1683), .Y(core__abc_21380_n1684) );
  AND2X2 AND2X2_1639 ( .A(core_v0_reg_23_), .B(core_v1_reg_23_), .Y(core__abc_21380_n1686) );
  AND2X2 AND2X2_164 ( .A(_abc_19068_n897_1_bF_buf3), .B(word0_reg_10_), .Y(_abc_19068_n1161_1) );
  AND2X2 AND2X2_1640 ( .A(core__abc_21380_n1685), .B(core__abc_21380_n1687), .Y(core__abc_21380_n1688) );
  AND2X2 AND2X2_1641 ( .A(core_v3_reg_23_), .B(core_v2_reg_23_), .Y(core__abc_21380_n1689) );
  AND2X2 AND2X2_1642 ( .A(core__abc_21380_n1690), .B(core__abc_21380_n1691), .Y(core__abc_21380_n1692) );
  AND2X2 AND2X2_1643 ( .A(core__abc_21380_n1696), .B(core__abc_21380_n1693), .Y(core__abc_21380_n1697) );
  AND2X2 AND2X2_1644 ( .A(core__abc_21380_n1699), .B(reset_n_bF_buf67), .Y(core__abc_21380_n1700) );
  AND2X2 AND2X2_1645 ( .A(core__abc_21380_n1698), .B(core__abc_21380_n1700), .Y(core_siphash_word1_reg_23__FF_INPUT) );
  AND2X2 AND2X2_1646 ( .A(core__abc_21380_n1702), .B(core__abc_21380_n1703), .Y(core__abc_21380_n1704) );
  AND2X2 AND2X2_1647 ( .A(core_v0_reg_24_), .B(core_v1_reg_24_), .Y(core__abc_21380_n1705) );
  AND2X2 AND2X2_1648 ( .A(core_v3_reg_24_), .B(core_v2_reg_24_), .Y(core__abc_21380_n1708) );
  AND2X2 AND2X2_1649 ( .A(core__abc_21380_n1709), .B(core__abc_21380_n1710), .Y(core__abc_21380_n1711) );
  AND2X2 AND2X2_165 ( .A(_abc_19068_n939_1_bF_buf4), .B(core_key_74_), .Y(_abc_19068_n1163) );
  AND2X2 AND2X2_1650 ( .A(core__abc_21380_n1712), .B(core__abc_21380_n1714), .Y(core__abc_21380_n1715) );
  AND2X2 AND2X2_1651 ( .A(core__abc_21380_n1717), .B(reset_n_bF_buf66), .Y(core__abc_21380_n1718) );
  AND2X2 AND2X2_1652 ( .A(core__abc_21380_n1716), .B(core__abc_21380_n1718), .Y(core_siphash_word1_reg_24__FF_INPUT) );
  AND2X2 AND2X2_1653 ( .A(core__abc_21380_n1720), .B(core__abc_21380_n1721), .Y(core__abc_21380_n1722) );
  AND2X2 AND2X2_1654 ( .A(core_v0_reg_25_), .B(core_v1_reg_25_), .Y(core__abc_21380_n1724) );
  AND2X2 AND2X2_1655 ( .A(core__abc_21380_n1723), .B(core__abc_21380_n1725), .Y(core__abc_21380_n1726) );
  AND2X2 AND2X2_1656 ( .A(core_v3_reg_25_), .B(core_v2_reg_25_), .Y(core__abc_21380_n1727) );
  AND2X2 AND2X2_1657 ( .A(core__abc_21380_n1728), .B(core__abc_21380_n1729), .Y(core__abc_21380_n1730) );
  AND2X2 AND2X2_1658 ( .A(core__abc_21380_n1734), .B(core__abc_21380_n1731), .Y(core__abc_21380_n1735) );
  AND2X2 AND2X2_1659 ( .A(core__abc_21380_n1737), .B(reset_n_bF_buf65), .Y(core__abc_21380_n1738) );
  AND2X2 AND2X2_166 ( .A(_abc_19068_n924_1_bF_buf4), .B(core_key_42_), .Y(_abc_19068_n1164_1) );
  AND2X2 AND2X2_1660 ( .A(core__abc_21380_n1736), .B(core__abc_21380_n1738), .Y(core_siphash_word1_reg_25__FF_INPUT) );
  AND2X2 AND2X2_1661 ( .A(core_v0_reg_26_), .B(core_v1_reg_26_), .Y(core__abc_21380_n1741) );
  AND2X2 AND2X2_1662 ( .A(core__abc_21380_n1742), .B(core__abc_21380_n1740), .Y(core__abc_21380_n1743) );
  AND2X2 AND2X2_1663 ( .A(core_v3_reg_26_), .B(core_v2_reg_26_), .Y(core__abc_21380_n1744) );
  AND2X2 AND2X2_1664 ( .A(core__abc_21380_n1745), .B(core__abc_21380_n1746), .Y(core__abc_21380_n1747) );
  AND2X2 AND2X2_1665 ( .A(core__abc_21380_n1751), .B(core__abc_21380_n1748), .Y(core__abc_21380_n1752) );
  AND2X2 AND2X2_1666 ( .A(core__abc_21380_n1754_1), .B(reset_n_bF_buf64), .Y(core__abc_21380_n1755) );
  AND2X2 AND2X2_1667 ( .A(core__abc_21380_n1753), .B(core__abc_21380_n1755), .Y(core_siphash_word1_reg_26__FF_INPUT) );
  AND2X2 AND2X2_1668 ( .A(core__abc_21380_n1757), .B(core__abc_21380_n1758), .Y(core__abc_21380_n1759) );
  AND2X2 AND2X2_1669 ( .A(core_v0_reg_27_), .B(core_v1_reg_27_), .Y(core__abc_21380_n1761) );
  AND2X2 AND2X2_167 ( .A(_abc_19068_n926_bF_buf4), .B(core_key_10_), .Y(_abc_19068_n1165_1) );
  AND2X2 AND2X2_1670 ( .A(core__abc_21380_n1760_1), .B(core__abc_21380_n1762), .Y(core__abc_21380_n1763) );
  AND2X2 AND2X2_1671 ( .A(core_v3_reg_27_), .B(core_v2_reg_27_), .Y(core__abc_21380_n1764) );
  AND2X2 AND2X2_1672 ( .A(core__abc_21380_n1765), .B(core__abc_21380_n1766), .Y(core__abc_21380_n1767) );
  AND2X2 AND2X2_1673 ( .A(core__abc_21380_n1771), .B(core__abc_21380_n1768), .Y(core__abc_21380_n1772) );
  AND2X2 AND2X2_1674 ( .A(core__abc_21380_n1774), .B(reset_n_bF_buf63), .Y(core__abc_21380_n1775) );
  AND2X2 AND2X2_1675 ( .A(core__abc_21380_n1773), .B(core__abc_21380_n1775), .Y(core_siphash_word1_reg_27__FF_INPUT) );
  AND2X2 AND2X2_1676 ( .A(core__abc_21380_n1777), .B(core__abc_21380_n1778), .Y(core__abc_21380_n1779) );
  AND2X2 AND2X2_1677 ( .A(core_v0_reg_28_), .B(core_v1_reg_28_), .Y(core__abc_21380_n1780) );
  AND2X2 AND2X2_1678 ( .A(core_v3_reg_28_), .B(core_v2_reg_28_), .Y(core__abc_21380_n1783) );
  AND2X2 AND2X2_1679 ( .A(core__abc_21380_n1784), .B(core__abc_21380_n1785), .Y(core__abc_21380_n1786_1) );
  AND2X2 AND2X2_168 ( .A(_abc_19068_n941_bF_buf4), .B(core_key_106_), .Y(_abc_19068_n1169) );
  AND2X2 AND2X2_1680 ( .A(core__abc_21380_n1787), .B(core__abc_21380_n1789), .Y(core__abc_21380_n1790) );
  AND2X2 AND2X2_1681 ( .A(core__abc_21380_n1792), .B(reset_n_bF_buf62), .Y(core__abc_21380_n1793) );
  AND2X2 AND2X2_1682 ( .A(core__abc_21380_n1791), .B(core__abc_21380_n1793), .Y(core_siphash_word1_reg_28__FF_INPUT) );
  AND2X2 AND2X2_1683 ( .A(core__abc_21380_n1795), .B(core__abc_21380_n1796), .Y(core__abc_21380_n1797) );
  AND2X2 AND2X2_1684 ( .A(core_v0_reg_29_), .B(core_v1_reg_29_), .Y(core__abc_21380_n1799) );
  AND2X2 AND2X2_1685 ( .A(core__abc_21380_n1798), .B(core__abc_21380_n1800), .Y(core__abc_21380_n1801) );
  AND2X2 AND2X2_1686 ( .A(core_v3_reg_29_), .B(core_v2_reg_29_), .Y(core__abc_21380_n1802) );
  AND2X2 AND2X2_1687 ( .A(core__abc_21380_n1803), .B(core__abc_21380_n1804), .Y(core__abc_21380_n1805) );
  AND2X2 AND2X2_1688 ( .A(core__abc_21380_n1809), .B(core__abc_21380_n1806), .Y(core__abc_21380_n1810) );
  AND2X2 AND2X2_1689 ( .A(core__abc_21380_n1812_1), .B(reset_n_bF_buf61), .Y(core__abc_21380_n1813) );
  AND2X2 AND2X2_169 ( .A(_abc_19068_n902_bF_buf3), .B(word2_reg_10_), .Y(_abc_19068_n1170_1) );
  AND2X2 AND2X2_1690 ( .A(core__abc_21380_n1811), .B(core__abc_21380_n1813), .Y(core_siphash_word1_reg_29__FF_INPUT) );
  AND2X2 AND2X2_1691 ( .A(core__abc_21380_n1815), .B(core__abc_21380_n1816_1), .Y(core__abc_21380_n1817) );
  AND2X2 AND2X2_1692 ( .A(core_v0_reg_30_), .B(core_v1_reg_30_), .Y(core__abc_21380_n1818) );
  AND2X2 AND2X2_1693 ( .A(core_v3_reg_30_), .B(core_v2_reg_30_), .Y(core__abc_21380_n1821) );
  AND2X2 AND2X2_1694 ( .A(core__abc_21380_n1822), .B(core__abc_21380_n1823), .Y(core__abc_21380_n1824) );
  AND2X2 AND2X2_1695 ( .A(core__abc_21380_n1825), .B(core__abc_21380_n1827), .Y(core__abc_21380_n1828) );
  AND2X2 AND2X2_1696 ( .A(core__abc_21380_n1830), .B(reset_n_bF_buf60), .Y(core__abc_21380_n1831) );
  AND2X2 AND2X2_1697 ( .A(core__abc_21380_n1829), .B(core__abc_21380_n1831), .Y(core_siphash_word1_reg_30__FF_INPUT) );
  AND2X2 AND2X2_1698 ( .A(core__abc_21380_n1833), .B(core__abc_21380_n1834), .Y(core__abc_21380_n1835) );
  AND2X2 AND2X2_1699 ( .A(core_v0_reg_31_), .B(core_v1_reg_31_), .Y(core__abc_21380_n1837) );
  AND2X2 AND2X2_17 ( .A(_abc_19068_n877_1), .B(_abc_19068_n895_1), .Y(_abc_19068_n896) );
  AND2X2 AND2X2_170 ( .A(_abc_19068_n899_bF_buf3), .B(word3_reg_10_), .Y(_abc_19068_n1171_1) );
  AND2X2 AND2X2_1700 ( .A(core__abc_21380_n1836), .B(core__abc_21380_n1838), .Y(core__abc_21380_n1839) );
  AND2X2 AND2X2_1701 ( .A(core_v3_reg_31_), .B(core_v2_reg_31_), .Y(core__abc_21380_n1840) );
  AND2X2 AND2X2_1702 ( .A(core__abc_21380_n1841), .B(core__abc_21380_n1842), .Y(core__abc_21380_n1843) );
  AND2X2 AND2X2_1703 ( .A(core__abc_21380_n1847), .B(core__abc_21380_n1844), .Y(core__abc_21380_n1848) );
  AND2X2 AND2X2_1704 ( .A(core__abc_21380_n1850), .B(reset_n_bF_buf59), .Y(core__abc_21380_n1851) );
  AND2X2 AND2X2_1705 ( .A(core__abc_21380_n1849), .B(core__abc_21380_n1851), .Y(core_siphash_word1_reg_31__FF_INPUT) );
  AND2X2 AND2X2_1706 ( .A(core__abc_21380_n1853), .B(core__abc_21380_n1854), .Y(core__abc_21380_n1855) );
  AND2X2 AND2X2_1707 ( .A(core_v0_reg_32_), .B(core_v1_reg_32_), .Y(core__abc_21380_n1856) );
  AND2X2 AND2X2_1708 ( .A(core_v3_reg_32_), .B(core_v2_reg_32_), .Y(core__abc_21380_n1859) );
  AND2X2 AND2X2_1709 ( .A(core__abc_21380_n1860), .B(core__abc_21380_n1861), .Y(core__abc_21380_n1862) );
  AND2X2 AND2X2_171 ( .A(_abc_19068_n945_1_bF_buf4), .B(core_mi_10_), .Y(_abc_19068_n1173_1) );
  AND2X2 AND2X2_1710 ( .A(core__abc_21380_n1863), .B(core__abc_21380_n1865), .Y(core__abc_21380_n1866) );
  AND2X2 AND2X2_1711 ( .A(core__abc_21380_n1868), .B(reset_n_bF_buf58), .Y(core__abc_21380_n1869) );
  AND2X2 AND2X2_1712 ( .A(core__abc_21380_n1867), .B(core__abc_21380_n1869), .Y(core_siphash_word1_reg_32__FF_INPUT) );
  AND2X2 AND2X2_1713 ( .A(core__abc_21380_n1871), .B(core__abc_21380_n1872), .Y(core__abc_21380_n1873) );
  AND2X2 AND2X2_1714 ( .A(core_v0_reg_33_), .B(core_v1_reg_33_), .Y(core__abc_21380_n1874) );
  AND2X2 AND2X2_1715 ( .A(core_v3_reg_33_), .B(core_v2_reg_33_), .Y(core__abc_21380_n1877) );
  AND2X2 AND2X2_1716 ( .A(core__abc_21380_n1878), .B(core__abc_21380_n1879), .Y(core__abc_21380_n1880) );
  AND2X2 AND2X2_1717 ( .A(core__abc_21380_n1881), .B(core__abc_21380_n1883), .Y(core__abc_21380_n1884) );
  AND2X2 AND2X2_1718 ( .A(core__abc_21380_n1886), .B(reset_n_bF_buf57), .Y(core__abc_21380_n1887) );
  AND2X2 AND2X2_1719 ( .A(core__abc_21380_n1885), .B(core__abc_21380_n1887), .Y(core_siphash_word1_reg_33__FF_INPUT) );
  AND2X2 AND2X2_172 ( .A(_abc_19068_n915_1_bF_buf3), .B(core_mi_42_), .Y(_abc_19068_n1174_1) );
  AND2X2 AND2X2_1720 ( .A(core__abc_21380_n1889), .B(core__abc_21380_n1890), .Y(core__abc_21380_n1891) );
  AND2X2 AND2X2_1721 ( .A(core_v0_reg_34_), .B(core_v1_reg_34_), .Y(core__abc_21380_n1892) );
  AND2X2 AND2X2_1722 ( .A(core_v3_reg_34_), .B(core_v2_reg_34_), .Y(core__abc_21380_n1895) );
  AND2X2 AND2X2_1723 ( .A(core__abc_21380_n1896), .B(core__abc_21380_n1897), .Y(core__abc_21380_n1898) );
  AND2X2 AND2X2_1724 ( .A(core__abc_21380_n1899), .B(core__abc_21380_n1901), .Y(core__abc_21380_n1902) );
  AND2X2 AND2X2_1725 ( .A(core__abc_21380_n1904), .B(reset_n_bF_buf56), .Y(core__abc_21380_n1905) );
  AND2X2 AND2X2_1726 ( .A(core__abc_21380_n1903), .B(core__abc_21380_n1905), .Y(core_siphash_word1_reg_34__FF_INPUT) );
  AND2X2 AND2X2_1727 ( .A(core__abc_21380_n1907), .B(core__abc_21380_n1908), .Y(core__abc_21380_n1909) );
  AND2X2 AND2X2_1728 ( .A(core_v0_reg_35_), .B(core_v1_reg_35_), .Y(core__abc_21380_n1911) );
  AND2X2 AND2X2_1729 ( .A(core__abc_21380_n1910), .B(core__abc_21380_n1912), .Y(core__abc_21380_n1913) );
  AND2X2 AND2X2_173 ( .A(_abc_19068_n923_bF_buf4), .B(_abc_19068_n1178), .Y(_auto_iopadmap_cc_313_execute_30317_10_) );
  AND2X2 AND2X2_1730 ( .A(core_v3_reg_35_), .B(core_v2_reg_35_), .Y(core__abc_21380_n1914) );
  AND2X2 AND2X2_1731 ( .A(core__abc_21380_n1915), .B(core__abc_21380_n1916), .Y(core__abc_21380_n1917) );
  AND2X2 AND2X2_1732 ( .A(core__abc_21380_n1921), .B(core__abc_21380_n1918), .Y(core__abc_21380_n1922) );
  AND2X2 AND2X2_1733 ( .A(core__abc_21380_n1924), .B(reset_n_bF_buf55), .Y(core__abc_21380_n1925) );
  AND2X2 AND2X2_1734 ( .A(core__abc_21380_n1923), .B(core__abc_21380_n1925), .Y(core_siphash_word1_reg_35__FF_INPUT) );
  AND2X2 AND2X2_1735 ( .A(core_v0_reg_36_), .B(core_v1_reg_36_), .Y(core__abc_21380_n1927) );
  AND2X2 AND2X2_1736 ( .A(core__abc_21380_n1928_1), .B(core__abc_21380_n1929), .Y(core__abc_21380_n1930) );
  AND2X2 AND2X2_1737 ( .A(core_v3_reg_36_), .B(core_v2_reg_36_), .Y(core__abc_21380_n1932) );
  AND2X2 AND2X2_1738 ( .A(core__abc_21380_n1933), .B(core__abc_21380_n1934_1), .Y(core__abc_21380_n1935) );
  AND2X2 AND2X2_1739 ( .A(core__abc_21380_n1931), .B(core__abc_21380_n1935), .Y(core__abc_21380_n1936) );
  AND2X2 AND2X2_174 ( .A(_abc_19068_n939_1_bF_buf3), .B(core_key_75_), .Y(_abc_19068_n1180_1) );
  AND2X2 AND2X2_1740 ( .A(core__abc_21380_n1937), .B(core__abc_21380_n1938), .Y(core__abc_21380_n1939) );
  AND2X2 AND2X2_1741 ( .A(core__abc_21380_n1942), .B(reset_n_bF_buf54), .Y(core__abc_21380_n1943) );
  AND2X2 AND2X2_1742 ( .A(core__abc_21380_n1941), .B(core__abc_21380_n1943), .Y(core_siphash_word1_reg_36__FF_INPUT) );
  AND2X2 AND2X2_1743 ( .A(core_v0_reg_37_), .B(core_v1_reg_37_), .Y(core__abc_21380_n1945) );
  AND2X2 AND2X2_1744 ( .A(core__abc_21380_n1947), .B(core__abc_21380_n1948), .Y(core__abc_21380_n1949) );
  AND2X2 AND2X2_1745 ( .A(core__abc_21380_n1950), .B(core__abc_21380_n1946), .Y(core__abc_21380_n1951) );
  AND2X2 AND2X2_1746 ( .A(core_v3_reg_37_), .B(core_v2_reg_37_), .Y(core__abc_21380_n1952) );
  AND2X2 AND2X2_1747 ( .A(core__abc_21380_n1953), .B(core__abc_21380_n1954), .Y(core__abc_21380_n1955) );
  AND2X2 AND2X2_1748 ( .A(core__abc_21380_n1956), .B(core__abc_21380_n1951), .Y(core__abc_21380_n1957) );
  AND2X2 AND2X2_1749 ( .A(core__abc_21380_n1958), .B(core__abc_21380_n1955), .Y(core__abc_21380_n1959) );
  AND2X2 AND2X2_175 ( .A(_abc_19068_n926_bF_buf3), .B(core_key_11_), .Y(_abc_19068_n1181) );
  AND2X2 AND2X2_1750 ( .A(core__abc_21380_n1962), .B(reset_n_bF_buf53), .Y(core__abc_21380_n1963) );
  AND2X2 AND2X2_1751 ( .A(core__abc_21380_n1961_1), .B(core__abc_21380_n1963), .Y(core_siphash_word1_reg_37__FF_INPUT) );
  AND2X2 AND2X2_1752 ( .A(core__abc_21380_n1965_1), .B(core__abc_21380_n1966), .Y(core__abc_21380_n1967) );
  AND2X2 AND2X2_1753 ( .A(core_v0_reg_38_), .B(core_v1_reg_38_), .Y(core__abc_21380_n1968) );
  AND2X2 AND2X2_1754 ( .A(core_v3_reg_38_), .B(core_v2_reg_38_), .Y(core__abc_21380_n1971) );
  AND2X2 AND2X2_1755 ( .A(core__abc_21380_n1972), .B(core__abc_21380_n1973), .Y(core__abc_21380_n1974) );
  AND2X2 AND2X2_1756 ( .A(core__abc_21380_n1975), .B(core__abc_21380_n1977), .Y(core__abc_21380_n1978) );
  AND2X2 AND2X2_1757 ( .A(core__abc_21380_n1980), .B(reset_n_bF_buf52), .Y(core__abc_21380_n1981) );
  AND2X2 AND2X2_1758 ( .A(core__abc_21380_n1979), .B(core__abc_21380_n1981), .Y(core_siphash_word1_reg_38__FF_INPUT) );
  AND2X2 AND2X2_1759 ( .A(core__abc_21380_n1983), .B(core__abc_21380_n1984), .Y(core__abc_21380_n1985) );
  AND2X2 AND2X2_176 ( .A(_abc_19068_n924_1_bF_buf3), .B(core_key_43_), .Y(_abc_19068_n1182_1) );
  AND2X2 AND2X2_1760 ( .A(core_v0_reg_39_), .B(core_v1_reg_39_), .Y(core__abc_21380_n1987) );
  AND2X2 AND2X2_1761 ( .A(core__abc_21380_n1986), .B(core__abc_21380_n1988), .Y(core__abc_21380_n1989) );
  AND2X2 AND2X2_1762 ( .A(core_v3_reg_39_), .B(core_v2_reg_39_), .Y(core__abc_21380_n1990) );
  AND2X2 AND2X2_1763 ( .A(core__abc_21380_n1991), .B(core__abc_21380_n1992), .Y(core__abc_21380_n1993) );
  AND2X2 AND2X2_1764 ( .A(core__abc_21380_n1997), .B(core__abc_21380_n1994), .Y(core__abc_21380_n1998) );
  AND2X2 AND2X2_1765 ( .A(core__abc_21380_n2000), .B(reset_n_bF_buf51), .Y(core__abc_21380_n2001_1) );
  AND2X2 AND2X2_1766 ( .A(core__abc_21380_n1999), .B(core__abc_21380_n2001_1), .Y(core_siphash_word1_reg_39__FF_INPUT) );
  AND2X2 AND2X2_1767 ( .A(core_v0_reg_40_), .B(core_v1_reg_40_), .Y(core__abc_21380_n2003) );
  AND2X2 AND2X2_1768 ( .A(core__abc_21380_n2004), .B(core__abc_21380_n2005), .Y(core__abc_21380_n2006) );
  AND2X2 AND2X2_1769 ( .A(core_v3_reg_40_), .B(core_v2_reg_40_), .Y(core__abc_21380_n2009) );
  AND2X2 AND2X2_177 ( .A(_abc_19068_n881), .B(_abc_19068_n907_1), .Y(_abc_19068_n1185_1) );
  AND2X2 AND2X2_1770 ( .A(core__abc_21380_n2010), .B(core__abc_21380_n2011), .Y(core__abc_21380_n2012) );
  AND2X2 AND2X2_1771 ( .A(core__abc_21380_n2008), .B(core__abc_21380_n2013), .Y(core__abc_21380_n2014) );
  AND2X2 AND2X2_1772 ( .A(core__abc_21380_n2007), .B(core__abc_21380_n2012), .Y(core__abc_21380_n2015) );
  AND2X2 AND2X2_1773 ( .A(core__abc_21380_n2018), .B(reset_n_bF_buf50), .Y(core__abc_21380_n2019) );
  AND2X2 AND2X2_1774 ( .A(core__abc_21380_n2017), .B(core__abc_21380_n2019), .Y(core_siphash_word1_reg_40__FF_INPUT) );
  AND2X2 AND2X2_1775 ( .A(core_v0_reg_41_), .B(core_v1_reg_41_), .Y(core__abc_21380_n2021) );
  AND2X2 AND2X2_1776 ( .A(core__abc_21380_n2022), .B(core__abc_21380_n2023), .Y(core__abc_21380_n2024) );
  AND2X2 AND2X2_1777 ( .A(core_v3_reg_41_), .B(core_v2_reg_41_), .Y(core__abc_21380_n2026) );
  AND2X2 AND2X2_1778 ( .A(core__abc_21380_n2027), .B(core__abc_21380_n2028), .Y(core__abc_21380_n2029) );
  AND2X2 AND2X2_1779 ( .A(core__abc_21380_n2025), .B(core__abc_21380_n2029), .Y(core__abc_21380_n2030) );
  AND2X2 AND2X2_178 ( .A(_abc_19068_n899_bF_buf2), .B(word3_reg_11_), .Y(_abc_19068_n1186_1) );
  AND2X2 AND2X2_1780 ( .A(core__abc_21380_n2031), .B(core__abc_21380_n2032), .Y(core__abc_21380_n2033) );
  AND2X2 AND2X2_1781 ( .A(core__abc_21380_n2036), .B(reset_n_bF_buf49), .Y(core__abc_21380_n2037) );
  AND2X2 AND2X2_1782 ( .A(core__abc_21380_n2035_1), .B(core__abc_21380_n2037), .Y(core_siphash_word1_reg_41__FF_INPUT) );
  AND2X2 AND2X2_1783 ( .A(core__abc_21380_n2039_1), .B(core__abc_21380_n2040), .Y(core__abc_21380_n2041) );
  AND2X2 AND2X2_1784 ( .A(core_v0_reg_42_), .B(core_v1_reg_42_), .Y(core__abc_21380_n2042) );
  AND2X2 AND2X2_1785 ( .A(core_v3_reg_42_), .B(core_v2_reg_42_), .Y(core__abc_21380_n2045) );
  AND2X2 AND2X2_1786 ( .A(core__abc_21380_n2046), .B(core__abc_21380_n2047), .Y(core__abc_21380_n2048) );
  AND2X2 AND2X2_1787 ( .A(core__abc_21380_n2049), .B(core__abc_21380_n2051), .Y(core__abc_21380_n2052) );
  AND2X2 AND2X2_1788 ( .A(core__abc_21380_n2054), .B(reset_n_bF_buf48), .Y(core__abc_21380_n2055) );
  AND2X2 AND2X2_1789 ( .A(core__abc_21380_n2053), .B(core__abc_21380_n2055), .Y(core_siphash_word1_reg_42__FF_INPUT) );
  AND2X2 AND2X2_179 ( .A(_abc_19068_n902_bF_buf2), .B(word2_reg_11_), .Y(_abc_19068_n1188_1) );
  AND2X2 AND2X2_1790 ( .A(core__abc_21380_n2057), .B(core__abc_21380_n2058), .Y(core__abc_21380_n2059) );
  AND2X2 AND2X2_1791 ( .A(core_v0_reg_43_), .B(core_v1_reg_43_), .Y(core__abc_21380_n2061) );
  AND2X2 AND2X2_1792 ( .A(core__abc_21380_n2060), .B(core__abc_21380_n2062), .Y(core__abc_21380_n2063) );
  AND2X2 AND2X2_1793 ( .A(core_v3_reg_43_), .B(core_v2_reg_43_), .Y(core__abc_21380_n2065) );
  AND2X2 AND2X2_1794 ( .A(core__abc_21380_n2066), .B(core__abc_21380_n2064), .Y(core__abc_21380_n2067_1) );
  AND2X2 AND2X2_1795 ( .A(core__abc_21380_n2071), .B(core__abc_21380_n2068), .Y(core__abc_21380_n2072) );
  AND2X2 AND2X2_1796 ( .A(core__abc_21380_n2074), .B(reset_n_bF_buf47), .Y(core__abc_21380_n2075) );
  AND2X2 AND2X2_1797 ( .A(core__abc_21380_n2073_1), .B(core__abc_21380_n2075), .Y(core_siphash_word1_reg_43__FF_INPUT) );
  AND2X2 AND2X2_1798 ( .A(core_v0_reg_44_), .B(core_v1_reg_44_), .Y(core__abc_21380_n2077) );
  AND2X2 AND2X2_1799 ( .A(core__abc_21380_n2078), .B(core__abc_21380_n2079), .Y(core__abc_21380_n2080) );
  AND2X2 AND2X2_18 ( .A(_abc_19068_n894_1), .B(_abc_19068_n896), .Y(_abc_19068_n897_1) );
  AND2X2 AND2X2_180 ( .A(_abc_19068_n916_1_bF_buf2), .B(word1_reg_11_), .Y(_abc_19068_n1189_1) );
  AND2X2 AND2X2_1800 ( .A(core_v2_reg_44_), .B(core_v3_reg_44_), .Y(core__abc_21380_n2083) );
  AND2X2 AND2X2_1801 ( .A(core__abc_21380_n2084), .B(core__abc_21380_n2082), .Y(core__abc_21380_n2085) );
  AND2X2 AND2X2_1802 ( .A(core__abc_21380_n2081), .B(core__abc_21380_n2085), .Y(core__abc_21380_n2086) );
  AND2X2 AND2X2_1803 ( .A(core__abc_21380_n2087), .B(core__abc_21380_n2088), .Y(core__abc_21380_n2089) );
  AND2X2 AND2X2_1804 ( .A(core__abc_21380_n2092), .B(reset_n_bF_buf46), .Y(core__abc_21380_n2093) );
  AND2X2 AND2X2_1805 ( .A(core__abc_21380_n2091), .B(core__abc_21380_n2093), .Y(core_siphash_word1_reg_44__FF_INPUT) );
  AND2X2 AND2X2_1806 ( .A(core__abc_21380_n2095), .B(core__abc_21380_n2096), .Y(core__abc_21380_n2097) );
  AND2X2 AND2X2_1807 ( .A(core_v0_reg_45_), .B(core_v1_reg_45_), .Y(core__abc_21380_n2099_1) );
  AND2X2 AND2X2_1808 ( .A(core__abc_21380_n2098), .B(core__abc_21380_n2100), .Y(core__abc_21380_n2101) );
  AND2X2 AND2X2_1809 ( .A(core_v3_reg_45_), .B(core_v2_reg_45_), .Y(core__abc_21380_n2103_1) );
  AND2X2 AND2X2_181 ( .A(_abc_19068_n941_bF_buf3), .B(core_key_107_), .Y(_abc_19068_n1192_1) );
  AND2X2 AND2X2_1810 ( .A(core__abc_21380_n2104), .B(core__abc_21380_n2102), .Y(core__abc_21380_n2105) );
  AND2X2 AND2X2_1811 ( .A(core__abc_21380_n2109), .B(core__abc_21380_n2106), .Y(core__abc_21380_n2110) );
  AND2X2 AND2X2_1812 ( .A(core__abc_21380_n2112), .B(reset_n_bF_buf45), .Y(core__abc_21380_n2113) );
  AND2X2 AND2X2_1813 ( .A(core__abc_21380_n2111), .B(core__abc_21380_n2113), .Y(core_siphash_word1_reg_45__FF_INPUT) );
  AND2X2 AND2X2_1814 ( .A(core_v0_reg_46_), .B(core_v1_reg_46_), .Y(core__abc_21380_n2115) );
  AND2X2 AND2X2_1815 ( .A(core__abc_21380_n2116), .B(core__abc_21380_n2117), .Y(core__abc_21380_n2118) );
  AND2X2 AND2X2_1816 ( .A(core_v2_reg_46_), .B(core_v3_reg_46_), .Y(core__abc_21380_n2121) );
  AND2X2 AND2X2_1817 ( .A(core__abc_21380_n2122), .B(core__abc_21380_n2120), .Y(core__abc_21380_n2123) );
  AND2X2 AND2X2_1818 ( .A(core__abc_21380_n2119), .B(core__abc_21380_n2123), .Y(core__abc_21380_n2124) );
  AND2X2 AND2X2_1819 ( .A(core__abc_21380_n2125), .B(core__abc_21380_n2126), .Y(core__abc_21380_n2127) );
  AND2X2 AND2X2_182 ( .A(_abc_19068_n945_1_bF_buf3), .B(core_mi_11_), .Y(_abc_19068_n1193) );
  AND2X2 AND2X2_1820 ( .A(core__abc_21380_n2130), .B(reset_n_bF_buf44), .Y(core__abc_21380_n2131) );
  AND2X2 AND2X2_1821 ( .A(core__abc_21380_n2129), .B(core__abc_21380_n2131), .Y(core_siphash_word1_reg_46__FF_INPUT) );
  AND2X2 AND2X2_1822 ( .A(core_v0_reg_47_), .B(core_v1_reg_47_), .Y(core__abc_21380_n2133) );
  AND2X2 AND2X2_1823 ( .A(core__abc_21380_n2135), .B(core__abc_21380_n2136), .Y(core__abc_21380_n2137) );
  AND2X2 AND2X2_1824 ( .A(core__abc_21380_n2138), .B(core__abc_21380_n2134), .Y(core__abc_21380_n2139_1) );
  AND2X2 AND2X2_1825 ( .A(core_v2_reg_47_), .B(core_v3_reg_47_), .Y(core__abc_21380_n2142) );
  AND2X2 AND2X2_1826 ( .A(core__abc_21380_n2143_1), .B(core__abc_21380_n2141), .Y(core__abc_21380_n2144) );
  AND2X2 AND2X2_1827 ( .A(core__abc_21380_n2140), .B(core__abc_21380_n2144), .Y(core__abc_21380_n2145) );
  AND2X2 AND2X2_1828 ( .A(core__abc_21380_n2146), .B(core__abc_21380_n2139_1), .Y(core__abc_21380_n2147) );
  AND2X2 AND2X2_1829 ( .A(core__abc_21380_n2150), .B(reset_n_bF_buf43), .Y(core__abc_21380_n2151) );
  AND2X2 AND2X2_183 ( .A(_abc_19068_n915_1_bF_buf2), .B(core_mi_43_), .Y(_abc_19068_n1195_1) );
  AND2X2 AND2X2_1830 ( .A(core__abc_21380_n2149), .B(core__abc_21380_n2151), .Y(core_siphash_word1_reg_47__FF_INPUT) );
  AND2X2 AND2X2_1831 ( .A(core__abc_21380_n2153), .B(core__abc_21380_n2154), .Y(core__abc_21380_n2155) );
  AND2X2 AND2X2_1832 ( .A(core_v0_reg_48_), .B(core_v1_reg_48_), .Y(core__abc_21380_n2156) );
  AND2X2 AND2X2_1833 ( .A(core_v2_reg_48_), .B(core_v3_reg_48_), .Y(core__abc_21380_n2160) );
  AND2X2 AND2X2_1834 ( .A(core__abc_21380_n2161), .B(core__abc_21380_n2159), .Y(core__abc_21380_n2162) );
  AND2X2 AND2X2_1835 ( .A(core__abc_21380_n2163), .B(core__abc_21380_n2165), .Y(core__abc_21380_n2166) );
  AND2X2 AND2X2_1836 ( .A(core__abc_21380_n2168), .B(reset_n_bF_buf42), .Y(core__abc_21380_n2169) );
  AND2X2 AND2X2_1837 ( .A(core__abc_21380_n2167), .B(core__abc_21380_n2169), .Y(core_siphash_word1_reg_48__FF_INPUT) );
  AND2X2 AND2X2_1838 ( .A(core_v0_reg_49_), .B(core_v1_reg_49_), .Y(core__abc_21380_n2171) );
  AND2X2 AND2X2_1839 ( .A(core__abc_21380_n2172), .B(core__abc_21380_n2173), .Y(core__abc_21380_n2174) );
  AND2X2 AND2X2_184 ( .A(_abc_19068_n897_1_bF_buf2), .B(word0_reg_11_), .Y(_abc_19068_n1196) );
  AND2X2 AND2X2_1840 ( .A(core_v2_reg_49_), .B(core_v3_reg_49_), .Y(core__abc_21380_n2177) );
  AND2X2 AND2X2_1841 ( .A(core__abc_21380_n2178), .B(core__abc_21380_n2176), .Y(core__abc_21380_n2179_1) );
  AND2X2 AND2X2_1842 ( .A(core__abc_21380_n2175), .B(core__abc_21380_n2179_1), .Y(core__abc_21380_n2180) );
  AND2X2 AND2X2_1843 ( .A(core__abc_21380_n2181), .B(core__abc_21380_n2182), .Y(core__abc_21380_n2183) );
  AND2X2 AND2X2_1844 ( .A(core__abc_21380_n2186), .B(reset_n_bF_buf41), .Y(core__abc_21380_n2187) );
  AND2X2 AND2X2_1845 ( .A(core__abc_21380_n2185_1), .B(core__abc_21380_n2187), .Y(core_siphash_word1_reg_49__FF_INPUT) );
  AND2X2 AND2X2_1846 ( .A(core_v0_reg_50_), .B(core_v1_reg_50_), .Y(core__abc_21380_n2189) );
  AND2X2 AND2X2_1847 ( .A(core__abc_21380_n2190), .B(core__abc_21380_n2191), .Y(core__abc_21380_n2192) );
  AND2X2 AND2X2_1848 ( .A(core_v2_reg_50_), .B(core_v3_reg_50_), .Y(core__abc_21380_n2195) );
  AND2X2 AND2X2_1849 ( .A(core__abc_21380_n2196), .B(core__abc_21380_n2194), .Y(core__abc_21380_n2197) );
  AND2X2 AND2X2_185 ( .A(_abc_19068_n923_bF_buf3), .B(_abc_19068_n1200_1), .Y(_auto_iopadmap_cc_313_execute_30317_11_) );
  AND2X2 AND2X2_1850 ( .A(core__abc_21380_n2193), .B(core__abc_21380_n2197), .Y(core__abc_21380_n2198) );
  AND2X2 AND2X2_1851 ( .A(core__abc_21380_n2199), .B(core__abc_21380_n2200), .Y(core__abc_21380_n2201) );
  AND2X2 AND2X2_1852 ( .A(core__abc_21380_n2204), .B(reset_n_bF_buf40), .Y(core__abc_21380_n2205) );
  AND2X2 AND2X2_1853 ( .A(core__abc_21380_n2203), .B(core__abc_21380_n2205), .Y(core_siphash_word1_reg_50__FF_INPUT) );
  AND2X2 AND2X2_1854 ( .A(core_v0_reg_51_), .B(core_v1_reg_51_), .Y(core__abc_21380_n2207) );
  AND2X2 AND2X2_1855 ( .A(core__abc_21380_n2209), .B(core__abc_21380_n2210), .Y(core__abc_21380_n2211) );
  AND2X2 AND2X2_1856 ( .A(core__abc_21380_n2212), .B(core__abc_21380_n2208), .Y(core__abc_21380_n2213_1) );
  AND2X2 AND2X2_1857 ( .A(core_v3_reg_51_), .B(core_v2_reg_51_), .Y(core__abc_21380_n2216) );
  AND2X2 AND2X2_1858 ( .A(core__abc_21380_n2217), .B(core__abc_21380_n2215), .Y(core__abc_21380_n2218) );
  AND2X2 AND2X2_1859 ( .A(core__abc_21380_n2214), .B(core__abc_21380_n2218), .Y(core__abc_21380_n2219_1) );
  AND2X2 AND2X2_186 ( .A(_abc_19068_n916_1_bF_buf1), .B(word1_reg_12_), .Y(_abc_19068_n1202) );
  AND2X2 AND2X2_1860 ( .A(core__abc_21380_n2220), .B(core__abc_21380_n2213_1), .Y(core__abc_21380_n2221) );
  AND2X2 AND2X2_1861 ( .A(core__abc_21380_n2224), .B(reset_n_bF_buf39), .Y(core__abc_21380_n2225) );
  AND2X2 AND2X2_1862 ( .A(core__abc_21380_n2223), .B(core__abc_21380_n2225), .Y(core_siphash_word1_reg_51__FF_INPUT) );
  AND2X2 AND2X2_1863 ( .A(core_v0_reg_52_), .B(core_v1_reg_52_), .Y(core__abc_21380_n2228) );
  AND2X2 AND2X2_1864 ( .A(core__abc_21380_n2229), .B(core__abc_21380_n2227), .Y(core__abc_21380_n2230) );
  AND2X2 AND2X2_1865 ( .A(core_v3_reg_52_), .B(core_v2_reg_52_), .Y(core__abc_21380_n2232) );
  AND2X2 AND2X2_1866 ( .A(core__abc_21380_n2233), .B(core__abc_21380_n2231), .Y(core__abc_21380_n2234) );
  AND2X2 AND2X2_1867 ( .A(core__abc_21380_n2238), .B(core__abc_21380_n2235), .Y(core__abc_21380_n2239) );
  AND2X2 AND2X2_1868 ( .A(core__abc_21380_n2241), .B(reset_n_bF_buf38), .Y(core__abc_21380_n2242) );
  AND2X2 AND2X2_1869 ( .A(core__abc_21380_n2240), .B(core__abc_21380_n2242), .Y(core_siphash_word1_reg_52__FF_INPUT) );
  AND2X2 AND2X2_187 ( .A(_abc_19068_n897_1_bF_buf1), .B(word0_reg_12_), .Y(_abc_19068_n1203_1) );
  AND2X2 AND2X2_1870 ( .A(core_v0_reg_53_), .B(core_v1_reg_53_), .Y(core__abc_21380_n2244) );
  AND2X2 AND2X2_1871 ( .A(core__abc_21380_n2246), .B(core__abc_21380_n2247_1), .Y(core__abc_21380_n2248) );
  AND2X2 AND2X2_1872 ( .A(core__abc_21380_n2249), .B(core__abc_21380_n2245), .Y(core__abc_21380_n2250) );
  AND2X2 AND2X2_1873 ( .A(core_v3_reg_53_), .B(core_v2_reg_53_), .Y(core__abc_21380_n2253) );
  AND2X2 AND2X2_1874 ( .A(core__abc_21380_n2254), .B(core__abc_21380_n2252), .Y(core__abc_21380_n2255) );
  AND2X2 AND2X2_1875 ( .A(core__abc_21380_n2251), .B(core__abc_21380_n2255), .Y(core__abc_21380_n2256) );
  AND2X2 AND2X2_1876 ( .A(core__abc_21380_n2257), .B(core__abc_21380_n2250), .Y(core__abc_21380_n2258) );
  AND2X2 AND2X2_1877 ( .A(core__abc_21380_n2261), .B(reset_n_bF_buf37), .Y(core__abc_21380_n2262) );
  AND2X2 AND2X2_1878 ( .A(core__abc_21380_n2260), .B(core__abc_21380_n2262), .Y(core_siphash_word1_reg_53__FF_INPUT) );
  AND2X2 AND2X2_1879 ( .A(core__abc_21380_n2264), .B(core__abc_21380_n2265), .Y(core__abc_21380_n2266) );
  AND2X2 AND2X2_188 ( .A(_abc_19068_n915_1_bF_buf1), .B(core_mi_44_), .Y(_abc_19068_n1205) );
  AND2X2 AND2X2_1880 ( .A(core_v0_reg_54_), .B(core_v1_reg_54_), .Y(core__abc_21380_n2267) );
  AND2X2 AND2X2_1881 ( .A(core_v3_reg_54_), .B(core_v2_reg_54_), .Y(core__abc_21380_n2271) );
  AND2X2 AND2X2_1882 ( .A(core__abc_21380_n2272), .B(core__abc_21380_n2270), .Y(core__abc_21380_n2273) );
  AND2X2 AND2X2_1883 ( .A(core__abc_21380_n2274), .B(core__abc_21380_n2276), .Y(core__abc_21380_n2277) );
  AND2X2 AND2X2_1884 ( .A(core__abc_21380_n2279), .B(reset_n_bF_buf36), .Y(core__abc_21380_n2280) );
  AND2X2 AND2X2_1885 ( .A(core__abc_21380_n2278), .B(core__abc_21380_n2280), .Y(core_siphash_word1_reg_54__FF_INPUT) );
  AND2X2 AND2X2_1886 ( .A(core__abc_21380_n2282), .B(core__abc_21380_n2283), .Y(core__abc_21380_n2284) );
  AND2X2 AND2X2_1887 ( .A(core_v0_reg_55_), .B(core_v1_reg_55_), .Y(core__abc_21380_n2286) );
  AND2X2 AND2X2_1888 ( .A(core__abc_21380_n2285), .B(core__abc_21380_n2287), .Y(core__abc_21380_n2288) );
  AND2X2 AND2X2_1889 ( .A(core_v3_reg_55_), .B(core_v2_reg_55_), .Y(core__abc_21380_n2290) );
  AND2X2 AND2X2_189 ( .A(_abc_19068_n945_1_bF_buf2), .B(core_mi_12_), .Y(_abc_19068_n1206_1) );
  AND2X2 AND2X2_1890 ( .A(core__abc_21380_n2291), .B(core__abc_21380_n2289), .Y(core__abc_21380_n2292) );
  AND2X2 AND2X2_1891 ( .A(core__abc_21380_n2296), .B(core__abc_21380_n2293), .Y(core__abc_21380_n2297) );
  AND2X2 AND2X2_1892 ( .A(core__abc_21380_n2299), .B(reset_n_bF_buf35), .Y(core__abc_21380_n2300) );
  AND2X2 AND2X2_1893 ( .A(core__abc_21380_n2298_1), .B(core__abc_21380_n2300), .Y(core_siphash_word1_reg_55__FF_INPUT) );
  AND2X2 AND2X2_1894 ( .A(core__abc_21380_n2302), .B(core__abc_21380_n2303), .Y(core__abc_21380_n2304) );
  AND2X2 AND2X2_1895 ( .A(core_v0_reg_56_), .B(core_v1_reg_56_), .Y(core__abc_21380_n2305) );
  AND2X2 AND2X2_1896 ( .A(core_v2_reg_56_), .B(core_v3_reg_56_), .Y(core__abc_21380_n2309) );
  AND2X2 AND2X2_1897 ( .A(core__abc_21380_n2310), .B(core__abc_21380_n2308), .Y(core__abc_21380_n2311) );
  AND2X2 AND2X2_1898 ( .A(core__abc_21380_n2312), .B(core__abc_21380_n2314), .Y(core__abc_21380_n2315) );
  AND2X2 AND2X2_1899 ( .A(core__abc_21380_n2317), .B(reset_n_bF_buf34), .Y(core__abc_21380_n2318) );
  AND2X2 AND2X2_19 ( .A(_abc_19068_n893), .B(_abc_19068_n883_1), .Y(_abc_19068_n898_1) );
  AND2X2 AND2X2_190 ( .A(_abc_19068_n926_bF_buf2), .B(core_key_12_), .Y(_abc_19068_n1210_1) );
  AND2X2 AND2X2_1900 ( .A(core__abc_21380_n2316), .B(core__abc_21380_n2318), .Y(core_siphash_word1_reg_56__FF_INPUT) );
  AND2X2 AND2X2_1901 ( .A(core__abc_21380_n2320), .B(core__abc_21380_n2321), .Y(core__abc_21380_n2322) );
  AND2X2 AND2X2_1902 ( .A(core_v0_reg_57_), .B(core_v1_reg_57_), .Y(core__abc_21380_n2323) );
  AND2X2 AND2X2_1903 ( .A(core_v2_reg_57_), .B(core_v3_reg_57_), .Y(core__abc_21380_n2327) );
  AND2X2 AND2X2_1904 ( .A(core__abc_21380_n2328_1), .B(core__abc_21380_n2326), .Y(core__abc_21380_n2329) );
  AND2X2 AND2X2_1905 ( .A(core__abc_21380_n2330), .B(core__abc_21380_n2332_1), .Y(core__abc_21380_n2333) );
  AND2X2 AND2X2_1906 ( .A(core__abc_21380_n2335), .B(reset_n_bF_buf33), .Y(core__abc_21380_n2336) );
  AND2X2 AND2X2_1907 ( .A(core__abc_21380_n2334), .B(core__abc_21380_n2336), .Y(core_siphash_word1_reg_57__FF_INPUT) );
  AND2X2 AND2X2_1908 ( .A(core__abc_21380_n2338), .B(core__abc_21380_n2339), .Y(core__abc_21380_n2340) );
  AND2X2 AND2X2_1909 ( .A(core_v0_reg_58_), .B(core_v1_reg_58_), .Y(core__abc_21380_n2341) );
  AND2X2 AND2X2_191 ( .A(_abc_19068_n924_1_bF_buf2), .B(core_key_44_), .Y(_abc_19068_n1211) );
  AND2X2 AND2X2_1910 ( .A(core_v3_reg_58_), .B(core_v2_reg_58_), .Y(core__abc_21380_n2345) );
  AND2X2 AND2X2_1911 ( .A(core__abc_21380_n2346), .B(core__abc_21380_n2344), .Y(core__abc_21380_n2347) );
  AND2X2 AND2X2_1912 ( .A(core__abc_21380_n2348), .B(core__abc_21380_n2350), .Y(core__abc_21380_n2351) );
  AND2X2 AND2X2_1913 ( .A(core__abc_21380_n2353), .B(reset_n_bF_buf32), .Y(core__abc_21380_n2354) );
  AND2X2 AND2X2_1914 ( .A(core__abc_21380_n2352), .B(core__abc_21380_n2354), .Y(core_siphash_word1_reg_58__FF_INPUT) );
  AND2X2 AND2X2_1915 ( .A(core__abc_21380_n2356), .B(core__abc_21380_n2357), .Y(core__abc_21380_n2358) );
  AND2X2 AND2X2_1916 ( .A(core_v0_reg_59_), .B(core_v1_reg_59_), .Y(core__abc_21380_n2360) );
  AND2X2 AND2X2_1917 ( .A(core__abc_21380_n2359), .B(core__abc_21380_n2361), .Y(core__abc_21380_n2362) );
  AND2X2 AND2X2_1918 ( .A(core_v3_reg_59_), .B(core_v2_reg_59_), .Y(core__abc_21380_n2364) );
  AND2X2 AND2X2_1919 ( .A(core__abc_21380_n2365), .B(core__abc_21380_n2363_1), .Y(core__abc_21380_n2366) );
  AND2X2 AND2X2_192 ( .A(_abc_19068_n902_bF_buf1), .B(word2_reg_12_), .Y(_abc_19068_n1214) );
  AND2X2 AND2X2_1920 ( .A(core__abc_21380_n2370), .B(core__abc_21380_n2367), .Y(core__abc_21380_n2371) );
  AND2X2 AND2X2_1921 ( .A(core__abc_21380_n2373), .B(reset_n_bF_buf31), .Y(core__abc_21380_n2374) );
  AND2X2 AND2X2_1922 ( .A(core__abc_21380_n2372), .B(core__abc_21380_n2374), .Y(core_siphash_word1_reg_59__FF_INPUT) );
  AND2X2 AND2X2_1923 ( .A(core__abc_21380_n2376), .B(core__abc_21380_n2377), .Y(core__abc_21380_n2378) );
  AND2X2 AND2X2_1924 ( .A(core_v0_reg_60_), .B(core_v1_reg_60_), .Y(core__abc_21380_n2379) );
  AND2X2 AND2X2_1925 ( .A(core_v3_reg_60_), .B(core_v2_reg_60_), .Y(core__abc_21380_n2383) );
  AND2X2 AND2X2_1926 ( .A(core__abc_21380_n2384), .B(core__abc_21380_n2382), .Y(core__abc_21380_n2385) );
  AND2X2 AND2X2_1927 ( .A(core__abc_21380_n2386), .B(core__abc_21380_n2388), .Y(core__abc_21380_n2389) );
  AND2X2 AND2X2_1928 ( .A(core__abc_21380_n2391_1), .B(reset_n_bF_buf30), .Y(core__abc_21380_n2392) );
  AND2X2 AND2X2_1929 ( .A(core__abc_21380_n2390), .B(core__abc_21380_n2392), .Y(core_siphash_word1_reg_60__FF_INPUT) );
  AND2X2 AND2X2_193 ( .A(_abc_19068_n899_bF_buf1), .B(word3_reg_12_), .Y(_abc_19068_n1215_1) );
  AND2X2 AND2X2_1930 ( .A(core__abc_21380_n2394), .B(core__abc_21380_n2395_1), .Y(core__abc_21380_n2396) );
  AND2X2 AND2X2_1931 ( .A(core_v0_reg_61_), .B(core_v1_reg_61_), .Y(core__abc_21380_n2397) );
  AND2X2 AND2X2_1932 ( .A(core_v3_reg_61_), .B(core_v2_reg_61_), .Y(core__abc_21380_n2401) );
  AND2X2 AND2X2_1933 ( .A(core__abc_21380_n2402), .B(core__abc_21380_n2400), .Y(core__abc_21380_n2403) );
  AND2X2 AND2X2_1934 ( .A(core__abc_21380_n2404), .B(core__abc_21380_n2406), .Y(core__abc_21380_n2407) );
  AND2X2 AND2X2_1935 ( .A(core__abc_21380_n2409), .B(reset_n_bF_buf29), .Y(core__abc_21380_n2410) );
  AND2X2 AND2X2_1936 ( .A(core__abc_21380_n2408), .B(core__abc_21380_n2410), .Y(core_siphash_word1_reg_61__FF_INPUT) );
  AND2X2 AND2X2_1937 ( .A(core__abc_21380_n2412), .B(core__abc_21380_n2413), .Y(core__abc_21380_n2414) );
  AND2X2 AND2X2_1938 ( .A(core_v0_reg_62_), .B(core_v1_reg_62_), .Y(core__abc_21380_n2415) );
  AND2X2 AND2X2_1939 ( .A(core_v3_reg_62_), .B(core_v2_reg_62_), .Y(core__abc_21380_n2419) );
  AND2X2 AND2X2_194 ( .A(_abc_19068_n939_1_bF_buf2), .B(core_key_76_), .Y(_abc_19068_n1217) );
  AND2X2 AND2X2_1940 ( .A(core__abc_21380_n2420), .B(core__abc_21380_n2418), .Y(core__abc_21380_n2421) );
  AND2X2 AND2X2_1941 ( .A(core__abc_21380_n2422), .B(core__abc_21380_n2424_1), .Y(core__abc_21380_n2425) );
  AND2X2 AND2X2_1942 ( .A(core__abc_21380_n2427), .B(reset_n_bF_buf28), .Y(core__abc_21380_n2428) );
  AND2X2 AND2X2_1943 ( .A(core__abc_21380_n2426), .B(core__abc_21380_n2428), .Y(core_siphash_word1_reg_62__FF_INPUT) );
  AND2X2 AND2X2_1944 ( .A(core__abc_21380_n2431), .B(core__abc_21380_n2433), .Y(core__abc_21380_n2434) );
  AND2X2 AND2X2_1945 ( .A(core_v3_reg_63_), .B(core_v2_reg_63_), .Y(core__abc_21380_n2437) );
  AND2X2 AND2X2_1946 ( .A(core__abc_21380_n2438), .B(core__abc_21380_n2436), .Y(core__abc_21380_n2439) );
  AND2X2 AND2X2_1947 ( .A(core__abc_21380_n2435), .B(core__abc_21380_n2440), .Y(core__abc_21380_n2441) );
  AND2X2 AND2X2_1948 ( .A(core__abc_21380_n2434), .B(core__abc_21380_n2439), .Y(core__abc_21380_n2442) );
  AND2X2 AND2X2_1949 ( .A(core__abc_21380_n2445_1), .B(reset_n_bF_buf27), .Y(core__abc_21380_n2446) );
  AND2X2 AND2X2_195 ( .A(_abc_19068_n941_bF_buf2), .B(core_key_108_), .Y(_abc_19068_n1218_1) );
  AND2X2 AND2X2_1950 ( .A(core__abc_21380_n2444), .B(core__abc_21380_n2446), .Y(core_siphash_word1_reg_63__FF_INPUT) );
  AND2X2 AND2X2_1951 ( .A(core__abc_21380_n1142_1), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n2448) );
  AND2X2 AND2X2_1952 ( .A(core__abc_21380_n1136_1), .B(core__abc_21380_n2449), .Y(core__abc_21380_n2450) );
  AND2X2 AND2X2_1953 ( .A(core__abc_21380_n2448), .B(core__abc_21380_n2450), .Y(core__abc_21380_n2451_1) );
  AND2X2 AND2X2_1954 ( .A(core__abc_21380_n2454), .B(reset_n_bF_buf26), .Y(core__abc_21380_n2455) );
  AND2X2 AND2X2_1955 ( .A(core__abc_21380_n2455), .B(core__abc_21380_n2453), .Y(core_siphash_word0_reg_0__FF_INPUT) );
  AND2X2 AND2X2_1956 ( .A(core__abc_21380_n2458), .B(reset_n_bF_buf25), .Y(core__abc_21380_n2459) );
  AND2X2 AND2X2_1957 ( .A(core__abc_21380_n2459), .B(core__abc_21380_n2457), .Y(core_siphash_word0_reg_1__FF_INPUT) );
  AND2X2 AND2X2_1958 ( .A(core__abc_21380_n2462), .B(reset_n_bF_buf24), .Y(core__abc_21380_n2463) );
  AND2X2 AND2X2_1959 ( .A(core__abc_21380_n2463), .B(core__abc_21380_n2461), .Y(core_siphash_word0_reg_2__FF_INPUT) );
  AND2X2 AND2X2_196 ( .A(_abc_19068_n923_bF_buf2), .B(_abc_19068_n1222_1), .Y(_auto_iopadmap_cc_313_execute_30317_12_) );
  AND2X2 AND2X2_1960 ( .A(core__abc_21380_n1331), .B(core__abc_21380_n2451_1_bF_buf3), .Y(core__abc_21380_n2465) );
  AND2X2 AND2X2_1961 ( .A(core__abc_21380_n2452_bF_buf4), .B(core_siphash_word_3_), .Y(core__abc_21380_n2466) );
  AND2X2 AND2X2_1962 ( .A(core__abc_21380_n2467), .B(reset_n_bF_buf23), .Y(core_siphash_word0_reg_3__FF_INPUT) );
  AND2X2 AND2X2_1963 ( .A(core__abc_21380_n2470), .B(reset_n_bF_buf22), .Y(core__abc_21380_n2471_1) );
  AND2X2 AND2X2_1964 ( .A(core__abc_21380_n2471_1), .B(core__abc_21380_n2469), .Y(core_siphash_word0_reg_4__FF_INPUT) );
  AND2X2 AND2X2_1965 ( .A(core__abc_21380_n1368), .B(core__abc_21380_n2451_1_bF_buf1), .Y(core__abc_21380_n2473) );
  AND2X2 AND2X2_1966 ( .A(core__abc_21380_n2452_bF_buf2), .B(core_siphash_word_5_), .Y(core__abc_21380_n2474) );
  AND2X2 AND2X2_1967 ( .A(core__abc_21380_n2475), .B(reset_n_bF_buf21), .Y(core_siphash_word0_reg_5__FF_INPUT) );
  AND2X2 AND2X2_1968 ( .A(core__abc_21380_n2478), .B(reset_n_bF_buf20), .Y(core__abc_21380_n2479) );
  AND2X2 AND2X2_1969 ( .A(core__abc_21380_n2479), .B(core__abc_21380_n2477_1), .Y(core_siphash_word0_reg_6__FF_INPUT) );
  AND2X2 AND2X2_197 ( .A(_abc_19068_n941_bF_buf1), .B(core_key_109_), .Y(_abc_19068_n1224_1) );
  AND2X2 AND2X2_1970 ( .A(core__abc_21380_n2482), .B(reset_n_bF_buf19), .Y(core__abc_21380_n2483) );
  AND2X2 AND2X2_1971 ( .A(core__abc_21380_n2483), .B(core__abc_21380_n2481), .Y(core_siphash_word0_reg_7__FF_INPUT) );
  AND2X2 AND2X2_1972 ( .A(core__abc_21380_n1423), .B(core__abc_21380_n2451_1_bF_buf6), .Y(core__abc_21380_n2485) );
  AND2X2 AND2X2_1973 ( .A(core__abc_21380_n2452_bF_buf7), .B(core_siphash_word_8_), .Y(core__abc_21380_n2486) );
  AND2X2 AND2X2_1974 ( .A(core__abc_21380_n2487), .B(reset_n_bF_buf18), .Y(core_siphash_word0_reg_8__FF_INPUT) );
  AND2X2 AND2X2_1975 ( .A(core__abc_21380_n2490), .B(reset_n_bF_buf17), .Y(core__abc_21380_n2491) );
  AND2X2 AND2X2_1976 ( .A(core__abc_21380_n2489), .B(core__abc_21380_n2491), .Y(core_siphash_word0_reg_9__FF_INPUT) );
  AND2X2 AND2X2_1977 ( .A(core__abc_21380_n2494), .B(reset_n_bF_buf16), .Y(core__abc_21380_n2495) );
  AND2X2 AND2X2_1978 ( .A(core__abc_21380_n2495), .B(core__abc_21380_n2493_1), .Y(core_siphash_word0_reg_10__FF_INPUT) );
  AND2X2 AND2X2_1979 ( .A(core__abc_21380_n2498), .B(reset_n_bF_buf15), .Y(core__abc_21380_n2499) );
  AND2X2 AND2X2_198 ( .A(_abc_19068_n899_bF_buf0), .B(word3_reg_13_), .Y(_abc_19068_n1225_1) );
  AND2X2 AND2X2_1980 ( .A(core__abc_21380_n2499), .B(core__abc_21380_n2497_1), .Y(core_siphash_word0_reg_11__FF_INPUT) );
  AND2X2 AND2X2_1981 ( .A(core__abc_21380_n1495), .B(core__abc_21380_n2451_1_bF_buf2), .Y(core__abc_21380_n2501) );
  AND2X2 AND2X2_1982 ( .A(core__abc_21380_n2452_bF_buf3), .B(core_siphash_word_12_), .Y(core__abc_21380_n2502) );
  AND2X2 AND2X2_1983 ( .A(core__abc_21380_n2503), .B(reset_n_bF_buf14), .Y(core_siphash_word0_reg_12__FF_INPUT) );
  AND2X2 AND2X2_1984 ( .A(core__abc_21380_n2506), .B(reset_n_bF_buf13), .Y(core__abc_21380_n2507) );
  AND2X2 AND2X2_1985 ( .A(core__abc_21380_n2507), .B(core__abc_21380_n2505), .Y(core_siphash_word0_reg_13__FF_INPUT) );
  AND2X2 AND2X2_1986 ( .A(core__abc_21380_n2510), .B(reset_n_bF_buf12), .Y(core__abc_21380_n2511) );
  AND2X2 AND2X2_1987 ( .A(core__abc_21380_n2511), .B(core__abc_21380_n2509), .Y(core_siphash_word0_reg_14__FF_INPUT) );
  AND2X2 AND2X2_1988 ( .A(core__abc_21380_n2514), .B(reset_n_bF_buf11), .Y(core__abc_21380_n2515) );
  AND2X2 AND2X2_1989 ( .A(core__abc_21380_n2513), .B(core__abc_21380_n2515), .Y(core_siphash_word0_reg_15__FF_INPUT) );
  AND2X2 AND2X2_199 ( .A(_abc_19068_n902_bF_buf0), .B(word2_reg_13_), .Y(_abc_19068_n1226) );
  AND2X2 AND2X2_1990 ( .A(core__abc_21380_n1569), .B(core__abc_21380_n2451_1_bF_buf6), .Y(core__abc_21380_n2517) );
  AND2X2 AND2X2_1991 ( .A(core__abc_21380_n2452_bF_buf7), .B(core_siphash_word_16_), .Y(core__abc_21380_n2518) );
  AND2X2 AND2X2_1992 ( .A(core__abc_21380_n2519), .B(reset_n_bF_buf10), .Y(core_siphash_word0_reg_16__FF_INPUT) );
  AND2X2 AND2X2_1993 ( .A(core__abc_21380_n2522), .B(reset_n_bF_buf9), .Y(core__abc_21380_n2523) );
  AND2X2 AND2X2_1994 ( .A(core__abc_21380_n2521), .B(core__abc_21380_n2523), .Y(core_siphash_word0_reg_17__FF_INPUT) );
  AND2X2 AND2X2_1995 ( .A(core__abc_21380_n2526), .B(reset_n_bF_buf8), .Y(core__abc_21380_n2527) );
  AND2X2 AND2X2_1996 ( .A(core__abc_21380_n2527), .B(core__abc_21380_n2525), .Y(core_siphash_word0_reg_18__FF_INPUT) );
  AND2X2 AND2X2_1997 ( .A(core__abc_21380_n1623), .B(core__abc_21380_n2451_1_bF_buf3), .Y(core__abc_21380_n2529) );
  AND2X2 AND2X2_1998 ( .A(core__abc_21380_n2452_bF_buf4), .B(core_siphash_word_19_), .Y(core__abc_21380_n2530) );
  AND2X2 AND2X2_1999 ( .A(core__abc_21380_n2531), .B(reset_n_bF_buf7), .Y(core_siphash_word0_reg_19__FF_INPUT) );
  AND2X2 AND2X2_2 ( .A(_abc_19068_n872), .B(\addr[0] ), .Y(_abc_19068_n873_1) );
  AND2X2 AND2X2_20 ( .A(_abc_19068_n898_1), .B(_abc_19068_n896), .Y(_abc_19068_n899) );
  AND2X2 AND2X2_200 ( .A(_abc_19068_n915_1_bF_buf0), .B(core_mi_45_), .Y(_abc_19068_n1228_1) );
  AND2X2 AND2X2_2000 ( .A(core__abc_21380_n2534_1), .B(reset_n_bF_buf6), .Y(core__abc_21380_n2535) );
  AND2X2 AND2X2_2001 ( .A(core__abc_21380_n2535), .B(core__abc_21380_n2533), .Y(core_siphash_word0_reg_20__FF_INPUT) );
  AND2X2 AND2X2_2002 ( .A(core__abc_21380_n2538), .B(reset_n_bF_buf5), .Y(core__abc_21380_n2539) );
  AND2X2 AND2X2_2003 ( .A(core__abc_21380_n2539), .B(core__abc_21380_n2537), .Y(core_siphash_word0_reg_21__FF_INPUT) );
  AND2X2 AND2X2_2004 ( .A(core__abc_21380_n2542), .B(reset_n_bF_buf4), .Y(core__abc_21380_n2543) );
  AND2X2 AND2X2_2005 ( .A(core__abc_21380_n2543), .B(core__abc_21380_n2541), .Y(core_siphash_word0_reg_22__FF_INPUT) );
  AND2X2 AND2X2_2006 ( .A(core__abc_21380_n2546), .B(reset_n_bF_buf3), .Y(core__abc_21380_n2547) );
  AND2X2 AND2X2_2007 ( .A(core__abc_21380_n2545), .B(core__abc_21380_n2547), .Y(core_siphash_word0_reg_23__FF_INPUT) );
  AND2X2 AND2X2_2008 ( .A(core__abc_21380_n2550), .B(reset_n_bF_buf2), .Y(core__abc_21380_n2551_1) );
  AND2X2 AND2X2_2009 ( .A(core__abc_21380_n2551_1), .B(core__abc_21380_n2549), .Y(core_siphash_word0_reg_24__FF_INPUT) );
  AND2X2 AND2X2_201 ( .A(_abc_19068_n945_1_bF_buf1), .B(core_mi_13_), .Y(_abc_19068_n1229) );
  AND2X2 AND2X2_2010 ( .A(core__abc_21380_n2554), .B(reset_n_bF_buf1), .Y(core__abc_21380_n2555_1) );
  AND2X2 AND2X2_2011 ( .A(core__abc_21380_n2553), .B(core__abc_21380_n2555_1), .Y(core_siphash_word0_reg_25__FF_INPUT) );
  AND2X2 AND2X2_2012 ( .A(core__abc_21380_n2558), .B(reset_n_bF_buf0), .Y(core__abc_21380_n2559) );
  AND2X2 AND2X2_2013 ( .A(core__abc_21380_n2559), .B(core__abc_21380_n2557), .Y(core_siphash_word0_reg_26__FF_INPUT) );
  AND2X2 AND2X2_2014 ( .A(core__abc_21380_n2562), .B(reset_n_bF_buf84), .Y(core__abc_21380_n2563) );
  AND2X2 AND2X2_2015 ( .A(core__abc_21380_n2561), .B(core__abc_21380_n2563), .Y(core_siphash_word0_reg_27__FF_INPUT) );
  AND2X2 AND2X2_2016 ( .A(core__abc_21380_n2566), .B(reset_n_bF_buf83), .Y(core__abc_21380_n2567) );
  AND2X2 AND2X2_2017 ( .A(core__abc_21380_n2567), .B(core__abc_21380_n2565), .Y(core_siphash_word0_reg_28__FF_INPUT) );
  AND2X2 AND2X2_2018 ( .A(core__abc_21380_n2570), .B(reset_n_bF_buf82), .Y(core__abc_21380_n2571) );
  AND2X2 AND2X2_2019 ( .A(core__abc_21380_n2569), .B(core__abc_21380_n2571), .Y(core_siphash_word0_reg_29__FF_INPUT) );
  AND2X2 AND2X2_202 ( .A(_abc_19068_n926_bF_buf1), .B(core_key_13_), .Y(_abc_19068_n1233_1) );
  AND2X2 AND2X2_2020 ( .A(core__abc_21380_n2574), .B(reset_n_bF_buf81), .Y(core__abc_21380_n2575) );
  AND2X2 AND2X2_2021 ( .A(core__abc_21380_n2575), .B(core__abc_21380_n2573), .Y(core_siphash_word0_reg_30__FF_INPUT) );
  AND2X2 AND2X2_2022 ( .A(core__abc_21380_n2578_1), .B(reset_n_bF_buf80), .Y(core__abc_21380_n2579) );
  AND2X2 AND2X2_2023 ( .A(core__abc_21380_n2577), .B(core__abc_21380_n2579), .Y(core_siphash_word0_reg_31__FF_INPUT) );
  AND2X2 AND2X2_2024 ( .A(core__abc_21380_n2582_1), .B(reset_n_bF_buf79), .Y(core__abc_21380_n2583) );
  AND2X2 AND2X2_2025 ( .A(core__abc_21380_n2583), .B(core__abc_21380_n2581), .Y(core_siphash_word0_reg_32__FF_INPUT) );
  AND2X2 AND2X2_2026 ( .A(core__abc_21380_n2586), .B(reset_n_bF_buf78), .Y(core__abc_21380_n2587) );
  AND2X2 AND2X2_2027 ( .A(core__abc_21380_n2587), .B(core__abc_21380_n2585), .Y(core_siphash_word0_reg_33__FF_INPUT) );
  AND2X2 AND2X2_2028 ( .A(core__abc_21380_n2590), .B(reset_n_bF_buf77), .Y(core__abc_21380_n2591) );
  AND2X2 AND2X2_2029 ( .A(core__abc_21380_n2591), .B(core__abc_21380_n2589), .Y(core_siphash_word0_reg_34__FF_INPUT) );
  AND2X2 AND2X2_203 ( .A(_abc_19068_n924_1_bF_buf1), .B(core_key_45_), .Y(_abc_19068_n1234) );
  AND2X2 AND2X2_2030 ( .A(core__abc_21380_n2594), .B(reset_n_bF_buf76), .Y(core__abc_21380_n2595) );
  AND2X2 AND2X2_2031 ( .A(core__abc_21380_n2593), .B(core__abc_21380_n2595), .Y(core_siphash_word0_reg_35__FF_INPUT) );
  AND2X2 AND2X2_2032 ( .A(core__abc_21380_n2598), .B(reset_n_bF_buf75), .Y(core__abc_21380_n2599) );
  AND2X2 AND2X2_2033 ( .A(core__abc_21380_n2599), .B(core__abc_21380_n2597_1), .Y(core_siphash_word0_reg_36__FF_INPUT) );
  AND2X2 AND2X2_2034 ( .A(core__abc_21380_n1960), .B(core__abc_21380_n2451_1_bF_buf1), .Y(core__abc_21380_n2601) );
  AND2X2 AND2X2_2035 ( .A(core__abc_21380_n2452_bF_buf2), .B(core_siphash_word_37_), .Y(core__abc_21380_n2602) );
  AND2X2 AND2X2_2036 ( .A(core__abc_21380_n2603_1), .B(reset_n_bF_buf74), .Y(core_siphash_word0_reg_37__FF_INPUT) );
  AND2X2 AND2X2_2037 ( .A(core__abc_21380_n2606), .B(reset_n_bF_buf73), .Y(core__abc_21380_n2607) );
  AND2X2 AND2X2_2038 ( .A(core__abc_21380_n2607), .B(core__abc_21380_n2605), .Y(core_siphash_word0_reg_38__FF_INPUT) );
  AND2X2 AND2X2_2039 ( .A(core__abc_21380_n2610), .B(reset_n_bF_buf72), .Y(core__abc_21380_n2611) );
  AND2X2 AND2X2_204 ( .A(_abc_19068_n939_1_bF_buf1), .B(core_key_77_), .Y(_abc_19068_n1236) );
  AND2X2 AND2X2_2040 ( .A(core__abc_21380_n2609), .B(core__abc_21380_n2611), .Y(core_siphash_word0_reg_39__FF_INPUT) );
  AND2X2 AND2X2_2041 ( .A(core__abc_21380_n2016), .B(core__abc_21380_n2451_1_bF_buf6), .Y(core__abc_21380_n2613) );
  AND2X2 AND2X2_2042 ( .A(core__abc_21380_n2452_bF_buf7), .B(core_siphash_word_40_), .Y(core__abc_21380_n2614) );
  AND2X2 AND2X2_2043 ( .A(core__abc_21380_n2615), .B(reset_n_bF_buf71), .Y(core_siphash_word0_reg_40__FF_INPUT) );
  AND2X2 AND2X2_2044 ( .A(core__abc_21380_n2618), .B(reset_n_bF_buf70), .Y(core__abc_21380_n2619) );
  AND2X2 AND2X2_2045 ( .A(core__abc_21380_n2619), .B(core__abc_21380_n2617), .Y(core_siphash_word0_reg_41__FF_INPUT) );
  AND2X2 AND2X2_2046 ( .A(core__abc_21380_n2622), .B(reset_n_bF_buf69), .Y(core__abc_21380_n2623) );
  AND2X2 AND2X2_2047 ( .A(core__abc_21380_n2623), .B(core__abc_21380_n2621), .Y(core_siphash_word0_reg_42__FF_INPUT) );
  AND2X2 AND2X2_2048 ( .A(core__abc_21380_n2626), .B(reset_n_bF_buf68), .Y(core__abc_21380_n2627_1) );
  AND2X2 AND2X2_2049 ( .A(core__abc_21380_n2625), .B(core__abc_21380_n2627_1), .Y(core_siphash_word0_reg_43__FF_INPUT) );
  AND2X2 AND2X2_205 ( .A(_abc_19068_n897_1_bF_buf0), .B(word0_reg_13_), .Y(_abc_19068_n1238) );
  AND2X2 AND2X2_2050 ( .A(core__abc_21380_n2090), .B(core__abc_21380_n2451_1_bF_buf2), .Y(core__abc_21380_n2629) );
  AND2X2 AND2X2_2051 ( .A(core__abc_21380_n2452_bF_buf3), .B(core_siphash_word_44_), .Y(core__abc_21380_n2630) );
  AND2X2 AND2X2_2052 ( .A(core__abc_21380_n2631), .B(reset_n_bF_buf67), .Y(core_siphash_word0_reg_44__FF_INPUT) );
  AND2X2 AND2X2_2053 ( .A(core__abc_21380_n2634), .B(reset_n_bF_buf66), .Y(core__abc_21380_n2635) );
  AND2X2 AND2X2_2054 ( .A(core__abc_21380_n2633_1), .B(core__abc_21380_n2635), .Y(core_siphash_word0_reg_45__FF_INPUT) );
  AND2X2 AND2X2_2055 ( .A(core__abc_21380_n2128), .B(core__abc_21380_n2451_1_bF_buf0), .Y(core__abc_21380_n2637) );
  AND2X2 AND2X2_2056 ( .A(core__abc_21380_n2452_bF_buf1), .B(core_siphash_word_46_), .Y(core__abc_21380_n2638) );
  AND2X2 AND2X2_2057 ( .A(core__abc_21380_n2639), .B(reset_n_bF_buf65), .Y(core_siphash_word0_reg_46__FF_INPUT) );
  AND2X2 AND2X2_2058 ( .A(core__abc_21380_n2642), .B(reset_n_bF_buf64), .Y(core__abc_21380_n2643) );
  AND2X2 AND2X2_2059 ( .A(core__abc_21380_n2641), .B(core__abc_21380_n2643), .Y(core_siphash_word0_reg_47__FF_INPUT) );
  AND2X2 AND2X2_206 ( .A(_abc_19068_n916_1_bF_buf0), .B(word1_reg_13_), .Y(_abc_19068_n1239_1) );
  AND2X2 AND2X2_2060 ( .A(core__abc_21380_n2646), .B(reset_n_bF_buf63), .Y(core__abc_21380_n2647) );
  AND2X2 AND2X2_2061 ( .A(core__abc_21380_n2647), .B(core__abc_21380_n2645), .Y(core_siphash_word0_reg_48__FF_INPUT) );
  AND2X2 AND2X2_2062 ( .A(core__abc_21380_n2184), .B(core__abc_21380_n2451_1_bF_buf5), .Y(core__abc_21380_n2649) );
  AND2X2 AND2X2_2063 ( .A(core__abc_21380_n2452_bF_buf6), .B(core_siphash_word_49_), .Y(core__abc_21380_n2650) );
  AND2X2 AND2X2_2064 ( .A(core__abc_21380_n2651), .B(reset_n_bF_buf62), .Y(core_siphash_word0_reg_49__FF_INPUT) );
  AND2X2 AND2X2_2065 ( .A(core__abc_21380_n2202), .B(core__abc_21380_n2451_1_bF_buf4), .Y(core__abc_21380_n2653) );
  AND2X2 AND2X2_2066 ( .A(core__abc_21380_n2452_bF_buf5), .B(core_siphash_word_50_), .Y(core__abc_21380_n2654_1) );
  AND2X2 AND2X2_2067 ( .A(core__abc_21380_n2655), .B(reset_n_bF_buf61), .Y(core_siphash_word0_reg_50__FF_INPUT) );
  AND2X2 AND2X2_2068 ( .A(core__abc_21380_n2222), .B(core__abc_21380_n2451_1_bF_buf3), .Y(core__abc_21380_n2657) );
  AND2X2 AND2X2_2069 ( .A(core__abc_21380_n2452_bF_buf4), .B(core_siphash_word_51_), .Y(core__abc_21380_n2658) );
  AND2X2 AND2X2_207 ( .A(_abc_19068_n1243_1), .B(_abc_19068_n923_bF_buf1), .Y(_auto_iopadmap_cc_313_execute_30317_13_) );
  AND2X2 AND2X2_2070 ( .A(core__abc_21380_n2659), .B(reset_n_bF_buf60), .Y(core_siphash_word0_reg_51__FF_INPUT) );
  AND2X2 AND2X2_2071 ( .A(core__abc_21380_n2662), .B(reset_n_bF_buf59), .Y(core__abc_21380_n2663) );
  AND2X2 AND2X2_2072 ( .A(core__abc_21380_n2663), .B(core__abc_21380_n2661), .Y(core_siphash_word0_reg_52__FF_INPUT) );
  AND2X2 AND2X2_2073 ( .A(core__abc_21380_n2259), .B(core__abc_21380_n2451_1_bF_buf1), .Y(core__abc_21380_n2665) );
  AND2X2 AND2X2_2074 ( .A(core__abc_21380_n2452_bF_buf2), .B(core_siphash_word_53_), .Y(core__abc_21380_n2666) );
  AND2X2 AND2X2_2075 ( .A(core__abc_21380_n2667), .B(reset_n_bF_buf58), .Y(core_siphash_word0_reg_53__FF_INPUT) );
  AND2X2 AND2X2_2076 ( .A(core__abc_21380_n2670), .B(reset_n_bF_buf57), .Y(core__abc_21380_n2671) );
  AND2X2 AND2X2_2077 ( .A(core__abc_21380_n2671), .B(core__abc_21380_n2669), .Y(core_siphash_word0_reg_54__FF_INPUT) );
  AND2X2 AND2X2_2078 ( .A(core__abc_21380_n2674), .B(reset_n_bF_buf56), .Y(core__abc_21380_n2675) );
  AND2X2 AND2X2_2079 ( .A(core__abc_21380_n2673), .B(core__abc_21380_n2675), .Y(core_siphash_word0_reg_55__FF_INPUT) );
  AND2X2 AND2X2_208 ( .A(_abc_19068_n941_bF_buf0), .B(core_key_110_), .Y(_abc_19068_n1245_1) );
  AND2X2 AND2X2_2080 ( .A(core__abc_21380_n2678), .B(reset_n_bF_buf55), .Y(core__abc_21380_n2679) );
  AND2X2 AND2X2_2081 ( .A(core__abc_21380_n2679), .B(core__abc_21380_n2677), .Y(core_siphash_word0_reg_56__FF_INPUT) );
  AND2X2 AND2X2_2082 ( .A(core__abc_21380_n2682_1), .B(reset_n_bF_buf54), .Y(core__abc_21380_n2683) );
  AND2X2 AND2X2_2083 ( .A(core__abc_21380_n2683), .B(core__abc_21380_n2681), .Y(core_siphash_word0_reg_57__FF_INPUT) );
  AND2X2 AND2X2_2084 ( .A(core__abc_21380_n2686), .B(reset_n_bF_buf53), .Y(core__abc_21380_n2687) );
  AND2X2 AND2X2_2085 ( .A(core__abc_21380_n2687), .B(core__abc_21380_n2685), .Y(core_siphash_word0_reg_58__FF_INPUT) );
  AND2X2 AND2X2_2086 ( .A(core__abc_21380_n2690), .B(reset_n_bF_buf52), .Y(core__abc_21380_n2691) );
  AND2X2 AND2X2_2087 ( .A(core__abc_21380_n2689), .B(core__abc_21380_n2691), .Y(core_siphash_word0_reg_59__FF_INPUT) );
  AND2X2 AND2X2_2088 ( .A(core__abc_21380_n2694), .B(reset_n_bF_buf51), .Y(core__abc_21380_n2695) );
  AND2X2 AND2X2_2089 ( .A(core__abc_21380_n2695), .B(core__abc_21380_n2693), .Y(core_siphash_word0_reg_60__FF_INPUT) );
  AND2X2 AND2X2_209 ( .A(_abc_19068_n945_1_bF_buf0), .B(core_mi_14_), .Y(_abc_19068_n1246) );
  AND2X2 AND2X2_2090 ( .A(core__abc_21380_n2698), .B(reset_n_bF_buf50), .Y(core__abc_21380_n2699) );
  AND2X2 AND2X2_2091 ( .A(core__abc_21380_n2699), .B(core__abc_21380_n2697), .Y(core_siphash_word0_reg_61__FF_INPUT) );
  AND2X2 AND2X2_2092 ( .A(core__abc_21380_n2702), .B(reset_n_bF_buf49), .Y(core__abc_21380_n2703) );
  AND2X2 AND2X2_2093 ( .A(core__abc_21380_n2703), .B(core__abc_21380_n2701), .Y(core_siphash_word0_reg_62__FF_INPUT) );
  AND2X2 AND2X2_2094 ( .A(core__abc_21380_n2443), .B(core__abc_21380_n2451_1_bF_buf7), .Y(core__abc_21380_n2705) );
  AND2X2 AND2X2_2095 ( .A(core__abc_21380_n2452_bF_buf0), .B(core_siphash_word_63_), .Y(core__abc_21380_n2706) );
  AND2X2 AND2X2_2096 ( .A(core__abc_21380_n2707), .B(reset_n_bF_buf48), .Y(core_siphash_word0_reg_63__FF_INPUT) );
  AND2X2 AND2X2_2097 ( .A(core__abc_21380_n1142_1), .B(core__abc_21380_n1137_1), .Y(core__abc_21380_n2710) );
  AND2X2 AND2X2_2098 ( .A(core__abc_21380_n2712), .B(core_ready), .Y(core__abc_21380_n2713) );
  AND2X2 AND2X2_2099 ( .A(core__abc_21380_n1139), .B(core__abc_21380_n2449), .Y(core__abc_21380_n2716) );
  AND2X2 AND2X2_21 ( .A(_abc_19068_n886_1), .B(\addr[1] ), .Y(_abc_19068_n900_1) );
  AND2X2 AND2X2_210 ( .A(_abc_19068_n899_bF_buf4), .B(word3_reg_14_), .Y(_abc_19068_n1249_1) );
  AND2X2 AND2X2_2100 ( .A(core__abc_21380_n2717), .B(core__abc_21380_n1137_1), .Y(core__abc_21380_n2718) );
  AND2X2 AND2X2_2101 ( .A(core__abc_21380_n2715), .B(core__abc_21380_n2718), .Y(core__abc_21380_n2719) );
  AND2X2 AND2X2_2102 ( .A(core__abc_21380_n2721), .B(reset_n_bF_buf47), .Y(core__abc_21380_n2722) );
  AND2X2 AND2X2_2103 ( .A(core__abc_21380_n2720), .B(core__abc_21380_n2722), .Y(core_loop_ctr_reg_0__FF_INPUT) );
  AND2X2 AND2X2_2104 ( .A(core__abc_21380_n2719), .B(core_loop_ctr_reg_1_), .Y(core__abc_21380_n2724_1) );
  AND2X2 AND2X2_2105 ( .A(core_loop_ctr_reg_1_), .B(core_loop_ctr_reg_0_), .Y(core__abc_21380_n2725) );
  AND2X2 AND2X2_2106 ( .A(core__abc_21380_n2716), .B(core__abc_21380_n2726), .Y(core__abc_21380_n2727) );
  AND2X2 AND2X2_2107 ( .A(core__abc_21380_n2729), .B(reset_n_bF_buf46), .Y(core__abc_21380_n2730) );
  AND2X2 AND2X2_2108 ( .A(core__abc_21380_n2728_1), .B(core__abc_21380_n2730), .Y(core_loop_ctr_reg_1__FF_INPUT) );
  AND2X2 AND2X2_2109 ( .A(core__abc_21380_n2719), .B(core_loop_ctr_reg_2_), .Y(core__abc_21380_n2732) );
  AND2X2 AND2X2_211 ( .A(_abc_19068_n939_1_bF_buf0), .B(core_key_78_), .Y(_abc_19068_n1252) );
  AND2X2 AND2X2_2110 ( .A(core__abc_21380_n2725), .B(core_loop_ctr_reg_2_), .Y(core__abc_21380_n2733) );
  AND2X2 AND2X2_2111 ( .A(core__abc_21380_n2716), .B(core__abc_21380_n2734), .Y(core__abc_21380_n2735) );
  AND2X2 AND2X2_2112 ( .A(core__abc_21380_n2737), .B(reset_n_bF_buf45), .Y(core__abc_21380_n2738) );
  AND2X2 AND2X2_2113 ( .A(core__abc_21380_n2736), .B(core__abc_21380_n2738), .Y(core_loop_ctr_reg_2__FF_INPUT) );
  AND2X2 AND2X2_2114 ( .A(core__abc_21380_n2716), .B(core__abc_21380_n2733), .Y(core__abc_21380_n2742) );
  AND2X2 AND2X2_2115 ( .A(core__abc_21380_n2743), .B(reset_n_bF_buf44), .Y(core__abc_21380_n2744) );
  AND2X2 AND2X2_2116 ( .A(core__abc_21380_n2741), .B(core__abc_21380_n2744), .Y(core_loop_ctr_reg_3__FF_INPUT) );
  AND2X2 AND2X2_2117 ( .A(core__abc_21380_n1133_1), .B(core_compress), .Y(core__abc_21380_n2746) );
  AND2X2 AND2X2_2118 ( .A(core__abc_21380_n2746), .B(core__abc_21380_n1144_1), .Y(core__abc_21380_n2747) );
  AND2X2 AND2X2_2119 ( .A(core__abc_21380_n2747), .B(core__abc_21380_n1138_1), .Y(core__abc_21380_n2748) );
  AND2X2 AND2X2_212 ( .A(_abc_19068_n926_bF_buf0), .B(core_key_14_), .Y(_abc_19068_n1253_1) );
  AND2X2 AND2X2_2120 ( .A(core__abc_21380_n2448), .B(core__abc_21380_n2748), .Y(core__abc_21380_n2749) );
  AND2X2 AND2X2_2121 ( .A(core__abc_21380_n2750_bF_buf7), .B(core_mi_reg_0_), .Y(core__abc_21380_n2751) );
  AND2X2 AND2X2_2122 ( .A(core__abc_21380_n2749_bF_buf9), .B(core_mi_0_), .Y(core__abc_21380_n2752) );
  AND2X2 AND2X2_2123 ( .A(core__abc_21380_n2753), .B(reset_n_bF_buf43), .Y(core_mi_reg_0__FF_INPUT) );
  AND2X2 AND2X2_2124 ( .A(core__abc_21380_n2750_bF_buf6), .B(core_mi_reg_1_), .Y(core__abc_21380_n2755) );
  AND2X2 AND2X2_2125 ( .A(core__abc_21380_n2749_bF_buf8), .B(core_mi_1_), .Y(core__abc_21380_n2756) );
  AND2X2 AND2X2_2126 ( .A(core__abc_21380_n2757), .B(reset_n_bF_buf42), .Y(core_mi_reg_1__FF_INPUT) );
  AND2X2 AND2X2_2127 ( .A(core__abc_21380_n2750_bF_buf5), .B(core_mi_reg_2_), .Y(core__abc_21380_n2759) );
  AND2X2 AND2X2_2128 ( .A(core__abc_21380_n2749_bF_buf7), .B(core_mi_2_), .Y(core__abc_21380_n2760) );
  AND2X2 AND2X2_2129 ( .A(core__abc_21380_n2761), .B(reset_n_bF_buf41), .Y(core_mi_reg_2__FF_INPUT) );
  AND2X2 AND2X2_213 ( .A(_abc_19068_n924_1_bF_buf0), .B(core_key_46_), .Y(_abc_19068_n1254) );
  AND2X2 AND2X2_2130 ( .A(core__abc_21380_n2750_bF_buf4), .B(core_mi_reg_3_), .Y(core__abc_21380_n2763) );
  AND2X2 AND2X2_2131 ( .A(core__abc_21380_n2749_bF_buf6), .B(core_mi_3_), .Y(core__abc_21380_n2764) );
  AND2X2 AND2X2_2132 ( .A(core__abc_21380_n2765), .B(reset_n_bF_buf40), .Y(core_mi_reg_3__FF_INPUT) );
  AND2X2 AND2X2_2133 ( .A(core__abc_21380_n2750_bF_buf3), .B(core_mi_reg_4_), .Y(core__abc_21380_n2767) );
  AND2X2 AND2X2_2134 ( .A(core__abc_21380_n2749_bF_buf5), .B(core_mi_4_), .Y(core__abc_21380_n2768) );
  AND2X2 AND2X2_2135 ( .A(core__abc_21380_n2769), .B(reset_n_bF_buf39), .Y(core_mi_reg_4__FF_INPUT) );
  AND2X2 AND2X2_2136 ( .A(core__abc_21380_n2750_bF_buf2), .B(core_mi_reg_5_), .Y(core__abc_21380_n2771) );
  AND2X2 AND2X2_2137 ( .A(core__abc_21380_n2749_bF_buf4), .B(core_mi_5_), .Y(core__abc_21380_n2772) );
  AND2X2 AND2X2_2138 ( .A(core__abc_21380_n2773), .B(reset_n_bF_buf38), .Y(core_mi_reg_5__FF_INPUT) );
  AND2X2 AND2X2_2139 ( .A(core__abc_21380_n2750_bF_buf1), .B(core_mi_reg_6_), .Y(core__abc_21380_n2775) );
  AND2X2 AND2X2_214 ( .A(_abc_19068_n916_1_bF_buf4), .B(word1_reg_14_), .Y(_abc_19068_n1257_1) );
  AND2X2 AND2X2_2140 ( .A(core__abc_21380_n2749_bF_buf3), .B(core_mi_6_), .Y(core__abc_21380_n2776) );
  AND2X2 AND2X2_2141 ( .A(core__abc_21380_n2777), .B(reset_n_bF_buf37), .Y(core_mi_reg_6__FF_INPUT) );
  AND2X2 AND2X2_2142 ( .A(core__abc_21380_n2750_bF_buf0), .B(core_mi_reg_7_), .Y(core__abc_21380_n2779) );
  AND2X2 AND2X2_2143 ( .A(core__abc_21380_n2749_bF_buf2), .B(core_mi_7_), .Y(core__abc_21380_n2780) );
  AND2X2 AND2X2_2144 ( .A(core__abc_21380_n2781), .B(reset_n_bF_buf36), .Y(core_mi_reg_7__FF_INPUT) );
  AND2X2 AND2X2_2145 ( .A(core__abc_21380_n2750_bF_buf7), .B(core_mi_reg_8_), .Y(core__abc_21380_n2783) );
  AND2X2 AND2X2_2146 ( .A(core__abc_21380_n2749_bF_buf1), .B(core_mi_8_), .Y(core__abc_21380_n2784) );
  AND2X2 AND2X2_2147 ( .A(core__abc_21380_n2785), .B(reset_n_bF_buf35), .Y(core_mi_reg_8__FF_INPUT) );
  AND2X2 AND2X2_2148 ( .A(core__abc_21380_n2750_bF_buf6), .B(core_mi_reg_9_), .Y(core__abc_21380_n2787) );
  AND2X2 AND2X2_2149 ( .A(core__abc_21380_n2749_bF_buf0), .B(core_mi_9_), .Y(core__abc_21380_n2788) );
  AND2X2 AND2X2_215 ( .A(_abc_19068_n902_bF_buf4), .B(word2_reg_14_), .Y(_abc_19068_n1258) );
  AND2X2 AND2X2_2150 ( .A(core__abc_21380_n2789), .B(reset_n_bF_buf34), .Y(core_mi_reg_9__FF_INPUT) );
  AND2X2 AND2X2_2151 ( .A(core__abc_21380_n2750_bF_buf5), .B(core_mi_reg_10_), .Y(core__abc_21380_n2791) );
  AND2X2 AND2X2_2152 ( .A(core__abc_21380_n2749_bF_buf10), .B(core_mi_10_), .Y(core__abc_21380_n2792) );
  AND2X2 AND2X2_2153 ( .A(core__abc_21380_n2793), .B(reset_n_bF_buf33), .Y(core_mi_reg_10__FF_INPUT) );
  AND2X2 AND2X2_2154 ( .A(core__abc_21380_n2750_bF_buf4), .B(core_mi_reg_11_), .Y(core__abc_21380_n2795) );
  AND2X2 AND2X2_2155 ( .A(core__abc_21380_n2749_bF_buf9), .B(core_mi_11_), .Y(core__abc_21380_n2796) );
  AND2X2 AND2X2_2156 ( .A(core__abc_21380_n2797), .B(reset_n_bF_buf32), .Y(core_mi_reg_11__FF_INPUT) );
  AND2X2 AND2X2_2157 ( .A(core__abc_21380_n2750_bF_buf3), .B(core_mi_reg_12_), .Y(core__abc_21380_n2799) );
  AND2X2 AND2X2_2158 ( .A(core__abc_21380_n2749_bF_buf8), .B(core_mi_12_), .Y(core__abc_21380_n2800_1) );
  AND2X2 AND2X2_2159 ( .A(core__abc_21380_n2801), .B(reset_n_bF_buf31), .Y(core_mi_reg_12__FF_INPUT) );
  AND2X2 AND2X2_216 ( .A(_abc_19068_n915_1_bF_buf4), .B(core_mi_46_), .Y(_abc_19068_n1260) );
  AND2X2 AND2X2_2160 ( .A(core__abc_21380_n2750_bF_buf2), .B(core_mi_reg_13_), .Y(core__abc_21380_n2803) );
  AND2X2 AND2X2_2161 ( .A(core__abc_21380_n2749_bF_buf7), .B(core_mi_13_), .Y(core__abc_21380_n2804_1) );
  AND2X2 AND2X2_2162 ( .A(core__abc_21380_n2805), .B(reset_n_bF_buf30), .Y(core_mi_reg_13__FF_INPUT) );
  AND2X2 AND2X2_2163 ( .A(core__abc_21380_n2750_bF_buf1), .B(core_mi_reg_14_), .Y(core__abc_21380_n2807) );
  AND2X2 AND2X2_2164 ( .A(core__abc_21380_n2749_bF_buf6), .B(core_mi_14_), .Y(core__abc_21380_n2808) );
  AND2X2 AND2X2_2165 ( .A(core__abc_21380_n2809), .B(reset_n_bF_buf29), .Y(core_mi_reg_14__FF_INPUT) );
  AND2X2 AND2X2_2166 ( .A(core__abc_21380_n2750_bF_buf0), .B(core_mi_reg_15_), .Y(core__abc_21380_n2811) );
  AND2X2 AND2X2_2167 ( .A(core__abc_21380_n2749_bF_buf5), .B(core_mi_15_), .Y(core__abc_21380_n2812) );
  AND2X2 AND2X2_2168 ( .A(core__abc_21380_n2813), .B(reset_n_bF_buf28), .Y(core_mi_reg_15__FF_INPUT) );
  AND2X2 AND2X2_2169 ( .A(core__abc_21380_n2750_bF_buf7), .B(core_mi_reg_16_), .Y(core__abc_21380_n2815) );
  AND2X2 AND2X2_217 ( .A(_abc_19068_n897_1_bF_buf4), .B(word0_reg_14_), .Y(_abc_19068_n1261_1) );
  AND2X2 AND2X2_2170 ( .A(core__abc_21380_n2749_bF_buf4), .B(core_mi_16_), .Y(core__abc_21380_n2816) );
  AND2X2 AND2X2_2171 ( .A(core__abc_21380_n2817_1), .B(reset_n_bF_buf27), .Y(core_mi_reg_16__FF_INPUT) );
  AND2X2 AND2X2_2172 ( .A(core__abc_21380_n2750_bF_buf6), .B(core_mi_reg_17_), .Y(core__abc_21380_n2819) );
  AND2X2 AND2X2_2173 ( .A(core__abc_21380_n2749_bF_buf3), .B(core_mi_17_), .Y(core__abc_21380_n2820) );
  AND2X2 AND2X2_2174 ( .A(core__abc_21380_n2821), .B(reset_n_bF_buf26), .Y(core_mi_reg_17__FF_INPUT) );
  AND2X2 AND2X2_2175 ( .A(core__abc_21380_n2750_bF_buf5), .B(core_mi_reg_18_), .Y(core__abc_21380_n2823_1) );
  AND2X2 AND2X2_2176 ( .A(core__abc_21380_n2749_bF_buf2), .B(core_mi_18_), .Y(core__abc_21380_n2824) );
  AND2X2 AND2X2_2177 ( .A(core__abc_21380_n2825), .B(reset_n_bF_buf25), .Y(core_mi_reg_18__FF_INPUT) );
  AND2X2 AND2X2_2178 ( .A(core__abc_21380_n2750_bF_buf4), .B(core_mi_reg_19_), .Y(core__abc_21380_n2827) );
  AND2X2 AND2X2_2179 ( .A(core__abc_21380_n2749_bF_buf1), .B(core_mi_19_), .Y(core__abc_21380_n2828) );
  AND2X2 AND2X2_218 ( .A(_abc_19068_n923_bF_buf0), .B(_abc_19068_n1265_1), .Y(_auto_iopadmap_cc_313_execute_30317_14_) );
  AND2X2 AND2X2_2180 ( .A(core__abc_21380_n2829), .B(reset_n_bF_buf24), .Y(core_mi_reg_19__FF_INPUT) );
  AND2X2 AND2X2_2181 ( .A(core__abc_21380_n2750_bF_buf3), .B(core_mi_reg_20_), .Y(core__abc_21380_n2831) );
  AND2X2 AND2X2_2182 ( .A(core__abc_21380_n2749_bF_buf0), .B(core_mi_20_), .Y(core__abc_21380_n2832) );
  AND2X2 AND2X2_2183 ( .A(core__abc_21380_n2833), .B(reset_n_bF_buf23), .Y(core_mi_reg_20__FF_INPUT) );
  AND2X2 AND2X2_2184 ( .A(core__abc_21380_n2750_bF_buf2), .B(core_mi_reg_21_), .Y(core__abc_21380_n2835) );
  AND2X2 AND2X2_2185 ( .A(core__abc_21380_n2749_bF_buf10), .B(core_mi_21_), .Y(core__abc_21380_n2836) );
  AND2X2 AND2X2_2186 ( .A(core__abc_21380_n2837), .B(reset_n_bF_buf22), .Y(core_mi_reg_21__FF_INPUT) );
  AND2X2 AND2X2_2187 ( .A(core__abc_21380_n2750_bF_buf1), .B(core_mi_reg_22_), .Y(core__abc_21380_n2839_1) );
  AND2X2 AND2X2_2188 ( .A(core__abc_21380_n2749_bF_buf9), .B(core_mi_22_), .Y(core__abc_21380_n2840) );
  AND2X2 AND2X2_2189 ( .A(core__abc_21380_n2841), .B(reset_n_bF_buf21), .Y(core_mi_reg_22__FF_INPUT) );
  AND2X2 AND2X2_219 ( .A(_abc_19068_n916_1_bF_buf3), .B(word1_reg_15_), .Y(_abc_19068_n1267_1) );
  AND2X2 AND2X2_2190 ( .A(core__abc_21380_n2750_bF_buf0), .B(core_mi_reg_23_), .Y(core__abc_21380_n2843) );
  AND2X2 AND2X2_2191 ( .A(core__abc_21380_n2749_bF_buf8), .B(core_mi_23_), .Y(core__abc_21380_n2844) );
  AND2X2 AND2X2_2192 ( .A(core__abc_21380_n2845_1), .B(reset_n_bF_buf20), .Y(core_mi_reg_23__FF_INPUT) );
  AND2X2 AND2X2_2193 ( .A(core__abc_21380_n2750_bF_buf7), .B(core_mi_reg_24_), .Y(core__abc_21380_n2847) );
  AND2X2 AND2X2_2194 ( .A(core__abc_21380_n2749_bF_buf7), .B(core_mi_24_), .Y(core__abc_21380_n2848) );
  AND2X2 AND2X2_2195 ( .A(core__abc_21380_n2849), .B(reset_n_bF_buf19), .Y(core_mi_reg_24__FF_INPUT) );
  AND2X2 AND2X2_2196 ( .A(core__abc_21380_n2750_bF_buf6), .B(core_mi_reg_25_), .Y(core__abc_21380_n2851) );
  AND2X2 AND2X2_2197 ( .A(core__abc_21380_n2749_bF_buf6), .B(core_mi_25_), .Y(core__abc_21380_n2852) );
  AND2X2 AND2X2_2198 ( .A(core__abc_21380_n2853), .B(reset_n_bF_buf18), .Y(core_mi_reg_25__FF_INPUT) );
  AND2X2 AND2X2_2199 ( .A(core__abc_21380_n2750_bF_buf5), .B(core_mi_reg_26_), .Y(core__abc_21380_n2855) );
  AND2X2 AND2X2_22 ( .A(_abc_19068_n893), .B(_abc_19068_n900_1), .Y(_abc_19068_n901_1) );
  AND2X2 AND2X2_220 ( .A(_abc_19068_n897_1_bF_buf3), .B(word0_reg_15_), .Y(_abc_19068_n1268) );
  AND2X2 AND2X2_2200 ( .A(core__abc_21380_n2749_bF_buf5), .B(core_mi_26_), .Y(core__abc_21380_n2856) );
  AND2X2 AND2X2_2201 ( .A(core__abc_21380_n2857), .B(reset_n_bF_buf17), .Y(core_mi_reg_26__FF_INPUT) );
  AND2X2 AND2X2_2202 ( .A(core__abc_21380_n2750_bF_buf4), .B(core_mi_reg_27_), .Y(core__abc_21380_n2859) );
  AND2X2 AND2X2_2203 ( .A(core__abc_21380_n2749_bF_buf4), .B(core_mi_27_), .Y(core__abc_21380_n2860_1) );
  AND2X2 AND2X2_2204 ( .A(core__abc_21380_n2861), .B(reset_n_bF_buf16), .Y(core_mi_reg_27__FF_INPUT) );
  AND2X2 AND2X2_2205 ( .A(core__abc_21380_n2750_bF_buf3), .B(core_mi_reg_28_), .Y(core__abc_21380_n2863) );
  AND2X2 AND2X2_2206 ( .A(core__abc_21380_n2749_bF_buf3), .B(core_mi_28_), .Y(core__abc_21380_n2864_1) );
  AND2X2 AND2X2_2207 ( .A(core__abc_21380_n2865), .B(reset_n_bF_buf15), .Y(core_mi_reg_28__FF_INPUT) );
  AND2X2 AND2X2_2208 ( .A(core__abc_21380_n2750_bF_buf2), .B(core_mi_reg_29_), .Y(core__abc_21380_n2867) );
  AND2X2 AND2X2_2209 ( .A(core__abc_21380_n2749_bF_buf2), .B(core_mi_29_), .Y(core__abc_21380_n2868) );
  AND2X2 AND2X2_221 ( .A(_abc_19068_n941_bF_buf4), .B(core_key_111_), .Y(_abc_19068_n1270) );
  AND2X2 AND2X2_2210 ( .A(core__abc_21380_n2869), .B(reset_n_bF_buf14), .Y(core_mi_reg_29__FF_INPUT) );
  AND2X2 AND2X2_2211 ( .A(core__abc_21380_n2750_bF_buf1), .B(core_mi_reg_30_), .Y(core__abc_21380_n2871) );
  AND2X2 AND2X2_2212 ( .A(core__abc_21380_n2749_bF_buf1), .B(core_mi_30_), .Y(core__abc_21380_n2872) );
  AND2X2 AND2X2_2213 ( .A(core__abc_21380_n2873), .B(reset_n_bF_buf13), .Y(core_mi_reg_30__FF_INPUT) );
  AND2X2 AND2X2_2214 ( .A(core__abc_21380_n2750_bF_buf0), .B(core_mi_reg_31_), .Y(core__abc_21380_n2875) );
  AND2X2 AND2X2_2215 ( .A(core__abc_21380_n2749_bF_buf0), .B(core_mi_31_), .Y(core__abc_21380_n2876) );
  AND2X2 AND2X2_2216 ( .A(core__abc_21380_n2877), .B(reset_n_bF_buf12), .Y(core_mi_reg_31__FF_INPUT) );
  AND2X2 AND2X2_2217 ( .A(core__abc_21380_n2750_bF_buf7), .B(core_mi_reg_32_), .Y(core__abc_21380_n2879) );
  AND2X2 AND2X2_2218 ( .A(core__abc_21380_n2749_bF_buf10), .B(core_mi_32_), .Y(core__abc_21380_n2880) );
  AND2X2 AND2X2_2219 ( .A(core__abc_21380_n2881_1), .B(reset_n_bF_buf11), .Y(core_mi_reg_32__FF_INPUT) );
  AND2X2 AND2X2_222 ( .A(_abc_19068_n924_1_bF_buf4), .B(core_key_47_), .Y(_abc_19068_n1271_1) );
  AND2X2 AND2X2_2220 ( .A(core__abc_21380_n2750_bF_buf6), .B(core_mi_reg_33_), .Y(core__abc_21380_n2883) );
  AND2X2 AND2X2_2221 ( .A(core__abc_21380_n2749_bF_buf9), .B(core_mi_33_), .Y(core__abc_21380_n2884) );
  AND2X2 AND2X2_2222 ( .A(core__abc_21380_n2885_1), .B(reset_n_bF_buf10), .Y(core_mi_reg_33__FF_INPUT) );
  AND2X2 AND2X2_2223 ( .A(core__abc_21380_n2750_bF_buf5), .B(core_mi_reg_34_), .Y(core__abc_21380_n2887) );
  AND2X2 AND2X2_2224 ( .A(core__abc_21380_n2749_bF_buf8), .B(core_mi_34_), .Y(core__abc_21380_n2888) );
  AND2X2 AND2X2_2225 ( .A(core__abc_21380_n2889), .B(reset_n_bF_buf9), .Y(core_mi_reg_34__FF_INPUT) );
  AND2X2 AND2X2_2226 ( .A(core__abc_21380_n2750_bF_buf4), .B(core_mi_reg_35_), .Y(core__abc_21380_n2891) );
  AND2X2 AND2X2_2227 ( .A(core__abc_21380_n2749_bF_buf7), .B(core_mi_35_), .Y(core__abc_21380_n2892) );
  AND2X2 AND2X2_2228 ( .A(core__abc_21380_n2893), .B(reset_n_bF_buf8), .Y(core_mi_reg_35__FF_INPUT) );
  AND2X2 AND2X2_2229 ( .A(core__abc_21380_n2750_bF_buf3), .B(core_mi_reg_36_), .Y(core__abc_21380_n2895) );
  AND2X2 AND2X2_223 ( .A(_abc_19068_n926_bF_buf4), .B(core_key_15_), .Y(_abc_19068_n1272) );
  AND2X2 AND2X2_2230 ( .A(core__abc_21380_n2749_bF_buf6), .B(core_mi_36_), .Y(core__abc_21380_n2896) );
  AND2X2 AND2X2_2231 ( .A(core__abc_21380_n2897), .B(reset_n_bF_buf7), .Y(core_mi_reg_36__FF_INPUT) );
  AND2X2 AND2X2_2232 ( .A(core__abc_21380_n2750_bF_buf2), .B(core_mi_reg_37_), .Y(core__abc_21380_n2899) );
  AND2X2 AND2X2_2233 ( .A(core__abc_21380_n2749_bF_buf5), .B(core_mi_37_), .Y(core__abc_21380_n2900_1) );
  AND2X2 AND2X2_2234 ( .A(core__abc_21380_n2901), .B(reset_n_bF_buf6), .Y(core_mi_reg_37__FF_INPUT) );
  AND2X2 AND2X2_2235 ( .A(core__abc_21380_n2750_bF_buf1), .B(core_mi_reg_38_), .Y(core__abc_21380_n2903) );
  AND2X2 AND2X2_2236 ( .A(core__abc_21380_n2749_bF_buf4), .B(core_mi_38_), .Y(core__abc_21380_n2904_1) );
  AND2X2 AND2X2_2237 ( .A(core__abc_21380_n2905), .B(reset_n_bF_buf5), .Y(core_mi_reg_38__FF_INPUT) );
  AND2X2 AND2X2_2238 ( .A(core__abc_21380_n2750_bF_buf0), .B(core_mi_reg_39_), .Y(core__abc_21380_n2907) );
  AND2X2 AND2X2_2239 ( .A(core__abc_21380_n2749_bF_buf3), .B(core_mi_39_), .Y(core__abc_21380_n2908) );
  AND2X2 AND2X2_224 ( .A(_abc_19068_n939_1_bF_buf4), .B(core_key_79_), .Y(_abc_19068_n1276) );
  AND2X2 AND2X2_2240 ( .A(core__abc_21380_n2909), .B(reset_n_bF_buf4), .Y(core_mi_reg_39__FF_INPUT) );
  AND2X2 AND2X2_2241 ( .A(core__abc_21380_n2750_bF_buf7), .B(core_mi_reg_40_), .Y(core__abc_21380_n2911) );
  AND2X2 AND2X2_2242 ( .A(core__abc_21380_n2749_bF_buf2), .B(core_mi_40_), .Y(core__abc_21380_n2912) );
  AND2X2 AND2X2_2243 ( .A(core__abc_21380_n2913), .B(reset_n_bF_buf3), .Y(core_mi_reg_40__FF_INPUT) );
  AND2X2 AND2X2_2244 ( .A(core__abc_21380_n2750_bF_buf6), .B(core_mi_reg_41_), .Y(core__abc_21380_n2915) );
  AND2X2 AND2X2_2245 ( .A(core__abc_21380_n2749_bF_buf1), .B(core_mi_41_), .Y(core__abc_21380_n2916_1) );
  AND2X2 AND2X2_2246 ( .A(core__abc_21380_n2917), .B(reset_n_bF_buf2), .Y(core_mi_reg_41__FF_INPUT) );
  AND2X2 AND2X2_2247 ( .A(core__abc_21380_n2750_bF_buf5), .B(core_mi_reg_42_), .Y(core__abc_21380_n2919) );
  AND2X2 AND2X2_2248 ( .A(core__abc_21380_n2749_bF_buf0), .B(core_mi_42_), .Y(core__abc_21380_n2920) );
  AND2X2 AND2X2_2249 ( .A(core__abc_21380_n2921), .B(reset_n_bF_buf1), .Y(core_mi_reg_42__FF_INPUT) );
  AND2X2 AND2X2_225 ( .A(_abc_19068_n902_bF_buf3), .B(word2_reg_15_), .Y(_abc_19068_n1277_1) );
  AND2X2 AND2X2_2250 ( .A(core__abc_21380_n2750_bF_buf4), .B(core_mi_reg_43_), .Y(core__abc_21380_n2923) );
  AND2X2 AND2X2_2251 ( .A(core__abc_21380_n2749_bF_buf10), .B(core_mi_43_), .Y(core__abc_21380_n2924) );
  AND2X2 AND2X2_2252 ( .A(core__abc_21380_n2925), .B(reset_n_bF_buf0), .Y(core_mi_reg_43__FF_INPUT) );
  AND2X2 AND2X2_2253 ( .A(core__abc_21380_n2750_bF_buf3), .B(core_mi_reg_44_), .Y(core__abc_21380_n2927) );
  AND2X2 AND2X2_2254 ( .A(core__abc_21380_n2749_bF_buf9), .B(core_mi_44_), .Y(core__abc_21380_n2928) );
  AND2X2 AND2X2_2255 ( .A(core__abc_21380_n2929), .B(reset_n_bF_buf84), .Y(core_mi_reg_44__FF_INPUT) );
  AND2X2 AND2X2_2256 ( .A(core__abc_21380_n2750_bF_buf2), .B(core_mi_reg_45_), .Y(core__abc_21380_n2931) );
  AND2X2 AND2X2_2257 ( .A(core__abc_21380_n2749_bF_buf8), .B(core_mi_45_), .Y(core__abc_21380_n2932) );
  AND2X2 AND2X2_2258 ( .A(core__abc_21380_n2933), .B(reset_n_bF_buf83), .Y(core_mi_reg_45__FF_INPUT) );
  AND2X2 AND2X2_2259 ( .A(core__abc_21380_n2750_bF_buf1), .B(core_mi_reg_46_), .Y(core__abc_21380_n2935) );
  AND2X2 AND2X2_226 ( .A(_abc_19068_n899_bF_buf3), .B(word3_reg_15_), .Y(_abc_19068_n1278) );
  AND2X2 AND2X2_2260 ( .A(core__abc_21380_n2749_bF_buf7), .B(core_mi_46_), .Y(core__abc_21380_n2936) );
  AND2X2 AND2X2_2261 ( .A(core__abc_21380_n2937), .B(reset_n_bF_buf82), .Y(core_mi_reg_46__FF_INPUT) );
  AND2X2 AND2X2_2262 ( .A(core__abc_21380_n2750_bF_buf0), .B(core_mi_reg_47_), .Y(core__abc_21380_n2939) );
  AND2X2 AND2X2_2263 ( .A(core__abc_21380_n2749_bF_buf6), .B(core_mi_47_), .Y(core__abc_21380_n2940) );
  AND2X2 AND2X2_2264 ( .A(core__abc_21380_n2941), .B(reset_n_bF_buf81), .Y(core_mi_reg_47__FF_INPUT) );
  AND2X2 AND2X2_2265 ( .A(core__abc_21380_n2750_bF_buf7), .B(core_mi_reg_48_), .Y(core__abc_21380_n2943) );
  AND2X2 AND2X2_2266 ( .A(core__abc_21380_n2749_bF_buf5), .B(core_mi_48_), .Y(core__abc_21380_n2944) );
  AND2X2 AND2X2_2267 ( .A(core__abc_21380_n2945), .B(reset_n_bF_buf80), .Y(core_mi_reg_48__FF_INPUT) );
  AND2X2 AND2X2_2268 ( .A(core__abc_21380_n2750_bF_buf6), .B(core_mi_reg_49_), .Y(core__abc_21380_n2947) );
  AND2X2 AND2X2_2269 ( .A(core__abc_21380_n2749_bF_buf4), .B(core_mi_49_), .Y(core__abc_21380_n2948) );
  AND2X2 AND2X2_227 ( .A(_abc_19068_n945_1_bF_buf4), .B(core_mi_15_), .Y(_abc_19068_n1280) );
  AND2X2 AND2X2_2270 ( .A(core__abc_21380_n2949), .B(reset_n_bF_buf79), .Y(core_mi_reg_49__FF_INPUT) );
  AND2X2 AND2X2_2271 ( .A(core__abc_21380_n2750_bF_buf5), .B(core_mi_reg_50_), .Y(core__abc_21380_n2951) );
  AND2X2 AND2X2_2272 ( .A(core__abc_21380_n2749_bF_buf3), .B(core_mi_50_), .Y(core__abc_21380_n2952_1) );
  AND2X2 AND2X2_2273 ( .A(core__abc_21380_n2953), .B(reset_n_bF_buf78), .Y(core_mi_reg_50__FF_INPUT) );
  AND2X2 AND2X2_2274 ( .A(core__abc_21380_n2750_bF_buf4), .B(core_mi_reg_51_), .Y(core__abc_21380_n2955) );
  AND2X2 AND2X2_2275 ( .A(core__abc_21380_n2749_bF_buf2), .B(core_mi_51_), .Y(core__abc_21380_n2956_1) );
  AND2X2 AND2X2_2276 ( .A(core__abc_21380_n2957), .B(reset_n_bF_buf77), .Y(core_mi_reg_51__FF_INPUT) );
  AND2X2 AND2X2_2277 ( .A(core__abc_21380_n2750_bF_buf3), .B(core_mi_reg_52_), .Y(core__abc_21380_n2959) );
  AND2X2 AND2X2_2278 ( .A(core__abc_21380_n2749_bF_buf1), .B(core_mi_52_), .Y(core__abc_21380_n2960) );
  AND2X2 AND2X2_2279 ( .A(core__abc_21380_n2961), .B(reset_n_bF_buf76), .Y(core_mi_reg_52__FF_INPUT) );
  AND2X2 AND2X2_228 ( .A(_abc_19068_n915_1_bF_buf3), .B(core_mi_47_), .Y(_abc_19068_n1281_1) );
  AND2X2 AND2X2_2280 ( .A(core__abc_21380_n2750_bF_buf2), .B(core_mi_reg_53_), .Y(core__abc_21380_n2963) );
  AND2X2 AND2X2_2281 ( .A(core__abc_21380_n2749_bF_buf0), .B(core_mi_53_), .Y(core__abc_21380_n2964) );
  AND2X2 AND2X2_2282 ( .A(core__abc_21380_n2965_1), .B(reset_n_bF_buf75), .Y(core_mi_reg_53__FF_INPUT) );
  AND2X2 AND2X2_2283 ( .A(core__abc_21380_n2750_bF_buf1), .B(core_mi_reg_54_), .Y(core__abc_21380_n2967) );
  AND2X2 AND2X2_2284 ( .A(core__abc_21380_n2749_bF_buf10), .B(core_mi_54_), .Y(core__abc_21380_n2968) );
  AND2X2 AND2X2_2285 ( .A(core__abc_21380_n2969), .B(reset_n_bF_buf74), .Y(core_mi_reg_54__FF_INPUT) );
  AND2X2 AND2X2_2286 ( .A(core__abc_21380_n2750_bF_buf0), .B(core_mi_reg_55_), .Y(core__abc_21380_n2971_1) );
  AND2X2 AND2X2_2287 ( .A(core__abc_21380_n2749_bF_buf9), .B(core_mi_55_), .Y(core__abc_21380_n2972) );
  AND2X2 AND2X2_2288 ( .A(core__abc_21380_n2973), .B(reset_n_bF_buf73), .Y(core_mi_reg_55__FF_INPUT) );
  AND2X2 AND2X2_2289 ( .A(core__abc_21380_n2750_bF_buf7), .B(core_mi_reg_56_), .Y(core__abc_21380_n2975) );
  AND2X2 AND2X2_229 ( .A(_abc_19068_n923_bF_buf4), .B(_abc_19068_n1285_1), .Y(_auto_iopadmap_cc_313_execute_30317_15_) );
  AND2X2 AND2X2_2290 ( .A(core__abc_21380_n2749_bF_buf8), .B(core_mi_56_), .Y(core__abc_21380_n2976) );
  AND2X2 AND2X2_2291 ( .A(core__abc_21380_n2977), .B(reset_n_bF_buf72), .Y(core_mi_reg_56__FF_INPUT) );
  AND2X2 AND2X2_2292 ( .A(core__abc_21380_n2750_bF_buf6), .B(core_mi_reg_57_), .Y(core__abc_21380_n2979) );
  AND2X2 AND2X2_2293 ( .A(core__abc_21380_n2749_bF_buf7), .B(core_mi_57_), .Y(core__abc_21380_n2980) );
  AND2X2 AND2X2_2294 ( .A(core__abc_21380_n2981), .B(reset_n_bF_buf71), .Y(core_mi_reg_57__FF_INPUT) );
  AND2X2 AND2X2_2295 ( .A(core__abc_21380_n2750_bF_buf5), .B(core_mi_reg_58_), .Y(core__abc_21380_n2983) );
  AND2X2 AND2X2_2296 ( .A(core__abc_21380_n2749_bF_buf6), .B(core_mi_58_), .Y(core__abc_21380_n2984) );
  AND2X2 AND2X2_2297 ( .A(core__abc_21380_n2985), .B(reset_n_bF_buf70), .Y(core_mi_reg_58__FF_INPUT) );
  AND2X2 AND2X2_2298 ( .A(core__abc_21380_n2750_bF_buf4), .B(core_mi_reg_59_), .Y(core__abc_21380_n2987) );
  AND2X2 AND2X2_2299 ( .A(core__abc_21380_n2749_bF_buf5), .B(core_mi_59_), .Y(core__abc_21380_n2988_1) );
  AND2X2 AND2X2_23 ( .A(_abc_19068_n901_1), .B(_abc_19068_n896), .Y(_abc_19068_n902) );
  AND2X2 AND2X2_230 ( .A(_abc_19068_n899_bF_buf2), .B(word3_reg_16_), .Y(_abc_19068_n1287_1) );
  AND2X2 AND2X2_2300 ( .A(core__abc_21380_n2989), .B(reset_n_bF_buf69), .Y(core_mi_reg_59__FF_INPUT) );
  AND2X2 AND2X2_2301 ( .A(core__abc_21380_n2750_bF_buf3), .B(core_mi_reg_60_), .Y(core__abc_21380_n2991) );
  AND2X2 AND2X2_2302 ( .A(core__abc_21380_n2749_bF_buf4), .B(core_mi_60_), .Y(core__abc_21380_n2992) );
  AND2X2 AND2X2_2303 ( .A(core__abc_21380_n2993), .B(reset_n_bF_buf68), .Y(core_mi_reg_60__FF_INPUT) );
  AND2X2 AND2X2_2304 ( .A(core__abc_21380_n2750_bF_buf2), .B(core_mi_reg_61_), .Y(core__abc_21380_n2995) );
  AND2X2 AND2X2_2305 ( .A(core__abc_21380_n2749_bF_buf3), .B(core_mi_61_), .Y(core__abc_21380_n2996) );
  AND2X2 AND2X2_2306 ( .A(core__abc_21380_n2997), .B(reset_n_bF_buf67), .Y(core_mi_reg_61__FF_INPUT) );
  AND2X2 AND2X2_2307 ( .A(core__abc_21380_n2750_bF_buf1), .B(core_mi_reg_62_), .Y(core__abc_21380_n2999) );
  AND2X2 AND2X2_2308 ( .A(core__abc_21380_n2749_bF_buf2), .B(core_mi_62_), .Y(core__abc_21380_n3000) );
  AND2X2 AND2X2_2309 ( .A(core__abc_21380_n3001_1), .B(reset_n_bF_buf66), .Y(core_mi_reg_62__FF_INPUT) );
  AND2X2 AND2X2_231 ( .A(_abc_19068_n945_1_bF_buf3), .B(core_mi_16_), .Y(_abc_19068_n1289_1) );
  AND2X2 AND2X2_2310 ( .A(core__abc_21380_n2750_bF_buf0), .B(core_mi_reg_63_), .Y(core__abc_21380_n3003) );
  AND2X2 AND2X2_2311 ( .A(core__abc_21380_n2749_bF_buf1), .B(core_mi_63_), .Y(core__abc_21380_n3004) );
  AND2X2 AND2X2_2312 ( .A(core__abc_21380_n3005_1), .B(reset_n_bF_buf65), .Y(core_mi_reg_63__FF_INPUT) );
  AND2X2 AND2X2_2313 ( .A(core__abc_21380_n3008), .B(core__abc_21380_n2027), .Y(core__abc_21380_n3009) );
  AND2X2 AND2X2_2314 ( .A(core__abc_21380_n1329), .B(core__abc_21380_n1304), .Y(core__abc_21380_n3011) );
  AND2X2 AND2X2_2315 ( .A(core__abc_21380_n1286_1), .B(core__abc_21380_n1266_1), .Y(core__abc_21380_n3013) );
  AND2X2 AND2X2_2316 ( .A(core__abc_21380_n1309), .B(core__abc_21380_n1329), .Y(core__abc_21380_n3015) );
  AND2X2 AND2X2_2317 ( .A(core__abc_21380_n3014), .B(core__abc_21380_n3015), .Y(core__abc_21380_n3016) );
  AND2X2 AND2X2_2318 ( .A(core__abc_21380_n3017), .B(core__abc_21380_n3021), .Y(core__abc_21380_n3022) );
  AND2X2 AND2X2_2319 ( .A(core__abc_21380_n1403), .B(core__abc_21380_n1379), .Y(core__abc_21380_n3028) );
  AND2X2 AND2X2_232 ( .A(_abc_19068_n941_bF_buf3), .B(core_key_112_), .Y(_abc_19068_n1290) );
  AND2X2 AND2X2_2320 ( .A(core__abc_21380_n3030_1), .B(core__abc_21380_n3027), .Y(core__abc_21380_n3031) );
  AND2X2 AND2X2_2321 ( .A(core__abc_21380_n3023), .B(core__abc_21380_n3031), .Y(core__abc_21380_n3032) );
  AND2X2 AND2X2_2322 ( .A(core__abc_21380_n1527), .B(core__abc_21380_n1546), .Y(core__abc_21380_n3033) );
  AND2X2 AND2X2_2323 ( .A(core__abc_21380_n1491), .B(core__abc_21380_n1509), .Y(core__abc_21380_n3034) );
  AND2X2 AND2X2_2324 ( .A(core__abc_21380_n3033), .B(core__abc_21380_n3034), .Y(core__abc_21380_n3035) );
  AND2X2 AND2X2_2325 ( .A(core__abc_21380_n1418), .B(core__abc_21380_n1438), .Y(core__abc_21380_n3036) );
  AND2X2 AND2X2_2326 ( .A(core__abc_21380_n1455), .B(core__abc_21380_n1472), .Y(core__abc_21380_n3037) );
  AND2X2 AND2X2_2327 ( .A(core__abc_21380_n3036), .B(core__abc_21380_n3037), .Y(core__abc_21380_n3038) );
  AND2X2 AND2X2_2328 ( .A(core__abc_21380_n3035), .B(core__abc_21380_n3038), .Y(core__abc_21380_n3039) );
  AND2X2 AND2X2_2329 ( .A(core__abc_21380_n1416), .B(core__abc_21380_n1436), .Y(core__abc_21380_n3043) );
  AND2X2 AND2X2_233 ( .A(_abc_19068_n939_1_bF_buf3), .B(core_key_80_), .Y(_abc_19068_n1293_1) );
  AND2X2 AND2X2_2330 ( .A(core__abc_21380_n3045), .B(core__abc_21380_n3037), .Y(core__abc_21380_n3046) );
  AND2X2 AND2X2_2331 ( .A(core__abc_21380_n1471), .B(core__abc_21380_n1452), .Y(core__abc_21380_n3047) );
  AND2X2 AND2X2_2332 ( .A(core__abc_21380_n3049), .B(core__abc_21380_n3035), .Y(core__abc_21380_n3050) );
  AND2X2 AND2X2_2333 ( .A(core__abc_21380_n3051), .B(core__abc_21380_n1507), .Y(core__abc_21380_n3052) );
  AND2X2 AND2X2_2334 ( .A(core__abc_21380_n3053), .B(core__abc_21380_n3033), .Y(core__abc_21380_n3054) );
  AND2X2 AND2X2_2335 ( .A(core__abc_21380_n1545), .B(core__abc_21380_n1524), .Y(core__abc_21380_n3055_1) );
  AND2X2 AND2X2_2336 ( .A(core__abc_21380_n3041), .B(core__abc_21380_n3059), .Y(core__abc_21380_n3060) );
  AND2X2 AND2X2_2337 ( .A(core__abc_21380_n1824), .B(core__abc_21380_n1843), .Y(core__abc_21380_n3061_1) );
  AND2X2 AND2X2_2338 ( .A(core__abc_21380_n1786_1), .B(core__abc_21380_n1805), .Y(core__abc_21380_n3062) );
  AND2X2 AND2X2_2339 ( .A(core__abc_21380_n3061_1), .B(core__abc_21380_n3062), .Y(core__abc_21380_n3063) );
  AND2X2 AND2X2_234 ( .A(_abc_19068_n924_1_bF_buf3), .B(core_key_48_), .Y(_abc_19068_n1294) );
  AND2X2 AND2X2_2340 ( .A(core__abc_21380_n1747), .B(core__abc_21380_n1767), .Y(core__abc_21380_n3064) );
  AND2X2 AND2X2_2341 ( .A(core__abc_21380_n1711), .B(core__abc_21380_n1730), .Y(core__abc_21380_n3065) );
  AND2X2 AND2X2_2342 ( .A(core__abc_21380_n3064), .B(core__abc_21380_n3065), .Y(core__abc_21380_n3066) );
  AND2X2 AND2X2_2343 ( .A(core__abc_21380_n3063), .B(core__abc_21380_n3066), .Y(core__abc_21380_n3067) );
  AND2X2 AND2X2_2344 ( .A(core__abc_21380_n1673), .B(core__abc_21380_n1692), .Y(core__abc_21380_n3068) );
  AND2X2 AND2X2_2345 ( .A(core__abc_21380_n1637), .B(core__abc_21380_n1655_1), .Y(core__abc_21380_n3069) );
  AND2X2 AND2X2_2346 ( .A(core__abc_21380_n3068), .B(core__abc_21380_n3069), .Y(core__abc_21380_n3070) );
  AND2X2 AND2X2_2347 ( .A(core__abc_21380_n1565), .B(core__abc_21380_n1584), .Y(core__abc_21380_n3071) );
  AND2X2 AND2X2_2348 ( .A(core__abc_21380_n1601), .B(core__abc_21380_n1618), .Y(core__abc_21380_n3072) );
  AND2X2 AND2X2_2349 ( .A(core__abc_21380_n3071), .B(core__abc_21380_n3072), .Y(core__abc_21380_n3073_1) );
  AND2X2 AND2X2_235 ( .A(_abc_19068_n926_bF_buf3), .B(core_key_16_), .Y(_abc_19068_n1295_1) );
  AND2X2 AND2X2_2350 ( .A(core__abc_21380_n3070), .B(core__abc_21380_n3073_1), .Y(core__abc_21380_n3074) );
  AND2X2 AND2X2_2351 ( .A(core__abc_21380_n3067), .B(core__abc_21380_n3074), .Y(core__abc_21380_n3075) );
  AND2X2 AND2X2_2352 ( .A(core__abc_21380_n1563), .B(core__abc_21380_n1582), .Y(core__abc_21380_n3079) );
  AND2X2 AND2X2_2353 ( .A(core__abc_21380_n3081), .B(core__abc_21380_n3072), .Y(core__abc_21380_n3082) );
  AND2X2 AND2X2_2354 ( .A(core__abc_21380_n1617), .B(core__abc_21380_n1598), .Y(core__abc_21380_n3083) );
  AND2X2 AND2X2_2355 ( .A(core__abc_21380_n3085), .B(core__abc_21380_n3070), .Y(core__abc_21380_n3086) );
  AND2X2 AND2X2_2356 ( .A(core__abc_21380_n3087), .B(core__abc_21380_n1653), .Y(core__abc_21380_n3088) );
  AND2X2 AND2X2_2357 ( .A(core__abc_21380_n3089), .B(core__abc_21380_n3068), .Y(core__abc_21380_n3090) );
  AND2X2 AND2X2_2358 ( .A(core__abc_21380_n1691), .B(core__abc_21380_n1670), .Y(core__abc_21380_n3091_1) );
  AND2X2 AND2X2_2359 ( .A(core__abc_21380_n3094), .B(core__abc_21380_n3067), .Y(core__abc_21380_n3095_1) );
  AND2X2 AND2X2_236 ( .A(_abc_19068_n916_1_bF_buf2), .B(word1_reg_16_), .Y(_abc_19068_n1298_1) );
  AND2X2 AND2X2_2360 ( .A(core__abc_21380_n3096), .B(core__abc_21380_n1728), .Y(core__abc_21380_n3097) );
  AND2X2 AND2X2_2361 ( .A(core__abc_21380_n3098), .B(core__abc_21380_n3064), .Y(core__abc_21380_n3099) );
  AND2X2 AND2X2_2362 ( .A(core__abc_21380_n1766), .B(core__abc_21380_n1744), .Y(core__abc_21380_n3100) );
  AND2X2 AND2X2_2363 ( .A(core__abc_21380_n3102), .B(core__abc_21380_n3063), .Y(core__abc_21380_n3103) );
  AND2X2 AND2X2_2364 ( .A(core__abc_21380_n1842), .B(core__abc_21380_n1821), .Y(core__abc_21380_n3104_1) );
  AND2X2 AND2X2_2365 ( .A(core__abc_21380_n1784), .B(core__abc_21380_n1803), .Y(core__abc_21380_n3107) );
  AND2X2 AND2X2_2366 ( .A(core__abc_21380_n3109), .B(core__abc_21380_n3061_1), .Y(core__abc_21380_n3110_1) );
  AND2X2 AND2X2_2367 ( .A(core__abc_21380_n3077_1), .B(core__abc_21380_n3114), .Y(core__abc_21380_n3115) );
  AND2X2 AND2X2_2368 ( .A(core__abc_21380_n1974), .B(core__abc_21380_n1993), .Y(core__abc_21380_n3116) );
  AND2X2 AND2X2_2369 ( .A(core__abc_21380_n1935), .B(core__abc_21380_n1955), .Y(core__abc_21380_n3117) );
  AND2X2 AND2X2_237 ( .A(_abc_19068_n902_bF_buf2), .B(word2_reg_16_), .Y(_abc_19068_n1299) );
  AND2X2 AND2X2_2370 ( .A(core__abc_21380_n3116), .B(core__abc_21380_n3117), .Y(core__abc_21380_n3118) );
  AND2X2 AND2X2_2371 ( .A(core__abc_21380_n1862), .B(core__abc_21380_n1880), .Y(core__abc_21380_n3119) );
  AND2X2 AND2X2_2372 ( .A(core__abc_21380_n1898), .B(core__abc_21380_n1917), .Y(core__abc_21380_n3120) );
  AND2X2 AND2X2_2373 ( .A(core__abc_21380_n3119), .B(core__abc_21380_n3120), .Y(core__abc_21380_n3121) );
  AND2X2 AND2X2_2374 ( .A(core__abc_21380_n3118), .B(core__abc_21380_n3121), .Y(core__abc_21380_n3122_1) );
  AND2X2 AND2X2_2375 ( .A(core__abc_21380_n1860), .B(core__abc_21380_n1878), .Y(core__abc_21380_n3126) );
  AND2X2 AND2X2_2376 ( .A(core__abc_21380_n3128_1), .B(core__abc_21380_n3120), .Y(core__abc_21380_n3129) );
  AND2X2 AND2X2_2377 ( .A(core__abc_21380_n1916), .B(core__abc_21380_n1895), .Y(core__abc_21380_n3130) );
  AND2X2 AND2X2_2378 ( .A(core__abc_21380_n3132), .B(core__abc_21380_n3118), .Y(core__abc_21380_n3133) );
  AND2X2 AND2X2_2379 ( .A(core__abc_21380_n3134), .B(core__abc_21380_n1953), .Y(core__abc_21380_n3135) );
  AND2X2 AND2X2_238 ( .A(_abc_19068_n897_1_bF_buf2), .B(word0_reg_16_), .Y(_abc_19068_n1301) );
  AND2X2 AND2X2_2380 ( .A(core__abc_21380_n3136), .B(core__abc_21380_n3116), .Y(core__abc_21380_n3137) );
  AND2X2 AND2X2_2381 ( .A(core__abc_21380_n1992), .B(core__abc_21380_n1971), .Y(core__abc_21380_n3138) );
  AND2X2 AND2X2_2382 ( .A(core__abc_21380_n3124), .B(core__abc_21380_n3142), .Y(core__abc_21380_n3143) );
  AND2X2 AND2X2_2383 ( .A(core__abc_21380_n2012), .B(core__abc_21380_n2029), .Y(core__abc_21380_n3145_1) );
  AND2X2 AND2X2_2384 ( .A(core__abc_21380_n3144), .B(core__abc_21380_n3145_1), .Y(core__abc_21380_n3146) );
  AND2X2 AND2X2_2385 ( .A(core__abc_21380_n3147), .B(core__abc_21380_n2048), .Y(core__abc_21380_n3148) );
  AND2X2 AND2X2_2386 ( .A(core__abc_21380_n3149), .B(core__abc_21380_n2046), .Y(core__abc_21380_n3150) );
  AND2X2 AND2X2_2387 ( .A(core__abc_21380_n3150), .B(core__abc_21380_n2070), .Y(core__abc_21380_n3151) );
  AND2X2 AND2X2_2388 ( .A(core__abc_21380_n3152), .B(core__abc_21380_n3153), .Y(core__abc_21380_n3154) );
  AND2X2 AND2X2_2389 ( .A(core__abc_21380_n3158), .B(core__abc_21380_n3155), .Y(core__abc_21380_n3159) );
  AND2X2 AND2X2_239 ( .A(_abc_19068_n915_1_bF_buf2), .B(core_mi_48_), .Y(_abc_19068_n1302_1) );
  AND2X2 AND2X2_2390 ( .A(core__abc_21380_n2715), .B(core__abc_21380_n1142_1), .Y(core__abc_21380_n3160) );
  AND2X2 AND2X2_2391 ( .A(core__abc_21380_n1143), .B(core__abc_21380_n1144_1), .Y(core__abc_21380_n3162) );
  AND2X2 AND2X2_2392 ( .A(core__abc_21380_n3162), .B(core__abc_21380_n1255), .Y(core__abc_21380_n3163_1) );
  AND2X2 AND2X2_2393 ( .A(core__abc_21380_n3164), .B(core__abc_21380_n1136_1), .Y(core__abc_21380_n3165) );
  AND2X2 AND2X2_2394 ( .A(core__abc_21380_n3165), .B(core__abc_21380_n2711), .Y(core__abc_21380_n3166) );
  AND2X2 AND2X2_2395 ( .A(core__abc_21380_n3166), .B(core__abc_21380_n3161), .Y(core__abc_21380_n3167_1) );
  AND2X2 AND2X2_2396 ( .A(core__abc_21380_n1280_1), .B(core__abc_21380_n1260_1), .Y(core__abc_21380_n3168) );
  AND2X2 AND2X2_2397 ( .A(core__abc_21380_n3169), .B(core__abc_21380_n3171), .Y(core__abc_21380_n3172) );
  AND2X2 AND2X2_2398 ( .A(core__abc_21380_n3173), .B(core__abc_21380_n1301), .Y(core__abc_21380_n3174) );
  AND2X2 AND2X2_2399 ( .A(core__abc_21380_n1378), .B(core__abc_21380_n1397), .Y(core__abc_21380_n3177_1) );
  AND2X2 AND2X2_24 ( .A(_abc_19068_n894_1), .B(_abc_19068_n881), .Y(_abc_19068_n906_1) );
  AND2X2 AND2X2_240 ( .A(_abc_19068_n923_bF_buf3), .B(_abc_19068_n1306_1), .Y(_auto_iopadmap_cc_313_execute_30317_16_) );
  AND2X2 AND2X2_2400 ( .A(core__abc_21380_n1359), .B(core__abc_21380_n1339), .Y(core__abc_21380_n3178) );
  AND2X2 AND2X2_2401 ( .A(core__abc_21380_n3177_1), .B(core__abc_21380_n3178), .Y(core__abc_21380_n3179) );
  AND2X2 AND2X2_2402 ( .A(core__abc_21380_n3176), .B(core__abc_21380_n3179), .Y(core__abc_21380_n3180) );
  AND2X2 AND2X2_2403 ( .A(core__abc_21380_n3182), .B(core__abc_21380_n3181_1), .Y(core__abc_21380_n3183) );
  AND2X2 AND2X2_2404 ( .A(core__abc_21380_n3177_1), .B(core__abc_21380_n3183), .Y(core__abc_21380_n3184) );
  AND2X2 AND2X2_2405 ( .A(core__abc_21380_n3185), .B(core__abc_21380_n1376), .Y(core__abc_21380_n3186) );
  AND2X2 AND2X2_2406 ( .A(core__abc_21380_n1523), .B(core__abc_21380_n1542), .Y(core__abc_21380_n3190) );
  AND2X2 AND2X2_2407 ( .A(core__abc_21380_n3192), .B(core__abc_21380_n3190), .Y(core__abc_21380_n3193) );
  AND2X2 AND2X2_2408 ( .A(core__abc_21380_n1434), .B(core__abc_21380_n1414), .Y(core__abc_21380_n3194_1) );
  AND2X2 AND2X2_2409 ( .A(core__abc_21380_n1451), .B(core__abc_21380_n1468), .Y(core__abc_21380_n3195) );
  AND2X2 AND2X2_241 ( .A(_abc_19068_n915_1_bF_buf1), .B(core_mi_49_), .Y(_abc_19068_n1308_1) );
  AND2X2 AND2X2_2410 ( .A(core__abc_21380_n3194_1), .B(core__abc_21380_n3195), .Y(core__abc_21380_n3196) );
  AND2X2 AND2X2_2411 ( .A(core__abc_21380_n3193), .B(core__abc_21380_n3196), .Y(core__abc_21380_n3197) );
  AND2X2 AND2X2_2412 ( .A(core__abc_21380_n3189), .B(core__abc_21380_n3197), .Y(core__abc_21380_n3198) );
  AND2X2 AND2X2_2413 ( .A(core__abc_21380_n3199), .B(core__abc_21380_n1433), .Y(core__abc_21380_n3200_1) );
  AND2X2 AND2X2_2414 ( .A(core__abc_21380_n3195), .B(core__abc_21380_n3200_1), .Y(core__abc_21380_n3201) );
  AND2X2 AND2X2_2415 ( .A(core__abc_21380_n1465), .B(core__abc_21380_n1449), .Y(core__abc_21380_n3202) );
  AND2X2 AND2X2_2416 ( .A(core__abc_21380_n3204), .B(core__abc_21380_n3193), .Y(core__abc_21380_n3205) );
  AND2X2 AND2X2_2417 ( .A(core__abc_21380_n3209), .B(core__abc_21380_n3190), .Y(core__abc_21380_n3210) );
  AND2X2 AND2X2_2418 ( .A(core__abc_21380_n1539), .B(core__abc_21380_n1521), .Y(core__abc_21380_n3211_1) );
  AND2X2 AND2X2_2419 ( .A(core__abc_21380_n1820), .B(core__abc_21380_n1839), .Y(core__abc_21380_n3216) );
  AND2X2 AND2X2_242 ( .A(_abc_19068_n897_1_bF_buf1), .B(word0_reg_17_), .Y(_abc_19068_n1309) );
  AND2X2 AND2X2_2420 ( .A(core__abc_21380_n1782_1), .B(core__abc_21380_n1801), .Y(core__abc_21380_n3217) );
  AND2X2 AND2X2_2421 ( .A(core__abc_21380_n3216), .B(core__abc_21380_n3217), .Y(core__abc_21380_n3218) );
  AND2X2 AND2X2_2422 ( .A(core__abc_21380_n1707), .B(core__abc_21380_n1726), .Y(core__abc_21380_n3219) );
  AND2X2 AND2X2_2423 ( .A(core__abc_21380_n1763), .B(core__abc_21380_n1743), .Y(core__abc_21380_n3220) );
  AND2X2 AND2X2_2424 ( .A(core__abc_21380_n3219), .B(core__abc_21380_n3220), .Y(core__abc_21380_n3221) );
  AND2X2 AND2X2_2425 ( .A(core__abc_21380_n3218), .B(core__abc_21380_n3221), .Y(core__abc_21380_n3222) );
  AND2X2 AND2X2_2426 ( .A(core__abc_21380_n1669), .B(core__abc_21380_n1688), .Y(core__abc_21380_n3223) );
  AND2X2 AND2X2_2427 ( .A(core__abc_21380_n3225), .B(core__abc_21380_n3223), .Y(core__abc_21380_n3226) );
  AND2X2 AND2X2_2428 ( .A(core__abc_21380_n1561), .B(core__abc_21380_n1580), .Y(core__abc_21380_n3227) );
  AND2X2 AND2X2_2429 ( .A(core__abc_21380_n1597), .B(core__abc_21380_n1614), .Y(core__abc_21380_n3228) );
  AND2X2 AND2X2_243 ( .A(_abc_19068_n916_1_bF_buf1), .B(word1_reg_17_), .Y(_abc_19068_n1311) );
  AND2X2 AND2X2_2430 ( .A(core__abc_21380_n3227), .B(core__abc_21380_n3228), .Y(core__abc_21380_n3229) );
  AND2X2 AND2X2_2431 ( .A(core__abc_21380_n3226), .B(core__abc_21380_n3229), .Y(core__abc_21380_n3230_1) );
  AND2X2 AND2X2_2432 ( .A(core__abc_21380_n3230_1), .B(core__abc_21380_n3222), .Y(core__abc_21380_n3231) );
  AND2X2 AND2X2_2433 ( .A(core__abc_21380_n3215_1), .B(core__abc_21380_n3231), .Y(core__abc_21380_n3232) );
  AND2X2 AND2X2_2434 ( .A(core__abc_21380_n3233), .B(core__abc_21380_n1579), .Y(core__abc_21380_n3234) );
  AND2X2 AND2X2_2435 ( .A(core__abc_21380_n3228), .B(core__abc_21380_n3234), .Y(core__abc_21380_n3235) );
  AND2X2 AND2X2_2436 ( .A(core__abc_21380_n1613), .B(core__abc_21380_n1595), .Y(core__abc_21380_n3236_1) );
  AND2X2 AND2X2_2437 ( .A(core__abc_21380_n3238), .B(core__abc_21380_n3226), .Y(core__abc_21380_n3239) );
  AND2X2 AND2X2_2438 ( .A(core__abc_21380_n3243), .B(core__abc_21380_n3223), .Y(core__abc_21380_n3244) );
  AND2X2 AND2X2_2439 ( .A(core__abc_21380_n1685), .B(core__abc_21380_n1667), .Y(core__abc_21380_n3245_1) );
  AND2X2 AND2X2_244 ( .A(_abc_19068_n939_1_bF_buf2), .B(core_key_81_), .Y(_abc_19068_n1314_1) );
  AND2X2 AND2X2_2440 ( .A(core__abc_21380_n3248), .B(core__abc_21380_n3222), .Y(core__abc_21380_n3249) );
  AND2X2 AND2X2_2441 ( .A(core__abc_21380_n3250), .B(core__abc_21380_n1725), .Y(core__abc_21380_n3251_1) );
  AND2X2 AND2X2_2442 ( .A(core__abc_21380_n3253), .B(core__abc_21380_n3220), .Y(core__abc_21380_n3254) );
  AND2X2 AND2X2_2443 ( .A(core__abc_21380_n1760_1), .B(core__abc_21380_n1741), .Y(core__abc_21380_n3255) );
  AND2X2 AND2X2_2444 ( .A(core__abc_21380_n3257), .B(core__abc_21380_n3218), .Y(core__abc_21380_n3258) );
  AND2X2 AND2X2_2445 ( .A(core__abc_21380_n1836), .B(core__abc_21380_n1818), .Y(core__abc_21380_n3259) );
  AND2X2 AND2X2_2446 ( .A(core__abc_21380_n3261), .B(core__abc_21380_n1800), .Y(core__abc_21380_n3262_1) );
  AND2X2 AND2X2_2447 ( .A(core__abc_21380_n3264), .B(core__abc_21380_n3216), .Y(core__abc_21380_n3265) );
  AND2X2 AND2X2_2448 ( .A(core__abc_21380_n3269), .B(core__abc_21380_n1858), .Y(core__abc_21380_n3270) );
  AND2X2 AND2X2_2449 ( .A(core__abc_21380_n3271), .B(core__abc_21380_n1279), .Y(core__abc_21380_n3272) );
  AND2X2 AND2X2_245 ( .A(_abc_19068_n924_1_bF_buf2), .B(core_key_49_), .Y(_abc_19068_n1315) );
  AND2X2 AND2X2_2450 ( .A(core__abc_21380_n3273), .B(core__abc_21380_n3274), .Y(core__abc_21380_n3275) );
  AND2X2 AND2X2_2451 ( .A(core__abc_21380_n3277_1), .B(core__abc_21380_n3278), .Y(core__abc_21380_n3279) );
  AND2X2 AND2X2_2452 ( .A(core__abc_21380_n3281_1), .B(core__abc_21380_n3282), .Y(core__abc_21380_n3283) );
  AND2X2 AND2X2_2453 ( .A(core__abc_21380_n3285), .B(core__abc_21380_n3286), .Y(core__abc_21380_n3287) );
  AND2X2 AND2X2_2454 ( .A(core__abc_21380_n3287), .B(core__abc_21380_n1857), .Y(core__abc_21380_n3288) );
  AND2X2 AND2X2_2455 ( .A(core__abc_21380_n1267), .B(core_v3_reg_48_), .Y(core__abc_21380_n3291) );
  AND2X2 AND2X2_2456 ( .A(core__abc_21380_n3292), .B(core__abc_21380_n3293), .Y(core__abc_21380_n3294) );
  AND2X2 AND2X2_2457 ( .A(core__abc_21380_n3290), .B(core__abc_21380_n3295), .Y(core__abc_21380_n3296) );
  AND2X2 AND2X2_2458 ( .A(core__abc_21380_n3289), .B(core__abc_21380_n3294), .Y(core__abc_21380_n3297) );
  AND2X2 AND2X2_2459 ( .A(core__abc_21380_n3298), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf3), .Y(core__abc_21380_n3299) );
  AND2X2 AND2X2_246 ( .A(_abc_19068_n926_bF_buf2), .B(core_key_17_), .Y(_abc_19068_n1316_1) );
  AND2X2 AND2X2_2460 ( .A(core__abc_21380_n3157), .B(core_v3_reg_27_), .Y(core__abc_21380_n3301) );
  AND2X2 AND2X2_2461 ( .A(core__abc_21380_n3154), .B(core__abc_21380_n3007), .Y(core__abc_21380_n3302) );
  AND2X2 AND2X2_2462 ( .A(core__abc_21380_n3304), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf3), .Y(core__abc_21380_n3305) );
  AND2X2 AND2X2_2463 ( .A(core__abc_21380_n3306), .B(core__abc_21380_n3300), .Y(core__abc_21380_n3307) );
  AND2X2 AND2X2_2464 ( .A(core__abc_21380_n3162), .B(core__abc_21380_n1132_1), .Y(core__abc_21380_n3308) );
  AND2X2 AND2X2_2465 ( .A(core__abc_21380_n1241_1), .B(core__abc_21380_n1138_1), .Y(core__abc_21380_n3309) );
  AND2X2 AND2X2_2466 ( .A(core__abc_21380_n3309), .B(core__abc_21380_n1142_1), .Y(core__abc_21380_n3310) );
  AND2X2 AND2X2_2467 ( .A(core__abc_21380_n3160), .B(core__abc_21380_n1137_1), .Y(core__abc_21380_n3312) );
  AND2X2 AND2X2_2468 ( .A(core__abc_21380_n3312), .B(core__abc_21380_n3165), .Y(core__abc_21380_n3313) );
  AND2X2 AND2X2_2469 ( .A(core__abc_21380_n3315), .B(core__abc_21380_n2750_bF_buf7), .Y(core__abc_21380_n3316) );
  AND2X2 AND2X2_247 ( .A(_abc_19068_n941_bF_buf2), .B(core_key_113_), .Y(_abc_19068_n1319) );
  AND2X2 AND2X2_2470 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n3318), .Y(core__abc_21380_n3319) );
  AND2X2 AND2X2_2471 ( .A(core_v3_reg_0_), .B(core_mi_0_), .Y(core__abc_21380_n3321) );
  AND2X2 AND2X2_2472 ( .A(core__abc_21380_n3322), .B(core__abc_21380_n3320), .Y(core__abc_21380_n3323) );
  AND2X2 AND2X2_2473 ( .A(core__abc_21380_n2749_bF_buf0), .B(core__abc_21380_n3323), .Y(core__abc_21380_n3324) );
  AND2X2 AND2X2_2474 ( .A(core__abc_21380_n3329), .B(reset_n_bF_buf64), .Y(core__abc_21380_n3330) );
  AND2X2 AND2X2_2475 ( .A(core__abc_21380_n3327), .B(core__abc_21380_n3330), .Y(core_v3_reg_0__FF_INPUT) );
  AND2X2 AND2X2_2476 ( .A(core__abc_21380_n1876), .B(core__abc_21380_n1856), .Y(core__abc_21380_n3332) );
  AND2X2 AND2X2_2477 ( .A(core__abc_21380_n1858), .B(core__abc_21380_n1876), .Y(core__abc_21380_n3336) );
  AND2X2 AND2X2_2478 ( .A(core__abc_21380_n3269), .B(core__abc_21380_n3336), .Y(core__abc_21380_n3337) );
  AND2X2 AND2X2_2479 ( .A(core__abc_21380_n3335), .B(core__abc_21380_n3338), .Y(core__abc_21380_n3339) );
  AND2X2 AND2X2_248 ( .A(_abc_19068_n945_1_bF_buf2), .B(core_mi_17_), .Y(_abc_19068_n1320_1) );
  AND2X2 AND2X2_2480 ( .A(core__abc_21380_n3339), .B(core__abc_21380_n3333), .Y(core__abc_21380_n3340) );
  AND2X2 AND2X2_2481 ( .A(core__abc_21380_n1285_1), .B(core__abc_21380_n3342), .Y(core__abc_21380_n3343) );
  AND2X2 AND2X2_2482 ( .A(core__abc_21380_n3346), .B(core__abc_21380_n3347), .Y(core__abc_21380_n3348) );
  AND2X2 AND2X2_2483 ( .A(core__abc_21380_n3340), .B(core__abc_21380_n3349), .Y(core__abc_21380_n3350) );
  AND2X2 AND2X2_2484 ( .A(core__abc_21380_n3351), .B(core__abc_21380_n3352), .Y(core__abc_21380_n3353) );
  AND2X2 AND2X2_2485 ( .A(core__abc_21380_n3353), .B(core__abc_21380_n3296), .Y(core__abc_21380_n3354) );
  AND2X2 AND2X2_2486 ( .A(core__abc_21380_n3357), .B(core__abc_21380_n1876), .Y(core__abc_21380_n3358) );
  AND2X2 AND2X2_2487 ( .A(core__abc_21380_n3359), .B(core__abc_21380_n3348), .Y(core__abc_21380_n3360) );
  AND2X2 AND2X2_2488 ( .A(core__abc_21380_n3361), .B(core__abc_21380_n3355), .Y(core__abc_21380_n3362) );
  AND2X2 AND2X2_2489 ( .A(core__abc_21380_n2048), .B(core__abc_21380_n2067_1), .Y(core__abc_21380_n3366) );
  AND2X2 AND2X2_249 ( .A(_abc_19068_n899_bF_buf1), .B(word3_reg_17_), .Y(_abc_19068_n1322_1) );
  AND2X2 AND2X2_2490 ( .A(core__abc_21380_n3010), .B(core__abc_21380_n3366), .Y(core__abc_21380_n3367) );
  AND2X2 AND2X2_2491 ( .A(core__abc_21380_n2064), .B(core__abc_21380_n2045), .Y(core__abc_21380_n3368) );
  AND2X2 AND2X2_2492 ( .A(core__abc_21380_n3145_1), .B(core__abc_21380_n3366), .Y(core__abc_21380_n3372) );
  AND2X2 AND2X2_2493 ( .A(core__abc_21380_n3374), .B(core__abc_21380_n3371), .Y(core__abc_21380_n3375) );
  AND2X2 AND2X2_2494 ( .A(core__abc_21380_n3376), .B(core__abc_21380_n2085), .Y(core__abc_21380_n3377) );
  AND2X2 AND2X2_2495 ( .A(core__abc_21380_n3375), .B(core__abc_21380_n2088), .Y(core__abc_21380_n3378) );
  AND2X2 AND2X2_2496 ( .A(core__abc_21380_n3381), .B(core__abc_21380_n3382), .Y(core__abc_21380_n3383) );
  AND2X2 AND2X2_2497 ( .A(core__abc_21380_n3386), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n3387) );
  AND2X2 AND2X2_2498 ( .A(core__abc_21380_n3387), .B(core__abc_21380_n3385), .Y(core__abc_21380_n3388) );
  AND2X2 AND2X2_2499 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n3389), .Y(core__abc_21380_n3390) );
  AND2X2 AND2X2_25 ( .A(_abc_19068_n893), .B(_abc_19068_n873_1), .Y(_abc_19068_n907_1) );
  AND2X2 AND2X2_250 ( .A(_abc_19068_n902_bF_buf1), .B(word2_reg_17_), .Y(_abc_19068_n1323) );
  AND2X2 AND2X2_2500 ( .A(core_v3_reg_1_), .B(core_mi_1_), .Y(core__abc_21380_n3392) );
  AND2X2 AND2X2_2501 ( .A(core__abc_21380_n3393), .B(core__abc_21380_n3391), .Y(core__abc_21380_n3394) );
  AND2X2 AND2X2_2502 ( .A(core__abc_21380_n2749_bF_buf10), .B(core__abc_21380_n3394), .Y(core__abc_21380_n3395) );
  AND2X2 AND2X2_2503 ( .A(core__abc_21380_n3399), .B(reset_n_bF_buf63), .Y(core__abc_21380_n3400) );
  AND2X2 AND2X2_2504 ( .A(core__abc_21380_n3398), .B(core__abc_21380_n3400), .Y(core_v3_reg_1__FF_INPUT) );
  AND2X2 AND2X2_2505 ( .A(core__abc_21380_n3402), .B(core__abc_21380_n3351), .Y(core__abc_21380_n3403) );
  AND2X2 AND2X2_2506 ( .A(core__abc_21380_n3406), .B(core__abc_21380_n1893), .Y(core__abc_21380_n3407) );
  AND2X2 AND2X2_2507 ( .A(core__abc_21380_n3405), .B(core__abc_21380_n1894_1), .Y(core__abc_21380_n3408) );
  AND2X2 AND2X2_2508 ( .A(core__abc_21380_n3014), .B(core__abc_21380_n1309), .Y(core__abc_21380_n3412) );
  AND2X2 AND2X2_2509 ( .A(core__abc_21380_n3413), .B(core__abc_21380_n1308), .Y(core__abc_21380_n3414) );
  AND2X2 AND2X2_251 ( .A(_abc_19068_n923_bF_buf2), .B(_abc_19068_n1327), .Y(_auto_iopadmap_cc_313_execute_30317_17_) );
  AND2X2 AND2X2_2510 ( .A(core__abc_21380_n3417), .B(core__abc_21380_n3418), .Y(core__abc_21380_n3419) );
  AND2X2 AND2X2_2511 ( .A(core__abc_21380_n3410), .B(core__abc_21380_n3420), .Y(core__abc_21380_n3421) );
  AND2X2 AND2X2_2512 ( .A(core__abc_21380_n3409), .B(core__abc_21380_n3419), .Y(core__abc_21380_n3422) );
  AND2X2 AND2X2_2513 ( .A(core__abc_21380_n3403), .B(core__abc_21380_n3423), .Y(core__abc_21380_n3424) );
  AND2X2 AND2X2_2514 ( .A(core__abc_21380_n3425), .B(core__abc_21380_n3426), .Y(core__abc_21380_n3427) );
  AND2X2 AND2X2_2515 ( .A(core__abc_21380_n3431), .B(core__abc_21380_n2108), .Y(core__abc_21380_n3432) );
  AND2X2 AND2X2_2516 ( .A(core__abc_21380_n3430), .B(core__abc_21380_n2105), .Y(core__abc_21380_n3433) );
  AND2X2 AND2X2_2517 ( .A(core__abc_21380_n3434), .B(core__abc_21380_n3429), .Y(core__abc_21380_n3435) );
  AND2X2 AND2X2_2518 ( .A(core__abc_21380_n3436), .B(core_v3_reg_29_), .Y(core__abc_21380_n3437) );
  AND2X2 AND2X2_2519 ( .A(core__abc_21380_n3441), .B(core__abc_21380_n3442), .Y(core__abc_21380_n3443) );
  AND2X2 AND2X2_252 ( .A(_abc_19068_n939_1_bF_buf1), .B(core_key_82_), .Y(_abc_19068_n1329) );
  AND2X2 AND2X2_2520 ( .A(core__abc_21380_n3444), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n3445) );
  AND2X2 AND2X2_2521 ( .A(core__abc_21380_n3445), .B(core__abc_21380_n3439), .Y(core__abc_21380_n3446) );
  AND2X2 AND2X2_2522 ( .A(core__abc_21380_n3313_bF_buf9), .B(core_key_66_), .Y(core__abc_21380_n3447) );
  AND2X2 AND2X2_2523 ( .A(core_v3_reg_2_), .B(core_mi_2_), .Y(core__abc_21380_n3449) );
  AND2X2 AND2X2_2524 ( .A(core__abc_21380_n3450), .B(core__abc_21380_n3448), .Y(core__abc_21380_n3451) );
  AND2X2 AND2X2_2525 ( .A(core__abc_21380_n2749_bF_buf9), .B(core__abc_21380_n3451), .Y(core__abc_21380_n3452) );
  AND2X2 AND2X2_2526 ( .A(core__abc_21380_n3456), .B(reset_n_bF_buf62), .Y(core__abc_21380_n3457) );
  AND2X2 AND2X2_2527 ( .A(core__abc_21380_n3455), .B(core__abc_21380_n3457), .Y(core_v3_reg_2__FF_INPUT) );
  AND2X2 AND2X2_2528 ( .A(core__abc_21380_n3460), .B(core__abc_21380_n1919), .Y(core__abc_21380_n3461) );
  AND2X2 AND2X2_2529 ( .A(core__abc_21380_n3459), .B(core__abc_21380_n1913), .Y(core__abc_21380_n3462) );
  AND2X2 AND2X2_253 ( .A(_abc_19068_n926_bF_buf1), .B(core_key_18_), .Y(_abc_19068_n1330_1) );
  AND2X2 AND2X2_2530 ( .A(core__abc_21380_n3465), .B(core__abc_21380_n3464), .Y(core__abc_21380_n3466) );
  AND2X2 AND2X2_2531 ( .A(core__abc_21380_n3467), .B(core__abc_21380_n1327), .Y(core__abc_21380_n3468) );
  AND2X2 AND2X2_2532 ( .A(core__abc_21380_n3466), .B(core__abc_21380_n1329), .Y(core__abc_21380_n3469) );
  AND2X2 AND2X2_2533 ( .A(core__abc_21380_n3472), .B(core__abc_21380_n3474), .Y(core__abc_21380_n3475) );
  AND2X2 AND2X2_2534 ( .A(core__abc_21380_n3479), .B(core__abc_21380_n3476), .Y(core__abc_21380_n3480) );
  AND2X2 AND2X2_2535 ( .A(core__abc_21380_n3483_1), .B(core__abc_21380_n3482), .Y(core__abc_21380_n3484) );
  AND2X2 AND2X2_2536 ( .A(core__abc_21380_n3484), .B(core__abc_21380_n3481), .Y(core__abc_21380_n3485_1) );
  AND2X2 AND2X2_2537 ( .A(core__abc_21380_n2085), .B(core__abc_21380_n2105), .Y(core__abc_21380_n3490_1) );
  AND2X2 AND2X2_2538 ( .A(core__abc_21380_n2084), .B(core__abc_21380_n2104), .Y(core__abc_21380_n3494) );
  AND2X2 AND2X2_2539 ( .A(core__abc_21380_n3492), .B(core__abc_21380_n3495), .Y(core__abc_21380_n3496) );
  AND2X2 AND2X2_254 ( .A(_abc_19068_n924_1_bF_buf1), .B(core_key_50_), .Y(_abc_19068_n1331) );
  AND2X2 AND2X2_2540 ( .A(core__abc_21380_n3496), .B(core__abc_21380_n2126), .Y(core__abc_21380_n3497) );
  AND2X2 AND2X2_2541 ( .A(core__abc_21380_n3498), .B(core__abc_21380_n2123), .Y(core__abc_21380_n3499) );
  AND2X2 AND2X2_2542 ( .A(core__abc_21380_n3502), .B(core__abc_21380_n3504), .Y(core__abc_21380_n3505_1) );
  AND2X2 AND2X2_2543 ( .A(core__abc_21380_n3508), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n3509) );
  AND2X2 AND2X2_2544 ( .A(core__abc_21380_n3509), .B(core__abc_21380_n3506), .Y(core__abc_21380_n3510) );
  AND2X2 AND2X2_2545 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_67_), .Y(core__abc_21380_n3511) );
  AND2X2 AND2X2_2546 ( .A(core_v3_reg_3_), .B(core_mi_3_), .Y(core__abc_21380_n3513) );
  AND2X2 AND2X2_2547 ( .A(core__abc_21380_n3514), .B(core__abc_21380_n3512), .Y(core__abc_21380_n3515) );
  AND2X2 AND2X2_2548 ( .A(core__abc_21380_n2749_bF_buf8), .B(core__abc_21380_n3515), .Y(core__abc_21380_n3516) );
  AND2X2 AND2X2_2549 ( .A(core__abc_21380_n3520), .B(reset_n_bF_buf61), .Y(core__abc_21380_n3521) );
  AND2X2 AND2X2_255 ( .A(_abc_19068_n899_bF_buf0), .B(word3_reg_18_), .Y(_abc_19068_n1334_1) );
  AND2X2 AND2X2_2550 ( .A(core__abc_21380_n3519), .B(core__abc_21380_n3521), .Y(core_v3_reg_3__FF_INPUT) );
  AND2X2 AND2X2_2551 ( .A(core__abc_21380_n1894_1), .B(core__abc_21380_n1913), .Y(core__abc_21380_n3523) );
  AND2X2 AND2X2_2552 ( .A(core__abc_21380_n3404), .B(core__abc_21380_n3523), .Y(core__abc_21380_n3524) );
  AND2X2 AND2X2_2553 ( .A(core__abc_21380_n1910), .B(core__abc_21380_n1892), .Y(core__abc_21380_n3525) );
  AND2X2 AND2X2_2554 ( .A(core__abc_21380_n3336), .B(core__abc_21380_n3523), .Y(core__abc_21380_n3528) );
  AND2X2 AND2X2_2555 ( .A(core__abc_21380_n3269), .B(core__abc_21380_n3528), .Y(core__abc_21380_n3529) );
  AND2X2 AND2X2_2556 ( .A(core__abc_21380_n3530), .B(core__abc_21380_n1937), .Y(core__abc_21380_n3531_1) );
  AND2X2 AND2X2_2557 ( .A(core__abc_21380_n3534), .B(core__abc_21380_n3532), .Y(core__abc_21380_n3535_1) );
  AND2X2 AND2X2_2558 ( .A(core__abc_21380_n3535_1), .B(core__abc_21380_n1931), .Y(core__abc_21380_n3536) );
  AND2X2 AND2X2_2559 ( .A(core__abc_21380_n3017), .B(core__abc_21380_n1345), .Y(core__abc_21380_n3540) );
  AND2X2 AND2X2_256 ( .A(_abc_19068_n902_bF_buf0), .B(word2_reg_18_), .Y(_abc_19068_n1336_1) );
  AND2X2 AND2X2_2560 ( .A(core__abc_21380_n3541), .B(core__abc_21380_n1344), .Y(core__abc_21380_n3542) );
  AND2X2 AND2X2_2561 ( .A(core__abc_21380_n3543), .B(core__abc_21380_n3539), .Y(core__abc_21380_n3544) );
  AND2X2 AND2X2_2562 ( .A(core__abc_21380_n3545), .B(core_v3_reg_52_), .Y(core__abc_21380_n3546) );
  AND2X2 AND2X2_2563 ( .A(core__abc_21380_n3538), .B(core__abc_21380_n3548_1), .Y(core__abc_21380_n3549) );
  AND2X2 AND2X2_2564 ( .A(core__abc_21380_n3537), .B(core__abc_21380_n3547), .Y(core__abc_21380_n3550) );
  AND2X2 AND2X2_2565 ( .A(core__abc_21380_n3476), .B(core__abc_21380_n3482), .Y(core__abc_21380_n3553) );
  AND2X2 AND2X2_2566 ( .A(core__abc_21380_n3555), .B(core__abc_21380_n3479), .Y(core__abc_21380_n3556) );
  AND2X2 AND2X2_2567 ( .A(core__abc_21380_n3556), .B(core__abc_21380_n3552_1), .Y(core__abc_21380_n3557) );
  AND2X2 AND2X2_2568 ( .A(core__abc_21380_n3483_1), .B(core__abc_21380_n3553), .Y(core__abc_21380_n3559) );
  AND2X2 AND2X2_2569 ( .A(core__abc_21380_n3560), .B(core__abc_21380_n3551), .Y(core__abc_21380_n3561_1) );
  AND2X2 AND2X2_257 ( .A(_abc_19068_n916_1_bF_buf0), .B(word1_reg_18_), .Y(_abc_19068_n1337) );
  AND2X2 AND2X2_2570 ( .A(core__abc_21380_n3564), .B(core__abc_21380_n2122), .Y(core__abc_21380_n3565) );
  AND2X2 AND2X2_2571 ( .A(core__abc_21380_n3565), .B(core__abc_21380_n2146), .Y(core__abc_21380_n3566) );
  AND2X2 AND2X2_2572 ( .A(core__abc_21380_n3567), .B(core__abc_21380_n2144), .Y(core__abc_21380_n3568) );
  AND2X2 AND2X2_2573 ( .A(core__abc_21380_n3569_1), .B(core_v3_reg_31_), .Y(core__abc_21380_n3570) );
  AND2X2 AND2X2_2574 ( .A(core__abc_21380_n3572), .B(core__abc_21380_n3573), .Y(core__abc_21380_n3574) );
  AND2X2 AND2X2_2575 ( .A(core__abc_21380_n3574), .B(core__abc_21380_n3571), .Y(core__abc_21380_n3575) );
  AND2X2 AND2X2_2576 ( .A(core__abc_21380_n3579), .B(core__abc_21380_n3578), .Y(core__abc_21380_n3580) );
  AND2X2 AND2X2_2577 ( .A(core__abc_21380_n3581_1), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n3582) );
  AND2X2 AND2X2_2578 ( .A(core__abc_21380_n3582), .B(core__abc_21380_n3577), .Y(core__abc_21380_n3583) );
  AND2X2 AND2X2_2579 ( .A(core__abc_21380_n3313_bF_buf7), .B(core__abc_21380_n3584), .Y(core__abc_21380_n3585) );
  AND2X2 AND2X2_258 ( .A(_abc_19068_n941_bF_buf1), .B(core_key_114_), .Y(_abc_19068_n1340_1) );
  AND2X2 AND2X2_2580 ( .A(core_v3_reg_4_), .B(core_mi_4_), .Y(core__abc_21380_n3587) );
  AND2X2 AND2X2_2581 ( .A(core__abc_21380_n3588), .B(core__abc_21380_n3586), .Y(core__abc_21380_n3589_1) );
  AND2X2 AND2X2_2582 ( .A(core__abc_21380_n2749_bF_buf7), .B(core__abc_21380_n3589_1), .Y(core__abc_21380_n3590) );
  AND2X2 AND2X2_2583 ( .A(core__abc_21380_n3594), .B(reset_n_bF_buf60), .Y(core__abc_21380_n3595) );
  AND2X2 AND2X2_2584 ( .A(core__abc_21380_n3593), .B(core__abc_21380_n3595), .Y(core_v3_reg_4__FF_INPUT) );
  AND2X2 AND2X2_2585 ( .A(core__abc_21380_n3600_1), .B(core__abc_21380_n1958), .Y(core__abc_21380_n3601) );
  AND2X2 AND2X2_2586 ( .A(core__abc_21380_n3599), .B(core__abc_21380_n1951), .Y(core__abc_21380_n3602) );
  AND2X2 AND2X2_2587 ( .A(core__abc_21380_n3607), .B(core__abc_21380_n1364), .Y(core__abc_21380_n3608) );
  AND2X2 AND2X2_2588 ( .A(core__abc_21380_n3606), .B(core__abc_21380_n1366), .Y(core__abc_21380_n3609) );
  AND2X2 AND2X2_2589 ( .A(core__abc_21380_n3610), .B(core__abc_21380_n3605), .Y(core__abc_21380_n3611) );
  AND2X2 AND2X2_259 ( .A(_abc_19068_n945_1_bF_buf1), .B(core_mi_18_), .Y(_abc_19068_n1341) );
  AND2X2 AND2X2_2590 ( .A(core__abc_21380_n3612), .B(core_v3_reg_53_), .Y(core__abc_21380_n3613) );
  AND2X2 AND2X2_2591 ( .A(core__abc_21380_n3604_1), .B(core__abc_21380_n3615), .Y(core__abc_21380_n3616) );
  AND2X2 AND2X2_2592 ( .A(core__abc_21380_n3603), .B(core__abc_21380_n3614), .Y(core__abc_21380_n3617) );
  AND2X2 AND2X2_2593 ( .A(core__abc_21380_n3598), .B(core__abc_21380_n3618), .Y(core__abc_21380_n3619_1) );
  AND2X2 AND2X2_2594 ( .A(core__abc_21380_n3597), .B(core__abc_21380_n3620), .Y(core__abc_21380_n3621) );
  AND2X2 AND2X2_2595 ( .A(core__abc_21380_n2123), .B(core__abc_21380_n2144), .Y(core__abc_21380_n3625) );
  AND2X2 AND2X2_2596 ( .A(core__abc_21380_n3490_1), .B(core__abc_21380_n3625), .Y(core__abc_21380_n3626) );
  AND2X2 AND2X2_2597 ( .A(core__abc_21380_n3370), .B(core__abc_21380_n3626), .Y(core__abc_21380_n3627) );
  AND2X2 AND2X2_2598 ( .A(core__abc_21380_n3628), .B(core__abc_21380_n3625), .Y(core__abc_21380_n3629) );
  AND2X2 AND2X2_2599 ( .A(core__abc_21380_n2141), .B(core__abc_21380_n2121), .Y(core__abc_21380_n3630) );
  AND2X2 AND2X2_26 ( .A(_abc_19068_n908), .B(_abc_19068_n881), .Y(_abc_19068_n909_1) );
  AND2X2 AND2X2_260 ( .A(_abc_19068_n915_1_bF_buf0), .B(core_mi_50_), .Y(_abc_19068_n1343) );
  AND2X2 AND2X2_2600 ( .A(core__abc_21380_n3144), .B(core__abc_21380_n3372), .Y(core__abc_21380_n3634) );
  AND2X2 AND2X2_2601 ( .A(core__abc_21380_n3634), .B(core__abc_21380_n3626), .Y(core__abc_21380_n3635) );
  AND2X2 AND2X2_2602 ( .A(core__abc_21380_n3636_1), .B(core__abc_21380_n2162), .Y(core__abc_21380_n3637) );
  AND2X2 AND2X2_2603 ( .A(core__abc_21380_n3640), .B(core__abc_21380_n3638), .Y(core__abc_21380_n3641) );
  AND2X2 AND2X2_2604 ( .A(core__abc_21380_n3641), .B(core__abc_21380_n2164), .Y(core__abc_21380_n3642) );
  AND2X2 AND2X2_2605 ( .A(core__abc_21380_n3645), .B(core__abc_21380_n3646), .Y(core__abc_21380_n3647_1) );
  AND2X2 AND2X2_2606 ( .A(core__abc_21380_n3650), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n3651_1) );
  AND2X2 AND2X2_2607 ( .A(core__abc_21380_n3651_1), .B(core__abc_21380_n3649), .Y(core__abc_21380_n3652) );
  AND2X2 AND2X2_2608 ( .A(core__abc_21380_n3313_bF_buf6), .B(core__abc_21380_n3653), .Y(core__abc_21380_n3654) );
  AND2X2 AND2X2_2609 ( .A(core_v3_reg_5_), .B(core_mi_5_), .Y(core__abc_21380_n3656) );
  AND2X2 AND2X2_261 ( .A(_abc_19068_n897_1_bF_buf0), .B(word0_reg_18_), .Y(_abc_19068_n1344_1) );
  AND2X2 AND2X2_2610 ( .A(core__abc_21380_n3657), .B(core__abc_21380_n3655), .Y(core__abc_21380_n3658) );
  AND2X2 AND2X2_2611 ( .A(core__abc_21380_n2749_bF_buf6), .B(core__abc_21380_n3658), .Y(core__abc_21380_n3659_1) );
  AND2X2 AND2X2_2612 ( .A(core__abc_21380_n3663_1), .B(reset_n_bF_buf59), .Y(core__abc_21380_n3664) );
  AND2X2 AND2X2_2613 ( .A(core__abc_21380_n3662), .B(core__abc_21380_n3664), .Y(core_v3_reg_5__FF_INPUT) );
  AND2X2 AND2X2_2614 ( .A(core__abc_21380_n3669), .B(core__abc_21380_n3668), .Y(core__abc_21380_n3670) );
  AND2X2 AND2X2_2615 ( .A(core__abc_21380_n3667), .B(core__abc_21380_n3671), .Y(core__abc_21380_n3672) );
  AND2X2 AND2X2_2616 ( .A(core__abc_21380_n1937), .B(core__abc_21380_n1951), .Y(core__abc_21380_n3674) );
  AND2X2 AND2X2_2617 ( .A(core__abc_21380_n3677), .B(core__abc_21380_n1946), .Y(core__abc_21380_n3678) );
  AND2X2 AND2X2_2618 ( .A(core__abc_21380_n3676_1), .B(core__abc_21380_n3679), .Y(core__abc_21380_n3680) );
  AND2X2 AND2X2_2619 ( .A(core__abc_21380_n3680), .B(core__abc_21380_n1969), .Y(core__abc_21380_n3681_1) );
  AND2X2 AND2X2_262 ( .A(_abc_19068_n923_bF_buf1), .B(_abc_19068_n1348_1), .Y(_auto_iopadmap_cc_313_execute_30317_18_) );
  AND2X2 AND2X2_2620 ( .A(core__abc_21380_n3530), .B(core__abc_21380_n3674), .Y(core__abc_21380_n3682) );
  AND2X2 AND2X2_2621 ( .A(core__abc_21380_n3684), .B(core__abc_21380_n1970), .Y(core__abc_21380_n3685) );
  AND2X2 AND2X2_2622 ( .A(core__abc_21380_n3688_1), .B(core__abc_21380_n3026), .Y(core__abc_21380_n3689) );
  AND2X2 AND2X2_2623 ( .A(core__abc_21380_n3689), .B(core__abc_21380_n1383), .Y(core__abc_21380_n3690) );
  AND2X2 AND2X2_2624 ( .A(core__abc_21380_n3695), .B(core__abc_21380_n3696), .Y(core__abc_21380_n3697) );
  AND2X2 AND2X2_2625 ( .A(core__abc_21380_n3686), .B(core__abc_21380_n3697), .Y(core__abc_21380_n3700) );
  AND2X2 AND2X2_2626 ( .A(core__abc_21380_n3673), .B(core__abc_21380_n3702), .Y(core__abc_21380_n3703_1) );
  AND2X2 AND2X2_2627 ( .A(core__abc_21380_n3672), .B(core__abc_21380_n3701), .Y(core__abc_21380_n3704) );
  AND2X2 AND2X2_2628 ( .A(core__abc_21380_n2182), .B(core__abc_21380_n2161), .Y(core__abc_21380_n3709) );
  AND2X2 AND2X2_2629 ( .A(core__abc_21380_n3708_1), .B(core__abc_21380_n3709), .Y(core__abc_21380_n3710) );
  AND2X2 AND2X2_263 ( .A(_abc_19068_n899_bF_buf4), .B(word3_reg_19_), .Y(_abc_19068_n1350_1) );
  AND2X2 AND2X2_2630 ( .A(core__abc_21380_n2179_1), .B(core__abc_21380_n2160), .Y(core__abc_21380_n3711) );
  AND2X2 AND2X2_2631 ( .A(core__abc_21380_n2162), .B(core__abc_21380_n2179_1), .Y(core__abc_21380_n3712) );
  AND2X2 AND2X2_2632 ( .A(core__abc_21380_n3636_1), .B(core__abc_21380_n3712), .Y(core__abc_21380_n3713) );
  AND2X2 AND2X2_2633 ( .A(core__abc_21380_n3715), .B(core__abc_21380_n3707), .Y(core__abc_21380_n3716_1) );
  AND2X2 AND2X2_2634 ( .A(core__abc_21380_n3717), .B(core_v3_reg_33_), .Y(core__abc_21380_n3718) );
  AND2X2 AND2X2_2635 ( .A(core__abc_21380_n3722), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n3723) );
  AND2X2 AND2X2_2636 ( .A(core__abc_21380_n3723), .B(core__abc_21380_n3721), .Y(core__abc_21380_n3724) );
  AND2X2 AND2X2_2637 ( .A(core__abc_21380_n3313_bF_buf5), .B(core__abc_21380_n3725), .Y(core__abc_21380_n3726) );
  AND2X2 AND2X2_2638 ( .A(core_v3_reg_6_), .B(core_mi_6_), .Y(core__abc_21380_n3728) );
  AND2X2 AND2X2_2639 ( .A(core__abc_21380_n3729), .B(core__abc_21380_n3727), .Y(core__abc_21380_n3730) );
  AND2X2 AND2X2_264 ( .A(_abc_19068_n945_1_bF_buf0), .B(core_mi_19_), .Y(_abc_19068_n1352_1) );
  AND2X2 AND2X2_2640 ( .A(core__abc_21380_n2749_bF_buf5), .B(core__abc_21380_n3730), .Y(core__abc_21380_n3731) );
  AND2X2 AND2X2_2641 ( .A(core__abc_21380_n3735), .B(reset_n_bF_buf58), .Y(core__abc_21380_n3736) );
  AND2X2 AND2X2_2642 ( .A(core__abc_21380_n3734), .B(core__abc_21380_n3736), .Y(core_v3_reg_6__FF_INPUT) );
  AND2X2 AND2X2_2643 ( .A(core__abc_21380_n3741), .B(core__abc_21380_n3740_1), .Y(core__abc_21380_n3742) );
  AND2X2 AND2X2_2644 ( .A(core__abc_21380_n3742), .B(core__abc_21380_n1995_1), .Y(core__abc_21380_n3743) );
  AND2X2 AND2X2_2645 ( .A(core__abc_21380_n3744), .B(core__abc_21380_n1989), .Y(core__abc_21380_n3745_1) );
  AND2X2 AND2X2_2646 ( .A(core__abc_21380_n3749), .B(core__abc_21380_n1402), .Y(core__abc_21380_n3750) );
  AND2X2 AND2X2_2647 ( .A(core__abc_21380_n3748), .B(core__abc_21380_n1403), .Y(core__abc_21380_n3751) );
  AND2X2 AND2X2_2648 ( .A(core__abc_21380_n3752_1), .B(core__abc_21380_n3747), .Y(core__abc_21380_n3753) );
  AND2X2 AND2X2_2649 ( .A(core__abc_21380_n3754), .B(core_v3_reg_55_), .Y(core__abc_21380_n3755) );
  AND2X2 AND2X2_265 ( .A(_abc_19068_n941_bF_buf0), .B(core_key_115_), .Y(_abc_19068_n1353) );
  AND2X2 AND2X2_2650 ( .A(core__abc_21380_n3759), .B(core__abc_21380_n3758), .Y(core__abc_21380_n3760) );
  AND2X2 AND2X2_2651 ( .A(core__abc_21380_n3757), .B(core__abc_21380_n3762), .Y(core__abc_21380_n3763) );
  AND2X2 AND2X2_2652 ( .A(core__abc_21380_n3739), .B(core__abc_21380_n3764), .Y(core__abc_21380_n3765) );
  AND2X2 AND2X2_2653 ( .A(core__abc_21380_n3738), .B(core__abc_21380_n3763), .Y(core__abc_21380_n3766) );
  AND2X2 AND2X2_2654 ( .A(core__abc_21380_n3771), .B(core__abc_21380_n2197), .Y(core__abc_21380_n3772_1) );
  AND2X2 AND2X2_2655 ( .A(core__abc_21380_n3773), .B(core__abc_21380_n3774), .Y(core__abc_21380_n3775) );
  AND2X2 AND2X2_2656 ( .A(core__abc_21380_n3778), .B(core__abc_21380_n3776), .Y(core__abc_21380_n3779_1) );
  AND2X2 AND2X2_2657 ( .A(core__abc_21380_n3782), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n3783_1) );
  AND2X2 AND2X2_2658 ( .A(core__abc_21380_n3783_1), .B(core__abc_21380_n3781), .Y(core__abc_21380_n3784) );
  AND2X2 AND2X2_2659 ( .A(core__abc_21380_n3313_bF_buf4), .B(core_key_71_), .Y(core__abc_21380_n3785) );
  AND2X2 AND2X2_266 ( .A(_abc_19068_n939_1_bF_buf0), .B(core_key_83_), .Y(_abc_19068_n1356_1) );
  AND2X2 AND2X2_2660 ( .A(core_v3_reg_7_), .B(core_mi_7_), .Y(core__abc_21380_n3787) );
  AND2X2 AND2X2_2661 ( .A(core__abc_21380_n3788), .B(core__abc_21380_n3786), .Y(core__abc_21380_n3789) );
  AND2X2 AND2X2_2662 ( .A(core__abc_21380_n2749_bF_buf4), .B(core__abc_21380_n3789), .Y(core__abc_21380_n3790) );
  AND2X2 AND2X2_2663 ( .A(core__abc_21380_n3794), .B(reset_n_bF_buf57), .Y(core__abc_21380_n3795) );
  AND2X2 AND2X2_2664 ( .A(core__abc_21380_n3793), .B(core__abc_21380_n3795), .Y(core_v3_reg_7__FF_INPUT) );
  AND2X2 AND2X2_2665 ( .A(core__abc_21380_n1970), .B(core__abc_21380_n1989), .Y(core__abc_21380_n3797_1) );
  AND2X2 AND2X2_2666 ( .A(core__abc_21380_n3674), .B(core__abc_21380_n3797_1), .Y(core__abc_21380_n3798) );
  AND2X2 AND2X2_2667 ( .A(core__abc_21380_n3527), .B(core__abc_21380_n3798), .Y(core__abc_21380_n3799) );
  AND2X2 AND2X2_2668 ( .A(core__abc_21380_n3683), .B(core__abc_21380_n3797_1), .Y(core__abc_21380_n3800) );
  AND2X2 AND2X2_2669 ( .A(core__abc_21380_n1986), .B(core__abc_21380_n1968), .Y(core__abc_21380_n3801_1) );
  AND2X2 AND2X2_267 ( .A(_abc_19068_n924_1_bF_buf0), .B(core_key_51_), .Y(_abc_19068_n1357) );
  AND2X2 AND2X2_2670 ( .A(core__abc_21380_n3528), .B(core__abc_21380_n3798), .Y(core__abc_21380_n3805) );
  AND2X2 AND2X2_2671 ( .A(core__abc_21380_n3269), .B(core__abc_21380_n3805), .Y(core__abc_21380_n3806) );
  AND2X2 AND2X2_2672 ( .A(core__abc_21380_n3807), .B(core__abc_21380_n2008), .Y(core__abc_21380_n3808) );
  AND2X2 AND2X2_2673 ( .A(core__abc_21380_n3811), .B(core__abc_21380_n3809_1), .Y(core__abc_21380_n3812) );
  AND2X2 AND2X2_2674 ( .A(core__abc_21380_n3812), .B(core__abc_21380_n2007), .Y(core__abc_21380_n3813) );
  AND2X2 AND2X2_2675 ( .A(core__abc_21380_n3032), .B(core__abc_21380_n1419), .Y(core__abc_21380_n3817) );
  AND2X2 AND2X2_2676 ( .A(core__abc_21380_n3818), .B(core__abc_21380_n1418), .Y(core__abc_21380_n3819) );
  AND2X2 AND2X2_2677 ( .A(core__abc_21380_n3822), .B(core__abc_21380_n3823_1), .Y(core__abc_21380_n3824) );
  AND2X2 AND2X2_2678 ( .A(core__abc_21380_n3815), .B(core__abc_21380_n3825), .Y(core__abc_21380_n3826) );
  AND2X2 AND2X2_2679 ( .A(core__abc_21380_n3814_1), .B(core__abc_21380_n3824), .Y(core__abc_21380_n3827) );
  AND2X2 AND2X2_268 ( .A(_abc_19068_n926_bF_buf0), .B(core_key_19_), .Y(_abc_19068_n1358_1) );
  AND2X2 AND2X2_2680 ( .A(core__abc_21380_n3746), .B(core__abc_21380_n3756_1), .Y(core__abc_21380_n3829) );
  AND2X2 AND2X2_2681 ( .A(core__abc_21380_n3830), .B(core__abc_21380_n3757), .Y(core__abc_21380_n3831) );
  AND2X2 AND2X2_2682 ( .A(core__abc_21380_n3831), .B(core__abc_21380_n3671), .Y(core__abc_21380_n3832) );
  AND2X2 AND2X2_2683 ( .A(core__abc_21380_n3667), .B(core__abc_21380_n3832), .Y(core__abc_21380_n3833) );
  AND2X2 AND2X2_2684 ( .A(core__abc_21380_n3757), .B(core__abc_21380_n3700), .Y(core__abc_21380_n3834_1) );
  AND2X2 AND2X2_2685 ( .A(core__abc_21380_n3836), .B(core__abc_21380_n3828_1), .Y(core__abc_21380_n3837) );
  AND2X2 AND2X2_2686 ( .A(core__abc_21380_n3763), .B(core__abc_21380_n3702), .Y(core__abc_21380_n3840) );
  AND2X2 AND2X2_2687 ( .A(core__abc_21380_n3840), .B(core__abc_21380_n3670), .Y(core__abc_21380_n3841) );
  AND2X2 AND2X2_2688 ( .A(core__abc_21380_n3556), .B(core__abc_21380_n3843), .Y(core__abc_21380_n3844) );
  AND2X2 AND2X2_2689 ( .A(core__abc_21380_n3844), .B(core__abc_21380_n3840), .Y(core__abc_21380_n3845) );
  AND2X2 AND2X2_269 ( .A(_abc_19068_n916_1_bF_buf4), .B(word1_reg_19_), .Y(_abc_19068_n1361) );
  AND2X2 AND2X2_2690 ( .A(core__abc_21380_n3846), .B(core__abc_21380_n3838_1), .Y(core__abc_21380_n3847) );
  AND2X2 AND2X2_2691 ( .A(core__abc_21380_n3773), .B(core__abc_21380_n2196), .Y(core__abc_21380_n3851) );
  AND2X2 AND2X2_2692 ( .A(core__abc_21380_n3851), .B(core__abc_21380_n2220), .Y(core__abc_21380_n3852) );
  AND2X2 AND2X2_2693 ( .A(core__abc_21380_n3853_1), .B(core__abc_21380_n3854), .Y(core__abc_21380_n3855) );
  AND2X2 AND2X2_2694 ( .A(core__abc_21380_n3855), .B(core__abc_21380_n3850), .Y(core__abc_21380_n3858) );
  AND2X2 AND2X2_2695 ( .A(core__abc_21380_n3861), .B(core__abc_21380_n3856), .Y(core__abc_21380_n3862) );
  AND2X2 AND2X2_2696 ( .A(core__abc_21380_n3863), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n3864_1) );
  AND2X2 AND2X2_2697 ( .A(core__abc_21380_n3864_1), .B(core__abc_21380_n3860), .Y(core__abc_21380_n3865) );
  AND2X2 AND2X2_2698 ( .A(core__abc_21380_n3313_bF_buf3), .B(core__abc_21380_n3866), .Y(core__abc_21380_n3867) );
  AND2X2 AND2X2_2699 ( .A(core_v3_reg_8_), .B(core_mi_8_), .Y(core__abc_21380_n3869_1) );
  AND2X2 AND2X2_27 ( .A(_abc_19068_n879_1), .B(\addr[4] ), .Y(_abc_19068_n911) );
  AND2X2 AND2X2_270 ( .A(_abc_19068_n902_bF_buf4), .B(word2_reg_19_), .Y(_abc_19068_n1362) );
  AND2X2 AND2X2_2700 ( .A(core__abc_21380_n3870), .B(core__abc_21380_n3868), .Y(core__abc_21380_n3871) );
  AND2X2 AND2X2_2701 ( .A(core__abc_21380_n2749_bF_buf3), .B(core__abc_21380_n3871), .Y(core__abc_21380_n3872) );
  AND2X2 AND2X2_2702 ( .A(core__abc_21380_n3876), .B(reset_n_bF_buf56), .Y(core__abc_21380_n3877) );
  AND2X2 AND2X2_2703 ( .A(core__abc_21380_n3875), .B(core__abc_21380_n3877), .Y(core_v3_reg_8__FF_INPUT) );
  AND2X2 AND2X2_2704 ( .A(core__abc_21380_n3880), .B(core__abc_21380_n3879), .Y(core__abc_21380_n3881_1) );
  AND2X2 AND2X2_2705 ( .A(core__abc_21380_n2031), .B(core__abc_21380_n2003), .Y(core__abc_21380_n3883) );
  AND2X2 AND2X2_2706 ( .A(core__abc_21380_n3885), .B(core__abc_21380_n2025), .Y(core__abc_21380_n3886_1) );
  AND2X2 AND2X2_2707 ( .A(core__abc_21380_n2008), .B(core__abc_21380_n2031), .Y(core__abc_21380_n3887) );
  AND2X2 AND2X2_2708 ( .A(core__abc_21380_n3807), .B(core__abc_21380_n3887), .Y(core__abc_21380_n3888) );
  AND2X2 AND2X2_2709 ( .A(core__abc_21380_n3893_1), .B(core__abc_21380_n1439), .Y(core__abc_21380_n3894) );
  AND2X2 AND2X2_271 ( .A(_abc_19068_n897_1_bF_buf4), .B(word0_reg_19_), .Y(_abc_19068_n1364) );
  AND2X2 AND2X2_2710 ( .A(core__abc_21380_n3892), .B(core__abc_21380_n1438), .Y(core__abc_21380_n3895) );
  AND2X2 AND2X2_2711 ( .A(core__abc_21380_n3896), .B(core__abc_21380_n3891), .Y(core__abc_21380_n3897) );
  AND2X2 AND2X2_2712 ( .A(core__abc_21380_n3898_1), .B(core_v3_reg_57_), .Y(core__abc_21380_n3899) );
  AND2X2 AND2X2_2713 ( .A(core__abc_21380_n3890), .B(core__abc_21380_n3900), .Y(core__abc_21380_n3902) );
  AND2X2 AND2X2_2714 ( .A(core__abc_21380_n3903), .B(core__abc_21380_n3901), .Y(core__abc_21380_n3904) );
  AND2X2 AND2X2_2715 ( .A(core__abc_21380_n3882), .B(core__abc_21380_n3905), .Y(core__abc_21380_n3906) );
  AND2X2 AND2X2_2716 ( .A(core__abc_21380_n3881_1), .B(core__abc_21380_n3904), .Y(core__abc_21380_n3907) );
  AND2X2 AND2X2_2717 ( .A(core__abc_21380_n2197), .B(core__abc_21380_n2218), .Y(core__abc_21380_n3910_1) );
  AND2X2 AND2X2_2718 ( .A(core__abc_21380_n3712), .B(core__abc_21380_n3910_1), .Y(core__abc_21380_n3911) );
  AND2X2 AND2X2_2719 ( .A(core__abc_21380_n3770), .B(core__abc_21380_n3910_1), .Y(core__abc_21380_n3914_1) );
  AND2X2 AND2X2_272 ( .A(_abc_19068_n915_1_bF_buf4), .B(core_mi_51_), .Y(_abc_19068_n1365_1) );
  AND2X2 AND2X2_2720 ( .A(core__abc_21380_n2215), .B(core__abc_21380_n2195), .Y(core__abc_21380_n3915) );
  AND2X2 AND2X2_2721 ( .A(core__abc_21380_n3913), .B(core__abc_21380_n3918), .Y(core__abc_21380_n3919) );
  AND2X2 AND2X2_2722 ( .A(core__abc_21380_n3920), .B(core__abc_21380_n2234), .Y(core__abc_21380_n3921) );
  AND2X2 AND2X2_2723 ( .A(core__abc_21380_n3919), .B(core__abc_21380_n2237), .Y(core__abc_21380_n3922_1) );
  AND2X2 AND2X2_2724 ( .A(core__abc_21380_n3925), .B(core__abc_21380_n3926), .Y(core__abc_21380_n3927_1) );
  AND2X2 AND2X2_2725 ( .A(core__abc_21380_n3931), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n3932) );
  AND2X2 AND2X2_2726 ( .A(core__abc_21380_n3932), .B(core__abc_21380_n3929), .Y(core__abc_21380_n3933) );
  AND2X2 AND2X2_2727 ( .A(core__abc_21380_n3313_bF_buf2), .B(core_key_73_), .Y(core__abc_21380_n3934) );
  AND2X2 AND2X2_2728 ( .A(core_v3_reg_9_), .B(core_mi_9_), .Y(core__abc_21380_n3936) );
  AND2X2 AND2X2_2729 ( .A(core__abc_21380_n3937_1), .B(core__abc_21380_n3935), .Y(core__abc_21380_n3938) );
  AND2X2 AND2X2_273 ( .A(_abc_19068_n923_bF_buf0), .B(_abc_19068_n1369_1), .Y(_auto_iopadmap_cc_313_execute_30317_19_) );
  AND2X2 AND2X2_2730 ( .A(core__abc_21380_n2749_bF_buf2), .B(core__abc_21380_n3938), .Y(core__abc_21380_n3939) );
  AND2X2 AND2X2_2731 ( .A(core__abc_21380_n3943), .B(reset_n_bF_buf55), .Y(core__abc_21380_n3944) );
  AND2X2 AND2X2_2732 ( .A(core__abc_21380_n3942_1), .B(core__abc_21380_n3944), .Y(core_v3_reg_9__FF_INPUT) );
  AND2X2 AND2X2_2733 ( .A(core__abc_21380_n3947), .B(core__abc_21380_n2044), .Y(core__abc_21380_n3948_1) );
  AND2X2 AND2X2_2734 ( .A(core__abc_21380_n3949), .B(core__abc_21380_n2043), .Y(core__abc_21380_n3950) );
  AND2X2 AND2X2_2735 ( .A(core__abc_21380_n3818), .B(core__abc_21380_n3036), .Y(core__abc_21380_n3954) );
  AND2X2 AND2X2_2736 ( .A(core__abc_21380_n3955_1), .B(core__abc_21380_n3044_1), .Y(core__abc_21380_n3956) );
  AND2X2 AND2X2_2737 ( .A(core__abc_21380_n3956), .B(core__abc_21380_n1458), .Y(core__abc_21380_n3957) );
  AND2X2 AND2X2_2738 ( .A(core__abc_21380_n3962), .B(core__abc_21380_n3963), .Y(core__abc_21380_n3964) );
  AND2X2 AND2X2_2739 ( .A(core__abc_21380_n3952_1), .B(core__abc_21380_n3965_1), .Y(core__abc_21380_n3966) );
  AND2X2 AND2X2_274 ( .A(_abc_19068_n939_1_bF_buf4), .B(core_key_84_), .Y(_abc_19068_n1371_1) );
  AND2X2 AND2X2_2740 ( .A(core__abc_21380_n3951), .B(core__abc_21380_n3964), .Y(core__abc_21380_n3967) );
  AND2X2 AND2X2_2741 ( .A(core__abc_21380_n3901), .B(core__abc_21380_n3879), .Y(core__abc_21380_n3970) );
  AND2X2 AND2X2_2742 ( .A(core__abc_21380_n3880), .B(core__abc_21380_n3970), .Y(core__abc_21380_n3971) );
  AND2X2 AND2X2_2743 ( .A(core__abc_21380_n3973), .B(core__abc_21380_n3969_1), .Y(core__abc_21380_n3974_1) );
  AND2X2 AND2X2_2744 ( .A(core__abc_21380_n3972), .B(core__abc_21380_n3968), .Y(core__abc_21380_n3975) );
  AND2X2 AND2X2_2745 ( .A(core__abc_21380_n3980), .B(core__abc_21380_n2257), .Y(core__abc_21380_n3981) );
  AND2X2 AND2X2_2746 ( .A(core__abc_21380_n3979_1), .B(core__abc_21380_n2255), .Y(core__abc_21380_n3982_1) );
  AND2X2 AND2X2_2747 ( .A(core__abc_21380_n3983), .B(core__abc_21380_n3978), .Y(core__abc_21380_n3984) );
  AND2X2 AND2X2_2748 ( .A(core__abc_21380_n3985), .B(core_v3_reg_37_), .Y(core__abc_21380_n3986_1) );
  AND2X2 AND2X2_2749 ( .A(core__abc_21380_n3990), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n3991) );
  AND2X2 AND2X2_275 ( .A(_abc_19068_n926_bF_buf4), .B(core_key_20_), .Y(_abc_19068_n1372) );
  AND2X2 AND2X2_2750 ( .A(core__abc_21380_n3991), .B(core__abc_21380_n3989), .Y(core__abc_21380_n3992_1) );
  AND2X2 AND2X2_2751 ( .A(core__abc_21380_n3313_bF_buf1), .B(core__abc_21380_n3993), .Y(core__abc_21380_n3994) );
  AND2X2 AND2X2_2752 ( .A(core_v3_reg_10_), .B(core_mi_10_), .Y(core__abc_21380_n3996) );
  AND2X2 AND2X2_2753 ( .A(core__abc_21380_n3997), .B(core__abc_21380_n3995_1), .Y(core__abc_21380_n3998) );
  AND2X2 AND2X2_2754 ( .A(core__abc_21380_n2749_bF_buf1), .B(core__abc_21380_n3998), .Y(core__abc_21380_n3999) );
  AND2X2 AND2X2_2755 ( .A(core__abc_21380_n4003_1), .B(reset_n_bF_buf54), .Y(core__abc_21380_n4004) );
  AND2X2 AND2X2_2756 ( .A(core__abc_21380_n4002), .B(core__abc_21380_n4004), .Y(core_v3_reg_10__FF_INPUT) );
  AND2X2 AND2X2_2757 ( .A(core__abc_21380_n4008_1), .B(core__abc_21380_n2069), .Y(core__abc_21380_n4009) );
  AND2X2 AND2X2_2758 ( .A(core__abc_21380_n4007), .B(core__abc_21380_n2063), .Y(core__abc_21380_n4010) );
  AND2X2 AND2X2_2759 ( .A(core__abc_21380_n3958), .B(core__abc_21380_n1453), .Y(core__abc_21380_n4013) );
  AND2X2 AND2X2_276 ( .A(_abc_19068_n924_1_bF_buf4), .B(core_key_52_), .Y(_abc_19068_n1373_1) );
  AND2X2 AND2X2_2760 ( .A(core__abc_21380_n4013), .B(core__abc_21380_n1475), .Y(core__abc_21380_n4014) );
  AND2X2 AND2X2_2761 ( .A(core__abc_21380_n4015), .B(core__abc_21380_n4016_1), .Y(core__abc_21380_n4017) );
  AND2X2 AND2X2_2762 ( .A(core__abc_21380_n4018_1), .B(core__abc_21380_n4012_1), .Y(core__abc_21380_n4019) );
  AND2X2 AND2X2_2763 ( .A(core__abc_21380_n4017), .B(core_v3_reg_59_), .Y(core__abc_21380_n4020) );
  AND2X2 AND2X2_2764 ( .A(core__abc_21380_n4011), .B(core__abc_21380_n4021), .Y(core__abc_21380_n4023_1) );
  AND2X2 AND2X2_2765 ( .A(core__abc_21380_n4024), .B(core__abc_21380_n4022), .Y(core__abc_21380_n4025) );
  AND2X2 AND2X2_2766 ( .A(core__abc_21380_n4006), .B(core__abc_21380_n4025), .Y(core__abc_21380_n4026_1) );
  AND2X2 AND2X2_2767 ( .A(core__abc_21380_n4027), .B(core__abc_21380_n4028), .Y(core__abc_21380_n4029) );
  AND2X2 AND2X2_2768 ( .A(core__abc_21380_n2234), .B(core__abc_21380_n2255), .Y(core__abc_21380_n4031_1) );
  AND2X2 AND2X2_2769 ( .A(core__abc_21380_n2233), .B(core__abc_21380_n2254), .Y(core__abc_21380_n4035) );
  AND2X2 AND2X2_277 ( .A(_abc_19068_n899_bF_buf3), .B(word3_reg_20_), .Y(_abc_19068_n1376) );
  AND2X2 AND2X2_2770 ( .A(core__abc_21380_n4033), .B(core__abc_21380_n4036), .Y(core__abc_21380_n4037) );
  AND2X2 AND2X2_2771 ( .A(core__abc_21380_n4038), .B(core__abc_21380_n2273), .Y(core__abc_21380_n4039_1) );
  AND2X2 AND2X2_2772 ( .A(core__abc_21380_n4037), .B(core__abc_21380_n2275), .Y(core__abc_21380_n4040) );
  AND2X2 AND2X2_2773 ( .A(core__abc_21380_n4043_1), .B(core__abc_21380_n4045), .Y(core__abc_21380_n4046) );
  AND2X2 AND2X2_2774 ( .A(core__abc_21380_n4049), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n4050_1) );
  AND2X2 AND2X2_2775 ( .A(core__abc_21380_n4050_1), .B(core__abc_21380_n4048), .Y(core__abc_21380_n4051) );
  AND2X2 AND2X2_2776 ( .A(core__abc_21380_n3313_bF_buf0), .B(core_key_75_), .Y(core__abc_21380_n4052) );
  AND2X2 AND2X2_2777 ( .A(core_v3_reg_11_), .B(core_mi_11_), .Y(core__abc_21380_n4054_1) );
  AND2X2 AND2X2_2778 ( .A(core__abc_21380_n4055), .B(core__abc_21380_n4053), .Y(core__abc_21380_n4056) );
  AND2X2 AND2X2_2779 ( .A(core__abc_21380_n2749_bF_buf0), .B(core__abc_21380_n4056), .Y(core__abc_21380_n4057_1) );
  AND2X2 AND2X2_278 ( .A(_abc_19068_n902_bF_buf3), .B(word2_reg_20_), .Y(_abc_19068_n1378) );
  AND2X2 AND2X2_2780 ( .A(core__abc_21380_n4061), .B(reset_n_bF_buf53), .Y(core__abc_21380_n4062_1) );
  AND2X2 AND2X2_2781 ( .A(core__abc_21380_n4060), .B(core__abc_21380_n4062_1), .Y(core_v3_reg_11__FF_INPUT) );
  AND2X2 AND2X2_2782 ( .A(core__abc_21380_n3904), .B(core__abc_21380_n3838_1), .Y(core__abc_21380_n4064) );
  AND2X2 AND2X2_2783 ( .A(core__abc_21380_n4025), .B(core__abc_21380_n3969_1), .Y(core__abc_21380_n4065) );
  AND2X2 AND2X2_2784 ( .A(core__abc_21380_n4065), .B(core__abc_21380_n4064), .Y(core__abc_21380_n4066) );
  AND2X2 AND2X2_2785 ( .A(core__abc_21380_n4070), .B(core__abc_21380_n4071), .Y(core__abc_21380_n4072_1) );
  AND2X2 AND2X2_2786 ( .A(core__abc_21380_n4072_1), .B(core__abc_21380_n4073), .Y(core__abc_21380_n4074) );
  AND2X2 AND2X2_2787 ( .A(core__abc_21380_n4024), .B(core__abc_21380_n3966), .Y(core__abc_21380_n4078) );
  AND2X2 AND2X2_2788 ( .A(core__abc_21380_n4077), .B(core__abc_21380_n4080_1), .Y(core__abc_21380_n4081) );
  AND2X2 AND2X2_2789 ( .A(core__abc_21380_n4068), .B(core__abc_21380_n4081), .Y(core__abc_21380_n4082_1) );
  AND2X2 AND2X2_279 ( .A(_abc_19068_n916_1_bF_buf3), .B(word1_reg_20_), .Y(_abc_19068_n1379_1) );
  AND2X2 AND2X2_2790 ( .A(core__abc_21380_n2044), .B(core__abc_21380_n2063), .Y(core__abc_21380_n4084) );
  AND2X2 AND2X2_2791 ( .A(core__abc_21380_n3946), .B(core__abc_21380_n4084), .Y(core__abc_21380_n4085) );
  AND2X2 AND2X2_2792 ( .A(core__abc_21380_n2060), .B(core__abc_21380_n2042), .Y(core__abc_21380_n4086) );
  AND2X2 AND2X2_2793 ( .A(core__abc_21380_n3887), .B(core__abc_21380_n4084), .Y(core__abc_21380_n4089) );
  AND2X2 AND2X2_2794 ( .A(core__abc_21380_n3807), .B(core__abc_21380_n4089), .Y(core__abc_21380_n4090) );
  AND2X2 AND2X2_2795 ( .A(core__abc_21380_n4091_1), .B(core__abc_21380_n2087), .Y(core__abc_21380_n4092) );
  AND2X2 AND2X2_2796 ( .A(core__abc_21380_n4095_1), .B(core__abc_21380_n4093), .Y(core__abc_21380_n4096) );
  AND2X2 AND2X2_2797 ( .A(core__abc_21380_n4096), .B(core__abc_21380_n2081), .Y(core__abc_21380_n4097) );
  AND2X2 AND2X2_2798 ( .A(core__abc_21380_n3818), .B(core__abc_21380_n3038), .Y(core__abc_21380_n4101) );
  AND2X2 AND2X2_2799 ( .A(core__abc_21380_n4102_1), .B(core__abc_21380_n1491), .Y(core__abc_21380_n4103) );
  AND2X2 AND2X2_28 ( .A(_abc_19068_n877_1), .B(_abc_19068_n911), .Y(_abc_19068_n912_1) );
  AND2X2 AND2X2_280 ( .A(_abc_19068_n941_bF_buf4), .B(core_key_116_), .Y(_abc_19068_n1382) );
  AND2X2 AND2X2_2800 ( .A(core__abc_21380_n4104), .B(core__abc_21380_n1492), .Y(core__abc_21380_n4105) );
  AND2X2 AND2X2_2801 ( .A(core__abc_21380_n4108), .B(core__abc_21380_n4109), .Y(core__abc_21380_n4110) );
  AND2X2 AND2X2_2802 ( .A(core__abc_21380_n4099), .B(core__abc_21380_n4111_1), .Y(core__abc_21380_n4112) );
  AND2X2 AND2X2_2803 ( .A(core__abc_21380_n4098_1), .B(core__abc_21380_n4110), .Y(core__abc_21380_n4113) );
  AND2X2 AND2X2_2804 ( .A(core__abc_21380_n4083), .B(core__abc_21380_n4115_1), .Y(core__abc_21380_n4116) );
  AND2X2 AND2X2_2805 ( .A(core__abc_21380_n4082_1), .B(core__abc_21380_n4114), .Y(core__abc_21380_n4117) );
  AND2X2 AND2X2_2806 ( .A(core__abc_21380_n4120_1), .B(core__abc_21380_n2272), .Y(core__abc_21380_n4121) );
  AND2X2 AND2X2_2807 ( .A(core__abc_21380_n4121), .B(core__abc_21380_n2295), .Y(core__abc_21380_n4122) );
  AND2X2 AND2X2_2808 ( .A(core__abc_21380_n4123), .B(core__abc_21380_n2292), .Y(core__abc_21380_n4124_1) );
  AND2X2 AND2X2_2809 ( .A(core__abc_21380_n4125), .B(core_v3_reg_39_), .Y(core__abc_21380_n4126) );
  AND2X2 AND2X2_281 ( .A(_abc_19068_n945_1_bF_buf4), .B(core_mi_20_), .Y(_abc_19068_n1383_1) );
  AND2X2 AND2X2_2810 ( .A(core__abc_21380_n4128), .B(core__abc_21380_n4129_1), .Y(core__abc_21380_n4130) );
  AND2X2 AND2X2_2811 ( .A(core__abc_21380_n4130), .B(core__abc_21380_n4127), .Y(core__abc_21380_n4131) );
  AND2X2 AND2X2_2812 ( .A(core__abc_21380_n4135), .B(core__abc_21380_n4134), .Y(core__abc_21380_n4136) );
  AND2X2 AND2X2_2813 ( .A(core__abc_21380_n4137), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n4138_1) );
  AND2X2 AND2X2_2814 ( .A(core__abc_21380_n4138_1), .B(core__abc_21380_n4133_1), .Y(core__abc_21380_n4139) );
  AND2X2 AND2X2_2815 ( .A(core__abc_21380_n3313_bF_buf12), .B(core_key_76_), .Y(core__abc_21380_n4140) );
  AND2X2 AND2X2_2816 ( .A(core_v3_reg_12_), .B(core_mi_12_), .Y(core__abc_21380_n4142) );
  AND2X2 AND2X2_2817 ( .A(core__abc_21380_n4143), .B(core__abc_21380_n4141_1), .Y(core__abc_21380_n4144) );
  AND2X2 AND2X2_2818 ( .A(core__abc_21380_n2749_bF_buf10), .B(core__abc_21380_n4144), .Y(core__abc_21380_n4145_1) );
  AND2X2 AND2X2_2819 ( .A(core__abc_21380_n4149_1), .B(reset_n_bF_buf52), .Y(core__abc_21380_n4150) );
  AND2X2 AND2X2_282 ( .A(_abc_19068_n915_1_bF_buf3), .B(core_mi_52_), .Y(_abc_19068_n1385_1) );
  AND2X2 AND2X2_2820 ( .A(core__abc_21380_n4148), .B(core__abc_21380_n4150), .Y(core_v3_reg_12__FF_INPUT) );
  AND2X2 AND2X2_2821 ( .A(core__abc_21380_n4153_1), .B(core__abc_21380_n4152), .Y(core__abc_21380_n4154) );
  AND2X2 AND2X2_2822 ( .A(core__abc_21380_n4156), .B(core__abc_21380_n2101), .Y(core__abc_21380_n4158) );
  AND2X2 AND2X2_2823 ( .A(core__abc_21380_n4159), .B(core__abc_21380_n4157_1), .Y(core__abc_21380_n4160) );
  AND2X2 AND2X2_2824 ( .A(core__abc_21380_n4163), .B(core__abc_21380_n1511), .Y(core__abc_21380_n4164) );
  AND2X2 AND2X2_2825 ( .A(core__abc_21380_n4162), .B(core__abc_21380_n1509), .Y(core__abc_21380_n4165_1) );
  AND2X2 AND2X2_2826 ( .A(core__abc_21380_n4166), .B(core__abc_21380_n4161_1), .Y(core__abc_21380_n4167) );
  AND2X2 AND2X2_2827 ( .A(core__abc_21380_n4168), .B(core_v3_reg_61_), .Y(core__abc_21380_n4169) );
  AND2X2 AND2X2_2828 ( .A(core__abc_21380_n4160), .B(core__abc_21380_n4171), .Y(core__abc_21380_n4172) );
  AND2X2 AND2X2_2829 ( .A(core__abc_21380_n4174), .B(core__abc_21380_n4170_1), .Y(core__abc_21380_n4175) );
  AND2X2 AND2X2_283 ( .A(_abc_19068_n897_1_bF_buf3), .B(word0_reg_20_), .Y(_abc_19068_n1386) );
  AND2X2 AND2X2_2830 ( .A(core__abc_21380_n4176), .B(core__abc_21380_n4173_1), .Y(core__abc_21380_n4177) );
  AND2X2 AND2X2_2831 ( .A(core__abc_21380_n4155), .B(core__abc_21380_n4178_1), .Y(core__abc_21380_n4179) );
  AND2X2 AND2X2_2832 ( .A(core__abc_21380_n4154), .B(core__abc_21380_n4177), .Y(core__abc_21380_n4180) );
  AND2X2 AND2X2_2833 ( .A(core__abc_21380_n2273), .B(core__abc_21380_n2292), .Y(core__abc_21380_n4183) );
  AND2X2 AND2X2_2834 ( .A(core__abc_21380_n4031_1), .B(core__abc_21380_n4183), .Y(core__abc_21380_n4184) );
  AND2X2 AND2X2_2835 ( .A(core__abc_21380_n3917), .B(core__abc_21380_n4184), .Y(core__abc_21380_n4185) );
  AND2X2 AND2X2_2836 ( .A(core__abc_21380_n4186_1), .B(core__abc_21380_n4183), .Y(core__abc_21380_n4187) );
  AND2X2 AND2X2_2837 ( .A(core__abc_21380_n2289), .B(core__abc_21380_n2271), .Y(core__abc_21380_n4188) );
  AND2X2 AND2X2_2838 ( .A(core__abc_21380_n3636_1), .B(core__abc_21380_n3911), .Y(core__abc_21380_n4192) );
  AND2X2 AND2X2_2839 ( .A(core__abc_21380_n4192), .B(core__abc_21380_n4184), .Y(core__abc_21380_n4193) );
  AND2X2 AND2X2_284 ( .A(_abc_19068_n923_bF_buf4), .B(_abc_19068_n1390), .Y(_auto_iopadmap_cc_313_execute_30317_20_) );
  AND2X2 AND2X2_2840 ( .A(core__abc_21380_n4195), .B(core__abc_21380_n2313), .Y(core__abc_21380_n4196) );
  AND2X2 AND2X2_2841 ( .A(core__abc_21380_n4194_1), .B(core__abc_21380_n2311), .Y(core__abc_21380_n4197) );
  AND2X2 AND2X2_2842 ( .A(core__abc_21380_n4200), .B(core__abc_21380_n4201), .Y(core__abc_21380_n4202) );
  AND2X2 AND2X2_2843 ( .A(core__abc_21380_n4206_1), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n4207) );
  AND2X2 AND2X2_2844 ( .A(core__abc_21380_n4207), .B(core__abc_21380_n4204), .Y(core__abc_21380_n4208) );
  AND2X2 AND2X2_2845 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n4209), .Y(core__abc_21380_n4210_1) );
  AND2X2 AND2X2_2846 ( .A(core_v3_reg_13_), .B(core_mi_13_), .Y(core__abc_21380_n4212) );
  AND2X2 AND2X2_2847 ( .A(core__abc_21380_n4213), .B(core__abc_21380_n4211), .Y(core__abc_21380_n4214) );
  AND2X2 AND2X2_2848 ( .A(core__abc_21380_n2749_bF_buf9), .B(core__abc_21380_n4214), .Y(core__abc_21380_n4215) );
  AND2X2 AND2X2_2849 ( .A(core__abc_21380_n4219), .B(reset_n_bF_buf51), .Y(core__abc_21380_n4220) );
  AND2X2 AND2X2_285 ( .A(_abc_19068_n945_1_bF_buf3), .B(core_mi_21_), .Y(_abc_19068_n1392) );
  AND2X2 AND2X2_2850 ( .A(core__abc_21380_n4218_1), .B(core__abc_21380_n4220), .Y(core_v3_reg_13__FF_INPUT) );
  AND2X2 AND2X2_2851 ( .A(core__abc_21380_n2087), .B(core__abc_21380_n2101), .Y(core__abc_21380_n4222) );
  AND2X2 AND2X2_2852 ( .A(core__abc_21380_n4225), .B(core__abc_21380_n2100), .Y(core__abc_21380_n4226) );
  AND2X2 AND2X2_2853 ( .A(core__abc_21380_n4224_1), .B(core__abc_21380_n4227), .Y(core__abc_21380_n4228) );
  AND2X2 AND2X2_2854 ( .A(core__abc_21380_n4228), .B(core__abc_21380_n2119), .Y(core__abc_21380_n4229) );
  AND2X2 AND2X2_2855 ( .A(core__abc_21380_n4091_1), .B(core__abc_21380_n4222), .Y(core__abc_21380_n4230_1) );
  AND2X2 AND2X2_2856 ( .A(core__abc_21380_n4232), .B(core__abc_21380_n2125), .Y(core__abc_21380_n4233) );
  AND2X2 AND2X2_2857 ( .A(core__abc_21380_n4102_1), .B(core__abc_21380_n3034), .Y(core__abc_21380_n4237_1) );
  AND2X2 AND2X2_2858 ( .A(core__abc_21380_n4239), .B(core__abc_21380_n1529), .Y(core__abc_21380_n4240) );
  AND2X2 AND2X2_2859 ( .A(core__abc_21380_n4238), .B(core__abc_21380_n1527), .Y(core__abc_21380_n4241) );
  AND2X2 AND2X2_286 ( .A(_abc_19068_n915_1_bF_buf2), .B(core_mi_53_), .Y(_abc_19068_n1393_1) );
  AND2X2 AND2X2_2860 ( .A(core__abc_21380_n4244), .B(core__abc_21380_n4245), .Y(core__abc_21380_n4246) );
  AND2X2 AND2X2_2861 ( .A(core__abc_21380_n4235), .B(core__abc_21380_n4247), .Y(core__abc_21380_n4248) );
  AND2X2 AND2X2_2862 ( .A(core__abc_21380_n4234), .B(core__abc_21380_n4246), .Y(core__abc_21380_n4249_1) );
  AND2X2 AND2X2_2863 ( .A(core__abc_21380_n4173_1), .B(core__abc_21380_n4152), .Y(core__abc_21380_n4251) );
  AND2X2 AND2X2_2864 ( .A(core__abc_21380_n4177), .B(core__abc_21380_n4115_1), .Y(core__abc_21380_n4253) );
  AND2X2 AND2X2_2865 ( .A(core__abc_21380_n4255_1), .B(core__abc_21380_n4252), .Y(core__abc_21380_n4256) );
  AND2X2 AND2X2_2866 ( .A(core__abc_21380_n4256), .B(core__abc_21380_n4250), .Y(core__abc_21380_n4257) );
  AND2X2 AND2X2_2867 ( .A(core__abc_21380_n2329), .B(core__abc_21380_n2309), .Y(core__abc_21380_n4262_1) );
  AND2X2 AND2X2_2868 ( .A(core__abc_21380_n2331), .B(core__abc_21380_n2310), .Y(core__abc_21380_n4264) );
  AND2X2 AND2X2_2869 ( .A(core__abc_21380_n4263), .B(core__abc_21380_n4264), .Y(core__abc_21380_n4265) );
  AND2X2 AND2X2_287 ( .A(_abc_19068_n899_bF_buf2), .B(word3_reg_21_), .Y(_abc_19068_n1395_1) );
  AND2X2 AND2X2_2870 ( .A(core__abc_21380_n4197), .B(core__abc_21380_n2329), .Y(core__abc_21380_n4266) );
  AND2X2 AND2X2_2871 ( .A(core__abc_21380_n4268), .B(core__abc_21380_n4261), .Y(core__abc_21380_n4269) );
  AND2X2 AND2X2_2872 ( .A(core__abc_21380_n4270), .B(core_v3_reg_41_), .Y(core__abc_21380_n4271) );
  AND2X2 AND2X2_2873 ( .A(core__abc_21380_n4276), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf2), .Y(core__abc_21380_n4277) );
  AND2X2 AND2X2_2874 ( .A(core__abc_21380_n4277), .B(core__abc_21380_n4273_1), .Y(core__abc_21380_n4278_1) );
  AND2X2 AND2X2_2875 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n4279), .Y(core__abc_21380_n4280) );
  AND2X2 AND2X2_2876 ( .A(core_v3_reg_14_), .B(core_mi_14_), .Y(core__abc_21380_n4282) );
  AND2X2 AND2X2_2877 ( .A(core__abc_21380_n4283), .B(core__abc_21380_n4281), .Y(core__abc_21380_n4284_1) );
  AND2X2 AND2X2_2878 ( .A(core__abc_21380_n2749_bF_buf8), .B(core__abc_21380_n4284_1), .Y(core__abc_21380_n4285) );
  AND2X2 AND2X2_2879 ( .A(core__abc_21380_n4289_1), .B(reset_n_bF_buf50), .Y(core__abc_21380_n4290) );
  AND2X2 AND2X2_288 ( .A(_abc_19068_n902_bF_buf2), .B(word2_reg_21_), .Y(_abc_19068_n1396) );
  AND2X2 AND2X2_2880 ( .A(core__abc_21380_n4288), .B(core__abc_21380_n4290), .Y(core_v3_reg_14__FF_INPUT) );
  AND2X2 AND2X2_2881 ( .A(core__abc_21380_n4258), .B(core__abc_21380_n4292), .Y(core__abc_21380_n4293) );
  AND2X2 AND2X2_2882 ( .A(core__abc_21380_n4295), .B(core__abc_21380_n4294_1), .Y(core__abc_21380_n4296) );
  AND2X2 AND2X2_2883 ( .A(core__abc_21380_n4296), .B(core__abc_21380_n2140), .Y(core__abc_21380_n4297) );
  AND2X2 AND2X2_2884 ( .A(core__abc_21380_n4298), .B(core__abc_21380_n2139_1), .Y(core__abc_21380_n4299_1) );
  AND2X2 AND2X2_2885 ( .A(core__abc_21380_n4303), .B(core__abc_21380_n1549), .Y(core__abc_21380_n4304_1) );
  AND2X2 AND2X2_2886 ( .A(core__abc_21380_n4302), .B(core__abc_21380_n1546), .Y(core__abc_21380_n4305) );
  AND2X2 AND2X2_2887 ( .A(core__abc_21380_n4306), .B(core__abc_21380_n4301), .Y(core__abc_21380_n4307) );
  AND2X2 AND2X2_2888 ( .A(core__abc_21380_n4308), .B(core_v3_reg_63_), .Y(core__abc_21380_n4309_1) );
  AND2X2 AND2X2_2889 ( .A(core__abc_21380_n4314_1), .B(core__abc_21380_n4313), .Y(core__abc_21380_n4315) );
  AND2X2 AND2X2_289 ( .A(_abc_19068_n926_bF_buf3), .B(core_key_21_), .Y(_abc_19068_n1399_1) );
  AND2X2 AND2X2_2890 ( .A(core__abc_21380_n4312), .B(core__abc_21380_n4316), .Y(core__abc_21380_n4317) );
  AND2X2 AND2X2_2891 ( .A(core__abc_21380_n4293), .B(core__abc_21380_n4317), .Y(core__abc_21380_n4318) );
  AND2X2 AND2X2_2892 ( .A(core__abc_21380_n4319_1), .B(core__abc_21380_n4320), .Y(core__abc_21380_n4321) );
  AND2X2 AND2X2_2893 ( .A(core__abc_21380_n4324_1), .B(core__abc_21380_n2347), .Y(core__abc_21380_n4325) );
  AND2X2 AND2X2_2894 ( .A(core__abc_21380_n4326), .B(core__abc_21380_n4327), .Y(core__abc_21380_n4328) );
  AND2X2 AND2X2_2895 ( .A(core__abc_21380_n4332), .B(core__abc_21380_n4329_1), .Y(core__abc_21380_n4333) );
  AND2X2 AND2X2_2896 ( .A(core__abc_21380_n4336), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf2), .Y(core__abc_21380_n4337) );
  AND2X2 AND2X2_2897 ( .A(core__abc_21380_n4337), .B(core__abc_21380_n4335), .Y(core__abc_21380_n4338) );
  AND2X2 AND2X2_2898 ( .A(core__abc_21380_n3313_bF_buf9), .B(core_key_79_), .Y(core__abc_21380_n4339_1) );
  AND2X2 AND2X2_2899 ( .A(core_v3_reg_15_), .B(core_mi_15_), .Y(core__abc_21380_n4341) );
  AND2X2 AND2X2_29 ( .A(_abc_19068_n913_1), .B(_abc_19068_n912_1), .Y(_abc_19068_n914) );
  AND2X2 AND2X2_290 ( .A(_abc_19068_n924_1_bF_buf3), .B(core_key_53_), .Y(_abc_19068_n1400) );
  AND2X2 AND2X2_2900 ( .A(core__abc_21380_n4342), .B(core__abc_21380_n4340), .Y(core__abc_21380_n4343) );
  AND2X2 AND2X2_2901 ( .A(core__abc_21380_n2749_bF_buf7), .B(core__abc_21380_n4343), .Y(core__abc_21380_n4344_1) );
  AND2X2 AND2X2_2902 ( .A(core__abc_21380_n4348), .B(reset_n_bF_buf49), .Y(core__abc_21380_n4349_1) );
  AND2X2 AND2X2_2903 ( .A(core__abc_21380_n4347), .B(core__abc_21380_n4349_1), .Y(core_v3_reg_15__FF_INPUT) );
  AND2X2 AND2X2_2904 ( .A(core__abc_21380_n3846), .B(core__abc_21380_n4066), .Y(core__abc_21380_n4351) );
  AND2X2 AND2X2_2905 ( .A(core__abc_21380_n4353), .B(core__abc_21380_n4354), .Y(core__abc_21380_n4355_1) );
  AND2X2 AND2X2_2906 ( .A(core__abc_21380_n4355_1), .B(core__abc_21380_n4352), .Y(core__abc_21380_n4356) );
  AND2X2 AND2X2_2907 ( .A(core__abc_21380_n4356), .B(core__abc_21380_n4253), .Y(core__abc_21380_n4357) );
  AND2X2 AND2X2_2908 ( .A(core__abc_21380_n4351), .B(core__abc_21380_n4357), .Y(core__abc_21380_n4358) );
  AND2X2 AND2X2_2909 ( .A(core__abc_21380_n4065), .B(core__abc_21380_n4359), .Y(core__abc_21380_n4360) );
  AND2X2 AND2X2_291 ( .A(_abc_19068_n941_bF_buf3), .B(core_key_117_), .Y(_abc_19068_n1402) );
  AND2X2 AND2X2_2910 ( .A(core__abc_21380_n4357), .B(core__abc_21380_n4361_1), .Y(core__abc_21380_n4362) );
  AND2X2 AND2X2_2911 ( .A(core__abc_21380_n4356), .B(core__abc_21380_n4363), .Y(core__abc_21380_n4364) );
  AND2X2 AND2X2_2912 ( .A(core__abc_21380_n4354), .B(core__abc_21380_n4248), .Y(core__abc_21380_n4366_1) );
  AND2X2 AND2X2_2913 ( .A(core__abc_21380_n2125), .B(core__abc_21380_n2139_1), .Y(core__abc_21380_n4371_1) );
  AND2X2 AND2X2_2914 ( .A(core__abc_21380_n4222), .B(core__abc_21380_n4371_1), .Y(core__abc_21380_n4372) );
  AND2X2 AND2X2_2915 ( .A(core__abc_21380_n4089), .B(core__abc_21380_n4372), .Y(core__abc_21380_n4373) );
  AND2X2 AND2X2_2916 ( .A(core__abc_21380_n3805), .B(core__abc_21380_n4373), .Y(core__abc_21380_n4374) );
  AND2X2 AND2X2_2917 ( .A(core__abc_21380_n3269), .B(core__abc_21380_n4374), .Y(core__abc_21380_n4375) );
  AND2X2 AND2X2_2918 ( .A(core__abc_21380_n3804), .B(core__abc_21380_n4373), .Y(core__abc_21380_n4376_1) );
  AND2X2 AND2X2_2919 ( .A(core__abc_21380_n4088), .B(core__abc_21380_n4372), .Y(core__abc_21380_n4377) );
  AND2X2 AND2X2_292 ( .A(_abc_19068_n939_1_bF_buf3), .B(core_key_85_), .Y(_abc_19068_n1403_1) );
  AND2X2 AND2X2_2920 ( .A(core__abc_21380_n4231), .B(core__abc_21380_n4371_1), .Y(core__abc_21380_n4378) );
  AND2X2 AND2X2_2921 ( .A(core__abc_21380_n2138), .B(core__abc_21380_n2115), .Y(core__abc_21380_n4379) );
  AND2X2 AND2X2_2922 ( .A(core__abc_21380_n4384), .B(core__abc_21380_n2158), .Y(core__abc_21380_n4385) );
  AND2X2 AND2X2_2923 ( .A(core__abc_21380_n4387), .B(core__abc_21380_n4388), .Y(core__abc_21380_n4389) );
  AND2X2 AND2X2_2924 ( .A(core__abc_21380_n4389), .B(core__abc_21380_n2157), .Y(core__abc_21380_n4390) );
  AND2X2 AND2X2_2925 ( .A(core__abc_21380_n3060), .B(core__abc_21380_n1566), .Y(core__abc_21380_n4393) );
  AND2X2 AND2X2_2926 ( .A(core__abc_21380_n4394), .B(core__abc_21380_n1565), .Y(core__abc_21380_n4395) );
  AND2X2 AND2X2_2927 ( .A(core__abc_21380_n4398), .B(core__abc_21380_n4399), .Y(core__abc_21380_n4400) );
  AND2X2 AND2X2_2928 ( .A(core__abc_21380_n4392_1), .B(core__abc_21380_n4400), .Y(core__abc_21380_n4401) );
  AND2X2 AND2X2_2929 ( .A(core__abc_21380_n4402_1), .B(core__abc_21380_n4391), .Y(core__abc_21380_n4403) );
  AND2X2 AND2X2_293 ( .A(_abc_19068_n897_1_bF_buf2), .B(word0_reg_21_), .Y(_abc_19068_n1406) );
  AND2X2 AND2X2_2930 ( .A(core__abc_21380_n4370), .B(core__abc_21380_n4405), .Y(core__abc_21380_n4406) );
  AND2X2 AND2X2_2931 ( .A(core__abc_21380_n4411), .B(core__abc_21380_n4412_1), .Y(core__abc_21380_n4413) );
  AND2X2 AND2X2_2932 ( .A(core__abc_21380_n4410), .B(core__abc_21380_n4413), .Y(core__abc_21380_n4414) );
  AND2X2 AND2X2_2933 ( .A(core__abc_21380_n4414), .B(core__abc_21380_n4409), .Y(core__abc_21380_n4415) );
  AND2X2 AND2X2_2934 ( .A(core__abc_21380_n4415), .B(core__abc_21380_n4404), .Y(core__abc_21380_n4416) );
  AND2X2 AND2X2_2935 ( .A(core__abc_21380_n4326), .B(core__abc_21380_n2346), .Y(core__abc_21380_n4418) );
  AND2X2 AND2X2_2936 ( .A(core__abc_21380_n4418), .B(core__abc_21380_n2369_1), .Y(core__abc_21380_n4419) );
  AND2X2 AND2X2_2937 ( .A(core__abc_21380_n4420), .B(core__abc_21380_n4421), .Y(core__abc_21380_n4422_1) );
  AND2X2 AND2X2_2938 ( .A(core__abc_21380_n4422_1), .B(core_v3_reg_43_), .Y(core__abc_21380_n4425) );
  AND2X2 AND2X2_2939 ( .A(core__abc_21380_n4429), .B(core__abc_21380_n4423), .Y(core__abc_21380_n4430) );
  AND2X2 AND2X2_294 ( .A(_abc_19068_n916_1_bF_buf2), .B(word1_reg_21_), .Y(_abc_19068_n1407_1) );
  AND2X2 AND2X2_2940 ( .A(core__abc_21380_n4431), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n4432_1) );
  AND2X2 AND2X2_2941 ( .A(core__abc_21380_n4432_1), .B(core__abc_21380_n4427_1), .Y(core__abc_21380_n4433) );
  AND2X2 AND2X2_2942 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_80_), .Y(core__abc_21380_n4434) );
  AND2X2 AND2X2_2943 ( .A(core_v3_reg_16_), .B(core_mi_16_), .Y(core__abc_21380_n4436) );
  AND2X2 AND2X2_2944 ( .A(core__abc_21380_n4437), .B(core__abc_21380_n4435), .Y(core__abc_21380_n4438_1) );
  AND2X2 AND2X2_2945 ( .A(core__abc_21380_n2749_bF_buf6), .B(core__abc_21380_n4438_1), .Y(core__abc_21380_n4439) );
  AND2X2 AND2X2_2946 ( .A(core__abc_21380_n4443_1), .B(reset_n_bF_buf48), .Y(core__abc_21380_n4444) );
  AND2X2 AND2X2_2947 ( .A(core__abc_21380_n4442), .B(core__abc_21380_n4444), .Y(core_v3_reg_16__FF_INPUT) );
  AND2X2 AND2X2_2948 ( .A(core__abc_21380_n4447), .B(core__abc_21380_n4446), .Y(core__abc_21380_n4448_1) );
  AND2X2 AND2X2_2949 ( .A(core__abc_21380_n2175), .B(core__abc_21380_n4451), .Y(core__abc_21380_n4452) );
  AND2X2 AND2X2_295 ( .A(_abc_19068_n1411_1), .B(_abc_19068_n923_bF_buf3), .Y(_auto_iopadmap_cc_313_execute_30317_21_) );
  AND2X2 AND2X2_2950 ( .A(core__abc_21380_n4450), .B(core__abc_21380_n4452), .Y(core__abc_21380_n4453) );
  AND2X2 AND2X2_2951 ( .A(core__abc_21380_n2181), .B(core__abc_21380_n2156), .Y(core__abc_21380_n4455) );
  AND2X2 AND2X2_2952 ( .A(core__abc_21380_n2158), .B(core__abc_21380_n2181), .Y(core__abc_21380_n4457) );
  AND2X2 AND2X2_2953 ( .A(core__abc_21380_n4384), .B(core__abc_21380_n4457), .Y(core__abc_21380_n4458) );
  AND2X2 AND2X2_2954 ( .A(core__abc_21380_n4459_1), .B(core__abc_21380_n4456), .Y(core__abc_21380_n4460) );
  AND2X2 AND2X2_2955 ( .A(core__abc_21380_n4454_1), .B(core__abc_21380_n4460), .Y(core__abc_21380_n4461) );
  AND2X2 AND2X2_2956 ( .A(core__abc_21380_n4463), .B(core__abc_21380_n1585), .Y(core__abc_21380_n4464_1) );
  AND2X2 AND2X2_2957 ( .A(core__abc_21380_n4462), .B(core__abc_21380_n1584), .Y(core__abc_21380_n4465) );
  AND2X2 AND2X2_2958 ( .A(core__abc_21380_n4466), .B(core__abc_21380_n1282_1), .Y(core__abc_21380_n4467) );
  AND2X2 AND2X2_2959 ( .A(core__abc_21380_n4468), .B(core_v3_reg_1_), .Y(core__abc_21380_n4469_1) );
  AND2X2 AND2X2_296 ( .A(_abc_19068_n899_bF_buf1), .B(word3_reg_22_), .Y(_abc_19068_n1413_1) );
  AND2X2 AND2X2_2960 ( .A(core__abc_21380_n4471), .B(core__abc_21380_n4461), .Y(core__abc_21380_n4472) );
  AND2X2 AND2X2_2961 ( .A(core__abc_21380_n4470), .B(core__abc_21380_n4474_1), .Y(core__abc_21380_n4475) );
  AND2X2 AND2X2_2962 ( .A(core__abc_21380_n4473), .B(core__abc_21380_n4476), .Y(core__abc_21380_n4477) );
  AND2X2 AND2X2_2963 ( .A(core__abc_21380_n4478), .B(core__abc_21380_n4480_1), .Y(core__abc_21380_n4481) );
  AND2X2 AND2X2_2964 ( .A(core__abc_21380_n4325), .B(core__abc_21380_n2366), .Y(core__abc_21380_n4483) );
  AND2X2 AND2X2_2965 ( .A(core__abc_21380_n2366), .B(core__abc_21380_n2345), .Y(core__abc_21380_n4484) );
  AND2X2 AND2X2_2966 ( .A(core__abc_21380_n4487), .B(core__abc_21380_n2387), .Y(core__abc_21380_n4488) );
  AND2X2 AND2X2_2967 ( .A(core__abc_21380_n4486), .B(core__abc_21380_n2385), .Y(core__abc_21380_n4489) );
  AND2X2 AND2X2_2968 ( .A(core__abc_21380_n4492), .B(core__abc_21380_n4494), .Y(core__abc_21380_n4495) );
  AND2X2 AND2X2_2969 ( .A(core__abc_21380_n4498), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n4499) );
  AND2X2 AND2X2_297 ( .A(_abc_19068_n945_1_bF_buf2), .B(core_mi_22_), .Y(_abc_19068_n1415_1) );
  AND2X2 AND2X2_2970 ( .A(core__abc_21380_n4499), .B(core__abc_21380_n4497), .Y(core__abc_21380_n4500) );
  AND2X2 AND2X2_2971 ( .A(core__abc_21380_n3313_bF_buf7), .B(core_key_81_), .Y(core__abc_21380_n4501_1) );
  AND2X2 AND2X2_2972 ( .A(core_v3_reg_17_), .B(core_mi_17_), .Y(core__abc_21380_n4503) );
  AND2X2 AND2X2_2973 ( .A(core__abc_21380_n4504), .B(core__abc_21380_n4502), .Y(core__abc_21380_n4505) );
  AND2X2 AND2X2_2974 ( .A(core__abc_21380_n2749_bF_buf5), .B(core__abc_21380_n4505), .Y(core__abc_21380_n4506_1) );
  AND2X2 AND2X2_2975 ( .A(core__abc_21380_n4510), .B(reset_n_bF_buf47), .Y(core__abc_21380_n4511_1) );
  AND2X2 AND2X2_2976 ( .A(core__abc_21380_n4509), .B(core__abc_21380_n4511_1), .Y(core_v3_reg_17__FF_INPUT) );
  AND2X2 AND2X2_2977 ( .A(core__abc_21380_n4473), .B(core__abc_21380_n4513), .Y(core__abc_21380_n4514) );
  AND2X2 AND2X2_2978 ( .A(core__abc_21380_n4477), .B(core__abc_21380_n4405), .Y(core__abc_21380_n4516_1) );
  AND2X2 AND2X2_2979 ( .A(core__abc_21380_n4370), .B(core__abc_21380_n4516_1), .Y(core__abc_21380_n4517) );
  AND2X2 AND2X2_298 ( .A(_abc_19068_n941_bF_buf2), .B(core_key_118_), .Y(_abc_19068_n1416) );
  AND2X2 AND2X2_2980 ( .A(core__abc_21380_n4522_1), .B(core__abc_21380_n2193), .Y(core__abc_21380_n4523) );
  AND2X2 AND2X2_2981 ( .A(core__abc_21380_n4521), .B(core__abc_21380_n2199), .Y(core__abc_21380_n4524) );
  AND2X2 AND2X2_2982 ( .A(core__abc_21380_n4528), .B(core__abc_21380_n3080), .Y(core__abc_21380_n4529) );
  AND2X2 AND2X2_2983 ( .A(core__abc_21380_n4529), .B(core__abc_21380_n1604), .Y(core__abc_21380_n4530) );
  AND2X2 AND2X2_2984 ( .A(core__abc_21380_n4535), .B(core__abc_21380_n4536), .Y(core__abc_21380_n4537_1) );
  AND2X2 AND2X2_2985 ( .A(core__abc_21380_n4526), .B(core__abc_21380_n4538), .Y(core__abc_21380_n4539) );
  AND2X2 AND2X2_2986 ( .A(core__abc_21380_n4525), .B(core__abc_21380_n4537_1), .Y(core__abc_21380_n4540) );
  AND2X2 AND2X2_2987 ( .A(core__abc_21380_n4519), .B(core__abc_21380_n4541), .Y(core__abc_21380_n4542_1) );
  AND2X2 AND2X2_2988 ( .A(core__abc_21380_n4518), .B(core__abc_21380_n4543), .Y(core__abc_21380_n4544) );
  AND2X2 AND2X2_2989 ( .A(core__abc_21380_n4546), .B(core__abc_21380_n2405), .Y(core__abc_21380_n4547_1) );
  AND2X2 AND2X2_299 ( .A(_abc_19068_n939_1_bF_buf2), .B(core_key_86_), .Y(_abc_19068_n1419_1) );
  AND2X2 AND2X2_2990 ( .A(core__abc_21380_n4548), .B(core__abc_21380_n2403), .Y(core__abc_21380_n4549) );
  AND2X2 AND2X2_2991 ( .A(core__abc_21380_n4550), .B(core_v3_reg_45_), .Y(core__abc_21380_n4551) );
  AND2X2 AND2X2_2992 ( .A(core__abc_21380_n4552_1), .B(core__abc_21380_n4553), .Y(core__abc_21380_n4554) );
  AND2X2 AND2X2_2993 ( .A(core__abc_21380_n4558), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n4559) );
  AND2X2 AND2X2_2994 ( .A(core__abc_21380_n4559), .B(core__abc_21380_n4556), .Y(core__abc_21380_n4560_1) );
  AND2X2 AND2X2_2995 ( .A(core__abc_21380_n3313_bF_buf6), .B(core__abc_21380_n4561), .Y(core__abc_21380_n4562) );
  AND2X2 AND2X2_2996 ( .A(core_v3_reg_18_), .B(core_mi_18_), .Y(core__abc_21380_n4564) );
  AND2X2 AND2X2_2997 ( .A(core__abc_21380_n4565_1), .B(core__abc_21380_n4563), .Y(core__abc_21380_n4566) );
  AND2X2 AND2X2_2998 ( .A(core__abc_21380_n2749_bF_buf4), .B(core__abc_21380_n4566), .Y(core__abc_21380_n4567) );
  AND2X2 AND2X2_2999 ( .A(core__abc_21380_n4571_1), .B(reset_n_bF_buf46), .Y(core__abc_21380_n4572) );
  AND2X2 AND2X2_3 ( .A(_abc_19068_n871_1), .B(_abc_19068_n873_1), .Y(_abc_19068_n874_1) );
  AND2X2 AND2X2_30 ( .A(_abc_19068_n912_1), .B(_abc_19068_n874_1), .Y(_abc_19068_n915_1) );
  AND2X2 AND2X2_300 ( .A(_abc_19068_n924_1_bF_buf2), .B(core_key_54_), .Y(_abc_19068_n1420) );
  AND2X2 AND2X2_3000 ( .A(core__abc_21380_n4570), .B(core__abc_21380_n4572), .Y(core_v3_reg_18__FF_INPUT) );
  AND2X2 AND2X2_3001 ( .A(core__abc_21380_n4548), .B(core__abc_21380_n2402), .Y(core__abc_21380_n4576_1) );
  AND2X2 AND2X2_3002 ( .A(core__abc_21380_n4578), .B(core__abc_21380_n2421), .Y(core__abc_21380_n4579) );
  AND2X2 AND2X2_3003 ( .A(core__abc_21380_n4577), .B(core__abc_21380_n2423), .Y(core__abc_21380_n4580) );
  AND2X2 AND2X2_3004 ( .A(core__abc_21380_n4581), .B(core__abc_21380_n4574), .Y(core__abc_21380_n4582_1) );
  AND2X2 AND2X2_3005 ( .A(core__abc_21380_n4583), .B(core_v3_reg_46_), .Y(core__abc_21380_n4584) );
  AND2X2 AND2X2_3006 ( .A(core__abc_21380_n4587_1), .B(core__abc_21380_n4586), .Y(core__abc_21380_n4588) );
  AND2X2 AND2X2_3007 ( .A(core__abc_21380_n4590), .B(core__abc_21380_n2213_1), .Y(core__abc_21380_n4592_1) );
  AND2X2 AND2X2_3008 ( .A(core__abc_21380_n4593), .B(core__abc_21380_n4591), .Y(core__abc_21380_n4594) );
  AND2X2 AND2X2_3009 ( .A(core__abc_21380_n4531), .B(core__abc_21380_n1599), .Y(core__abc_21380_n4595) );
  AND2X2 AND2X2_301 ( .A(_abc_19068_n926_bF_buf2), .B(core_key_22_), .Y(_abc_19068_n1421_1) );
  AND2X2 AND2X2_3010 ( .A(core__abc_21380_n4595), .B(core__abc_21380_n1619), .Y(core__abc_21380_n4596) );
  AND2X2 AND2X2_3011 ( .A(core__abc_21380_n4597_1), .B(core__abc_21380_n4598), .Y(core__abc_21380_n4599) );
  AND2X2 AND2X2_3012 ( .A(core__abc_21380_n4600), .B(core__abc_21380_n1325), .Y(core__abc_21380_n4601) );
  AND2X2 AND2X2_3013 ( .A(core__abc_21380_n4599), .B(core_v3_reg_3_), .Y(core__abc_21380_n4602) );
  AND2X2 AND2X2_3014 ( .A(core__abc_21380_n4604), .B(core__abc_21380_n4594), .Y(core__abc_21380_n4605) );
  AND2X2 AND2X2_3015 ( .A(core__abc_21380_n4606), .B(core__abc_21380_n4603_1), .Y(core__abc_21380_n4607) );
  AND2X2 AND2X2_3016 ( .A(core__abc_21380_n4610), .B(core__abc_21380_n4611), .Y(core__abc_21380_n4612) );
  AND2X2 AND2X2_3017 ( .A(core__abc_21380_n4613), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n4614_1) );
  AND2X2 AND2X2_3018 ( .A(core__abc_21380_n4612), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n4617) );
  AND2X2 AND2X2_3019 ( .A(core__abc_21380_n4615), .B(core__abc_21380_n4618), .Y(core__abc_21380_n4619_1) );
  AND2X2 AND2X2_302 ( .A(_abc_19068_n916_1_bF_buf1), .B(word1_reg_22_), .Y(_abc_19068_n1424) );
  AND2X2 AND2X2_3020 ( .A(core__abc_21380_n3313_bF_buf5), .B(core_key_83_), .Y(core__abc_21380_n4620) );
  AND2X2 AND2X2_3021 ( .A(core_v3_reg_19_), .B(core_mi_19_), .Y(core__abc_21380_n4621) );
  AND2X2 AND2X2_3022 ( .A(core__abc_21380_n4622), .B(core__abc_21380_n4623), .Y(core__abc_21380_n4624_1) );
  AND2X2 AND2X2_3023 ( .A(core__abc_21380_n2749_bF_buf3), .B(core__abc_21380_n4624_1), .Y(core__abc_21380_n4625) );
  AND2X2 AND2X2_3024 ( .A(core__abc_21380_n4629_1), .B(reset_n_bF_buf45), .Y(core__abc_21380_n4630) );
  AND2X2 AND2X2_3025 ( .A(core__abc_21380_n4628), .B(core__abc_21380_n4630), .Y(core_v3_reg_19__FF_INPUT) );
  AND2X2 AND2X2_3026 ( .A(core__abc_21380_n2199), .B(core__abc_21380_n2213_1), .Y(core__abc_21380_n4632) );
  AND2X2 AND2X2_3027 ( .A(core__abc_21380_n4520), .B(core__abc_21380_n4632), .Y(core__abc_21380_n4633) );
  AND2X2 AND2X2_3028 ( .A(core__abc_21380_n2212), .B(core__abc_21380_n2189), .Y(core__abc_21380_n4634_1) );
  AND2X2 AND2X2_3029 ( .A(core__abc_21380_n4457), .B(core__abc_21380_n4632), .Y(core__abc_21380_n4637) );
  AND2X2 AND2X2_303 ( .A(_abc_19068_n902_bF_buf1), .B(word2_reg_22_), .Y(_abc_19068_n1425_1) );
  AND2X2 AND2X2_3030 ( .A(core__abc_21380_n4384), .B(core__abc_21380_n4637), .Y(core__abc_21380_n4638) );
  AND2X2 AND2X2_3031 ( .A(core__abc_21380_n4640), .B(core__abc_21380_n2236), .Y(core__abc_21380_n4641) );
  AND2X2 AND2X2_3032 ( .A(core__abc_21380_n4639_1), .B(core__abc_21380_n2230), .Y(core__abc_21380_n4642) );
  AND2X2 AND2X2_3033 ( .A(core__abc_21380_n4394), .B(core__abc_21380_n3073_1), .Y(core__abc_21380_n4645) );
  AND2X2 AND2X2_3034 ( .A(core__abc_21380_n4646), .B(core__abc_21380_n1637), .Y(core__abc_21380_n4647) );
  AND2X2 AND2X2_3035 ( .A(core__abc_21380_n4648), .B(core__abc_21380_n1639), .Y(core__abc_21380_n4649) );
  AND2X2 AND2X2_3036 ( .A(core__abc_21380_n4652), .B(core__abc_21380_n4653), .Y(core__abc_21380_n4654) );
  AND2X2 AND2X2_3037 ( .A(core__abc_21380_n4655_1), .B(core__abc_21380_n4644_1), .Y(core__abc_21380_n4656) );
  AND2X2 AND2X2_3038 ( .A(core__abc_21380_n4654), .B(core__abc_21380_n4643), .Y(core__abc_21380_n4657) );
  AND2X2 AND2X2_3039 ( .A(core__abc_21380_n4659), .B(core__abc_21380_n4586), .Y(core__abc_21380_n4660_1) );
  AND2X2 AND2X2_304 ( .A(_abc_19068_n897_1_bF_buf1), .B(word0_reg_22_), .Y(_abc_19068_n1427) );
  AND2X2 AND2X2_3040 ( .A(core__abc_21380_n4609), .B(core__abc_21380_n4543), .Y(core__abc_21380_n4663) );
  AND2X2 AND2X2_3041 ( .A(core__abc_21380_n4663), .B(core__abc_21380_n4515), .Y(core__abc_21380_n4664) );
  AND2X2 AND2X2_3042 ( .A(core__abc_21380_n4663), .B(core__abc_21380_n4516_1), .Y(core__abc_21380_n4667) );
  AND2X2 AND2X2_3043 ( .A(core__abc_21380_n4669), .B(core__abc_21380_n4666_1), .Y(core__abc_21380_n4670) );
  AND2X2 AND2X2_3044 ( .A(core__abc_21380_n4670), .B(core__abc_21380_n4658), .Y(core__abc_21380_n4671_1) );
  AND2X2 AND2X2_3045 ( .A(core__abc_21380_n4677), .B(core__abc_21380_n2440), .Y(core__abc_21380_n4678) );
  AND2X2 AND2X2_3046 ( .A(core__abc_21380_n4676_1), .B(core__abc_21380_n2439), .Y(core__abc_21380_n4679) );
  AND2X2 AND2X2_3047 ( .A(core__abc_21380_n4680), .B(core__abc_21380_n4675), .Y(core__abc_21380_n4681_1) );
  AND2X2 AND2X2_3048 ( .A(core__abc_21380_n4682), .B(core_v3_reg_47_), .Y(core__abc_21380_n4683) );
  AND2X2 AND2X2_3049 ( .A(core__abc_21380_n4687), .B(core__abc_21380_n4688), .Y(core__abc_21380_n4689) );
  AND2X2 AND2X2_305 ( .A(_abc_19068_n915_1_bF_buf1), .B(core_mi_54_), .Y(_abc_19068_n1428_1) );
  AND2X2 AND2X2_3050 ( .A(core__abc_21380_n4690), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n4691_1) );
  AND2X2 AND2X2_3051 ( .A(core__abc_21380_n4691_1), .B(core__abc_21380_n4685), .Y(core__abc_21380_n4692) );
  AND2X2 AND2X2_3052 ( .A(core__abc_21380_n3313_bF_buf4), .B(core__abc_21380_n4693), .Y(core__abc_21380_n4694) );
  AND2X2 AND2X2_3053 ( .A(core_v3_reg_20_), .B(core_mi_20_), .Y(core__abc_21380_n4696_1) );
  AND2X2 AND2X2_3054 ( .A(core__abc_21380_n4697), .B(core__abc_21380_n4695), .Y(core__abc_21380_n4698) );
  AND2X2 AND2X2_3055 ( .A(core__abc_21380_n2749_bF_buf2), .B(core__abc_21380_n4698), .Y(core__abc_21380_n4699) );
  AND2X2 AND2X2_3056 ( .A(core__abc_21380_n4703), .B(reset_n_bF_buf44), .Y(core__abc_21380_n4704) );
  AND2X2 AND2X2_3057 ( .A(core__abc_21380_n4702), .B(core__abc_21380_n4704), .Y(core_v3_reg_20__FF_INPUT) );
  AND2X2 AND2X2_3058 ( .A(core__abc_21380_n4707_1), .B(core__abc_21380_n2251), .Y(core__abc_21380_n4708) );
  AND2X2 AND2X2_3059 ( .A(core__abc_21380_n4706), .B(core__abc_21380_n2250), .Y(core__abc_21380_n4709) );
  AND2X2 AND2X2_306 ( .A(_abc_19068_n923_bF_buf2), .B(_abc_19068_n1432_1), .Y(_auto_iopadmap_cc_313_execute_30317_22_) );
  AND2X2 AND2X2_3060 ( .A(core__abc_21380_n4713), .B(core__abc_21380_n1657), .Y(core__abc_21380_n4714) );
  AND2X2 AND2X2_3061 ( .A(core__abc_21380_n4712_1), .B(core__abc_21380_n1655_1), .Y(core__abc_21380_n4715) );
  AND2X2 AND2X2_3062 ( .A(core__abc_21380_n4716), .B(core__abc_21380_n1362), .Y(core__abc_21380_n4717_1) );
  AND2X2 AND2X2_3063 ( .A(core__abc_21380_n4718), .B(core_v3_reg_5_), .Y(core__abc_21380_n4719) );
  AND2X2 AND2X2_3064 ( .A(core__abc_21380_n4721), .B(core__abc_21380_n4711), .Y(core__abc_21380_n4722_1) );
  AND2X2 AND2X2_3065 ( .A(core__abc_21380_n4720), .B(core__abc_21380_n4710), .Y(core__abc_21380_n4723) );
  AND2X2 AND2X2_3066 ( .A(core__abc_21380_n4672), .B(core__abc_21380_n4725), .Y(core__abc_21380_n4726) );
  AND2X2 AND2X2_3067 ( .A(core__abc_21380_n4726), .B(core__abc_21380_n4724), .Y(core__abc_21380_n4727_1) );
  AND2X2 AND2X2_3068 ( .A(core__abc_21380_n4733), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n4734) );
  AND2X2 AND2X2_3069 ( .A(core__abc_21380_n4734), .B(core__abc_21380_n4732_1), .Y(core__abc_21380_n4735) );
  AND2X2 AND2X2_307 ( .A(_abc_19068_n916_1_bF_buf0), .B(word1_reg_23_), .Y(_abc_19068_n1434_1) );
  AND2X2 AND2X2_3070 ( .A(core__abc_21380_n3313_bF_buf3), .B(core__abc_21380_n4736), .Y(core__abc_21380_n4737_1) );
  AND2X2 AND2X2_3071 ( .A(core_v3_reg_21_), .B(core_mi_21_), .Y(core__abc_21380_n4739) );
  AND2X2 AND2X2_3072 ( .A(core__abc_21380_n4740), .B(core__abc_21380_n4738), .Y(core__abc_21380_n4741) );
  AND2X2 AND2X2_3073 ( .A(core__abc_21380_n2749_bF_buf1), .B(core__abc_21380_n4741), .Y(core__abc_21380_n4742_1) );
  AND2X2 AND2X2_3074 ( .A(core__abc_21380_n4746), .B(reset_n_bF_buf43), .Y(core__abc_21380_n4747_1) );
  AND2X2 AND2X2_3075 ( .A(core__abc_21380_n4745), .B(core__abc_21380_n4747_1), .Y(core_v3_reg_21__FF_INPUT) );
  AND2X2 AND2X2_3076 ( .A(core__abc_21380_n4751), .B(core__abc_21380_n4725), .Y(core__abc_21380_n4752_1) );
  AND2X2 AND2X2_3077 ( .A(core__abc_21380_n4750), .B(core__abc_21380_n4753), .Y(core__abc_21380_n4754) );
  AND2X2 AND2X2_3078 ( .A(core__abc_21380_n2229), .B(core__abc_21380_n2245), .Y(core__abc_21380_n4755) );
  AND2X2 AND2X2_3079 ( .A(core__abc_21380_n2250), .B(core__abc_21380_n2230), .Y(core__abc_21380_n4758) );
  AND2X2 AND2X2_308 ( .A(_abc_19068_n897_1_bF_buf0), .B(word0_reg_23_), .Y(_abc_19068_n1435) );
  AND2X2 AND2X2_3080 ( .A(core__abc_21380_n4639_1), .B(core__abc_21380_n4758), .Y(core__abc_21380_n4759) );
  AND2X2 AND2X2_3081 ( .A(core__abc_21380_n4761), .B(core__abc_21380_n2268), .Y(core__abc_21380_n4762_1) );
  AND2X2 AND2X2_3082 ( .A(core__abc_21380_n4760), .B(core__abc_21380_n2269), .Y(core__abc_21380_n4763) );
  AND2X2 AND2X2_3083 ( .A(core__abc_21380_n4646), .B(core__abc_21380_n3069), .Y(core__abc_21380_n4766) );
  AND2X2 AND2X2_3084 ( .A(core__abc_21380_n4768), .B(core__abc_21380_n1675), .Y(core__abc_21380_n4769) );
  AND2X2 AND2X2_3085 ( .A(core__abc_21380_n4767_1), .B(core__abc_21380_n1673), .Y(core__abc_21380_n4770) );
  AND2X2 AND2X2_3086 ( .A(core__abc_21380_n4773), .B(core__abc_21380_n4774), .Y(core__abc_21380_n4775) );
  AND2X2 AND2X2_3087 ( .A(core__abc_21380_n4776), .B(core__abc_21380_n4765), .Y(core__abc_21380_n4777_1) );
  AND2X2 AND2X2_3088 ( .A(core__abc_21380_n4775), .B(core__abc_21380_n4764), .Y(core__abc_21380_n4778) );
  AND2X2 AND2X2_3089 ( .A(core__abc_21380_n4754), .B(core__abc_21380_n4779), .Y(core__abc_21380_n4780) );
  AND2X2 AND2X2_309 ( .A(_abc_19068_n941_bF_buf1), .B(core_key_119_), .Y(_abc_19068_n1437) );
  AND2X2 AND2X2_3090 ( .A(core__abc_21380_n4786), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n4787) );
  AND2X2 AND2X2_3091 ( .A(core__abc_21380_n4787), .B(core__abc_21380_n4785), .Y(core__abc_21380_n4788_1) );
  AND2X2 AND2X2_3092 ( .A(core__abc_21380_n3313_bF_buf2), .B(core__abc_21380_n4789), .Y(core__abc_21380_n4790) );
  AND2X2 AND2X2_3093 ( .A(core_v3_reg_22_), .B(core_mi_22_), .Y(core__abc_21380_n4792) );
  AND2X2 AND2X2_3094 ( .A(core__abc_21380_n4793_1), .B(core__abc_21380_n4791), .Y(core__abc_21380_n4794) );
  AND2X2 AND2X2_3095 ( .A(core__abc_21380_n2749_bF_buf0), .B(core__abc_21380_n4794), .Y(core__abc_21380_n4795) );
  AND2X2 AND2X2_3096 ( .A(core__abc_21380_n4799), .B(reset_n_bF_buf42), .Y(core__abc_21380_n4800) );
  AND2X2 AND2X2_3097 ( .A(core__abc_21380_n4798_1), .B(core__abc_21380_n4800), .Y(core_v3_reg_22__FF_INPUT) );
  AND2X2 AND2X2_3098 ( .A(core__abc_21380_n4781), .B(core__abc_21380_n4802), .Y(core__abc_21380_n4803_1) );
  AND2X2 AND2X2_3099 ( .A(core__abc_21380_n4806), .B(core__abc_21380_n2294_1), .Y(core__abc_21380_n4807) );
  AND2X2 AND2X2_31 ( .A(_abc_19068_n907_1), .B(_abc_19068_n896), .Y(_abc_19068_n916_1) );
  AND2X2 AND2X2_310 ( .A(_abc_19068_n924_1_bF_buf1), .B(core_key_55_), .Y(_abc_19068_n1438_1) );
  AND2X2 AND2X2_3100 ( .A(core__abc_21380_n4805), .B(core__abc_21380_n2288), .Y(core__abc_21380_n4808_1) );
  AND2X2 AND2X2_3101 ( .A(core__abc_21380_n4811), .B(core__abc_21380_n1695), .Y(core__abc_21380_n4812) );
  AND2X2 AND2X2_3102 ( .A(core__abc_21380_n4810), .B(core__abc_21380_n1692), .Y(core__abc_21380_n4813) );
  AND2X2 AND2X2_3103 ( .A(core__abc_21380_n4814_1), .B(core__abc_21380_n1399), .Y(core__abc_21380_n4815) );
  AND2X2 AND2X2_3104 ( .A(core__abc_21380_n4820_1), .B(core__abc_21380_n4821), .Y(core__abc_21380_n4822) );
  AND2X2 AND2X2_3105 ( .A(core__abc_21380_n4823), .B(core__abc_21380_n4816), .Y(core__abc_21380_n4824) );
  AND2X2 AND2X2_3106 ( .A(core__abc_21380_n4825_1), .B(core__abc_21380_n4819), .Y(core__abc_21380_n4826) );
  AND2X2 AND2X2_3107 ( .A(core__abc_21380_n4822), .B(core__abc_21380_n4824), .Y(core__abc_21380_n4828) );
  AND2X2 AND2X2_3108 ( .A(core__abc_21380_n4818), .B(core__abc_21380_n4809), .Y(core__abc_21380_n4829) );
  AND2X2 AND2X2_3109 ( .A(core__abc_21380_n4827), .B(core__abc_21380_n4831), .Y(core__abc_21380_n4832) );
  AND2X2 AND2X2_311 ( .A(_abc_19068_n926_bF_buf1), .B(core_key_23_), .Y(_abc_19068_n1439) );
  AND2X2 AND2X2_3110 ( .A(core__abc_21380_n4835_1), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n4836) );
  AND2X2 AND2X2_3111 ( .A(core__abc_21380_n4836), .B(core__abc_21380_n4833), .Y(core__abc_21380_n4837) );
  AND2X2 AND2X2_3112 ( .A(core__abc_21380_n3313_bF_buf1), .B(core_key_87_), .Y(core__abc_21380_n4838) );
  AND2X2 AND2X2_3113 ( .A(core_v3_reg_23_), .B(core_mi_23_), .Y(core__abc_21380_n4840_1) );
  AND2X2 AND2X2_3114 ( .A(core__abc_21380_n4841), .B(core__abc_21380_n4839), .Y(core__abc_21380_n4842) );
  AND2X2 AND2X2_3115 ( .A(core__abc_21380_n2749_bF_buf10), .B(core__abc_21380_n4842), .Y(core__abc_21380_n4843) );
  AND2X2 AND2X2_3116 ( .A(core__abc_21380_n4847), .B(reset_n_bF_buf41), .Y(core__abc_21380_n4848) );
  AND2X2 AND2X2_3117 ( .A(core__abc_21380_n4846), .B(core__abc_21380_n4848), .Y(core_v3_reg_23__FF_INPUT) );
  AND2X2 AND2X2_3118 ( .A(core__abc_21380_n4826), .B(core__abc_21380_n4851_1), .Y(core__abc_21380_n4852) );
  AND2X2 AND2X2_3119 ( .A(core__abc_21380_n4852), .B(core__abc_21380_n4850), .Y(core__abc_21380_n4853) );
  AND2X2 AND2X2_312 ( .A(_abc_19068_n939_1_bF_buf1), .B(core_key_87_), .Y(_abc_19068_n1443) );
  AND2X2 AND2X2_3120 ( .A(core__abc_21380_n4853), .B(core__abc_21380_n4667), .Y(core__abc_21380_n4854) );
  AND2X2 AND2X2_3121 ( .A(core__abc_21380_n4825_1), .B(core__abc_21380_n4777_1), .Y(core__abc_21380_n4861) );
  AND2X2 AND2X2_3122 ( .A(core__abc_21380_n4860), .B(core__abc_21380_n4863), .Y(core__abc_21380_n4864) );
  AND2X2 AND2X2_3123 ( .A(core__abc_21380_n4859), .B(core__abc_21380_n4864), .Y(core__abc_21380_n4865) );
  AND2X2 AND2X2_3124 ( .A(core__abc_21380_n4856), .B(core__abc_21380_n4865), .Y(core__abc_21380_n4866) );
  AND2X2 AND2X2_3125 ( .A(core__abc_21380_n2269), .B(core__abc_21380_n2288), .Y(core__abc_21380_n4868) );
  AND2X2 AND2X2_3126 ( .A(core__abc_21380_n4868), .B(core__abc_21380_n4758), .Y(core__abc_21380_n4869) );
  AND2X2 AND2X2_3127 ( .A(core__abc_21380_n4637), .B(core__abc_21380_n4869), .Y(core__abc_21380_n4870) );
  AND2X2 AND2X2_3128 ( .A(core__abc_21380_n4636), .B(core__abc_21380_n4869), .Y(core__abc_21380_n4873_1) );
  AND2X2 AND2X2_3129 ( .A(core__abc_21380_n4757_1), .B(core__abc_21380_n4868), .Y(core__abc_21380_n4874) );
  AND2X2 AND2X2_313 ( .A(_abc_19068_n902_bF_buf0), .B(word2_reg_23_), .Y(_abc_19068_n1444_1) );
  AND2X2 AND2X2_3130 ( .A(core__abc_21380_n2285), .B(core__abc_21380_n2267), .Y(core__abc_21380_n4875) );
  AND2X2 AND2X2_3131 ( .A(core__abc_21380_n4872), .B(core__abc_21380_n4879), .Y(core__abc_21380_n4880) );
  AND2X2 AND2X2_3132 ( .A(core__abc_21380_n4880), .B(core__abc_21380_n2306), .Y(core__abc_21380_n4881) );
  AND2X2 AND2X2_3133 ( .A(core__abc_21380_n4384), .B(core__abc_21380_n4870), .Y(core__abc_21380_n4882) );
  AND2X2 AND2X2_3134 ( .A(core__abc_21380_n4883_1), .B(core__abc_21380_n2307), .Y(core__abc_21380_n4884) );
  AND2X2 AND2X2_3135 ( .A(core__abc_21380_n4890), .B(core__abc_21380_n4888_1), .Y(core__abc_21380_n4891) );
  AND2X2 AND2X2_3136 ( .A(core__abc_21380_n4891), .B(core__abc_21380_n1713), .Y(core__abc_21380_n4892_1) );
  AND2X2 AND2X2_3137 ( .A(core__abc_21380_n4893_1), .B(core__abc_21380_n1711), .Y(core__abc_21380_n4894) );
  AND2X2 AND2X2_3138 ( .A(core__abc_21380_n4897), .B(core__abc_21380_n4898_1), .Y(core__abc_21380_n4899) );
  AND2X2 AND2X2_3139 ( .A(core__abc_21380_n4900_1), .B(core__abc_21380_n4886), .Y(core__abc_21380_n4901) );
  AND2X2 AND2X2_314 ( .A(_abc_19068_n899_bF_buf0), .B(word3_reg_23_), .Y(_abc_19068_n1445) );
  AND2X2 AND2X2_3140 ( .A(core__abc_21380_n4899), .B(core__abc_21380_n4885), .Y(core__abc_21380_n4902_1) );
  AND2X2 AND2X2_3141 ( .A(core__abc_21380_n4867_1), .B(core__abc_21380_n4904), .Y(core__abc_21380_n4905) );
  AND2X2 AND2X2_3142 ( .A(core__abc_21380_n4866), .B(core__abc_21380_n4903), .Y(core__abc_21380_n4906) );
  AND2X2 AND2X2_3143 ( .A(core__abc_21380_n4910), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n4911) );
  AND2X2 AND2X2_3144 ( .A(core__abc_21380_n4911), .B(core__abc_21380_n4909), .Y(core__abc_21380_n4912) );
  AND2X2 AND2X2_3145 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n4913), .Y(core__abc_21380_n4914) );
  AND2X2 AND2X2_3146 ( .A(core_v3_reg_24_), .B(core_mi_24_), .Y(core__abc_21380_n4916) );
  AND2X2 AND2X2_3147 ( .A(core__abc_21380_n4917), .B(core__abc_21380_n4915), .Y(core__abc_21380_n4918) );
  AND2X2 AND2X2_3148 ( .A(core__abc_21380_n2749_bF_buf9), .B(core__abc_21380_n4918), .Y(core__abc_21380_n4919) );
  AND2X2 AND2X2_3149 ( .A(core__abc_21380_n4923), .B(reset_n_bF_buf40), .Y(core__abc_21380_n4924) );
  AND2X2 AND2X2_315 ( .A(_abc_19068_n945_1_bF_buf1), .B(core_mi_23_), .Y(_abc_19068_n1447) );
  AND2X2 AND2X2_3150 ( .A(core__abc_21380_n4922), .B(core__abc_21380_n4924), .Y(core_v3_reg_24__FF_INPUT) );
  AND2X2 AND2X2_3151 ( .A(core__abc_21380_n4927), .B(core__abc_21380_n4926), .Y(core__abc_21380_n4928) );
  AND2X2 AND2X2_3152 ( .A(core__abc_21380_n2325), .B(core__abc_21380_n2305), .Y(core__abc_21380_n4929) );
  AND2X2 AND2X2_3153 ( .A(core__abc_21380_n4931), .B(core__abc_21380_n2324), .Y(core__abc_21380_n4932) );
  AND2X2 AND2X2_3154 ( .A(core__abc_21380_n2307), .B(core__abc_21380_n2325), .Y(core__abc_21380_n4933) );
  AND2X2 AND2X2_3155 ( .A(core__abc_21380_n4883_1), .B(core__abc_21380_n4933), .Y(core__abc_21380_n4934) );
  AND2X2 AND2X2_3156 ( .A(core__abc_21380_n4939), .B(core__abc_21380_n1733), .Y(core__abc_21380_n4940) );
  AND2X2 AND2X2_3157 ( .A(core__abc_21380_n4938), .B(core__abc_21380_n1730), .Y(core__abc_21380_n4941) );
  AND2X2 AND2X2_3158 ( .A(core__abc_21380_n4942), .B(core__abc_21380_n4937), .Y(core__abc_21380_n4943) );
  AND2X2 AND2X2_3159 ( .A(core__abc_21380_n4944), .B(core_v3_reg_9_), .Y(core__abc_21380_n4945) );
  AND2X2 AND2X2_316 ( .A(_abc_19068_n915_1_bF_buf0), .B(core_mi_55_), .Y(_abc_19068_n1448_1) );
  AND2X2 AND2X2_3160 ( .A(core__abc_21380_n4936), .B(core__abc_21380_n4946), .Y(core__abc_21380_n4948) );
  AND2X2 AND2X2_3161 ( .A(core__abc_21380_n4949), .B(core__abc_21380_n4947), .Y(core__abc_21380_n4950) );
  AND2X2 AND2X2_3162 ( .A(core__abc_21380_n4954), .B(core__abc_21380_n4951), .Y(core__abc_21380_n4955) );
  AND2X2 AND2X2_3163 ( .A(core__abc_21380_n4958), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n4959) );
  AND2X2 AND2X2_3164 ( .A(core__abc_21380_n4959), .B(core__abc_21380_n4957), .Y(core__abc_21380_n4960) );
  AND2X2 AND2X2_3165 ( .A(core__abc_21380_n3313_bF_buf12), .B(core_key_89_), .Y(core__abc_21380_n4961) );
  AND2X2 AND2X2_3166 ( .A(core_v3_reg_25_), .B(core_mi_25_), .Y(core__abc_21380_n4963) );
  AND2X2 AND2X2_3167 ( .A(core__abc_21380_n4964), .B(core__abc_21380_n4962), .Y(core__abc_21380_n4965) );
  AND2X2 AND2X2_3168 ( .A(core__abc_21380_n2749_bF_buf8), .B(core__abc_21380_n4965), .Y(core__abc_21380_n4966) );
  AND2X2 AND2X2_3169 ( .A(core__abc_21380_n4970), .B(reset_n_bF_buf39), .Y(core__abc_21380_n4971) );
  AND2X2 AND2X2_317 ( .A(_abc_19068_n923_bF_buf1), .B(_abc_19068_n1452_1), .Y(_auto_iopadmap_cc_313_execute_30317_23_) );
  AND2X2 AND2X2_3170 ( .A(core__abc_21380_n4969), .B(core__abc_21380_n4971), .Y(core_v3_reg_25__FF_INPUT) );
  AND2X2 AND2X2_3171 ( .A(core__abc_21380_n4974), .B(core__abc_21380_n2343), .Y(core__abc_21380_n4975) );
  AND2X2 AND2X2_3172 ( .A(core__abc_21380_n4976), .B(core__abc_21380_n2342), .Y(core__abc_21380_n4977) );
  AND2X2 AND2X2_3173 ( .A(core__abc_21380_n4893_1), .B(core__abc_21380_n3065), .Y(core__abc_21380_n4981) );
  AND2X2 AND2X2_3174 ( .A(core__abc_21380_n4983), .B(core__abc_21380_n1750), .Y(core__abc_21380_n4984) );
  AND2X2 AND2X2_3175 ( .A(core__abc_21380_n4982), .B(core__abc_21380_n1747), .Y(core__abc_21380_n4985) );
  AND2X2 AND2X2_3176 ( .A(core__abc_21380_n4988), .B(core__abc_21380_n4989), .Y(core__abc_21380_n4990) );
  AND2X2 AND2X2_3177 ( .A(core__abc_21380_n4991), .B(core__abc_21380_n4979), .Y(core__abc_21380_n4992) );
  AND2X2 AND2X2_3178 ( .A(core__abc_21380_n4990), .B(core__abc_21380_n4978), .Y(core__abc_21380_n4993) );
  AND2X2 AND2X2_3179 ( .A(core__abc_21380_n4947), .B(core__abc_21380_n4926), .Y(core__abc_21380_n4995) );
  AND2X2 AND2X2_318 ( .A(_abc_19068_n899_bF_buf4), .B(word3_reg_24_), .Y(_abc_19068_n1454_1) );
  AND2X2 AND2X2_3180 ( .A(core__abc_21380_n4950), .B(core__abc_21380_n4904), .Y(core__abc_21380_n4997) );
  AND2X2 AND2X2_3181 ( .A(core__abc_21380_n4999), .B(core__abc_21380_n4996), .Y(core__abc_21380_n5000) );
  AND2X2 AND2X2_3182 ( .A(core__abc_21380_n5000), .B(core__abc_21380_n4994), .Y(core__abc_21380_n5001) );
  AND2X2 AND2X2_3183 ( .A(core__abc_21380_n5007), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n5008) );
  AND2X2 AND2X2_3184 ( .A(core__abc_21380_n5008), .B(core__abc_21380_n5005), .Y(core__abc_21380_n5009) );
  AND2X2 AND2X2_3185 ( .A(core__abc_21380_n3313_bF_buf11), .B(core_key_90_), .Y(core__abc_21380_n5010) );
  AND2X2 AND2X2_3186 ( .A(core_v3_reg_26_), .B(core_mi_26_), .Y(core__abc_21380_n5012) );
  AND2X2 AND2X2_3187 ( .A(core__abc_21380_n5013), .B(core__abc_21380_n5011), .Y(core__abc_21380_n5014) );
  AND2X2 AND2X2_3188 ( .A(core__abc_21380_n2749_bF_buf7), .B(core__abc_21380_n5014), .Y(core__abc_21380_n5015) );
  AND2X2 AND2X2_3189 ( .A(core__abc_21380_n5019), .B(reset_n_bF_buf38), .Y(core__abc_21380_n5020) );
  AND2X2 AND2X2_319 ( .A(_abc_19068_n945_1_bF_buf0), .B(core_mi_24_), .Y(_abc_19068_n1456_1) );
  AND2X2 AND2X2_3190 ( .A(core__abc_21380_n5018), .B(core__abc_21380_n5020), .Y(core_v3_reg_26__FF_INPUT) );
  AND2X2 AND2X2_3191 ( .A(core__abc_21380_n5002), .B(core__abc_21380_n5023), .Y(core__abc_21380_n5024) );
  AND2X2 AND2X2_3192 ( .A(core__abc_21380_n5026), .B(core__abc_21380_n2368), .Y(core__abc_21380_n5027) );
  AND2X2 AND2X2_3193 ( .A(core__abc_21380_n5025), .B(core__abc_21380_n2362), .Y(core__abc_21380_n5029) );
  AND2X2 AND2X2_3194 ( .A(core__abc_21380_n5028), .B(core__abc_21380_n5030), .Y(core__abc_21380_n5031) );
  AND2X2 AND2X2_3195 ( .A(core__abc_21380_n5034), .B(core__abc_21380_n1770), .Y(core__abc_21380_n5035) );
  AND2X2 AND2X2_3196 ( .A(core__abc_21380_n5033), .B(core__abc_21380_n1767), .Y(core__abc_21380_n5036) );
  AND2X2 AND2X2_3197 ( .A(core__abc_21380_n5037), .B(core__abc_21380_n5032), .Y(core__abc_21380_n5038) );
  AND2X2 AND2X2_3198 ( .A(core__abc_21380_n5039), .B(core__abc_21380_n5040), .Y(core__abc_21380_n5041) );
  AND2X2 AND2X2_3199 ( .A(core__abc_21380_n5031), .B(core__abc_21380_n5041), .Y(core__abc_21380_n5042) );
  AND2X2 AND2X2_32 ( .A(_abc_19068_n921_1), .B(cs), .Y(_abc_19068_n922_1) );
  AND2X2 AND2X2_320 ( .A(_abc_19068_n941_bF_buf0), .B(core_key_120_), .Y(_abc_19068_n1457) );
  AND2X2 AND2X2_3200 ( .A(core__abc_21380_n5045), .B(core__abc_21380_n5043), .Y(core__abc_21380_n5046) );
  AND2X2 AND2X2_3201 ( .A(core__abc_21380_n5051), .B(core__abc_21380_n5050), .Y(core__abc_21380_n5052) );
  AND2X2 AND2X2_3202 ( .A(core__abc_21380_n5053), .B(core__abc_21380_n5048), .Y(core__abc_21380_n5054) );
  AND2X2 AND2X2_3203 ( .A(core__abc_21380_n5057), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n5058) );
  AND2X2 AND2X2_3204 ( .A(core__abc_21380_n5058), .B(core__abc_21380_n5055), .Y(core__abc_21380_n5059) );
  AND2X2 AND2X2_3205 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n5060), .Y(core__abc_21380_n5061) );
  AND2X2 AND2X2_3206 ( .A(core_v3_reg_27_), .B(core_mi_27_), .Y(core__abc_21380_n5063) );
  AND2X2 AND2X2_3207 ( .A(core__abc_21380_n5064), .B(core__abc_21380_n5062), .Y(core__abc_21380_n5065) );
  AND2X2 AND2X2_3208 ( .A(core__abc_21380_n2749_bF_buf6), .B(core__abc_21380_n5065), .Y(core__abc_21380_n5066) );
  AND2X2 AND2X2_3209 ( .A(core__abc_21380_n5070), .B(reset_n_bF_buf37), .Y(core__abc_21380_n5071) );
  AND2X2 AND2X2_321 ( .A(_abc_19068_n939_1_bF_buf0), .B(core_key_88_), .Y(_abc_19068_n1460_1) );
  AND2X2 AND2X2_3210 ( .A(core__abc_21380_n5069), .B(core__abc_21380_n5071), .Y(core_v3_reg_27__FF_INPUT) );
  AND2X2 AND2X2_3211 ( .A(core__abc_21380_n5052), .B(core__abc_21380_n5074), .Y(core__abc_21380_n5075) );
  AND2X2 AND2X2_3212 ( .A(core__abc_21380_n5075), .B(core__abc_21380_n5073), .Y(core__abc_21380_n5076) );
  AND2X2 AND2X2_3213 ( .A(core__abc_21380_n5051), .B(core__abc_21380_n4992), .Y(core__abc_21380_n5077) );
  AND2X2 AND2X2_3214 ( .A(core__abc_21380_n5075), .B(core__abc_21380_n4997), .Y(core__abc_21380_n5080) );
  AND2X2 AND2X2_3215 ( .A(core__abc_21380_n4867_1), .B(core__abc_21380_n5080), .Y(core__abc_21380_n5081) );
  AND2X2 AND2X2_3216 ( .A(core__abc_21380_n2343), .B(core__abc_21380_n2362), .Y(core__abc_21380_n5084) );
  AND2X2 AND2X2_3217 ( .A(core__abc_21380_n4933), .B(core__abc_21380_n5084), .Y(core__abc_21380_n5085) );
  AND2X2 AND2X2_3218 ( .A(core__abc_21380_n4883_1), .B(core__abc_21380_n5085), .Y(core__abc_21380_n5086) );
  AND2X2 AND2X2_3219 ( .A(core__abc_21380_n4973), .B(core__abc_21380_n5084), .Y(core__abc_21380_n5087) );
  AND2X2 AND2X2_322 ( .A(_abc_19068_n924_1_bF_buf0), .B(core_key_56_), .Y(_abc_19068_n1461) );
  AND2X2 AND2X2_3220 ( .A(core__abc_21380_n2359), .B(core__abc_21380_n2341), .Y(core__abc_21380_n5088) );
  AND2X2 AND2X2_3221 ( .A(core__abc_21380_n5091), .B(core__abc_21380_n2381), .Y(core__abc_21380_n5092) );
  AND2X2 AND2X2_3222 ( .A(core__abc_21380_n5094), .B(core__abc_21380_n5095), .Y(core__abc_21380_n5096) );
  AND2X2 AND2X2_3223 ( .A(core__abc_21380_n5096), .B(core__abc_21380_n2380), .Y(core__abc_21380_n5097) );
  AND2X2 AND2X2_3224 ( .A(core__abc_21380_n5103), .B(core__abc_21380_n5101), .Y(core__abc_21380_n5104) );
  AND2X2 AND2X2_3225 ( .A(core__abc_21380_n5105), .B(core__abc_21380_n1786_1), .Y(core__abc_21380_n5106) );
  AND2X2 AND2X2_3226 ( .A(core__abc_21380_n5104), .B(core__abc_21380_n1788), .Y(core__abc_21380_n5107) );
  AND2X2 AND2X2_3227 ( .A(core__abc_21380_n5110), .B(core__abc_21380_n5111), .Y(core__abc_21380_n5112) );
  AND2X2 AND2X2_3228 ( .A(core__abc_21380_n5113), .B(core__abc_21380_n5099), .Y(core__abc_21380_n5114) );
  AND2X2 AND2X2_3229 ( .A(core__abc_21380_n5112), .B(core__abc_21380_n5098), .Y(core__abc_21380_n5115) );
  AND2X2 AND2X2_323 ( .A(_abc_19068_n926_bF_buf0), .B(core_key_24_), .Y(_abc_19068_n1462_1) );
  AND2X2 AND2X2_3230 ( .A(core__abc_21380_n5083), .B(core__abc_21380_n5116), .Y(core__abc_21380_n5117) );
  AND2X2 AND2X2_3231 ( .A(core__abc_21380_n5082), .B(core__abc_21380_n5118), .Y(core__abc_21380_n5119) );
  AND2X2 AND2X2_3232 ( .A(core__abc_21380_n5123), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n5124) );
  AND2X2 AND2X2_3233 ( .A(core__abc_21380_n5124), .B(core__abc_21380_n5121), .Y(core__abc_21380_n5125) );
  AND2X2 AND2X2_3234 ( .A(core__abc_21380_n3313_bF_buf9), .B(core__abc_21380_n5126), .Y(core__abc_21380_n5127) );
  AND2X2 AND2X2_3235 ( .A(core_v3_reg_28_), .B(core_mi_28_), .Y(core__abc_21380_n5129) );
  AND2X2 AND2X2_3236 ( .A(core__abc_21380_n5130), .B(core__abc_21380_n5128), .Y(core__abc_21380_n5131) );
  AND2X2 AND2X2_3237 ( .A(core__abc_21380_n2749_bF_buf5), .B(core__abc_21380_n5131), .Y(core__abc_21380_n5132) );
  AND2X2 AND2X2_3238 ( .A(core__abc_21380_n5136), .B(reset_n_bF_buf36), .Y(core__abc_21380_n5137) );
  AND2X2 AND2X2_3239 ( .A(core__abc_21380_n5135), .B(core__abc_21380_n5137), .Y(core_v3_reg_28__FF_INPUT) );
  AND2X2 AND2X2_324 ( .A(_abc_19068_n916_1_bF_buf4), .B(word1_reg_24_), .Y(_abc_19068_n1465) );
  AND2X2 AND2X2_3240 ( .A(core__abc_21380_n2399), .B(core__abc_21380_n2379), .Y(core__abc_21380_n5141) );
  AND2X2 AND2X2_3241 ( .A(core__abc_21380_n2381), .B(core__abc_21380_n2399), .Y(core__abc_21380_n5142) );
  AND2X2 AND2X2_3242 ( .A(core__abc_21380_n5091), .B(core__abc_21380_n5142), .Y(core__abc_21380_n5143) );
  AND2X2 AND2X2_3243 ( .A(core__abc_21380_n5152), .B(core__abc_21380_n1808), .Y(core__abc_21380_n5153) );
  AND2X2 AND2X2_3244 ( .A(core__abc_21380_n5151), .B(core__abc_21380_n1805), .Y(core__abc_21380_n5154) );
  AND2X2 AND2X2_3245 ( .A(core__abc_21380_n5155), .B(core__abc_21380_n5150), .Y(core__abc_21380_n5156) );
  AND2X2 AND2X2_3246 ( .A(core__abc_21380_n5157), .B(core__abc_21380_n5158), .Y(core__abc_21380_n5159) );
  AND2X2 AND2X2_3247 ( .A(core__abc_21380_n5159), .B(core__abc_21380_n5149), .Y(core__abc_21380_n5160) );
  AND2X2 AND2X2_3248 ( .A(core__abc_21380_n5162), .B(core__abc_21380_n5148), .Y(core__abc_21380_n5163) );
  AND2X2 AND2X2_3249 ( .A(core__abc_21380_n5164), .B(core__abc_21380_n5140), .Y(core__abc_21380_n5165) );
  AND2X2 AND2X2_325 ( .A(_abc_19068_n902_bF_buf4), .B(word2_reg_24_), .Y(_abc_19068_n1466_1) );
  AND2X2 AND2X2_3250 ( .A(core__abc_21380_n5139), .B(core__abc_21380_n5165), .Y(core__abc_21380_n5166) );
  AND2X2 AND2X2_3251 ( .A(core__abc_21380_n5169), .B(core__abc_21380_n5170), .Y(core__abc_21380_n5171) );
  AND2X2 AND2X2_3252 ( .A(core__abc_21380_n5171), .B(core__abc_21380_n5118), .Y(core__abc_21380_n5172) );
  AND2X2 AND2X2_3253 ( .A(core__abc_21380_n5082), .B(core__abc_21380_n5172), .Y(core__abc_21380_n5173) );
  AND2X2 AND2X2_3254 ( .A(core__abc_21380_n5174), .B(core__abc_21380_n5168), .Y(core__abc_21380_n5175) );
  AND2X2 AND2X2_3255 ( .A(core__abc_21380_n5167), .B(core__abc_21380_n5175), .Y(core__abc_21380_n5176) );
  AND2X2 AND2X2_3256 ( .A(core__abc_21380_n5179), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf1), .Y(core__abc_21380_n5180) );
  AND2X2 AND2X2_3257 ( .A(core__abc_21380_n5180), .B(core__abc_21380_n5177), .Y(core__abc_21380_n5181) );
  AND2X2 AND2X2_3258 ( .A(core__abc_21380_n3313_bF_buf8), .B(core__abc_21380_n5182), .Y(core__abc_21380_n5183) );
  AND2X2 AND2X2_3259 ( .A(core_v3_reg_29_), .B(core_mi_29_), .Y(core__abc_21380_n5185) );
  AND2X2 AND2X2_326 ( .A(_abc_19068_n897_1_bF_buf4), .B(word0_reg_24_), .Y(_abc_19068_n1468_1) );
  AND2X2 AND2X2_3260 ( .A(core__abc_21380_n5186), .B(core__abc_21380_n5184), .Y(core__abc_21380_n5187) );
  AND2X2 AND2X2_3261 ( .A(core__abc_21380_n2749_bF_buf4), .B(core__abc_21380_n5187), .Y(core__abc_21380_n5188) );
  AND2X2 AND2X2_3262 ( .A(core__abc_21380_n5192), .B(reset_n_bF_buf35), .Y(core__abc_21380_n5193) );
  AND2X2 AND2X2_3263 ( .A(core__abc_21380_n5191), .B(core__abc_21380_n5193), .Y(core_v3_reg_29__FF_INPUT) );
  AND2X2 AND2X2_3264 ( .A(core__abc_21380_n5168), .B(core__abc_21380_n5169), .Y(core__abc_21380_n5196) );
  AND2X2 AND2X2_3265 ( .A(core__abc_21380_n5174), .B(core__abc_21380_n5196), .Y(core__abc_21380_n5197) );
  AND2X2 AND2X2_3266 ( .A(core__abc_21380_n5199), .B(core__abc_21380_n5201), .Y(core__abc_21380_n5202) );
  AND2X2 AND2X2_3267 ( .A(core__abc_21380_n5202), .B(core__abc_21380_n2416), .Y(core__abc_21380_n5203) );
  AND2X2 AND2X2_3268 ( .A(core__abc_21380_n5204), .B(core__abc_21380_n2417), .Y(core__abc_21380_n5205) );
  AND2X2 AND2X2_3269 ( .A(core__abc_21380_n5209), .B(core__abc_21380_n3108), .Y(core__abc_21380_n5210) );
  AND2X2 AND2X2_327 ( .A(_abc_19068_n915_1_bF_buf4), .B(core_mi_56_), .Y(_abc_19068_n1469) );
  AND2X2 AND2X2_3270 ( .A(core__abc_21380_n5210), .B(core__abc_21380_n1826), .Y(core__abc_21380_n5211) );
  AND2X2 AND2X2_3271 ( .A(core__abc_21380_n5216), .B(core__abc_21380_n5218), .Y(core__abc_21380_n5219) );
  AND2X2 AND2X2_3272 ( .A(core__abc_21380_n5207), .B(core__abc_21380_n5219), .Y(core__abc_21380_n5220) );
  AND2X2 AND2X2_3273 ( .A(core__abc_21380_n5221), .B(core__abc_21380_n5206), .Y(core__abc_21380_n5222) );
  AND2X2 AND2X2_3274 ( .A(core__abc_21380_n5197), .B(core__abc_21380_n5223), .Y(core__abc_21380_n5224) );
  AND2X2 AND2X2_3275 ( .A(core__abc_21380_n5230), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf1), .Y(core__abc_21380_n5231) );
  AND2X2 AND2X2_3276 ( .A(core__abc_21380_n5231), .B(core__abc_21380_n5229), .Y(core__abc_21380_n5232) );
  AND2X2 AND2X2_3277 ( .A(core__abc_21380_n3313_bF_buf7), .B(core__abc_21380_n5233), .Y(core__abc_21380_n5234) );
  AND2X2 AND2X2_3278 ( .A(core_v3_reg_30_), .B(core_mi_30_), .Y(core__abc_21380_n5236) );
  AND2X2 AND2X2_3279 ( .A(core__abc_21380_n5237), .B(core__abc_21380_n5235), .Y(core__abc_21380_n5238) );
  AND2X2 AND2X2_328 ( .A(_abc_19068_n923_bF_buf0), .B(_abc_19068_n1473), .Y(_auto_iopadmap_cc_313_execute_30317_24_) );
  AND2X2 AND2X2_3280 ( .A(core__abc_21380_n2749_bF_buf3), .B(core__abc_21380_n5238), .Y(core__abc_21380_n5239) );
  AND2X2 AND2X2_3281 ( .A(core__abc_21380_n5243), .B(reset_n_bF_buf34), .Y(core__abc_21380_n5244) );
  AND2X2 AND2X2_3282 ( .A(core__abc_21380_n5242), .B(core__abc_21380_n5244), .Y(core_v3_reg_30__FF_INPUT) );
  AND2X2 AND2X2_3283 ( .A(core__abc_21380_n5225), .B(core__abc_21380_n5246), .Y(core__abc_21380_n5247) );
  AND2X2 AND2X2_3284 ( .A(core__abc_21380_n5250), .B(core__abc_21380_n5249), .Y(core__abc_21380_n5251) );
  AND2X2 AND2X2_3285 ( .A(core__abc_21380_n5251), .B(core__abc_21380_n2434), .Y(core__abc_21380_n5252) );
  AND2X2 AND2X2_3286 ( .A(core__abc_21380_n5253), .B(core__abc_21380_n2435), .Y(core__abc_21380_n5254) );
  AND2X2 AND2X2_3287 ( .A(core__abc_21380_n5212), .B(core__abc_21380_n1822), .Y(core__abc_21380_n5257) );
  AND2X2 AND2X2_3288 ( .A(core__abc_21380_n5257), .B(core__abc_21380_n1846_1), .Y(core__abc_21380_n5258) );
  AND2X2 AND2X2_3289 ( .A(core__abc_21380_n5261), .B(core__abc_21380_n5256), .Y(core__abc_21380_n5262) );
  AND2X2 AND2X2_329 ( .A(_abc_19068_n899_bF_buf3), .B(word3_reg_25_), .Y(_abc_19068_n1475) );
  AND2X2 AND2X2_3290 ( .A(core__abc_21380_n5263), .B(core__abc_21380_n5259), .Y(core__abc_21380_n5264) );
  AND2X2 AND2X2_3291 ( .A(core__abc_21380_n5264), .B(core_v3_reg_15_), .Y(core__abc_21380_n5265) );
  AND2X2 AND2X2_3292 ( .A(core__abc_21380_n5269), .B(core__abc_21380_n5268), .Y(core__abc_21380_n5270) );
  AND2X2 AND2X2_3293 ( .A(core__abc_21380_n5272), .B(core__abc_21380_n5271), .Y(core__abc_21380_n5273) );
  AND2X2 AND2X2_3294 ( .A(core__abc_21380_n5267), .B(core__abc_21380_n5274), .Y(core__abc_21380_n5275) );
  AND2X2 AND2X2_3295 ( .A(core__abc_21380_n5277), .B(core__abc_21380_n5278), .Y(core__abc_21380_n5279) );
  AND2X2 AND2X2_3296 ( .A(core__abc_21380_n5276), .B(core__abc_21380_n5280), .Y(core__abc_21380_n5281) );
  AND2X2 AND2X2_3297 ( .A(core__abc_21380_n5284), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n5285) );
  AND2X2 AND2X2_3298 ( .A(core__abc_21380_n5285), .B(core__abc_21380_n5282), .Y(core__abc_21380_n5286) );
  AND2X2 AND2X2_3299 ( .A(core__abc_21380_n3313_bF_buf6), .B(core_key_95_), .Y(core__abc_21380_n5287) );
  AND2X2 AND2X2_33 ( .A(_abc_19068_n920), .B(_abc_19068_n922_1), .Y(_abc_19068_n923) );
  AND2X2 AND2X2_330 ( .A(_abc_19068_n945_1_bF_buf4), .B(core_mi_25_), .Y(_abc_19068_n1477) );
  AND2X2 AND2X2_3300 ( .A(core_v3_reg_31_), .B(core_mi_31_), .Y(core__abc_21380_n5289) );
  AND2X2 AND2X2_3301 ( .A(core__abc_21380_n5290), .B(core__abc_21380_n5288), .Y(core__abc_21380_n5291) );
  AND2X2 AND2X2_3302 ( .A(core__abc_21380_n2749_bF_buf2), .B(core__abc_21380_n5291), .Y(core__abc_21380_n5292) );
  AND2X2 AND2X2_3303 ( .A(core__abc_21380_n5296), .B(reset_n_bF_buf33), .Y(core__abc_21380_n5297) );
  AND2X2 AND2X2_3304 ( .A(core__abc_21380_n5295), .B(core__abc_21380_n5297), .Y(core_v3_reg_31__FF_INPUT) );
  AND2X2 AND2X2_3305 ( .A(core__abc_21380_n5307), .B(core__abc_21380_n5308), .Y(core__abc_21380_n5309) );
  AND2X2 AND2X2_3306 ( .A(core__abc_21380_n5274), .B(core__abc_21380_n5220), .Y(core__abc_21380_n5313) );
  AND2X2 AND2X2_3307 ( .A(core__abc_21380_n5311), .B(core__abc_21380_n5315), .Y(core__abc_21380_n5316) );
  AND2X2 AND2X2_3308 ( .A(core__abc_21380_n5310), .B(core__abc_21380_n5316), .Y(core__abc_21380_n5317) );
  AND2X2 AND2X2_3309 ( .A(core__abc_21380_n5305), .B(core__abc_21380_n5317), .Y(core__abc_21380_n5318) );
  AND2X2 AND2X2_331 ( .A(_abc_19068_n941_bF_buf4), .B(core_key_121_), .Y(_abc_19068_n1478_1) );
  AND2X2 AND2X2_3310 ( .A(core__abc_21380_n5304), .B(core__abc_21380_n5318), .Y(core__abc_21380_n5319) );
  AND2X2 AND2X2_3311 ( .A(core__abc_21380_n5321), .B(core__abc_21380_n1862), .Y(core__abc_21380_n5322) );
  AND2X2 AND2X2_3312 ( .A(core__abc_21380_n3115), .B(core__abc_21380_n1864), .Y(core__abc_21380_n5323) );
  AND2X2 AND2X2_3313 ( .A(core__abc_21380_n5326), .B(core__abc_21380_n5327), .Y(core__abc_21380_n5328) );
  AND2X2 AND2X2_3314 ( .A(core__abc_21380_n5329), .B(core__abc_21380_n1262_1), .Y(core__abc_21380_n5330) );
  AND2X2 AND2X2_3315 ( .A(core__abc_21380_n5328), .B(core__abc_21380_n1270_1), .Y(core__abc_21380_n5331) );
  AND2X2 AND2X2_3316 ( .A(core__abc_21380_n5319), .B(core__abc_21380_n5332), .Y(core__abc_21380_n5333) );
  AND2X2 AND2X2_3317 ( .A(core__abc_21380_n4370), .B(core__abc_21380_n4854), .Y(core__abc_21380_n5334) );
  AND2X2 AND2X2_3318 ( .A(core__abc_21380_n5275), .B(core__abc_21380_n5335), .Y(core__abc_21380_n5336) );
  AND2X2 AND2X2_3319 ( .A(core__abc_21380_n5336), .B(core__abc_21380_n5172), .Y(core__abc_21380_n5337) );
  AND2X2 AND2X2_332 ( .A(_abc_19068_n939_1_bF_buf4), .B(core_key_89_), .Y(_abc_19068_n1481) );
  AND2X2 AND2X2_3320 ( .A(core__abc_21380_n5337), .B(core__abc_21380_n5080), .Y(core__abc_21380_n5338) );
  AND2X2 AND2X2_3321 ( .A(core__abc_21380_n5334), .B(core__abc_21380_n5338), .Y(core__abc_21380_n5339) );
  AND2X2 AND2X2_3322 ( .A(core__abc_21380_n4853), .B(core__abc_21380_n4665), .Y(core__abc_21380_n5340) );
  AND2X2 AND2X2_3323 ( .A(core__abc_21380_n4852), .B(core__abc_21380_n5341), .Y(core__abc_21380_n5342) );
  AND2X2 AND2X2_3324 ( .A(core__abc_21380_n5344), .B(core__abc_21380_n5338), .Y(core__abc_21380_n5345) );
  AND2X2 AND2X2_3325 ( .A(core__abc_21380_n5337), .B(core__abc_21380_n5079), .Y(core__abc_21380_n5346) );
  AND2X2 AND2X2_3326 ( .A(core__abc_21380_n5171), .B(core__abc_21380_n5114), .Y(core__abc_21380_n5347) );
  AND2X2 AND2X2_3327 ( .A(core__abc_21380_n5336), .B(core__abc_21380_n5348), .Y(core__abc_21380_n5349) );
  AND2X2 AND2X2_3328 ( .A(core__abc_21380_n5353), .B(core__abc_21380_n5354), .Y(core__abc_21380_n5355) );
  AND2X2 AND2X2_3329 ( .A(core__abc_21380_n5359), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n5360) );
  AND2X2 AND2X2_333 ( .A(_abc_19068_n924_1_bF_buf4), .B(core_key_57_), .Y(_abc_19068_n1482_1) );
  AND2X2 AND2X2_3330 ( .A(core__abc_21380_n5360), .B(core__abc_21380_n5357), .Y(core__abc_21380_n5361) );
  AND2X2 AND2X2_3331 ( .A(core__abc_21380_n3313_bF_buf5), .B(core_key_96_), .Y(core__abc_21380_n5362) );
  AND2X2 AND2X2_3332 ( .A(core_v3_reg_32_), .B(core_mi_32_), .Y(core__abc_21380_n5364) );
  AND2X2 AND2X2_3333 ( .A(core__abc_21380_n5365), .B(core__abc_21380_n5363), .Y(core__abc_21380_n5366) );
  AND2X2 AND2X2_3334 ( .A(core__abc_21380_n2749_bF_buf1), .B(core__abc_21380_n5366), .Y(core__abc_21380_n5367) );
  AND2X2 AND2X2_3335 ( .A(core__abc_21380_n5371), .B(reset_n_bF_buf32), .Y(core__abc_21380_n5372) );
  AND2X2 AND2X2_3336 ( .A(core__abc_21380_n5370), .B(core__abc_21380_n5372), .Y(core_v3_reg_32__FF_INPUT) );
  AND2X2 AND2X2_3337 ( .A(core__abc_21380_n1291), .B(core__abc_21380_n1261_1), .Y(core__abc_21380_n5374) );
  AND2X2 AND2X2_3338 ( .A(core__abc_21380_n5379), .B(core__abc_21380_n1882), .Y(core__abc_21380_n5380) );
  AND2X2 AND2X2_3339 ( .A(core__abc_21380_n5378), .B(core__abc_21380_n1880), .Y(core__abc_21380_n5381) );
  AND2X2 AND2X2_334 ( .A(_abc_19068_n926_bF_buf4), .B(core_key_25_), .Y(_abc_19068_n1483) );
  AND2X2 AND2X2_3340 ( .A(core__abc_21380_n5382), .B(core__abc_21380_n5377), .Y(core__abc_21380_n5383) );
  AND2X2 AND2X2_3341 ( .A(core__abc_21380_n5384), .B(core_v3_reg_17_), .Y(core__abc_21380_n5385) );
  AND2X2 AND2X2_3342 ( .A(core__abc_21380_n5387), .B(core__abc_21380_n5376), .Y(core__abc_21380_n5388) );
  AND2X2 AND2X2_3343 ( .A(core__abc_21380_n5386), .B(core__abc_21380_n5375), .Y(core__abc_21380_n5389) );
  AND2X2 AND2X2_3344 ( .A(core__abc_21380_n5392), .B(core__abc_21380_n5391), .Y(core__abc_21380_n5393) );
  AND2X2 AND2X2_3345 ( .A(core__abc_21380_n5393), .B(core__abc_21380_n5390), .Y(core__abc_21380_n5394) );
  AND2X2 AND2X2_3346 ( .A(core__abc_21380_n5400), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n5401) );
  AND2X2 AND2X2_3347 ( .A(core__abc_21380_n5401), .B(core__abc_21380_n5399), .Y(core__abc_21380_n5402) );
  AND2X2 AND2X2_3348 ( .A(core__abc_21380_n3313_bF_buf4), .B(core__abc_21380_n5403), .Y(core__abc_21380_n5404) );
  AND2X2 AND2X2_3349 ( .A(core_v3_reg_33_), .B(core_mi_33_), .Y(core__abc_21380_n5406) );
  AND2X2 AND2X2_335 ( .A(_abc_19068_n916_1_bF_buf3), .B(word1_reg_25_), .Y(_abc_19068_n1486_1) );
  AND2X2 AND2X2_3350 ( .A(core__abc_21380_n5407), .B(core__abc_21380_n5405), .Y(core__abc_21380_n5408) );
  AND2X2 AND2X2_3351 ( .A(core__abc_21380_n2749_bF_buf0), .B(core__abc_21380_n5408), .Y(core__abc_21380_n5409) );
  AND2X2 AND2X2_3352 ( .A(core__abc_21380_n5413), .B(reset_n_bF_buf31), .Y(core__abc_21380_n5414) );
  AND2X2 AND2X2_3353 ( .A(core__abc_21380_n5412), .B(core__abc_21380_n5414), .Y(core_v3_reg_33__FF_INPUT) );
  AND2X2 AND2X2_3354 ( .A(core__abc_21380_n5416), .B(core__abc_21380_n5354), .Y(core__abc_21380_n5417) );
  AND2X2 AND2X2_3355 ( .A(core__abc_21380_n5353), .B(core__abc_21380_n5417), .Y(core__abc_21380_n5418) );
  AND2X2 AND2X2_3356 ( .A(core__abc_21380_n5416), .B(core__abc_21380_n5330), .Y(core__abc_21380_n5420) );
  AND2X2 AND2X2_3357 ( .A(core__abc_21380_n5419), .B(core__abc_21380_n5422), .Y(core__abc_21380_n5423) );
  AND2X2 AND2X2_3358 ( .A(core__abc_21380_n3169), .B(core__abc_21380_n1303), .Y(core__abc_21380_n5424) );
  AND2X2 AND2X2_3359 ( .A(core__abc_21380_n3272), .B(core__abc_21380_n1302), .Y(core__abc_21380_n5425) );
  AND2X2 AND2X2_336 ( .A(_abc_19068_n902_bF_buf3), .B(word2_reg_25_), .Y(_abc_19068_n1487) );
  AND2X2 AND2X2_3360 ( .A(core__abc_21380_n5430), .B(core__abc_21380_n3127), .Y(core__abc_21380_n5431) );
  AND2X2 AND2X2_3361 ( .A(core__abc_21380_n5431), .B(core__abc_21380_n1900), .Y(core__abc_21380_n5432) );
  AND2X2 AND2X2_3362 ( .A(core__abc_21380_n5437), .B(core__abc_21380_n5438), .Y(core__abc_21380_n5439) );
  AND2X2 AND2X2_3363 ( .A(core__abc_21380_n5440), .B(core__abc_21380_n5427), .Y(core__abc_21380_n5441) );
  AND2X2 AND2X2_3364 ( .A(core__abc_21380_n5439), .B(core__abc_21380_n5426), .Y(core__abc_21380_n5442) );
  AND2X2 AND2X2_3365 ( .A(core__abc_21380_n5423), .B(core__abc_21380_n5443), .Y(core__abc_21380_n5444) );
  AND2X2 AND2X2_3366 ( .A(core__abc_21380_n5450), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n5451) );
  AND2X2 AND2X2_3367 ( .A(core__abc_21380_n5451), .B(core__abc_21380_n5448), .Y(core__abc_21380_n5452) );
  AND2X2 AND2X2_3368 ( .A(core__abc_21380_n3313_bF_buf3), .B(core_key_98_), .Y(core__abc_21380_n5453) );
  AND2X2 AND2X2_3369 ( .A(core_v3_reg_34_), .B(core_mi_34_), .Y(core__abc_21380_n5455) );
  AND2X2 AND2X2_337 ( .A(_abc_19068_n897_1_bF_buf3), .B(word0_reg_25_), .Y(_abc_19068_n1489) );
  AND2X2 AND2X2_3370 ( .A(core__abc_21380_n5456), .B(core__abc_21380_n5454), .Y(core__abc_21380_n5457) );
  AND2X2 AND2X2_3371 ( .A(core__abc_21380_n2749_bF_buf10), .B(core__abc_21380_n5457), .Y(core__abc_21380_n5458) );
  AND2X2 AND2X2_3372 ( .A(core__abc_21380_n5462), .B(reset_n_bF_buf30), .Y(core__abc_21380_n5463) );
  AND2X2 AND2X2_3373 ( .A(core__abc_21380_n5461), .B(core__abc_21380_n5463), .Y(core_v3_reg_34__FF_INPUT) );
  AND2X2 AND2X2_3374 ( .A(core__abc_21380_n5445), .B(core__abc_21380_n5465), .Y(core__abc_21380_n5466) );
  AND2X2 AND2X2_3375 ( .A(core__abc_21380_n5469), .B(core__abc_21380_n1321), .Y(core__abc_21380_n5470) );
  AND2X2 AND2X2_3376 ( .A(core__abc_21380_n5468), .B(core__abc_21380_n1322), .Y(core__abc_21380_n5471) );
  AND2X2 AND2X2_3377 ( .A(core__abc_21380_n5433), .B(core__abc_21380_n1896), .Y(core__abc_21380_n5475) );
  AND2X2 AND2X2_3378 ( .A(core__abc_21380_n5475), .B(core__abc_21380_n1920), .Y(core__abc_21380_n5476) );
  AND2X2 AND2X2_3379 ( .A(core__abc_21380_n5477), .B(core__abc_21380_n5478), .Y(core__abc_21380_n5479) );
  AND2X2 AND2X2_338 ( .A(_abc_19068_n915_1_bF_buf3), .B(core_mi_57_), .Y(_abc_19068_n1490_1) );
  AND2X2 AND2X2_3380 ( .A(core__abc_21380_n5480), .B(core__abc_21380_n5474), .Y(core__abc_21380_n5481) );
  AND2X2 AND2X2_3381 ( .A(core__abc_21380_n5479), .B(core_v3_reg_19_), .Y(core__abc_21380_n5482) );
  AND2X2 AND2X2_3382 ( .A(core__abc_21380_n5484), .B(core__abc_21380_n5473), .Y(core__abc_21380_n5485) );
  AND2X2 AND2X2_3383 ( .A(core__abc_21380_n5483), .B(core__abc_21380_n5472), .Y(core__abc_21380_n5486) );
  AND2X2 AND2X2_3384 ( .A(core__abc_21380_n5489), .B(core__abc_21380_n5490), .Y(core__abc_21380_n5491) );
  AND2X2 AND2X2_3385 ( .A(core__abc_21380_n5494), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n5495) );
  AND2X2 AND2X2_3386 ( .A(core__abc_21380_n5495), .B(core__abc_21380_n5492), .Y(core__abc_21380_n5496) );
  AND2X2 AND2X2_3387 ( .A(core__abc_21380_n3313_bF_buf2), .B(core_key_99_), .Y(core__abc_21380_n5497) );
  AND2X2 AND2X2_3388 ( .A(core_v3_reg_35_), .B(core_mi_35_), .Y(core__abc_21380_n5499) );
  AND2X2 AND2X2_3389 ( .A(core__abc_21380_n5500), .B(core__abc_21380_n5498), .Y(core__abc_21380_n5501) );
  AND2X2 AND2X2_339 ( .A(_abc_19068_n923_bF_buf4), .B(_abc_19068_n1494), .Y(_auto_iopadmap_cc_313_execute_30317_25_) );
  AND2X2 AND2X2_3390 ( .A(core__abc_21380_n2749_bF_buf9), .B(core__abc_21380_n5501), .Y(core__abc_21380_n5502) );
  AND2X2 AND2X2_3391 ( .A(core__abc_21380_n5506), .B(reset_n_bF_buf29), .Y(core__abc_21380_n5507) );
  AND2X2 AND2X2_3392 ( .A(core__abc_21380_n5505), .B(core__abc_21380_n5507), .Y(core_v3_reg_35__FF_INPUT) );
  AND2X2 AND2X2_3393 ( .A(core__abc_21380_n5510), .B(core__abc_21380_n5421), .Y(core__abc_21380_n5511) );
  AND2X2 AND2X2_3394 ( .A(core__abc_21380_n5512), .B(core__abc_21380_n5513), .Y(core__abc_21380_n5514) );
  AND2X2 AND2X2_3395 ( .A(core__abc_21380_n5510), .B(core__abc_21380_n5417), .Y(core__abc_21380_n5517) );
  AND2X2 AND2X2_3396 ( .A(core__abc_21380_n5353), .B(core__abc_21380_n5517), .Y(core__abc_21380_n5518) );
  AND2X2 AND2X2_3397 ( .A(core__abc_21380_n3176), .B(core__abc_21380_n1339), .Y(core__abc_21380_n5520) );
  AND2X2 AND2X2_3398 ( .A(core__abc_21380_n3275), .B(core__abc_21380_n1347), .Y(core__abc_21380_n5521) );
  AND2X2 AND2X2_3399 ( .A(core__abc_21380_n5321), .B(core__abc_21380_n3121), .Y(core__abc_21380_n5525) );
  AND2X2 AND2X2_34 ( .A(_abc_19068_n912_1), .B(_abc_19068_n907_1), .Y(_abc_19068_n924_1) );
  AND2X2 AND2X2_340 ( .A(_abc_19068_n916_1_bF_buf2), .B(word1_reg_26_), .Y(_abc_19068_n1496) );
  AND2X2 AND2X2_3400 ( .A(core__abc_21380_n5526), .B(core__abc_21380_n1935), .Y(core__abc_21380_n5527) );
  AND2X2 AND2X2_3401 ( .A(core__abc_21380_n5528), .B(core__abc_21380_n1938), .Y(core__abc_21380_n5529) );
  AND2X2 AND2X2_3402 ( .A(core__abc_21380_n5532), .B(core__abc_21380_n5533), .Y(core__abc_21380_n5534) );
  AND2X2 AND2X2_3403 ( .A(core__abc_21380_n5535), .B(core__abc_21380_n5523), .Y(core__abc_21380_n5536) );
  AND2X2 AND2X2_3404 ( .A(core__abc_21380_n5534), .B(core__abc_21380_n5522), .Y(core__abc_21380_n5537) );
  AND2X2 AND2X2_3405 ( .A(core__abc_21380_n5519), .B(core__abc_21380_n5539), .Y(core__abc_21380_n5540) );
  AND2X2 AND2X2_3406 ( .A(core__abc_21380_n5541), .B(core__abc_21380_n5538), .Y(core__abc_21380_n5542) );
  AND2X2 AND2X2_3407 ( .A(core__abc_21380_n5546), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n5547) );
  AND2X2 AND2X2_3408 ( .A(core__abc_21380_n5547), .B(core__abc_21380_n5544), .Y(core__abc_21380_n5548) );
  AND2X2 AND2X2_3409 ( .A(core__abc_21380_n3313_bF_buf1), .B(core_key_100_), .Y(core__abc_21380_n5549) );
  AND2X2 AND2X2_341 ( .A(_abc_19068_n897_1_bF_buf2), .B(word0_reg_26_), .Y(_abc_19068_n1497_1) );
  AND2X2 AND2X2_3410 ( .A(core_v3_reg_36_), .B(core_mi_36_), .Y(core__abc_21380_n5551) );
  AND2X2 AND2X2_3411 ( .A(core__abc_21380_n5552), .B(core__abc_21380_n5550), .Y(core__abc_21380_n5553) );
  AND2X2 AND2X2_3412 ( .A(core__abc_21380_n2749_bF_buf8), .B(core__abc_21380_n5553), .Y(core__abc_21380_n5554) );
  AND2X2 AND2X2_3413 ( .A(core__abc_21380_n5558), .B(reset_n_bF_buf28), .Y(core__abc_21380_n5559) );
  AND2X2 AND2X2_3414 ( .A(core__abc_21380_n5557), .B(core__abc_21380_n5559), .Y(core_v3_reg_36__FF_INPUT) );
  AND2X2 AND2X2_3415 ( .A(core__abc_21380_n5563), .B(core__abc_21380_n1358), .Y(core__abc_21380_n5564) );
  AND2X2 AND2X2_3416 ( .A(core__abc_21380_n5562), .B(core__abc_21380_n1359), .Y(core__abc_21380_n5565) );
  AND2X2 AND2X2_3417 ( .A(core__abc_21380_n5569), .B(core__abc_21380_n1956), .Y(core__abc_21380_n5570) );
  AND2X2 AND2X2_3418 ( .A(core__abc_21380_n5568), .B(core__abc_21380_n1955), .Y(core__abc_21380_n5571) );
  AND2X2 AND2X2_3419 ( .A(core__abc_21380_n5572), .B(core_v3_reg_21_), .Y(core__abc_21380_n5573) );
  AND2X2 AND2X2_342 ( .A(_abc_19068_n939_1_bF_buf3), .B(core_key_90_), .Y(_abc_19068_n1499_1) );
  AND2X2 AND2X2_3420 ( .A(core__abc_21380_n5574), .B(core__abc_21380_n5575), .Y(core__abc_21380_n5576) );
  AND2X2 AND2X2_3421 ( .A(core__abc_21380_n5577), .B(core__abc_21380_n5567), .Y(core__abc_21380_n5578) );
  AND2X2 AND2X2_3422 ( .A(core__abc_21380_n5576), .B(core__abc_21380_n5566), .Y(core__abc_21380_n5580) );
  AND2X2 AND2X2_3423 ( .A(core__abc_21380_n5579), .B(core__abc_21380_n5581), .Y(core__abc_21380_n5582) );
  AND2X2 AND2X2_3424 ( .A(core__abc_21380_n5586), .B(core__abc_21380_n5583), .Y(core__abc_21380_n5587) );
  AND2X2 AND2X2_3425 ( .A(core__abc_21380_n5590), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n5591) );
  AND2X2 AND2X2_3426 ( .A(core__abc_21380_n5591), .B(core__abc_21380_n5589), .Y(core__abc_21380_n5592) );
  AND2X2 AND2X2_3427 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n5593), .Y(core__abc_21380_n5594) );
  AND2X2 AND2X2_3428 ( .A(core_v3_reg_37_), .B(core_mi_37_), .Y(core__abc_21380_n5596) );
  AND2X2 AND2X2_3429 ( .A(core__abc_21380_n5597), .B(core__abc_21380_n5595), .Y(core__abc_21380_n5598) );
  AND2X2 AND2X2_343 ( .A(_abc_19068_n924_1_bF_buf3), .B(core_key_58_), .Y(_abc_19068_n1500) );
  AND2X2 AND2X2_3430 ( .A(core__abc_21380_n2749_bF_buf7), .B(core__abc_21380_n5598), .Y(core__abc_21380_n5599) );
  AND2X2 AND2X2_3431 ( .A(core__abc_21380_n5603), .B(reset_n_bF_buf27), .Y(core__abc_21380_n5604) );
  AND2X2 AND2X2_3432 ( .A(core__abc_21380_n5602), .B(core__abc_21380_n5604), .Y(core_v3_reg_37__FF_INPUT) );
  AND2X2 AND2X2_3433 ( .A(core__abc_21380_n5606), .B(core__abc_21380_n5581), .Y(core__abc_21380_n5607) );
  AND2X2 AND2X2_3434 ( .A(core__abc_21380_n5582), .B(core__abc_21380_n5539), .Y(core__abc_21380_n5608) );
  AND2X2 AND2X2_3435 ( .A(core__abc_21380_n5519), .B(core__abc_21380_n5608), .Y(core__abc_21380_n5609) );
  AND2X2 AND2X2_3436 ( .A(core__abc_21380_n3176), .B(core__abc_21380_n3178), .Y(core__abc_21380_n5612) );
  AND2X2 AND2X2_3437 ( .A(core__abc_21380_n5613), .B(core__abc_21380_n1378), .Y(core__abc_21380_n5614) );
  AND2X2 AND2X2_3438 ( .A(core__abc_21380_n5615), .B(core__abc_21380_n5616), .Y(core__abc_21380_n5617) );
  AND2X2 AND2X2_3439 ( .A(core__abc_21380_n5526), .B(core__abc_21380_n3117), .Y(core__abc_21380_n5618) );
  AND2X2 AND2X2_344 ( .A(_abc_19068_n926_bF_buf3), .B(core_key_26_), .Y(_abc_19068_n1501_1) );
  AND2X2 AND2X2_3440 ( .A(core__abc_21380_n5620), .B(core__abc_21380_n1976), .Y(core__abc_21380_n5621) );
  AND2X2 AND2X2_3441 ( .A(core__abc_21380_n5619), .B(core__abc_21380_n1974), .Y(core__abc_21380_n5622) );
  AND2X2 AND2X2_3442 ( .A(core__abc_21380_n5625), .B(core__abc_21380_n5627), .Y(core__abc_21380_n5628) );
  AND2X2 AND2X2_3443 ( .A(core__abc_21380_n5628), .B(core__abc_21380_n5617), .Y(core__abc_21380_n5629) );
  AND2X2 AND2X2_3444 ( .A(core__abc_21380_n5631), .B(core__abc_21380_n5630), .Y(core__abc_21380_n5632) );
  AND2X2 AND2X2_3445 ( .A(core__abc_21380_n5611), .B(core__abc_21380_n5633), .Y(core__abc_21380_n5634) );
  AND2X2 AND2X2_3446 ( .A(core__abc_21380_n5610), .B(core__abc_21380_n5635), .Y(core__abc_21380_n5636) );
  AND2X2 AND2X2_3447 ( .A(core__abc_21380_n5640), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n5641) );
  AND2X2 AND2X2_3448 ( .A(core__abc_21380_n5641), .B(core__abc_21380_n5638), .Y(core__abc_21380_n5642) );
  AND2X2 AND2X2_3449 ( .A(core__abc_21380_n3313_bF_buf12), .B(core__abc_21380_n5643), .Y(core__abc_21380_n5644) );
  AND2X2 AND2X2_345 ( .A(_abc_19068_n941_bF_buf3), .B(core_key_122_), .Y(_abc_19068_n1505_1) );
  AND2X2 AND2X2_3450 ( .A(core_v3_reg_38_), .B(core_mi_38_), .Y(core__abc_21380_n5646) );
  AND2X2 AND2X2_3451 ( .A(core__abc_21380_n5647), .B(core__abc_21380_n5645), .Y(core__abc_21380_n5648) );
  AND2X2 AND2X2_3452 ( .A(core__abc_21380_n2749_bF_buf6), .B(core__abc_21380_n5648), .Y(core__abc_21380_n5649) );
  AND2X2 AND2X2_3453 ( .A(core__abc_21380_n5653), .B(reset_n_bF_buf26), .Y(core__abc_21380_n5654) );
  AND2X2 AND2X2_3454 ( .A(core__abc_21380_n5652), .B(core__abc_21380_n5654), .Y(core_v3_reg_38__FF_INPUT) );
  AND2X2 AND2X2_3455 ( .A(core__abc_21380_n5615), .B(core__abc_21380_n5657), .Y(core__abc_21380_n5658) );
  AND2X2 AND2X2_3456 ( .A(core__abc_21380_n5658), .B(core__abc_21380_n1396), .Y(core__abc_21380_n5659) );
  AND2X2 AND2X2_3457 ( .A(core__abc_21380_n5660), .B(core__abc_21380_n5661), .Y(core__abc_21380_n5662) );
  AND2X2 AND2X2_3458 ( .A(core__abc_21380_n5665), .B(core__abc_21380_n1996), .Y(core__abc_21380_n5666) );
  AND2X2 AND2X2_3459 ( .A(core__abc_21380_n5664), .B(core__abc_21380_n1993), .Y(core__abc_21380_n5667) );
  AND2X2 AND2X2_346 ( .A(_abc_19068_n902_bF_buf2), .B(word2_reg_26_), .Y(_abc_19068_n1506) );
  AND2X2 AND2X2_3460 ( .A(core__abc_21380_n5668), .B(core__abc_21380_n5663), .Y(core__abc_21380_n5669) );
  AND2X2 AND2X2_3461 ( .A(core__abc_21380_n5670), .B(core__abc_21380_n5671), .Y(core__abc_21380_n5672) );
  AND2X2 AND2X2_3462 ( .A(core__abc_21380_n5672), .B(core__abc_21380_n5662), .Y(core__abc_21380_n5673) );
  AND2X2 AND2X2_3463 ( .A(core__abc_21380_n5674), .B(core__abc_21380_n5675), .Y(core__abc_21380_n5676) );
  AND2X2 AND2X2_3464 ( .A(core__abc_21380_n5681), .B(core__abc_21380_n5679), .Y(core__abc_21380_n5682) );
  AND2X2 AND2X2_3465 ( .A(core__abc_21380_n5684), .B(core__abc_21380_n5677), .Y(core__abc_21380_n5685) );
  AND2X2 AND2X2_3466 ( .A(core__abc_21380_n5688), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n5689) );
  AND2X2 AND2X2_3467 ( .A(core__abc_21380_n5689), .B(core__abc_21380_n5686), .Y(core__abc_21380_n5690) );
  AND2X2 AND2X2_3468 ( .A(core__abc_21380_n3313_bF_buf11), .B(core_key_103_), .Y(core__abc_21380_n5691) );
  AND2X2 AND2X2_3469 ( .A(core_v3_reg_39_), .B(core_mi_39_), .Y(core__abc_21380_n5693) );
  AND2X2 AND2X2_347 ( .A(_abc_19068_n899_bF_buf2), .B(word3_reg_26_), .Y(_abc_19068_n1507_1) );
  AND2X2 AND2X2_3470 ( .A(core__abc_21380_n5694), .B(core__abc_21380_n5692), .Y(core__abc_21380_n5695) );
  AND2X2 AND2X2_3471 ( .A(core__abc_21380_n2749_bF_buf5), .B(core__abc_21380_n5695), .Y(core__abc_21380_n5696) );
  AND2X2 AND2X2_3472 ( .A(core__abc_21380_n5700), .B(reset_n_bF_buf25), .Y(core__abc_21380_n5701) );
  AND2X2 AND2X2_3473 ( .A(core__abc_21380_n5699), .B(core__abc_21380_n5701), .Y(core_v3_reg_39__FF_INPUT) );
  AND2X2 AND2X2_3474 ( .A(core__abc_21380_n5676), .B(core__abc_21380_n5635), .Y(core__abc_21380_n5703) );
  AND2X2 AND2X2_3475 ( .A(core__abc_21380_n5703), .B(core__abc_21380_n5608), .Y(core__abc_21380_n5704) );
  AND2X2 AND2X2_3476 ( .A(core__abc_21380_n5704), .B(core__abc_21380_n5516), .Y(core__abc_21380_n5705) );
  AND2X2 AND2X2_3477 ( .A(core__abc_21380_n5703), .B(core__abc_21380_n5607), .Y(core__abc_21380_n5706) );
  AND2X2 AND2X2_3478 ( .A(core__abc_21380_n5675), .B(core__abc_21380_n5629), .Y(core__abc_21380_n5707) );
  AND2X2 AND2X2_3479 ( .A(core__abc_21380_n5704), .B(core__abc_21380_n5517), .Y(core__abc_21380_n5711) );
  AND2X2 AND2X2_348 ( .A(_abc_19068_n945_1_bF_buf3), .B(core_mi_26_), .Y(_abc_19068_n1509_1) );
  AND2X2 AND2X2_3480 ( .A(core__abc_21380_n5353), .B(core__abc_21380_n5711), .Y(core__abc_21380_n5712) );
  AND2X2 AND2X2_3481 ( .A(core__abc_21380_n3189), .B(core__abc_21380_n1414), .Y(core__abc_21380_n5714) );
  AND2X2 AND2X2_3482 ( .A(core__abc_21380_n3279), .B(core__abc_21380_n1421), .Y(core__abc_21380_n5715) );
  AND2X2 AND2X2_3483 ( .A(core__abc_21380_n3143), .B(core__abc_21380_n2013), .Y(core__abc_21380_n5719) );
  AND2X2 AND2X2_3484 ( .A(core__abc_21380_n3144), .B(core__abc_21380_n2012), .Y(core__abc_21380_n5720) );
  AND2X2 AND2X2_3485 ( .A(core__abc_21380_n5723), .B(core__abc_21380_n5724), .Y(core__abc_21380_n5725) );
  AND2X2 AND2X2_3486 ( .A(core__abc_21380_n5726), .B(core__abc_21380_n5717), .Y(core__abc_21380_n5727) );
  AND2X2 AND2X2_3487 ( .A(core__abc_21380_n5725), .B(core__abc_21380_n5716), .Y(core__abc_21380_n5728) );
  AND2X2 AND2X2_3488 ( .A(core__abc_21380_n5713), .B(core__abc_21380_n5730), .Y(core__abc_21380_n5731) );
  AND2X2 AND2X2_3489 ( .A(core__abc_21380_n5732), .B(core__abc_21380_n5729), .Y(core__abc_21380_n5733) );
  AND2X2 AND2X2_349 ( .A(_abc_19068_n915_1_bF_buf2), .B(core_mi_58_), .Y(_abc_19068_n1510) );
  AND2X2 AND2X2_3490 ( .A(core__abc_21380_n5737), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n5738) );
  AND2X2 AND2X2_3491 ( .A(core__abc_21380_n5738), .B(core__abc_21380_n5736), .Y(core__abc_21380_n5739) );
  AND2X2 AND2X2_3492 ( .A(core__abc_21380_n3313_bF_buf10), .B(core_key_104_), .Y(core__abc_21380_n5740) );
  AND2X2 AND2X2_3493 ( .A(core_v3_reg_40_), .B(core_mi_40_), .Y(core__abc_21380_n5742) );
  AND2X2 AND2X2_3494 ( .A(core__abc_21380_n5743), .B(core__abc_21380_n5741), .Y(core__abc_21380_n5744) );
  AND2X2 AND2X2_3495 ( .A(core__abc_21380_n2749_bF_buf4), .B(core__abc_21380_n5744), .Y(core__abc_21380_n5745) );
  AND2X2 AND2X2_3496 ( .A(core__abc_21380_n5749), .B(reset_n_bF_buf24), .Y(core__abc_21380_n5750) );
  AND2X2 AND2X2_3497 ( .A(core__abc_21380_n5748), .B(core__abc_21380_n5750), .Y(core_v3_reg_40__FF_INPUT) );
  AND2X2 AND2X2_3498 ( .A(core__abc_21380_n5753), .B(core__abc_21380_n5752), .Y(core__abc_21380_n5754) );
  AND2X2 AND2X2_3499 ( .A(core__abc_21380_n5756), .B(core__abc_21380_n1441), .Y(core__abc_21380_n5757) );
  AND2X2 AND2X2_35 ( .A(_abc_19068_n924_1_bF_buf4), .B(core_key_32_), .Y(_abc_19068_n925_1) );
  AND2X2 AND2X2_350 ( .A(_abc_19068_n923_bF_buf3), .B(_abc_19068_n1514), .Y(_auto_iopadmap_cc_313_execute_30317_26_) );
  AND2X2 AND2X2_3500 ( .A(core__abc_21380_n5755), .B(core__abc_21380_n1434), .Y(core__abc_21380_n5758) );
  AND2X2 AND2X2_3501 ( .A(core__abc_21380_n5763), .B(core__abc_21380_n2032), .Y(core__abc_21380_n5764) );
  AND2X2 AND2X2_3502 ( .A(core__abc_21380_n5762), .B(core__abc_21380_n2029), .Y(core__abc_21380_n5765) );
  AND2X2 AND2X2_3503 ( .A(core__abc_21380_n5766), .B(core__abc_21380_n5761), .Y(core__abc_21380_n5767) );
  AND2X2 AND2X2_3504 ( .A(core__abc_21380_n5768), .B(core_v3_reg_25_), .Y(core__abc_21380_n5769) );
  AND2X2 AND2X2_3505 ( .A(core__abc_21380_n5771), .B(core__abc_21380_n5760), .Y(core__abc_21380_n5772) );
  AND2X2 AND2X2_3506 ( .A(core__abc_21380_n5770), .B(core__abc_21380_n5759), .Y(core__abc_21380_n5774) );
  AND2X2 AND2X2_3507 ( .A(core__abc_21380_n5773), .B(core__abc_21380_n5775), .Y(core__abc_21380_n5776) );
  AND2X2 AND2X2_3508 ( .A(core__abc_21380_n5780), .B(core__abc_21380_n5777), .Y(core__abc_21380_n5781) );
  AND2X2 AND2X2_3509 ( .A(core__abc_21380_n5784), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n5785) );
  AND2X2 AND2X2_351 ( .A(_abc_19068_n916_1_bF_buf1), .B(word1_reg_27_), .Y(_abc_19068_n1516) );
  AND2X2 AND2X2_3510 ( .A(core__abc_21380_n5785), .B(core__abc_21380_n5783), .Y(core__abc_21380_n5786) );
  AND2X2 AND2X2_3511 ( .A(core__abc_21380_n3313_bF_buf9), .B(core_key_105_), .Y(core__abc_21380_n5787) );
  AND2X2 AND2X2_3512 ( .A(core_v3_reg_41_), .B(core_mi_41_), .Y(core__abc_21380_n5789) );
  AND2X2 AND2X2_3513 ( .A(core__abc_21380_n5790), .B(core__abc_21380_n5788), .Y(core__abc_21380_n5791) );
  AND2X2 AND2X2_3514 ( .A(core__abc_21380_n2749_bF_buf3), .B(core__abc_21380_n5791), .Y(core__abc_21380_n5792) );
  AND2X2 AND2X2_3515 ( .A(core__abc_21380_n5796), .B(reset_n_bF_buf23), .Y(core__abc_21380_n5797) );
  AND2X2 AND2X2_3516 ( .A(core__abc_21380_n5795), .B(core__abc_21380_n5797), .Y(core_v3_reg_41__FF_INPUT) );
  AND2X2 AND2X2_3517 ( .A(core__abc_21380_n3189), .B(core__abc_21380_n3194_1), .Y(core__abc_21380_n5799) );
  AND2X2 AND2X2_3518 ( .A(core__abc_21380_n5800), .B(core__abc_21380_n1451), .Y(core__abc_21380_n5801) );
  AND2X2 AND2X2_3519 ( .A(core__abc_21380_n5802), .B(core__abc_21380_n5803), .Y(core__abc_21380_n5804) );
  AND2X2 AND2X2_352 ( .A(_abc_19068_n897_1_bF_buf1), .B(word0_reg_27_), .Y(_abc_19068_n1517_1) );
  AND2X2 AND2X2_3520 ( .A(core__abc_21380_n3149), .B(core__abc_21380_n5806), .Y(core__abc_21380_n5807) );
  AND2X2 AND2X2_3521 ( .A(core__abc_21380_n5810), .B(core__abc_21380_n5808), .Y(core__abc_21380_n5811) );
  AND2X2 AND2X2_3522 ( .A(core__abc_21380_n5812), .B(core__abc_21380_n5804), .Y(core__abc_21380_n5813) );
  AND2X2 AND2X2_3523 ( .A(core__abc_21380_n5811), .B(core__abc_21380_n5814), .Y(core__abc_21380_n5815) );
  AND2X2 AND2X2_3524 ( .A(core__abc_21380_n5773), .B(core__abc_21380_n5752), .Y(core__abc_21380_n5817) );
  AND2X2 AND2X2_3525 ( .A(core__abc_21380_n5753), .B(core__abc_21380_n5817), .Y(core__abc_21380_n5818) );
  AND2X2 AND2X2_3526 ( .A(core__abc_21380_n5819), .B(core__abc_21380_n5816), .Y(core__abc_21380_n5820) );
  AND2X2 AND2X2_3527 ( .A(core__abc_21380_n5826), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n5827) );
  AND2X2 AND2X2_3528 ( .A(core__abc_21380_n5827), .B(core__abc_21380_n5824), .Y(core__abc_21380_n5828) );
  AND2X2 AND2X2_3529 ( .A(core__abc_21380_n3313_bF_buf8), .B(core__abc_21380_n5829), .Y(core__abc_21380_n5830) );
  AND2X2 AND2X2_353 ( .A(_abc_19068_n939_1_bF_buf2), .B(core_key_91_), .Y(_abc_19068_n1519_1) );
  AND2X2 AND2X2_3530 ( .A(core_v3_reg_42_), .B(core_mi_42_), .Y(core__abc_21380_n5832) );
  AND2X2 AND2X2_3531 ( .A(core__abc_21380_n5833), .B(core__abc_21380_n5831), .Y(core__abc_21380_n5834) );
  AND2X2 AND2X2_3532 ( .A(core__abc_21380_n2749_bF_buf2), .B(core__abc_21380_n5834), .Y(core__abc_21380_n5835) );
  AND2X2 AND2X2_3533 ( .A(core__abc_21380_n5839), .B(reset_n_bF_buf22), .Y(core__abc_21380_n5840) );
  AND2X2 AND2X2_3534 ( .A(core__abc_21380_n5838), .B(core__abc_21380_n5840), .Y(core_v3_reg_42__FF_INPUT) );
  AND2X2 AND2X2_3535 ( .A(core__abc_21380_n5821), .B(core__abc_21380_n5842), .Y(core__abc_21380_n5843) );
  AND2X2 AND2X2_3536 ( .A(core__abc_21380_n5802), .B(core__abc_21380_n1450), .Y(core__abc_21380_n5844) );
  AND2X2 AND2X2_3537 ( .A(core__abc_21380_n5844), .B(core__abc_21380_n1474), .Y(core__abc_21380_n5845) );
  AND2X2 AND2X2_3538 ( .A(core__abc_21380_n5846), .B(core__abc_21380_n5847), .Y(core__abc_21380_n5848) );
  AND2X2 AND2X2_3539 ( .A(core__abc_21380_n5851), .B(core__abc_21380_n5850), .Y(core__abc_21380_n5852) );
  AND2X2 AND2X2_354 ( .A(_abc_19068_n924_1_bF_buf2), .B(core_key_59_), .Y(_abc_19068_n1520) );
  AND2X2 AND2X2_3540 ( .A(core__abc_21380_n5843), .B(core__abc_21380_n5853), .Y(core__abc_21380_n5854) );
  AND2X2 AND2X2_3541 ( .A(core__abc_21380_n5855), .B(core__abc_21380_n5852), .Y(core__abc_21380_n5856) );
  AND2X2 AND2X2_3542 ( .A(core__abc_21380_n5860), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n5861) );
  AND2X2 AND2X2_3543 ( .A(core__abc_21380_n5861), .B(core__abc_21380_n5859), .Y(core__abc_21380_n5862) );
  AND2X2 AND2X2_3544 ( .A(core__abc_21380_n3313_bF_buf7), .B(core_key_107_), .Y(core__abc_21380_n5863) );
  AND2X2 AND2X2_3545 ( .A(core_v3_reg_43_), .B(core_mi_43_), .Y(core__abc_21380_n5865) );
  AND2X2 AND2X2_3546 ( .A(core__abc_21380_n5866), .B(core__abc_21380_n5864), .Y(core__abc_21380_n5867) );
  AND2X2 AND2X2_3547 ( .A(core__abc_21380_n2749_bF_buf1), .B(core__abc_21380_n5867), .Y(core__abc_21380_n5868) );
  AND2X2 AND2X2_3548 ( .A(core__abc_21380_n5872), .B(reset_n_bF_buf21), .Y(core__abc_21380_n5873) );
  AND2X2 AND2X2_3549 ( .A(core__abc_21380_n5871), .B(core__abc_21380_n5873), .Y(core_v3_reg_43__FF_INPUT) );
  AND2X2 AND2X2_355 ( .A(_abc_19068_n926_bF_buf2), .B(core_key_27_), .Y(_abc_19068_n1521_1) );
  AND2X2 AND2X2_3550 ( .A(core__abc_21380_n5852), .B(core__abc_21380_n5877), .Y(core__abc_21380_n5878) );
  AND2X2 AND2X2_3551 ( .A(core__abc_21380_n5878), .B(core__abc_21380_n5876), .Y(core__abc_21380_n5879) );
  AND2X2 AND2X2_3552 ( .A(core__abc_21380_n3159), .B(core__abc_21380_n5849), .Y(core__abc_21380_n5880) );
  AND2X2 AND2X2_3553 ( .A(core__abc_21380_n5881), .B(core__abc_21380_n5850), .Y(core__abc_21380_n5882) );
  AND2X2 AND2X2_3554 ( .A(core__abc_21380_n5776), .B(core__abc_21380_n5730), .Y(core__abc_21380_n5885) );
  AND2X2 AND2X2_3555 ( .A(core__abc_21380_n5878), .B(core__abc_21380_n5885), .Y(core__abc_21380_n5886) );
  AND2X2 AND2X2_3556 ( .A(core__abc_21380_n5713), .B(core__abc_21380_n5886), .Y(core__abc_21380_n5887) );
  AND2X2 AND2X2_3557 ( .A(core__abc_21380_n3189), .B(core__abc_21380_n3196), .Y(core__abc_21380_n5890) );
  AND2X2 AND2X2_3558 ( .A(core__abc_21380_n5892), .B(core__abc_21380_n1486), .Y(core__abc_21380_n5893) );
  AND2X2 AND2X2_3559 ( .A(core__abc_21380_n5891), .B(core__abc_21380_n1487), .Y(core__abc_21380_n5894) );
  AND2X2 AND2X2_356 ( .A(_abc_19068_n941_bF_buf2), .B(core_key_123_), .Y(_abc_19068_n1525_1) );
  AND2X2 AND2X2_3560 ( .A(core__abc_21380_n3384), .B(core__abc_21380_n5896), .Y(core__abc_21380_n5897) );
  AND2X2 AND2X2_3561 ( .A(core__abc_21380_n3383), .B(core__abc_21380_n5895), .Y(core__abc_21380_n5898) );
  AND2X2 AND2X2_3562 ( .A(core__abc_21380_n5889), .B(core__abc_21380_n5899), .Y(core__abc_21380_n5900) );
  AND2X2 AND2X2_3563 ( .A(core__abc_21380_n5888), .B(core__abc_21380_n5901), .Y(core__abc_21380_n5902) );
  AND2X2 AND2X2_3564 ( .A(core__abc_21380_n5906), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n5907) );
  AND2X2 AND2X2_3565 ( .A(core__abc_21380_n5907), .B(core__abc_21380_n5904), .Y(core__abc_21380_n5908) );
  AND2X2 AND2X2_3566 ( .A(core__abc_21380_n3313_bF_buf6), .B(core_key_108_), .Y(core__abc_21380_n5909) );
  AND2X2 AND2X2_3567 ( .A(core_v3_reg_44_), .B(core_mi_44_), .Y(core__abc_21380_n5911) );
  AND2X2 AND2X2_3568 ( .A(core__abc_21380_n5912), .B(core__abc_21380_n5910), .Y(core__abc_21380_n5913) );
  AND2X2 AND2X2_3569 ( .A(core__abc_21380_n2749_bF_buf0), .B(core__abc_21380_n5913), .Y(core__abc_21380_n5914) );
  AND2X2 AND2X2_357 ( .A(_abc_19068_n902_bF_buf1), .B(word2_reg_27_), .Y(_abc_19068_n1526) );
  AND2X2 AND2X2_3570 ( .A(core__abc_21380_n5918), .B(reset_n_bF_buf20), .Y(core__abc_21380_n5919) );
  AND2X2 AND2X2_3571 ( .A(core__abc_21380_n5917), .B(core__abc_21380_n5919), .Y(core_v3_reg_44__FF_INPUT) );
  AND2X2 AND2X2_3572 ( .A(core__abc_21380_n5922), .B(core__abc_21380_n1504), .Y(core__abc_21380_n5923) );
  AND2X2 AND2X2_3573 ( .A(core__abc_21380_n5921), .B(core__abc_21380_n1505), .Y(core__abc_21380_n5924) );
  AND2X2 AND2X2_3574 ( .A(core__abc_21380_n5926), .B(core__abc_21380_n5928), .Y(core__abc_21380_n5929) );
  AND2X2 AND2X2_3575 ( .A(core__abc_21380_n5932), .B(core__abc_21380_n5931), .Y(core__abc_21380_n5933) );
  AND2X2 AND2X2_3576 ( .A(core__abc_21380_n5933), .B(core__abc_21380_n5930), .Y(core__abc_21380_n5934) );
  AND2X2 AND2X2_3577 ( .A(core__abc_21380_n5940), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf0), .Y(core__abc_21380_n5941) );
  AND2X2 AND2X2_3578 ( .A(core__abc_21380_n5941), .B(core__abc_21380_n5939), .Y(core__abc_21380_n5942) );
  AND2X2 AND2X2_3579 ( .A(core__abc_21380_n3313_bF_buf5), .B(core__abc_21380_n5943), .Y(core__abc_21380_n5944) );
  AND2X2 AND2X2_358 ( .A(_abc_19068_n899_bF_buf1), .B(word3_reg_27_), .Y(_abc_19068_n1527_1) );
  AND2X2 AND2X2_3580 ( .A(core_v3_reg_45_), .B(core_mi_45_), .Y(core__abc_21380_n5946) );
  AND2X2 AND2X2_3581 ( .A(core__abc_21380_n5947), .B(core__abc_21380_n5945), .Y(core__abc_21380_n5948) );
  AND2X2 AND2X2_3582 ( .A(core__abc_21380_n2749_bF_buf10), .B(core__abc_21380_n5948), .Y(core__abc_21380_n5949) );
  AND2X2 AND2X2_3583 ( .A(core__abc_21380_n5953), .B(reset_n_bF_buf19), .Y(core__abc_21380_n5954) );
  AND2X2 AND2X2_3584 ( .A(core__abc_21380_n5952), .B(core__abc_21380_n5954), .Y(core_v3_reg_45__FF_INPUT) );
  AND2X2 AND2X2_3585 ( .A(core__abc_21380_n5929), .B(core__abc_21380_n5901), .Y(core__abc_21380_n5956) );
  AND2X2 AND2X2_3586 ( .A(core__abc_21380_n5888), .B(core__abc_21380_n5956), .Y(core__abc_21380_n5957) );
  AND2X2 AND2X2_3587 ( .A(core__abc_21380_n5929), .B(core__abc_21380_n5897), .Y(core__abc_21380_n5959) );
  AND2X2 AND2X2_3588 ( .A(core__abc_21380_n5891), .B(core__abc_21380_n3192), .Y(core__abc_21380_n5963) );
  AND2X2 AND2X2_3589 ( .A(core__abc_21380_n5964), .B(core__abc_21380_n1523), .Y(core__abc_21380_n5965) );
  AND2X2 AND2X2_359 ( .A(_abc_19068_n945_1_bF_buf2), .B(core_mi_27_), .Y(_abc_19068_n1529_1) );
  AND2X2 AND2X2_3590 ( .A(core__abc_21380_n5966), .B(core__abc_21380_n5967), .Y(core__abc_21380_n5968) );
  AND2X2 AND2X2_3591 ( .A(core__abc_21380_n3505_1), .B(core__abc_21380_n5968), .Y(core__abc_21380_n5969) );
  AND2X2 AND2X2_3592 ( .A(core__abc_21380_n3507), .B(core__abc_21380_n5970), .Y(core__abc_21380_n5971) );
  AND2X2 AND2X2_3593 ( .A(core__abc_21380_n5962), .B(core__abc_21380_n5972), .Y(core__abc_21380_n5973) );
  AND2X2 AND2X2_3594 ( .A(core__abc_21380_n5961), .B(core__abc_21380_n5974), .Y(core__abc_21380_n5975) );
  AND2X2 AND2X2_3595 ( .A(core__abc_21380_n5980), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf0), .Y(core__abc_21380_n5981) );
  AND2X2 AND2X2_3596 ( .A(core__abc_21380_n5981), .B(core__abc_21380_n5977), .Y(core__abc_21380_n5982) );
  AND2X2 AND2X2_3597 ( .A(core__abc_21380_n3313_bF_buf4), .B(core__abc_21380_n5983), .Y(core__abc_21380_n5984) );
  AND2X2 AND2X2_3598 ( .A(core_v3_reg_46_), .B(core_mi_46_), .Y(core__abc_21380_n5986) );
  AND2X2 AND2X2_3599 ( .A(core__abc_21380_n5987), .B(core__abc_21380_n5985), .Y(core__abc_21380_n5988) );
  AND2X2 AND2X2_36 ( .A(_abc_19068_n894_1), .B(_abc_19068_n912_1), .Y(_abc_19068_n926) );
  AND2X2 AND2X2_360 ( .A(_abc_19068_n915_1_bF_buf1), .B(core_mi_59_), .Y(_abc_19068_n1530) );
  AND2X2 AND2X2_3600 ( .A(core__abc_21380_n2749_bF_buf9), .B(core__abc_21380_n5988), .Y(core__abc_21380_n5989) );
  AND2X2 AND2X2_3601 ( .A(core__abc_21380_n5993), .B(reset_n_bF_buf18), .Y(core__abc_21380_n5994) );
  AND2X2 AND2X2_3602 ( .A(core__abc_21380_n5992), .B(core__abc_21380_n5994), .Y(core_v3_reg_46__FF_INPUT) );
  AND2X2 AND2X2_3603 ( .A(core__abc_21380_n5998), .B(core__abc_21380_n1548), .Y(core__abc_21380_n5999) );
  AND2X2 AND2X2_3604 ( .A(core__abc_21380_n5997), .B(core__abc_21380_n1542), .Y(core__abc_21380_n6000) );
  AND2X2 AND2X2_3605 ( .A(core__abc_21380_n3576), .B(core__abc_21380_n6002), .Y(core__abc_21380_n6003) );
  AND2X2 AND2X2_3606 ( .A(core__abc_21380_n3580), .B(core__abc_21380_n6001), .Y(core__abc_21380_n6004) );
  AND2X2 AND2X2_3607 ( .A(core__abc_21380_n6009), .B(core__abc_21380_n6008), .Y(core__abc_21380_n6010) );
  AND2X2 AND2X2_3608 ( .A(core__abc_21380_n6011), .B(core__abc_21380_n6006), .Y(core__abc_21380_n6012) );
  AND2X2 AND2X2_3609 ( .A(core__abc_21380_n6015), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n6016) );
  AND2X2 AND2X2_361 ( .A(_abc_19068_n923_bF_buf2), .B(_abc_19068_n1534), .Y(_auto_iopadmap_cc_313_execute_30317_27_) );
  AND2X2 AND2X2_3610 ( .A(core__abc_21380_n6016), .B(core__abc_21380_n6014), .Y(core__abc_21380_n6017) );
  AND2X2 AND2X2_3611 ( .A(core__abc_21380_n3313_bF_buf3), .B(core_key_111_), .Y(core__abc_21380_n6018) );
  AND2X2 AND2X2_3612 ( .A(core_v3_reg_47_), .B(core_mi_47_), .Y(core__abc_21380_n6020) );
  AND2X2 AND2X2_3613 ( .A(core__abc_21380_n6021), .B(core__abc_21380_n6019), .Y(core__abc_21380_n6022) );
  AND2X2 AND2X2_3614 ( .A(core__abc_21380_n2749_bF_buf8), .B(core__abc_21380_n6022), .Y(core__abc_21380_n6023) );
  AND2X2 AND2X2_3615 ( .A(core__abc_21380_n6027), .B(reset_n_bF_buf17), .Y(core__abc_21380_n6028) );
  AND2X2 AND2X2_3616 ( .A(core__abc_21380_n6026), .B(core__abc_21380_n6028), .Y(core_v3_reg_47__FF_INPUT) );
  AND2X2 AND2X2_3617 ( .A(core__abc_21380_n6010), .B(core__abc_21380_n5974), .Y(core__abc_21380_n6030) );
  AND2X2 AND2X2_3618 ( .A(core__abc_21380_n6030), .B(core__abc_21380_n5956), .Y(core__abc_21380_n6031) );
  AND2X2 AND2X2_3619 ( .A(core__abc_21380_n6031), .B(core__abc_21380_n5886), .Y(core__abc_21380_n6032) );
  AND2X2 AND2X2_362 ( .A(_abc_19068_n899_bF_buf0), .B(word3_reg_28_), .Y(_abc_19068_n1536) );
  AND2X2 AND2X2_3620 ( .A(core__abc_21380_n6032), .B(core__abc_21380_n5711), .Y(core__abc_21380_n6033) );
  AND2X2 AND2X2_3621 ( .A(core__abc_21380_n5353), .B(core__abc_21380_n6033), .Y(core__abc_21380_n6034) );
  AND2X2 AND2X2_3622 ( .A(core__abc_21380_n5710), .B(core__abc_21380_n6032), .Y(core__abc_21380_n6035) );
  AND2X2 AND2X2_3623 ( .A(core__abc_21380_n5884), .B(core__abc_21380_n6031), .Y(core__abc_21380_n6036) );
  AND2X2 AND2X2_3624 ( .A(core__abc_21380_n5960), .B(core__abc_21380_n6030), .Y(core__abc_21380_n6037) );
  AND2X2 AND2X2_3625 ( .A(core__abc_21380_n6039), .B(core__abc_21380_n6008), .Y(core__abc_21380_n6040) );
  AND2X2 AND2X2_3626 ( .A(core__abc_21380_n3215_1), .B(core__abc_21380_n1561), .Y(core__abc_21380_n6046) );
  AND2X2 AND2X2_3627 ( .A(core__abc_21380_n3283), .B(core__abc_21380_n1560), .Y(core__abc_21380_n6047) );
  AND2X2 AND2X2_3628 ( .A(core__abc_21380_n3648), .B(core__abc_21380_n6049), .Y(core__abc_21380_n6050) );
  AND2X2 AND2X2_3629 ( .A(core__abc_21380_n3647_1), .B(core__abc_21380_n6048), .Y(core__abc_21380_n6051) );
  AND2X2 AND2X2_363 ( .A(_abc_19068_n945_1_bF_buf1), .B(core_mi_28_), .Y(_abc_19068_n1538) );
  AND2X2 AND2X2_3630 ( .A(core__abc_21380_n6045), .B(core__abc_21380_n6053), .Y(core__abc_21380_n6054) );
  AND2X2 AND2X2_3631 ( .A(core__abc_21380_n6063), .B(core__abc_21380_n6064), .Y(core__abc_21380_n6065) );
  AND2X2 AND2X2_3632 ( .A(core__abc_21380_n6061), .B(core__abc_21380_n6065), .Y(core__abc_21380_n6066) );
  AND2X2 AND2X2_3633 ( .A(core__abc_21380_n6070), .B(core__abc_21380_n6069), .Y(core__abc_21380_n6071) );
  AND2X2 AND2X2_3634 ( .A(core__abc_21380_n6071), .B(core__abc_21380_n6068), .Y(core__abc_21380_n6072) );
  AND2X2 AND2X2_3635 ( .A(core__abc_21380_n6056), .B(core__abc_21380_n6072), .Y(core__abc_21380_n6073) );
  AND2X2 AND2X2_3636 ( .A(core__abc_21380_n6073), .B(core__abc_21380_n6052), .Y(core__abc_21380_n6074) );
  AND2X2 AND2X2_3637 ( .A(core__abc_21380_n6078), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n6079) );
  AND2X2 AND2X2_3638 ( .A(core__abc_21380_n6079), .B(core__abc_21380_n6077), .Y(core__abc_21380_n6080) );
  AND2X2 AND2X2_3639 ( .A(core__abc_21380_n3313_bF_buf2), .B(core__abc_21380_n6081), .Y(core__abc_21380_n6082) );
  AND2X2 AND2X2_364 ( .A(_abc_19068_n941_bF_buf1), .B(core_key_124_), .Y(_abc_19068_n1539_1) );
  AND2X2 AND2X2_3640 ( .A(core_v3_reg_48_), .B(core_mi_48_), .Y(core__abc_21380_n6084) );
  AND2X2 AND2X2_3641 ( .A(core__abc_21380_n6085), .B(core__abc_21380_n6083), .Y(core__abc_21380_n6086) );
  AND2X2 AND2X2_3642 ( .A(core__abc_21380_n2749_bF_buf7), .B(core__abc_21380_n6086), .Y(core__abc_21380_n6087) );
  AND2X2 AND2X2_3643 ( .A(core__abc_21380_n6091), .B(reset_n_bF_buf16), .Y(core__abc_21380_n6092) );
  AND2X2 AND2X2_3644 ( .A(core__abc_21380_n6090), .B(core__abc_21380_n6092), .Y(core_v3_reg_48__FF_INPUT) );
  AND2X2 AND2X2_3645 ( .A(core__abc_21380_n6095), .B(core__abc_21380_n6094), .Y(core__abc_21380_n6096) );
  AND2X2 AND2X2_3646 ( .A(core__abc_21380_n6099), .B(core__abc_21380_n1587), .Y(core__abc_21380_n6100) );
  AND2X2 AND2X2_3647 ( .A(core__abc_21380_n6098), .B(core__abc_21380_n1580), .Y(core__abc_21380_n6101) );
  AND2X2 AND2X2_3648 ( .A(core__abc_21380_n3720_1), .B(core__abc_21380_n6103), .Y(core__abc_21380_n6104) );
  AND2X2 AND2X2_3649 ( .A(core__abc_21380_n3719), .B(core__abc_21380_n6102), .Y(core__abc_21380_n6106) );
  AND2X2 AND2X2_365 ( .A(_abc_19068_n939_1_bF_buf1), .B(core_key_92_), .Y(_abc_19068_n1542) );
  AND2X2 AND2X2_3650 ( .A(core__abc_21380_n6105), .B(core__abc_21380_n6107), .Y(core__abc_21380_n6108) );
  AND2X2 AND2X2_3651 ( .A(core__abc_21380_n6109), .B(core__abc_21380_n6111), .Y(core__abc_21380_n6112) );
  AND2X2 AND2X2_3652 ( .A(core__abc_21380_n6115), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n6116) );
  AND2X2 AND2X2_3653 ( .A(core__abc_21380_n6116), .B(core__abc_21380_n6113), .Y(core__abc_21380_n6117) );
  AND2X2 AND2X2_3654 ( .A(core__abc_21380_n3313_bF_buf1), .B(core_key_113_), .Y(core__abc_21380_n6118) );
  AND2X2 AND2X2_3655 ( .A(core_v3_reg_49_), .B(core_mi_49_), .Y(core__abc_21380_n6120) );
  AND2X2 AND2X2_3656 ( .A(core__abc_21380_n6121), .B(core__abc_21380_n6119), .Y(core__abc_21380_n6122) );
  AND2X2 AND2X2_3657 ( .A(core__abc_21380_n2749_bF_buf6), .B(core__abc_21380_n6122), .Y(core__abc_21380_n6123) );
  AND2X2 AND2X2_3658 ( .A(core__abc_21380_n6127), .B(reset_n_bF_buf15), .Y(core__abc_21380_n6128) );
  AND2X2 AND2X2_3659 ( .A(core__abc_21380_n6126), .B(core__abc_21380_n6128), .Y(core_v3_reg_49__FF_INPUT) );
  AND2X2 AND2X2_366 ( .A(_abc_19068_n924_1_bF_buf1), .B(core_key_60_), .Y(_abc_19068_n1543_1) );
  AND2X2 AND2X2_3660 ( .A(core__abc_21380_n6105), .B(core__abc_21380_n6130), .Y(core__abc_21380_n6131) );
  AND2X2 AND2X2_3661 ( .A(core__abc_21380_n6108), .B(core__abc_21380_n6053), .Y(core__abc_21380_n6133) );
  AND2X2 AND2X2_3662 ( .A(core__abc_21380_n6045), .B(core__abc_21380_n6133), .Y(core__abc_21380_n6134) );
  AND2X2 AND2X2_3663 ( .A(core__abc_21380_n3215_1), .B(core__abc_21380_n3227), .Y(core__abc_21380_n6137) );
  AND2X2 AND2X2_3664 ( .A(core__abc_21380_n6138), .B(core__abc_21380_n1597), .Y(core__abc_21380_n6139) );
  AND2X2 AND2X2_3665 ( .A(core__abc_21380_n6140), .B(core__abc_21380_n6141), .Y(core__abc_21380_n6142) );
  AND2X2 AND2X2_3666 ( .A(core__abc_21380_n3780), .B(core__abc_21380_n6142), .Y(core__abc_21380_n6143) );
  AND2X2 AND2X2_3667 ( .A(core__abc_21380_n3779_1), .B(core__abc_21380_n6144), .Y(core__abc_21380_n6145) );
  AND2X2 AND2X2_3668 ( .A(core__abc_21380_n6136), .B(core__abc_21380_n6146), .Y(core__abc_21380_n6147) );
  AND2X2 AND2X2_3669 ( .A(core__abc_21380_n6135), .B(core__abc_21380_n6148), .Y(core__abc_21380_n6149) );
  AND2X2 AND2X2_367 ( .A(_abc_19068_n926_bF_buf1), .B(core_key_28_), .Y(_abc_19068_n1544) );
  AND2X2 AND2X2_3670 ( .A(core__abc_21380_n6153), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n6154) );
  AND2X2 AND2X2_3671 ( .A(core__abc_21380_n6154), .B(core__abc_21380_n6151), .Y(core__abc_21380_n6155) );
  AND2X2 AND2X2_3672 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n6156), .Y(core__abc_21380_n6157) );
  AND2X2 AND2X2_3673 ( .A(core_v3_reg_50_), .B(core_mi_50_), .Y(core__abc_21380_n6159) );
  AND2X2 AND2X2_3674 ( .A(core__abc_21380_n6160), .B(core__abc_21380_n6158), .Y(core__abc_21380_n6161) );
  AND2X2 AND2X2_3675 ( .A(core__abc_21380_n2749_bF_buf5), .B(core__abc_21380_n6161), .Y(core__abc_21380_n6162) );
  AND2X2 AND2X2_3676 ( .A(core__abc_21380_n6166), .B(reset_n_bF_buf14), .Y(core__abc_21380_n6167) );
  AND2X2 AND2X2_3677 ( .A(core__abc_21380_n6165), .B(core__abc_21380_n6167), .Y(core_v3_reg_50__FF_INPUT) );
  AND2X2 AND2X2_3678 ( .A(core__abc_21380_n6140), .B(core__abc_21380_n1596), .Y(core__abc_21380_n6170) );
  AND2X2 AND2X2_3679 ( .A(core__abc_21380_n6170), .B(core__abc_21380_n1621), .Y(core__abc_21380_n6171) );
  AND2X2 AND2X2_368 ( .A(_abc_19068_n916_1_bF_buf0), .B(word1_reg_28_), .Y(_abc_19068_n1547_1) );
  AND2X2 AND2X2_3680 ( .A(core__abc_21380_n6172), .B(core__abc_21380_n6173), .Y(core__abc_21380_n6174) );
  AND2X2 AND2X2_3681 ( .A(core__abc_21380_n6177), .B(core__abc_21380_n6176), .Y(core__abc_21380_n6178) );
  AND2X2 AND2X2_3682 ( .A(core__abc_21380_n3859), .B(core__abc_21380_n6174), .Y(core__abc_21380_n6181) );
  AND2X2 AND2X2_3683 ( .A(core__abc_21380_n3862), .B(core__abc_21380_n6175), .Y(core__abc_21380_n6182) );
  AND2X2 AND2X2_3684 ( .A(core__abc_21380_n6184), .B(core__abc_21380_n6179), .Y(core__abc_21380_n6185) );
  AND2X2 AND2X2_3685 ( .A(core__abc_21380_n6188), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n6189) );
  AND2X2 AND2X2_3686 ( .A(core__abc_21380_n6189), .B(core__abc_21380_n6187), .Y(core__abc_21380_n6190) );
  AND2X2 AND2X2_3687 ( .A(core__abc_21380_n3313_bF_buf12), .B(core_key_115_), .Y(core__abc_21380_n6191) );
  AND2X2 AND2X2_3688 ( .A(core_v3_reg_51_), .B(core_mi_51_), .Y(core__abc_21380_n6193) );
  AND2X2 AND2X2_3689 ( .A(core__abc_21380_n6194), .B(core__abc_21380_n6192), .Y(core__abc_21380_n6195) );
  AND2X2 AND2X2_369 ( .A(_abc_19068_n902_bF_buf0), .B(word2_reg_28_), .Y(_abc_19068_n1548) );
  AND2X2 AND2X2_3690 ( .A(core__abc_21380_n2749_bF_buf4), .B(core__abc_21380_n6195), .Y(core__abc_21380_n6196) );
  AND2X2 AND2X2_3691 ( .A(core__abc_21380_n6200), .B(reset_n_bF_buf13), .Y(core__abc_21380_n6201) );
  AND2X2 AND2X2_3692 ( .A(core__abc_21380_n6199), .B(core__abc_21380_n6201), .Y(core_v3_reg_51__FF_INPUT) );
  AND2X2 AND2X2_3693 ( .A(core__abc_21380_n6178), .B(core__abc_21380_n6148), .Y(core__abc_21380_n6203) );
  AND2X2 AND2X2_3694 ( .A(core__abc_21380_n6203), .B(core__abc_21380_n6132), .Y(core__abc_21380_n6204) );
  AND2X2 AND2X2_3695 ( .A(core__abc_21380_n6205), .B(core__abc_21380_n6177), .Y(core__abc_21380_n6206) );
  AND2X2 AND2X2_3696 ( .A(core__abc_21380_n6203), .B(core__abc_21380_n6133), .Y(core__abc_21380_n6208) );
  AND2X2 AND2X2_3697 ( .A(core__abc_21380_n6045), .B(core__abc_21380_n6208), .Y(core__abc_21380_n6209) );
  AND2X2 AND2X2_3698 ( .A(core__abc_21380_n3215_1), .B(core__abc_21380_n3229), .Y(core__abc_21380_n6212) );
  AND2X2 AND2X2_3699 ( .A(core__abc_21380_n6214), .B(core__abc_21380_n1632), .Y(core__abc_21380_n6215) );
  AND2X2 AND2X2_37 ( .A(_abc_19068_n926_bF_buf4), .B(core_key_0_), .Y(_abc_19068_n927_1) );
  AND2X2 AND2X2_370 ( .A(_abc_19068_n897_1_bF_buf0), .B(word0_reg_28_), .Y(_abc_19068_n1550) );
  AND2X2 AND2X2_3700 ( .A(core__abc_21380_n6213), .B(core__abc_21380_n1633), .Y(core__abc_21380_n6216) );
  AND2X2 AND2X2_3701 ( .A(core__abc_21380_n3928), .B(core__abc_21380_n6218), .Y(core__abc_21380_n6219) );
  AND2X2 AND2X2_3702 ( .A(core__abc_21380_n3927_1), .B(core__abc_21380_n6217), .Y(core__abc_21380_n6220) );
  AND2X2 AND2X2_3703 ( .A(core__abc_21380_n6211), .B(core__abc_21380_n6221), .Y(core__abc_21380_n6222) );
  AND2X2 AND2X2_3704 ( .A(core__abc_21380_n6210), .B(core__abc_21380_n6223), .Y(core__abc_21380_n6224) );
  AND2X2 AND2X2_3705 ( .A(core__abc_21380_n6228), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n6229) );
  AND2X2 AND2X2_3706 ( .A(core__abc_21380_n6229), .B(core__abc_21380_n6226), .Y(core__abc_21380_n6230) );
  AND2X2 AND2X2_3707 ( .A(core__abc_21380_n3313_bF_buf11), .B(core_key_116_), .Y(core__abc_21380_n6231) );
  AND2X2 AND2X2_3708 ( .A(core_v3_reg_52_), .B(core_mi_52_), .Y(core__abc_21380_n6233) );
  AND2X2 AND2X2_3709 ( .A(core__abc_21380_n6234), .B(core__abc_21380_n6232), .Y(core__abc_21380_n6235) );
  AND2X2 AND2X2_371 ( .A(_abc_19068_n915_1_bF_buf0), .B(core_mi_60_), .Y(_abc_19068_n1551_1) );
  AND2X2 AND2X2_3710 ( .A(core__abc_21380_n2749_bF_buf3), .B(core__abc_21380_n6235), .Y(core__abc_21380_n6236) );
  AND2X2 AND2X2_3711 ( .A(core__abc_21380_n6240), .B(reset_n_bF_buf12), .Y(core__abc_21380_n6241) );
  AND2X2 AND2X2_3712 ( .A(core__abc_21380_n6239), .B(core__abc_21380_n6241), .Y(core_v3_reg_52__FF_INPUT) );
  AND2X2 AND2X2_3713 ( .A(core__abc_21380_n6245), .B(core__abc_21380_n1650), .Y(core__abc_21380_n6246) );
  AND2X2 AND2X2_3714 ( .A(core__abc_21380_n6244), .B(core__abc_21380_n1651), .Y(core__abc_21380_n6247) );
  AND2X2 AND2X2_3715 ( .A(core__abc_21380_n3988_1), .B(core__abc_21380_n6249), .Y(core__abc_21380_n6250) );
  AND2X2 AND2X2_3716 ( .A(core__abc_21380_n3987), .B(core__abc_21380_n6248), .Y(core__abc_21380_n6251) );
  AND2X2 AND2X2_3717 ( .A(core__abc_21380_n6256), .B(core__abc_21380_n6254), .Y(core__abc_21380_n6257) );
  AND2X2 AND2X2_3718 ( .A(core__abc_21380_n6260), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n6261) );
  AND2X2 AND2X2_3719 ( .A(core__abc_21380_n6261), .B(core__abc_21380_n6258), .Y(core__abc_21380_n6262) );
  AND2X2 AND2X2_372 ( .A(_abc_19068_n923_bF_buf1), .B(_abc_19068_n1555_1), .Y(_auto_iopadmap_cc_313_execute_30317_28_) );
  AND2X2 AND2X2_3720 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n6263), .Y(core__abc_21380_n6264) );
  AND2X2 AND2X2_3721 ( .A(core_v3_reg_53_), .B(core_mi_53_), .Y(core__abc_21380_n6266) );
  AND2X2 AND2X2_3722 ( .A(core__abc_21380_n6267), .B(core__abc_21380_n6265), .Y(core__abc_21380_n6268) );
  AND2X2 AND2X2_3723 ( .A(core__abc_21380_n2749_bF_buf2), .B(core__abc_21380_n6268), .Y(core__abc_21380_n6269) );
  AND2X2 AND2X2_3724 ( .A(core__abc_21380_n6273), .B(reset_n_bF_buf11), .Y(core__abc_21380_n6274) );
  AND2X2 AND2X2_3725 ( .A(core__abc_21380_n6272), .B(core__abc_21380_n6274), .Y(core_v3_reg_53__FF_INPUT) );
  AND2X2 AND2X2_3726 ( .A(core__abc_21380_n6276), .B(core__abc_21380_n6278), .Y(core__abc_21380_n6279) );
  AND2X2 AND2X2_3727 ( .A(core__abc_21380_n6210), .B(core__abc_21380_n6282), .Y(core__abc_21380_n6283) );
  AND2X2 AND2X2_3728 ( .A(core__abc_21380_n6213), .B(core__abc_21380_n3225), .Y(core__abc_21380_n6286) );
  AND2X2 AND2X2_3729 ( .A(core__abc_21380_n6287), .B(core__abc_21380_n1669), .Y(core__abc_21380_n6288) );
  AND2X2 AND2X2_373 ( .A(_abc_19068_n945_1_bF_buf0), .B(core_mi_29_), .Y(_abc_19068_n1557) );
  AND2X2 AND2X2_3730 ( .A(core__abc_21380_n6289), .B(core__abc_21380_n6290), .Y(core__abc_21380_n6291) );
  AND2X2 AND2X2_3731 ( .A(core__abc_21380_n4046), .B(core__abc_21380_n6291), .Y(core__abc_21380_n6292) );
  AND2X2 AND2X2_3732 ( .A(core__abc_21380_n4047_1), .B(core__abc_21380_n6293), .Y(core__abc_21380_n6294) );
  AND2X2 AND2X2_3733 ( .A(core__abc_21380_n6285), .B(core__abc_21380_n6295), .Y(core__abc_21380_n6296) );
  AND2X2 AND2X2_3734 ( .A(core__abc_21380_n6284), .B(core__abc_21380_n6297), .Y(core__abc_21380_n6298) );
  AND2X2 AND2X2_3735 ( .A(core__abc_21380_n6302), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n6303) );
  AND2X2 AND2X2_3736 ( .A(core__abc_21380_n6303), .B(core__abc_21380_n6300), .Y(core__abc_21380_n6304) );
  AND2X2 AND2X2_3737 ( .A(core__abc_21380_n3313_bF_buf9), .B(core__abc_21380_n6305), .Y(core__abc_21380_n6306) );
  AND2X2 AND2X2_3738 ( .A(core_v3_reg_54_), .B(core_mi_54_), .Y(core__abc_21380_n6308) );
  AND2X2 AND2X2_3739 ( .A(core__abc_21380_n6309), .B(core__abc_21380_n6307), .Y(core__abc_21380_n6310) );
  AND2X2 AND2X2_374 ( .A(_abc_19068_n915_1_bF_buf4), .B(core_mi_61_), .Y(_abc_19068_n1558_1) );
  AND2X2 AND2X2_3740 ( .A(core__abc_21380_n2749_bF_buf1), .B(core__abc_21380_n6310), .Y(core__abc_21380_n6311) );
  AND2X2 AND2X2_3741 ( .A(core__abc_21380_n6315), .B(reset_n_bF_buf10), .Y(core__abc_21380_n6316) );
  AND2X2 AND2X2_3742 ( .A(core__abc_21380_n6314), .B(core__abc_21380_n6316), .Y(core_v3_reg_54__FF_INPUT) );
  AND2X2 AND2X2_3743 ( .A(core__abc_21380_n6319), .B(core__abc_21380_n1688), .Y(core__abc_21380_n6321) );
  AND2X2 AND2X2_3744 ( .A(core__abc_21380_n6322), .B(core__abc_21380_n6320), .Y(core__abc_21380_n6323) );
  AND2X2 AND2X2_3745 ( .A(core__abc_21380_n4132), .B(core__abc_21380_n6323), .Y(core__abc_21380_n6324) );
  AND2X2 AND2X2_3746 ( .A(core__abc_21380_n4136), .B(core__abc_21380_n6325), .Y(core__abc_21380_n6326) );
  AND2X2 AND2X2_3747 ( .A(core__abc_21380_n6331), .B(core__abc_21380_n6330), .Y(core__abc_21380_n6332) );
  AND2X2 AND2X2_3748 ( .A(core__abc_21380_n6333), .B(core__abc_21380_n6328), .Y(core__abc_21380_n6334) );
  AND2X2 AND2X2_3749 ( .A(core__abc_21380_n6337), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n6338) );
  AND2X2 AND2X2_375 ( .A(_abc_19068_n899_bF_buf4), .B(word3_reg_29_), .Y(_abc_19068_n1560) );
  AND2X2 AND2X2_3750 ( .A(core__abc_21380_n6338), .B(core__abc_21380_n6336), .Y(core__abc_21380_n6339) );
  AND2X2 AND2X2_3751 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_119_), .Y(core__abc_21380_n6340) );
  AND2X2 AND2X2_3752 ( .A(core_v3_reg_55_), .B(core_mi_55_), .Y(core__abc_21380_n6342) );
  AND2X2 AND2X2_3753 ( .A(core__abc_21380_n6343), .B(core__abc_21380_n6341), .Y(core__abc_21380_n6344) );
  AND2X2 AND2X2_3754 ( .A(core__abc_21380_n2749_bF_buf0), .B(core__abc_21380_n6344), .Y(core__abc_21380_n6345) );
  AND2X2 AND2X2_3755 ( .A(core__abc_21380_n6349), .B(reset_n_bF_buf9), .Y(core__abc_21380_n6350) );
  AND2X2 AND2X2_3756 ( .A(core__abc_21380_n6348), .B(core__abc_21380_n6350), .Y(core_v3_reg_55__FF_INPUT) );
  AND2X2 AND2X2_3757 ( .A(core__abc_21380_n6358), .B(core__abc_21380_n6359), .Y(core__abc_21380_n6360) );
  AND2X2 AND2X2_3758 ( .A(core__abc_21380_n6332), .B(core__abc_21380_n6297), .Y(core__abc_21380_n6362) );
  AND2X2 AND2X2_3759 ( .A(core__abc_21380_n6362), .B(core__abc_21380_n6280), .Y(core__abc_21380_n6363) );
  AND2X2 AND2X2_376 ( .A(_abc_19068_n902_bF_buf4), .B(word2_reg_29_), .Y(_abc_19068_n1561_1) );
  AND2X2 AND2X2_3760 ( .A(core__abc_21380_n6365), .B(core__abc_21380_n6330), .Y(core__abc_21380_n6366) );
  AND2X2 AND2X2_3761 ( .A(core__abc_21380_n6361), .B(core__abc_21380_n6369), .Y(core__abc_21380_n6370) );
  AND2X2 AND2X2_3762 ( .A(core__abc_21380_n6356), .B(core__abc_21380_n6370), .Y(core__abc_21380_n6371) );
  AND2X2 AND2X2_3763 ( .A(core__abc_21380_n3215_1), .B(core__abc_21380_n3230_1), .Y(core__abc_21380_n6372) );
  AND2X2 AND2X2_3764 ( .A(core__abc_21380_n6373), .B(core__abc_21380_n1707), .Y(core__abc_21380_n6374) );
  AND2X2 AND2X2_3765 ( .A(core__abc_21380_n6377), .B(core__abc_21380_n6375), .Y(core__abc_21380_n6378) );
  AND2X2 AND2X2_3766 ( .A(core__abc_21380_n6378), .B(core__abc_21380_n1706), .Y(core__abc_21380_n6379) );
  AND2X2 AND2X2_3767 ( .A(core__abc_21380_n4203_1), .B(core__abc_21380_n6381), .Y(core__abc_21380_n6382) );
  AND2X2 AND2X2_3768 ( .A(core__abc_21380_n4202), .B(core__abc_21380_n6380), .Y(core__abc_21380_n6383) );
  AND2X2 AND2X2_3769 ( .A(core__abc_21380_n6371), .B(core__abc_21380_n6384), .Y(core__abc_21380_n6385) );
  AND2X2 AND2X2_377 ( .A(_abc_19068_n926_bF_buf0), .B(core_key_29_), .Y(_abc_19068_n1564) );
  AND2X2 AND2X2_3770 ( .A(core__abc_21380_n6282), .B(core__abc_21380_n6362), .Y(core__abc_21380_n6386) );
  AND2X2 AND2X2_3771 ( .A(core__abc_21380_n6386), .B(core__abc_21380_n6208), .Y(core__abc_21380_n6387) );
  AND2X2 AND2X2_3772 ( .A(core__abc_21380_n6045), .B(core__abc_21380_n6387), .Y(core__abc_21380_n6388) );
  AND2X2 AND2X2_3773 ( .A(core__abc_21380_n6207), .B(core__abc_21380_n6386), .Y(core__abc_21380_n6389) );
  AND2X2 AND2X2_3774 ( .A(core__abc_21380_n6391), .B(core__abc_21380_n6392), .Y(core__abc_21380_n6393) );
  AND2X2 AND2X2_3775 ( .A(core__abc_21380_n6397), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n6398) );
  AND2X2 AND2X2_3776 ( .A(core__abc_21380_n6398), .B(core__abc_21380_n6396), .Y(core__abc_21380_n6399) );
  AND2X2 AND2X2_3777 ( .A(core__abc_21380_n3313_bF_buf7), .B(core_key_120_), .Y(core__abc_21380_n6400) );
  AND2X2 AND2X2_3778 ( .A(core_v3_reg_56_), .B(core_mi_56_), .Y(core__abc_21380_n6402) );
  AND2X2 AND2X2_3779 ( .A(core__abc_21380_n6403), .B(core__abc_21380_n6401), .Y(core__abc_21380_n6404) );
  AND2X2 AND2X2_378 ( .A(_abc_19068_n924_1_bF_buf0), .B(core_key_61_), .Y(_abc_19068_n1565_1) );
  AND2X2 AND2X2_3780 ( .A(core__abc_21380_n2749_bF_buf10), .B(core__abc_21380_n6404), .Y(core__abc_21380_n6405) );
  AND2X2 AND2X2_3781 ( .A(core__abc_21380_n6409), .B(reset_n_bF_buf8), .Y(core__abc_21380_n6410) );
  AND2X2 AND2X2_3782 ( .A(core__abc_21380_n6408), .B(core__abc_21380_n6410), .Y(core_v3_reg_56__FF_INPUT) );
  AND2X2 AND2X2_3783 ( .A(core__abc_21380_n6413), .B(core__abc_21380_n6412), .Y(core__abc_21380_n6414) );
  AND2X2 AND2X2_3784 ( .A(core__abc_21380_n6417), .B(core__abc_21380_n1732), .Y(core__abc_21380_n6418) );
  AND2X2 AND2X2_3785 ( .A(core__abc_21380_n6416), .B(core__abc_21380_n1726), .Y(core__abc_21380_n6419) );
  AND2X2 AND2X2_3786 ( .A(core__abc_21380_n4275), .B(core__abc_21380_n6421), .Y(core__abc_21380_n6422) );
  AND2X2 AND2X2_3787 ( .A(core__abc_21380_n4272), .B(core__abc_21380_n6420), .Y(core__abc_21380_n6424) );
  AND2X2 AND2X2_3788 ( .A(core__abc_21380_n6423), .B(core__abc_21380_n6425), .Y(core__abc_21380_n6426) );
  AND2X2 AND2X2_3789 ( .A(core__abc_21380_n6427), .B(core__abc_21380_n6429), .Y(core__abc_21380_n6430) );
  AND2X2 AND2X2_379 ( .A(_abc_19068_n941_bF_buf0), .B(core_key_125_), .Y(_abc_19068_n1567_1) );
  AND2X2 AND2X2_3790 ( .A(core__abc_21380_n6433), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n6434) );
  AND2X2 AND2X2_3791 ( .A(core__abc_21380_n6434), .B(core__abc_21380_n6431), .Y(core__abc_21380_n6435) );
  AND2X2 AND2X2_3792 ( .A(core__abc_21380_n3313_bF_buf6), .B(core_key_121_), .Y(core__abc_21380_n6436) );
  AND2X2 AND2X2_3793 ( .A(core_v3_reg_57_), .B(core_mi_57_), .Y(core__abc_21380_n6438) );
  AND2X2 AND2X2_3794 ( .A(core__abc_21380_n6439), .B(core__abc_21380_n6437), .Y(core__abc_21380_n6440) );
  AND2X2 AND2X2_3795 ( .A(core__abc_21380_n2749_bF_buf9), .B(core__abc_21380_n6440), .Y(core__abc_21380_n6441) );
  AND2X2 AND2X2_3796 ( .A(core__abc_21380_n6445), .B(reset_n_bF_buf7), .Y(core__abc_21380_n6446) );
  AND2X2 AND2X2_3797 ( .A(core__abc_21380_n6444), .B(core__abc_21380_n6446), .Y(core_v3_reg_57__FF_INPUT) );
  AND2X2 AND2X2_3798 ( .A(core__abc_21380_n6423), .B(core__abc_21380_n6448), .Y(core__abc_21380_n6449) );
  AND2X2 AND2X2_3799 ( .A(core__abc_21380_n6426), .B(core__abc_21380_n6392), .Y(core__abc_21380_n6451) );
  AND2X2 AND2X2_38 ( .A(_abc_19068_n882_1), .B(core_ready), .Y(_abc_19068_n929) );
  AND2X2 AND2X2_380 ( .A(_abc_19068_n939_1_bF_buf0), .B(core_key_93_), .Y(_abc_19068_n1568) );
  AND2X2 AND2X2_3800 ( .A(core__abc_21380_n6391), .B(core__abc_21380_n6451), .Y(core__abc_21380_n6452) );
  AND2X2 AND2X2_3801 ( .A(core__abc_21380_n6456), .B(core__abc_21380_n3252), .Y(core__abc_21380_n6457) );
  AND2X2 AND2X2_3802 ( .A(core__abc_21380_n6458), .B(core__abc_21380_n1743), .Y(core__abc_21380_n6459) );
  AND2X2 AND2X2_3803 ( .A(core__abc_21380_n6457), .B(core__abc_21380_n1749), .Y(core__abc_21380_n6460) );
  AND2X2 AND2X2_3804 ( .A(core__abc_21380_n4333), .B(core__abc_21380_n6462), .Y(core__abc_21380_n6463) );
  AND2X2 AND2X2_3805 ( .A(core__abc_21380_n4334_1), .B(core__abc_21380_n6461), .Y(core__abc_21380_n6464) );
  AND2X2 AND2X2_3806 ( .A(core__abc_21380_n6454), .B(core__abc_21380_n6465), .Y(core__abc_21380_n6466) );
  AND2X2 AND2X2_3807 ( .A(core__abc_21380_n6453), .B(core__abc_21380_n6467), .Y(core__abc_21380_n6468) );
  AND2X2 AND2X2_3808 ( .A(core__abc_21380_n6472), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n6473) );
  AND2X2 AND2X2_3809 ( .A(core__abc_21380_n6473), .B(core__abc_21380_n6471), .Y(core__abc_21380_n6474) );
  AND2X2 AND2X2_381 ( .A(_abc_19068_n897_1_bF_buf4), .B(word0_reg_29_), .Y(_abc_19068_n1571_1) );
  AND2X2 AND2X2_3810 ( .A(core__abc_21380_n3313_bF_buf5), .B(core__abc_21380_n6475), .Y(core__abc_21380_n6476) );
  AND2X2 AND2X2_3811 ( .A(core_v3_reg_58_), .B(core_mi_58_), .Y(core__abc_21380_n6478) );
  AND2X2 AND2X2_3812 ( .A(core__abc_21380_n6479), .B(core__abc_21380_n6477), .Y(core__abc_21380_n6480) );
  AND2X2 AND2X2_3813 ( .A(core__abc_21380_n2749_bF_buf8), .B(core__abc_21380_n6480), .Y(core__abc_21380_n6481) );
  AND2X2 AND2X2_3814 ( .A(core__abc_21380_n6485), .B(reset_n_bF_buf6), .Y(core__abc_21380_n6486) );
  AND2X2 AND2X2_3815 ( .A(core__abc_21380_n6484), .B(core__abc_21380_n6486), .Y(core_v3_reg_58__FF_INPUT) );
  AND2X2 AND2X2_3816 ( .A(core__abc_21380_n6490), .B(core__abc_21380_n1769), .Y(core__abc_21380_n6491) );
  AND2X2 AND2X2_3817 ( .A(core__abc_21380_n6489), .B(core__abc_21380_n1763), .Y(core__abc_21380_n6492) );
  AND2X2 AND2X2_3818 ( .A(core__abc_21380_n4430), .B(core__abc_21380_n6494), .Y(core__abc_21380_n6495) );
  AND2X2 AND2X2_3819 ( .A(core__abc_21380_n6496), .B(core__abc_21380_n6497), .Y(core__abc_21380_n6498) );
  AND2X2 AND2X2_382 ( .A(_abc_19068_n916_1_bF_buf4), .B(word1_reg_29_), .Y(_abc_19068_n1572) );
  AND2X2 AND2X2_3820 ( .A(core__abc_21380_n4426), .B(core__abc_21380_n6493), .Y(core__abc_21380_n6501) );
  AND2X2 AND2X2_3821 ( .A(core__abc_21380_n6503), .B(core__abc_21380_n6499), .Y(core__abc_21380_n6504) );
  AND2X2 AND2X2_3822 ( .A(core__abc_21380_n6507), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n6508) );
  AND2X2 AND2X2_3823 ( .A(core__abc_21380_n6508), .B(core__abc_21380_n6506), .Y(core__abc_21380_n6509) );
  AND2X2 AND2X2_3824 ( .A(core__abc_21380_n3313_bF_buf4), .B(core_key_123_), .Y(core__abc_21380_n6510) );
  AND2X2 AND2X2_3825 ( .A(core_v3_reg_59_), .B(core_mi_59_), .Y(core__abc_21380_n6512) );
  AND2X2 AND2X2_3826 ( .A(core__abc_21380_n6513), .B(core__abc_21380_n6511), .Y(core__abc_21380_n6514) );
  AND2X2 AND2X2_3827 ( .A(core__abc_21380_n2749_bF_buf7), .B(core__abc_21380_n6514), .Y(core__abc_21380_n6515) );
  AND2X2 AND2X2_3828 ( .A(core__abc_21380_n6519), .B(reset_n_bF_buf5), .Y(core__abc_21380_n6520) );
  AND2X2 AND2X2_3829 ( .A(core__abc_21380_n6518), .B(core__abc_21380_n6520), .Y(core_v3_reg_59__FF_INPUT) );
  AND2X2 AND2X2_383 ( .A(_abc_19068_n1576), .B(_abc_19068_n923_bF_buf0), .Y(_auto_iopadmap_cc_313_execute_30317_29_) );
  AND2X2 AND2X2_3830 ( .A(core__abc_21380_n6498), .B(core__abc_21380_n6467), .Y(core__abc_21380_n6522) );
  AND2X2 AND2X2_3831 ( .A(core__abc_21380_n6522), .B(core__abc_21380_n6451), .Y(core__abc_21380_n6523) );
  AND2X2 AND2X2_3832 ( .A(core__abc_21380_n6391), .B(core__abc_21380_n6523), .Y(core__abc_21380_n6524) );
  AND2X2 AND2X2_3833 ( .A(core__abc_21380_n6522), .B(core__abc_21380_n6450), .Y(core__abc_21380_n6525) );
  AND2X2 AND2X2_3834 ( .A(core__abc_21380_n6496), .B(core__abc_21380_n6526), .Y(core__abc_21380_n6527) );
  AND2X2 AND2X2_3835 ( .A(core__abc_21380_n6373), .B(core__abc_21380_n3221), .Y(core__abc_21380_n6532) );
  AND2X2 AND2X2_3836 ( .A(core__abc_21380_n6534), .B(core__abc_21380_n1781), .Y(core__abc_21380_n6535) );
  AND2X2 AND2X2_3837 ( .A(core__abc_21380_n6533), .B(core__abc_21380_n1782_1), .Y(core__abc_21380_n6536) );
  AND2X2 AND2X2_3838 ( .A(core__abc_21380_n4496_1), .B(core__abc_21380_n6537), .Y(core__abc_21380_n6538) );
  AND2X2 AND2X2_3839 ( .A(core__abc_21380_n4495), .B(core__abc_21380_n6539), .Y(core__abc_21380_n6540) );
  AND2X2 AND2X2_384 ( .A(_abc_19068_n899_bF_buf3), .B(word3_reg_30_), .Y(_abc_19068_n1578) );
  AND2X2 AND2X2_3840 ( .A(core__abc_21380_n6531), .B(core__abc_21380_n6542), .Y(core__abc_21380_n6543) );
  AND2X2 AND2X2_3841 ( .A(core__abc_21380_n6548), .B(core__abc_21380_n6528), .Y(core__abc_21380_n6549) );
  AND2X2 AND2X2_3842 ( .A(core__abc_21380_n6547), .B(core__abc_21380_n6549), .Y(core__abc_21380_n6550) );
  AND2X2 AND2X2_3843 ( .A(core__abc_21380_n6550), .B(core__abc_21380_n6541), .Y(core__abc_21380_n6551) );
  AND2X2 AND2X2_3844 ( .A(core__abc_21380_n6555), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n6556) );
  AND2X2 AND2X2_3845 ( .A(core__abc_21380_n6556), .B(core__abc_21380_n6554), .Y(core__abc_21380_n6557) );
  AND2X2 AND2X2_3846 ( .A(core__abc_21380_n3313_bF_buf3), .B(core__abc_21380_n6558), .Y(core__abc_21380_n6559) );
  AND2X2 AND2X2_3847 ( .A(core_v3_reg_60_), .B(core_mi_60_), .Y(core__abc_21380_n6561) );
  AND2X2 AND2X2_3848 ( .A(core__abc_21380_n6562), .B(core__abc_21380_n6560), .Y(core__abc_21380_n6563) );
  AND2X2 AND2X2_3849 ( .A(core__abc_21380_n2749_bF_buf6), .B(core__abc_21380_n6563), .Y(core__abc_21380_n6564) );
  AND2X2 AND2X2_385 ( .A(_abc_19068_n945_1_bF_buf4), .B(core_mi_30_), .Y(_abc_19068_n1580_1) );
  AND2X2 AND2X2_3850 ( .A(core__abc_21380_n6568), .B(reset_n_bF_buf4), .Y(core__abc_21380_n6569) );
  AND2X2 AND2X2_3851 ( .A(core__abc_21380_n6567), .B(core__abc_21380_n6569), .Y(core_v3_reg_60__FF_INPUT) );
  AND2X2 AND2X2_3852 ( .A(core__abc_21380_n6573), .B(core__abc_21380_n1807), .Y(core__abc_21380_n6574) );
  AND2X2 AND2X2_3853 ( .A(core__abc_21380_n6572), .B(core__abc_21380_n1801), .Y(core__abc_21380_n6575) );
  AND2X2 AND2X2_3854 ( .A(core__abc_21380_n4554), .B(core__abc_21380_n6577), .Y(core__abc_21380_n6578) );
  AND2X2 AND2X2_3855 ( .A(core__abc_21380_n6584), .B(core__abc_21380_n6579), .Y(core__abc_21380_n6585) );
  AND2X2 AND2X2_3856 ( .A(core__abc_21380_n6586), .B(core__abc_21380_n6582), .Y(core__abc_21380_n6587) );
  AND2X2 AND2X2_3857 ( .A(core__abc_21380_n6590), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf3), .Y(core__abc_21380_n6591) );
  AND2X2 AND2X2_3858 ( .A(core__abc_21380_n6591), .B(core__abc_21380_n6589), .Y(core__abc_21380_n6592) );
  AND2X2 AND2X2_3859 ( .A(core__abc_21380_n3313_bF_buf2), .B(core__abc_21380_n6593), .Y(core__abc_21380_n6594) );
  AND2X2 AND2X2_386 ( .A(_abc_19068_n941_bF_buf4), .B(core_key_126_), .Y(_abc_19068_n1581) );
  AND2X2 AND2X2_3860 ( .A(core_v3_reg_61_), .B(core_mi_61_), .Y(core__abc_21380_n6596) );
  AND2X2 AND2X2_3861 ( .A(core__abc_21380_n6597), .B(core__abc_21380_n6595), .Y(core__abc_21380_n6598) );
  AND2X2 AND2X2_3862 ( .A(core__abc_21380_n2749_bF_buf5), .B(core__abc_21380_n6598), .Y(core__abc_21380_n6599) );
  AND2X2 AND2X2_3863 ( .A(core__abc_21380_n6603), .B(reset_n_bF_buf3), .Y(core__abc_21380_n6604) );
  AND2X2 AND2X2_3864 ( .A(core__abc_21380_n6602), .B(core__abc_21380_n6604), .Y(core_v3_reg_61__FF_INPUT) );
  AND2X2 AND2X2_3865 ( .A(core__abc_21380_n6585), .B(core__abc_21380_n6542), .Y(core__abc_21380_n6606) );
  AND2X2 AND2X2_3866 ( .A(core__abc_21380_n6531), .B(core__abc_21380_n6606), .Y(core__abc_21380_n6607) );
  AND2X2 AND2X2_3867 ( .A(core__abc_21380_n6585), .B(core__abc_21380_n6540), .Y(core__abc_21380_n6608) );
  AND2X2 AND2X2_3868 ( .A(core__abc_21380_n6533), .B(core__abc_21380_n3217), .Y(core__abc_21380_n6611) );
  AND2X2 AND2X2_3869 ( .A(core__abc_21380_n6612), .B(core__abc_21380_n1820), .Y(core__abc_21380_n6613) );
  AND2X2 AND2X2_387 ( .A(_abc_19068_n939_1_bF_buf4), .B(core_key_94_), .Y(_abc_19068_n1584) );
  AND2X2 AND2X2_3870 ( .A(core__abc_21380_n6614), .B(core__abc_21380_n6615), .Y(core__abc_21380_n6616) );
  AND2X2 AND2X2_3871 ( .A(core__abc_21380_n4616), .B(core__abc_21380_n6616), .Y(core__abc_21380_n6617) );
  AND2X2 AND2X2_3872 ( .A(core__abc_21380_n4585), .B(core__abc_21380_n6618), .Y(core__abc_21380_n6619) );
  AND2X2 AND2X2_3873 ( .A(core__abc_21380_n6625), .B(core__abc_21380_n6584), .Y(core__abc_21380_n6626) );
  AND2X2 AND2X2_3874 ( .A(core__abc_21380_n6624), .B(core__abc_21380_n6626), .Y(core__abc_21380_n6627) );
  AND2X2 AND2X2_3875 ( .A(core__abc_21380_n6628), .B(core__abc_21380_n6622), .Y(core__abc_21380_n6629) );
  AND2X2 AND2X2_3876 ( .A(core__abc_21380_n6632), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf3), .Y(core__abc_21380_n6633) );
  AND2X2 AND2X2_3877 ( .A(core__abc_21380_n6633), .B(core__abc_21380_n6631), .Y(core__abc_21380_n6634) );
  AND2X2 AND2X2_3878 ( .A(core__abc_21380_n3313_bF_buf1), .B(core__abc_21380_n6635), .Y(core__abc_21380_n6636) );
  AND2X2 AND2X2_3879 ( .A(core_v3_reg_62_), .B(core_mi_62_), .Y(core__abc_21380_n6638) );
  AND2X2 AND2X2_388 ( .A(_abc_19068_n924_1_bF_buf4), .B(core_key_62_), .Y(_abc_19068_n1585) );
  AND2X2 AND2X2_3880 ( .A(core__abc_21380_n6639), .B(core__abc_21380_n6637), .Y(core__abc_21380_n6640) );
  AND2X2 AND2X2_3881 ( .A(core__abc_21380_n2749_bF_buf4), .B(core__abc_21380_n6640), .Y(core__abc_21380_n6641) );
  AND2X2 AND2X2_3882 ( .A(core__abc_21380_n6645), .B(reset_n_bF_buf2), .Y(core__abc_21380_n6646) );
  AND2X2 AND2X2_3883 ( .A(core__abc_21380_n6644), .B(core__abc_21380_n6646), .Y(core_v3_reg_62__FF_INPUT) );
  AND2X2 AND2X2_3884 ( .A(core__abc_21380_n6610), .B(core__abc_21380_n6621), .Y(core__abc_21380_n6648) );
  AND2X2 AND2X2_3885 ( .A(core__abc_21380_n6650), .B(core__abc_21380_n1839), .Y(core__abc_21380_n6652) );
  AND2X2 AND2X2_3886 ( .A(core__abc_21380_n6653), .B(core__abc_21380_n6651), .Y(core__abc_21380_n6654) );
  AND2X2 AND2X2_3887 ( .A(core__abc_21380_n4684), .B(core__abc_21380_n6654), .Y(core__abc_21380_n6655) );
  AND2X2 AND2X2_3888 ( .A(core__abc_21380_n4689), .B(core__abc_21380_n6657), .Y(core__abc_21380_n6658) );
  AND2X2 AND2X2_3889 ( .A(core__abc_21380_n6656), .B(core__abc_21380_n6659), .Y(core__abc_21380_n6660) );
  AND2X2 AND2X2_389 ( .A(_abc_19068_n926_bF_buf4), .B(core_key_30_), .Y(_abc_19068_n1586) );
  AND2X2 AND2X2_3890 ( .A(core__abc_21380_n6628), .B(core__abc_21380_n6662), .Y(core__abc_21380_n6663) );
  AND2X2 AND2X2_3891 ( .A(core__abc_21380_n6665), .B(core__abc_21380_n6661), .Y(core__abc_21380_n6666) );
  AND2X2 AND2X2_3892 ( .A(core__abc_21380_n6669), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n6670) );
  AND2X2 AND2X2_3893 ( .A(core__abc_21380_n6670), .B(core__abc_21380_n6668), .Y(core__abc_21380_n6671) );
  AND2X2 AND2X2_3894 ( .A(core__abc_21380_n3313_bF_buf0), .B(core_key_127_), .Y(core__abc_21380_n6672) );
  AND2X2 AND2X2_3895 ( .A(core_v3_reg_63_), .B(core_mi_63_), .Y(core__abc_21380_n6674) );
  AND2X2 AND2X2_3896 ( .A(core__abc_21380_n6675), .B(core__abc_21380_n6673), .Y(core__abc_21380_n6676) );
  AND2X2 AND2X2_3897 ( .A(core__abc_21380_n2749_bF_buf3), .B(core__abc_21380_n6676), .Y(core__abc_21380_n6677) );
  AND2X2 AND2X2_3898 ( .A(core__abc_21380_n6681), .B(reset_n_bF_buf1), .Y(core__abc_21380_n6682) );
  AND2X2 AND2X2_3899 ( .A(core__abc_21380_n6680), .B(core__abc_21380_n6682), .Y(core_v3_reg_63__FF_INPUT) );
  AND2X2 AND2X2_39 ( .A(_abc_19068_n885_1), .B(core_compression_rounds_0_), .Y(_abc_19068_n930_1) );
  AND2X2 AND2X2_390 ( .A(_abc_19068_n916_1_bF_buf3), .B(word1_reg_30_), .Y(_abc_19068_n1589_1) );
  AND2X2 AND2X2_3900 ( .A(core__abc_21380_n6654), .B(core__abc_21380_n6684), .Y(core__abc_21380_n6686) );
  AND2X2 AND2X2_3901 ( .A(core__abc_21380_n6687), .B(core__abc_21380_n6685), .Y(core__abc_21380_n6688) );
  AND2X2 AND2X2_3902 ( .A(core__abc_21380_n6692), .B(core__abc_21380_n6689), .Y(core__abc_21380_n6693) );
  AND2X2 AND2X2_3903 ( .A(core__abc_21380_n6695), .B(core__abc_21380_n6694), .Y(core__abc_21380_n6696) );
  AND2X2 AND2X2_3904 ( .A(core__abc_21380_n6697), .B(core__abc_21380_n5215), .Y(core__abc_21380_n6698) );
  AND2X2 AND2X2_3905 ( .A(core__abc_21380_n6696), .B(core__abc_21380_n5214), .Y(core__abc_21380_n6699) );
  AND2X2 AND2X2_3906 ( .A(core__abc_21380_n6693), .B(core__abc_21380_n6701), .Y(core__abc_21380_n6702) );
  AND2X2 AND2X2_3907 ( .A(core__abc_21380_n6576), .B(core__abc_21380_n1558), .Y(core__abc_21380_n6704) );
  AND2X2 AND2X2_3908 ( .A(core__abc_21380_n6577), .B(core_v1_reg_16_), .Y(core__abc_21380_n6705) );
  AND2X2 AND2X2_3909 ( .A(core__abc_21380_n6707), .B(core__abc_21380_n6703), .Y(core__abc_21380_n6708) );
  AND2X2 AND2X2_391 ( .A(_abc_19068_n902_bF_buf3), .B(word2_reg_30_), .Y(_abc_19068_n1590) );
  AND2X2 AND2X2_3910 ( .A(core__abc_21380_n6706), .B(core__abc_21380_n5155), .Y(core__abc_21380_n6710) );
  AND2X2 AND2X2_3911 ( .A(core__abc_21380_n6709), .B(core__abc_21380_n6711), .Y(core__abc_21380_n6712) );
  AND2X2 AND2X2_3912 ( .A(core__abc_21380_n6713), .B(core__abc_21380_n6714), .Y(core__abc_21380_n6715) );
  AND2X2 AND2X2_3913 ( .A(core__abc_21380_n6716), .B(core__abc_21380_n5109), .Y(core__abc_21380_n6717) );
  AND2X2 AND2X2_3914 ( .A(core__abc_21380_n6715), .B(core__abc_21380_n5108), .Y(core__abc_21380_n6718) );
  AND2X2 AND2X2_3915 ( .A(core__abc_21380_n6712), .B(core__abc_21380_n6720), .Y(core__abc_21380_n6721) );
  AND2X2 AND2X2_3916 ( .A(core__abc_21380_n6702), .B(core__abc_21380_n6721), .Y(core__abc_21380_n6722) );
  AND2X2 AND2X2_3917 ( .A(core__abc_21380_n6493), .B(core_v1_reg_14_), .Y(core__abc_21380_n6723) );
  AND2X2 AND2X2_3918 ( .A(core__abc_21380_n6724), .B(core__abc_21380_n6725), .Y(core__abc_21380_n6726) );
  AND2X2 AND2X2_3919 ( .A(core__abc_21380_n6726), .B(core__abc_21380_n5037), .Y(core__abc_21380_n6728) );
  AND2X2 AND2X2_392 ( .A(_abc_19068_n897_1_bF_buf3), .B(word0_reg_30_), .Y(_abc_19068_n1592) );
  AND2X2 AND2X2_3920 ( .A(core__abc_21380_n6729), .B(core__abc_21380_n6727), .Y(core__abc_21380_n6730) );
  AND2X2 AND2X2_3921 ( .A(core__abc_21380_n6731), .B(core__abc_21380_n6732), .Y(core__abc_21380_n6733) );
  AND2X2 AND2X2_3922 ( .A(core__abc_21380_n6734), .B(core__abc_21380_n4987), .Y(core__abc_21380_n6735) );
  AND2X2 AND2X2_3923 ( .A(core__abc_21380_n6733), .B(core__abc_21380_n4986), .Y(core__abc_21380_n6736) );
  AND2X2 AND2X2_3924 ( .A(core__abc_21380_n6730), .B(core__abc_21380_n6738), .Y(core__abc_21380_n6739) );
  AND2X2 AND2X2_3925 ( .A(core__abc_21380_n6420), .B(core__abc_21380_n1484), .Y(core__abc_21380_n6740) );
  AND2X2 AND2X2_3926 ( .A(core__abc_21380_n6421), .B(core_v1_reg_12_), .Y(core__abc_21380_n6741) );
  AND2X2 AND2X2_3927 ( .A(core__abc_21380_n6742), .B(core__abc_21380_n4942), .Y(core__abc_21380_n6743) );
  AND2X2 AND2X2_3928 ( .A(core__abc_21380_n6745), .B(core__abc_21380_n4944), .Y(core__abc_21380_n6746) );
  AND2X2 AND2X2_3929 ( .A(core__abc_21380_n6749), .B(core__abc_21380_n6750), .Y(core__abc_21380_n6751) );
  AND2X2 AND2X2_393 ( .A(_abc_19068_n915_1_bF_buf3), .B(core_mi_62_), .Y(_abc_19068_n1593) );
  AND2X2 AND2X2_3930 ( .A(core__abc_21380_n6752), .B(core__abc_21380_n4896_1), .Y(core__abc_21380_n6753) );
  AND2X2 AND2X2_3931 ( .A(core__abc_21380_n6747), .B(core__abc_21380_n6754), .Y(core__abc_21380_n6755) );
  AND2X2 AND2X2_3932 ( .A(core__abc_21380_n6756), .B(core__abc_21380_n6744), .Y(core__abc_21380_n6757) );
  AND2X2 AND2X2_3933 ( .A(core__abc_21380_n6739), .B(core__abc_21380_n6757), .Y(core__abc_21380_n6758) );
  AND2X2 AND2X2_3934 ( .A(core__abc_21380_n6760), .B(core__abc_21380_n6727), .Y(core__abc_21380_n6761) );
  AND2X2 AND2X2_3935 ( .A(core__abc_21380_n6763), .B(core__abc_21380_n6722), .Y(core__abc_21380_n6764) );
  AND2X2 AND2X2_3936 ( .A(core__abc_21380_n6709), .B(core__abc_21380_n6765), .Y(core__abc_21380_n6766) );
  AND2X2 AND2X2_3937 ( .A(core__abc_21380_n6767), .B(core__abc_21380_n6711), .Y(core__abc_21380_n6768) );
  AND2X2 AND2X2_3938 ( .A(core__abc_21380_n6702), .B(core__abc_21380_n6768), .Y(core__abc_21380_n6769) );
  AND2X2 AND2X2_3939 ( .A(core__abc_21380_n6688), .B(core__abc_21380_n5261), .Y(core__abc_21380_n6770) );
  AND2X2 AND2X2_394 ( .A(_abc_19068_n923_bF_buf4), .B(_abc_19068_n1597), .Y(_auto_iopadmap_cc_313_execute_30317_30_) );
  AND2X2 AND2X2_3940 ( .A(core__abc_21380_n6772), .B(core__abc_21380_n6689), .Y(core__abc_21380_n6773) );
  AND2X2 AND2X2_3941 ( .A(core__abc_21380_n6747), .B(core__abc_21380_n6744), .Y(core__abc_21380_n6777) );
  AND2X2 AND2X2_3942 ( .A(core__abc_21380_n6751), .B(core__abc_21380_n4895), .Y(core__abc_21380_n6778) );
  AND2X2 AND2X2_3943 ( .A(core__abc_21380_n6777), .B(core__abc_21380_n6780), .Y(core__abc_21380_n6781) );
  AND2X2 AND2X2_3944 ( .A(core__abc_21380_n6739), .B(core__abc_21380_n6781), .Y(core__abc_21380_n6782) );
  AND2X2 AND2X2_3945 ( .A(core__abc_21380_n6722), .B(core__abc_21380_n6782), .Y(core__abc_21380_n6783) );
  AND2X2 AND2X2_3946 ( .A(core__abc_21380_n6323), .B(core__abc_21380_n6784), .Y(core__abc_21380_n6786) );
  AND2X2 AND2X2_3947 ( .A(core__abc_21380_n6787), .B(core__abc_21380_n6785), .Y(core__abc_21380_n6788) );
  AND2X2 AND2X2_3948 ( .A(core__abc_21380_n6325), .B(core_v1_reg_10_), .Y(core__abc_21380_n6791) );
  AND2X2 AND2X2_3949 ( .A(core__abc_21380_n6793), .B(core__abc_21380_n6789), .Y(core__abc_21380_n6794) );
  AND2X2 AND2X2_395 ( .A(_abc_19068_n916_1_bF_buf2), .B(word1_reg_31_), .Y(_abc_19068_n1599) );
  AND2X2 AND2X2_3950 ( .A(core__abc_21380_n6796), .B(core__abc_21380_n6795), .Y(core__abc_21380_n6797) );
  AND2X2 AND2X2_3951 ( .A(core__abc_21380_n6798), .B(core__abc_21380_n4772_1), .Y(core__abc_21380_n6799) );
  AND2X2 AND2X2_3952 ( .A(core__abc_21380_n6797), .B(core__abc_21380_n4771), .Y(core__abc_21380_n6800) );
  AND2X2 AND2X2_3953 ( .A(core__abc_21380_n6794), .B(core__abc_21380_n6802), .Y(core__abc_21380_n6803) );
  AND2X2 AND2X2_3954 ( .A(core__abc_21380_n6248), .B(core__abc_21380_n6804), .Y(core__abc_21380_n6805) );
  AND2X2 AND2X2_3955 ( .A(core__abc_21380_n6249), .B(core_v1_reg_8_), .Y(core__abc_21380_n6806) );
  AND2X2 AND2X2_3956 ( .A(core__abc_21380_n6808), .B(core__abc_21380_n4718), .Y(core__abc_21380_n6809) );
  AND2X2 AND2X2_3957 ( .A(core__abc_21380_n6807), .B(core__abc_21380_n4716), .Y(core__abc_21380_n6811) );
  AND2X2 AND2X2_3958 ( .A(core__abc_21380_n6810), .B(core__abc_21380_n6812), .Y(core__abc_21380_n6813) );
  AND2X2 AND2X2_3959 ( .A(core__abc_21380_n6814), .B(core__abc_21380_n6815), .Y(core__abc_21380_n6816) );
  AND2X2 AND2X2_396 ( .A(_abc_19068_n897_1_bF_buf2), .B(word0_reg_31_), .Y(_abc_19068_n1600) );
  AND2X2 AND2X2_3960 ( .A(core__abc_21380_n6817), .B(core__abc_21380_n4651), .Y(core__abc_21380_n6818) );
  AND2X2 AND2X2_3961 ( .A(core__abc_21380_n6816), .B(core__abc_21380_n4650_1), .Y(core__abc_21380_n6819) );
  AND2X2 AND2X2_3962 ( .A(core__abc_21380_n6813), .B(core__abc_21380_n6821), .Y(core__abc_21380_n6822) );
  AND2X2 AND2X2_3963 ( .A(core__abc_21380_n6803), .B(core__abc_21380_n6822), .Y(core__abc_21380_n6823) );
  AND2X2 AND2X2_3964 ( .A(core__abc_21380_n6175), .B(core_v1_reg_6_), .Y(core__abc_21380_n6824) );
  AND2X2 AND2X2_3965 ( .A(core__abc_21380_n6174), .B(core__abc_21380_n1374), .Y(core__abc_21380_n6825) );
  AND2X2 AND2X2_3966 ( .A(core__abc_21380_n6826), .B(core__abc_21380_n4599), .Y(core__abc_21380_n6827) );
  AND2X2 AND2X2_3967 ( .A(core__abc_21380_n6828), .B(core__abc_21380_n6829), .Y(core__abc_21380_n6830) );
  AND2X2 AND2X2_3968 ( .A(core__abc_21380_n6832), .B(core__abc_21380_n6831), .Y(core__abc_21380_n6833) );
  AND2X2 AND2X2_3969 ( .A(core__abc_21380_n6834), .B(core__abc_21380_n4534), .Y(core__abc_21380_n6835) );
  AND2X2 AND2X2_397 ( .A(_abc_19068_n939_1_bF_buf3), .B(core_key_95_), .Y(_abc_19068_n1602) );
  AND2X2 AND2X2_3970 ( .A(core__abc_21380_n6833), .B(core__abc_21380_n4533), .Y(core__abc_21380_n6836) );
  AND2X2 AND2X2_3971 ( .A(core__abc_21380_n6830), .B(core__abc_21380_n6838), .Y(core__abc_21380_n6839) );
  AND2X2 AND2X2_3972 ( .A(core__abc_21380_n6102), .B(core__abc_21380_n6840), .Y(core__abc_21380_n6841) );
  AND2X2 AND2X2_3973 ( .A(core__abc_21380_n6103), .B(core_v1_reg_4_), .Y(core__abc_21380_n6842) );
  AND2X2 AND2X2_3974 ( .A(core__abc_21380_n6844), .B(core__abc_21380_n4468), .Y(core__abc_21380_n6845) );
  AND2X2 AND2X2_3975 ( .A(core__abc_21380_n6846), .B(core__abc_21380_n6847), .Y(core__abc_21380_n6848) );
  AND2X2 AND2X2_3976 ( .A(core__abc_21380_n6849), .B(core__abc_21380_n4397_1), .Y(core__abc_21380_n6850) );
  AND2X2 AND2X2_3977 ( .A(core__abc_21380_n6843), .B(core__abc_21380_n4466), .Y(core__abc_21380_n6851) );
  AND2X2 AND2X2_3978 ( .A(core__abc_21380_n6852), .B(core__abc_21380_n6850), .Y(core__abc_21380_n6853) );
  AND2X2 AND2X2_3979 ( .A(core__abc_21380_n6839), .B(core__abc_21380_n6854), .Y(core__abc_21380_n6855) );
  AND2X2 AND2X2_398 ( .A(_abc_19068_n924_1_bF_buf3), .B(core_key_63_), .Y(_abc_19068_n1603) );
  AND2X2 AND2X2_3980 ( .A(core__abc_21380_n6828), .B(core__abc_21380_n6857), .Y(core__abc_21380_n6858) );
  AND2X2 AND2X2_3981 ( .A(core__abc_21380_n6823), .B(core__abc_21380_n6861), .Y(core__abc_21380_n6862) );
  AND2X2 AND2X2_3982 ( .A(core__abc_21380_n6810), .B(core__abc_21380_n6863), .Y(core__abc_21380_n6864) );
  AND2X2 AND2X2_3983 ( .A(core__abc_21380_n6865), .B(core__abc_21380_n6812), .Y(core__abc_21380_n6866) );
  AND2X2 AND2X2_3984 ( .A(core__abc_21380_n6803), .B(core__abc_21380_n6866), .Y(core__abc_21380_n6867) );
  AND2X2 AND2X2_3985 ( .A(core__abc_21380_n6788), .B(core__abc_21380_n4814_1), .Y(core__abc_21380_n6868) );
  AND2X2 AND2X2_3986 ( .A(core__abc_21380_n6870), .B(core__abc_21380_n6789), .Y(core__abc_21380_n6871) );
  AND2X2 AND2X2_3987 ( .A(core__abc_21380_n6001), .B(core_v1_reg_2_), .Y(core__abc_21380_n6875) );
  AND2X2 AND2X2_3988 ( .A(core__abc_21380_n6002), .B(core__abc_21380_n1299), .Y(core__abc_21380_n6876) );
  AND2X2 AND2X2_3989 ( .A(core__abc_21380_n6877), .B(core__abc_21380_n4308), .Y(core__abc_21380_n6878) );
  AND2X2 AND2X2_399 ( .A(_abc_19068_n926_bF_buf3), .B(core_key_31_), .Y(_abc_19068_n1604) );
  AND2X2 AND2X2_3990 ( .A(core__abc_21380_n6879), .B(core__abc_21380_n6880), .Y(core__abc_21380_n6881) );
  AND2X2 AND2X2_3991 ( .A(core__abc_21380_n6883), .B(core__abc_21380_n6882), .Y(core__abc_21380_n6884) );
  AND2X2 AND2X2_3992 ( .A(core__abc_21380_n6885), .B(core__abc_21380_n4243_1), .Y(core__abc_21380_n6886) );
  AND2X2 AND2X2_3993 ( .A(core__abc_21380_n6884), .B(core__abc_21380_n4242), .Y(core__abc_21380_n6887) );
  AND2X2 AND2X2_3994 ( .A(core__abc_21380_n6881), .B(core__abc_21380_n6889), .Y(core__abc_21380_n6890) );
  AND2X2 AND2X2_3995 ( .A(core__abc_21380_n5925), .B(core__abc_21380_n6891), .Y(core__abc_21380_n6892) );
  AND2X2 AND2X2_3996 ( .A(core__abc_21380_n5927), .B(core_v1_reg_0_), .Y(core__abc_21380_n6893) );
  AND2X2 AND2X2_3997 ( .A(core__abc_21380_n6894), .B(core__abc_21380_n4166), .Y(core__abc_21380_n6895) );
  AND2X2 AND2X2_3998 ( .A(core__abc_21380_n6896), .B(core__abc_21380_n4168), .Y(core__abc_21380_n6897) );
  AND2X2 AND2X2_3999 ( .A(core__abc_21380_n6899), .B(core__abc_21380_n6900), .Y(core__abc_21380_n6901) );
  AND2X2 AND2X2_4 ( .A(_abc_19068_n875), .B(_abc_19068_n876_1), .Y(_abc_19068_n877_1) );
  AND2X2 AND2X2_40 ( .A(_abc_19068_n902_bF_buf3), .B(word2_reg_0_), .Y(_abc_19068_n933_1) );
  AND2X2 AND2X2_400 ( .A(_abc_19068_n941_bF_buf3), .B(core_key_127_), .Y(_abc_19068_n1608) );
  AND2X2 AND2X2_4000 ( .A(core__abc_21380_n6902), .B(core__abc_21380_n4107), .Y(core__abc_21380_n6903) );
  AND2X2 AND2X2_4001 ( .A(core__abc_21380_n6898), .B(core__abc_21380_n6904), .Y(core__abc_21380_n6905) );
  AND2X2 AND2X2_4002 ( .A(core__abc_21380_n6890), .B(core__abc_21380_n6907), .Y(core__abc_21380_n6908) );
  AND2X2 AND2X2_4003 ( .A(core__abc_21380_n6909), .B(core__abc_21380_n6880), .Y(core__abc_21380_n6910) );
  AND2X2 AND2X2_4004 ( .A(core__abc_21380_n6898), .B(core__abc_21380_n6912), .Y(core__abc_21380_n6913) );
  AND2X2 AND2X2_4005 ( .A(core__abc_21380_n6901), .B(core__abc_21380_n4106_1), .Y(core__abc_21380_n6914) );
  AND2X2 AND2X2_4006 ( .A(core__abc_21380_n6913), .B(core__abc_21380_n6916), .Y(core__abc_21380_n6917) );
  AND2X2 AND2X2_4007 ( .A(core__abc_21380_n6890), .B(core__abc_21380_n6917), .Y(core__abc_21380_n6918) );
  AND2X2 AND2X2_4008 ( .A(core__abc_21380_n5848), .B(core__abc_21380_n2413), .Y(core__abc_21380_n6920) );
  AND2X2 AND2X2_4009 ( .A(core__abc_21380_n6921), .B(core__abc_21380_n6919), .Y(core__abc_21380_n6922) );
  AND2X2 AND2X2_401 ( .A(_abc_19068_n902_bF_buf2), .B(word2_reg_31_), .Y(_abc_19068_n1609) );
  AND2X2 AND2X2_4010 ( .A(core__abc_21380_n6922), .B(core__abc_21380_n4018_1), .Y(core__abc_21380_n6923) );
  AND2X2 AND2X2_4011 ( .A(core__abc_21380_n6925), .B(core__abc_21380_n6924), .Y(core__abc_21380_n6926) );
  AND2X2 AND2X2_4012 ( .A(core__abc_21380_n6927), .B(core__abc_21380_n3961_1), .Y(core__abc_21380_n6928) );
  AND2X2 AND2X2_4013 ( .A(core__abc_21380_n6930), .B(core__abc_21380_n6929), .Y(core__abc_21380_n6931) );
  AND2X2 AND2X2_4014 ( .A(core__abc_21380_n5759), .B(core__abc_21380_n2377), .Y(core__abc_21380_n6934) );
  AND2X2 AND2X2_4015 ( .A(core__abc_21380_n5760), .B(core_v1_reg_60_), .Y(core__abc_21380_n6935) );
  AND2X2 AND2X2_4016 ( .A(core__abc_21380_n6937), .B(core__abc_21380_n3898_1), .Y(core__abc_21380_n6938) );
  AND2X2 AND2X2_4017 ( .A(core__abc_21380_n6936), .B(core__abc_21380_n3896), .Y(core__abc_21380_n6940) );
  AND2X2 AND2X2_4018 ( .A(core__abc_21380_n6941), .B(core__abc_21380_n6942), .Y(core__abc_21380_n6943) );
  AND2X2 AND2X2_4019 ( .A(core__abc_21380_n6944), .B(core__abc_21380_n3821), .Y(core__abc_21380_n6945) );
  AND2X2 AND2X2_402 ( .A(_abc_19068_n899_bF_buf2), .B(word3_reg_31_), .Y(_abc_19068_n1610) );
  AND2X2 AND2X2_4020 ( .A(core__abc_21380_n6939), .B(core__abc_21380_n6947), .Y(core__abc_21380_n6948) );
  AND2X2 AND2X2_4021 ( .A(core__abc_21380_n6950), .B(core__abc_21380_n6930), .Y(core__abc_21380_n6951) );
  AND2X2 AND2X2_4022 ( .A(core__abc_21380_n6926), .B(core__abc_21380_n3960), .Y(core__abc_21380_n6952) );
  AND2X2 AND2X2_4023 ( .A(core__abc_21380_n6951), .B(core__abc_21380_n6954), .Y(core__abc_21380_n6955) );
  AND2X2 AND2X2_4024 ( .A(core__abc_21380_n6955), .B(core__abc_21380_n6949), .Y(core__abc_21380_n6956) );
  AND2X2 AND2X2_4025 ( .A(core__abc_21380_n5679), .B(core_v1_reg_58_), .Y(core__abc_21380_n6958) );
  AND2X2 AND2X2_4026 ( .A(core__abc_21380_n5662), .B(core__abc_21380_n2339), .Y(core__abc_21380_n6959) );
  AND2X2 AND2X2_4027 ( .A(core__abc_21380_n6960), .B(core__abc_21380_n3754), .Y(core__abc_21380_n6961) );
  AND2X2 AND2X2_4028 ( .A(core__abc_21380_n6962), .B(core__abc_21380_n3752_1), .Y(core__abc_21380_n6963) );
  AND2X2 AND2X2_4029 ( .A(core__abc_21380_n6966), .B(core__abc_21380_n6965), .Y(core__abc_21380_n6967) );
  AND2X2 AND2X2_403 ( .A(_abc_19068_n945_1_bF_buf3), .B(core_mi_31_), .Y(_abc_19068_n1612) );
  AND2X2 AND2X2_4030 ( .A(core__abc_21380_n6968), .B(core__abc_21380_n3694), .Y(core__abc_21380_n6969) );
  AND2X2 AND2X2_4031 ( .A(core__abc_21380_n6964), .B(core__abc_21380_n6969), .Y(core__abc_21380_n6970) );
  AND2X2 AND2X2_4032 ( .A(core__abc_21380_n6964), .B(core__abc_21380_n6972), .Y(core__abc_21380_n6973) );
  AND2X2 AND2X2_4033 ( .A(core__abc_21380_n6967), .B(core__abc_21380_n3693_1), .Y(core__abc_21380_n6974) );
  AND2X2 AND2X2_4034 ( .A(core__abc_21380_n6973), .B(core__abc_21380_n6976), .Y(core__abc_21380_n6977) );
  AND2X2 AND2X2_4035 ( .A(core__abc_21380_n5566), .B(core__abc_21380_n2303), .Y(core__abc_21380_n6978) );
  AND2X2 AND2X2_4036 ( .A(core__abc_21380_n5567), .B(core_v1_reg_56_), .Y(core__abc_21380_n6979) );
  AND2X2 AND2X2_4037 ( .A(core__abc_21380_n6981), .B(core__abc_21380_n3612), .Y(core__abc_21380_n6982) );
  AND2X2 AND2X2_4038 ( .A(core__abc_21380_n6980), .B(core__abc_21380_n3610), .Y(core__abc_21380_n6983) );
  AND2X2 AND2X2_4039 ( .A(core__abc_21380_n6986), .B(core__abc_21380_n6987), .Y(core__abc_21380_n6988) );
  AND2X2 AND2X2_404 ( .A(_abc_19068_n915_1_bF_buf2), .B(core_mi_63_), .Y(_abc_19068_n1613) );
  AND2X2 AND2X2_4040 ( .A(core__abc_21380_n6989), .B(core__abc_21380_n3545), .Y(core__abc_21380_n6990) );
  AND2X2 AND2X2_4041 ( .A(core__abc_21380_n5472), .B(core__abc_21380_n2265), .Y(core__abc_21380_n6991) );
  AND2X2 AND2X2_4042 ( .A(core__abc_21380_n5473), .B(core_v1_reg_54_), .Y(core__abc_21380_n6992) );
  AND2X2 AND2X2_4043 ( .A(core__abc_21380_n6993), .B(core__abc_21380_n3471), .Y(core__abc_21380_n6996) );
  AND2X2 AND2X2_4044 ( .A(core__abc_21380_n6997), .B(core__abc_21380_n6994), .Y(core__abc_21380_n6998) );
  AND2X2 AND2X2_4045 ( .A(core__abc_21380_n6999), .B(core__abc_21380_n7000), .Y(core__abc_21380_n7001) );
  AND2X2 AND2X2_4046 ( .A(core__abc_21380_n7002), .B(core__abc_21380_n3416), .Y(core__abc_21380_n7003) );
  AND2X2 AND2X2_4047 ( .A(core__abc_21380_n7005), .B(core__abc_21380_n7006), .Y(core__abc_21380_n7007) );
  AND2X2 AND2X2_4048 ( .A(core__abc_21380_n7008), .B(core__abc_21380_n3345), .Y(core__abc_21380_n7009) );
  AND2X2 AND2X2_4049 ( .A(core__abc_21380_n1270_1), .B(core_v1_reg_51_), .Y(core__abc_21380_n7010) );
  AND2X2 AND2X2_405 ( .A(_abc_19068_n923_bF_buf3), .B(_abc_19068_n1617), .Y(_auto_iopadmap_cc_313_execute_30317_31_) );
  AND2X2 AND2X2_4050 ( .A(core__abc_21380_n1262_1), .B(core__abc_21380_n2210), .Y(core__abc_21380_n7011) );
  AND2X2 AND2X2_4051 ( .A(core__abc_21380_n7012), .B(core__abc_21380_n1268_1), .Y(core__abc_21380_n7013) );
  AND2X2 AND2X2_4052 ( .A(core__abc_21380_n7007), .B(core__abc_21380_n3344), .Y(core__abc_21380_n7015) );
  AND2X2 AND2X2_4053 ( .A(core__abc_21380_n7014), .B(core__abc_21380_n7016), .Y(core__abc_21380_n7017) );
  AND2X2 AND2X2_4054 ( .A(core__abc_21380_n7017), .B(core__abc_21380_n7013), .Y(core__abc_21380_n7018) );
  AND2X2 AND2X2_4055 ( .A(core__abc_21380_n7001), .B(core__abc_21380_n3415), .Y(core__abc_21380_n7021) );
  AND2X2 AND2X2_4056 ( .A(core__abc_21380_n7020), .B(core__abc_21380_n7022), .Y(core__abc_21380_n7023) );
  AND2X2 AND2X2_4057 ( .A(core__abc_21380_n7019), .B(core__abc_21380_n7023), .Y(core__abc_21380_n7024) );
  AND2X2 AND2X2_4058 ( .A(core__abc_21380_n7025), .B(core__abc_21380_n6998), .Y(core__abc_21380_n7026) );
  AND2X2 AND2X2_4059 ( .A(core__abc_21380_n6988), .B(core__abc_21380_n3543), .Y(core__abc_21380_n7028) );
  AND2X2 AND2X2_406 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_96_), .Y(_abc_19068_n1619) );
  AND2X2 AND2X2_4060 ( .A(core__abc_21380_n7027), .B(core__abc_21380_n7030), .Y(core__abc_21380_n7031) );
  AND2X2 AND2X2_4061 ( .A(core__abc_21380_n7032), .B(core__abc_21380_n6985), .Y(core__abc_21380_n7033) );
  AND2X2 AND2X2_4062 ( .A(core__abc_21380_n7034), .B(core__abc_21380_n6977), .Y(core__abc_21380_n7035) );
  AND2X2 AND2X2_4063 ( .A(core__abc_21380_n6939), .B(core__abc_21380_n7037), .Y(core__abc_21380_n7038) );
  AND2X2 AND2X2_4064 ( .A(core__abc_21380_n6943), .B(core__abc_21380_n3820), .Y(core__abc_21380_n7039) );
  AND2X2 AND2X2_4065 ( .A(core__abc_21380_n7038), .B(core__abc_21380_n7041), .Y(core__abc_21380_n7042) );
  AND2X2 AND2X2_4066 ( .A(core__abc_21380_n6955), .B(core__abc_21380_n7042), .Y(core__abc_21380_n7043) );
  AND2X2 AND2X2_4067 ( .A(core__abc_21380_n7036), .B(core__abc_21380_n7043), .Y(core__abc_21380_n7044) );
  AND2X2 AND2X2_4068 ( .A(core__abc_21380_n7045), .B(core__abc_21380_n6918), .Y(core__abc_21380_n7046) );
  AND2X2 AND2X2_4069 ( .A(core__abc_21380_n7048), .B(core__abc_21380_n6852), .Y(core__abc_21380_n7049) );
  AND2X2 AND2X2_407 ( .A(_abc_19068_n1620_bF_buf10), .B(word3_reg_0_), .Y(_abc_19068_n1621) );
  AND2X2 AND2X2_4070 ( .A(core__abc_21380_n6848), .B(core__abc_21380_n4396), .Y(core__abc_21380_n7050) );
  AND2X2 AND2X2_4071 ( .A(core__abc_21380_n7049), .B(core__abc_21380_n7052), .Y(core__abc_21380_n7053) );
  AND2X2 AND2X2_4072 ( .A(core__abc_21380_n6839), .B(core__abc_21380_n7053), .Y(core__abc_21380_n7054) );
  AND2X2 AND2X2_4073 ( .A(core__abc_21380_n6823), .B(core__abc_21380_n7054), .Y(core__abc_21380_n7055) );
  AND2X2 AND2X2_4074 ( .A(core__abc_21380_n7047), .B(core__abc_21380_n7055), .Y(core__abc_21380_n7056) );
  AND2X2 AND2X2_4075 ( .A(core__abc_21380_n7057), .B(core__abc_21380_n6783), .Y(core__abc_21380_n7058) );
  AND2X2 AND2X2_4076 ( .A(core__abc_21380_n7062), .B(core__abc_21380_n7063), .Y(core__abc_21380_n7064) );
  AND2X2 AND2X2_4077 ( .A(core__abc_21380_n7065), .B(core__abc_21380_n5325), .Y(core__abc_21380_n7066) );
  AND2X2 AND2X2_4078 ( .A(core__abc_21380_n7064), .B(core__abc_21380_n5324), .Y(core__abc_21380_n7067) );
  AND2X2 AND2X2_4079 ( .A(core__abc_21380_n7060), .B(core__abc_21380_n7068), .Y(core__abc_21380_n7069) );
  AND2X2 AND2X2_408 ( .A(_abc_19068_n1622), .B(reset_n_bF_buf84), .Y(word3_reg_0__FF_INPUT) );
  AND2X2 AND2X2_4080 ( .A(core__abc_21380_n7059), .B(core__abc_21380_n7070), .Y(core__abc_21380_n7071) );
  AND2X2 AND2X2_4081 ( .A(core__abc_21380_n7073), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n7074) );
  AND2X2 AND2X2_4082 ( .A(core__abc_21380_n3315), .B(core__abc_21380_n3164), .Y(core__abc_21380_n7075) );
  AND2X2 AND2X2_4083 ( .A(core__abc_21380_n3313_bF_buf12), .B(core__abc_21380_n7077), .Y(core__abc_21380_n7078) );
  AND2X2 AND2X2_4084 ( .A(core__abc_21380_n7080), .B(core__abc_21380_n7081), .Y(core__abc_21380_n7082) );
  AND2X2 AND2X2_4085 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core__abc_21380_n7082), .Y(core__abc_21380_n7083) );
  AND2X2 AND2X2_4086 ( .A(core__abc_21380_n7088), .B(reset_n_bF_buf0), .Y(core__abc_21380_n7089) );
  AND2X2 AND2X2_4087 ( .A(core__abc_21380_n7086), .B(core__abc_21380_n7089), .Y(core_v2_reg_0__FF_INPUT) );
  AND2X2 AND2X2_4088 ( .A(core__abc_21380_n3340), .B(core__abc_21380_n1629), .Y(core__abc_21380_n7091) );
  AND2X2 AND2X2_4089 ( .A(core__abc_21380_n3359), .B(core_v1_reg_20_), .Y(core__abc_21380_n7092) );
  AND2X2 AND2X2_409 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_97_), .Y(_abc_19068_n1624) );
  AND2X2 AND2X2_4090 ( .A(core__abc_21380_n5384), .B(core__abc_21380_n7093), .Y(core__abc_21380_n7094) );
  AND2X2 AND2X2_4091 ( .A(core__abc_21380_n7095), .B(core__abc_21380_n5382), .Y(core__abc_21380_n7096) );
  AND2X2 AND2X2_4092 ( .A(core__abc_21380_n7099), .B(core__abc_21380_n7098), .Y(core__abc_21380_n7100) );
  AND2X2 AND2X2_4093 ( .A(core__abc_21380_n7100), .B(core__abc_21380_n7097), .Y(core__abc_21380_n7101) );
  AND2X2 AND2X2_4094 ( .A(core__abc_21380_n7105), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n7106) );
  AND2X2 AND2X2_4095 ( .A(core__abc_21380_n3313_bF_buf11), .B(core_key_1_), .Y(core__abc_21380_n7107) );
  AND2X2 AND2X2_4096 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core__abc_21380_n1283), .Y(core__abc_21380_n7108) );
  AND2X2 AND2X2_4097 ( .A(core__abc_21380_n7112), .B(reset_n_bF_buf84), .Y(core__abc_21380_n7113) );
  AND2X2 AND2X2_4098 ( .A(core__abc_21380_n7111), .B(core__abc_21380_n7113), .Y(core_v2_reg_1__FF_INPUT) );
  AND2X2 AND2X2_4099 ( .A(core__abc_21380_n7115), .B(core__abc_21380_n7070), .Y(core__abc_21380_n7116) );
  AND2X2 AND2X2_41 ( .A(_abc_19068_n915_1_bF_buf3), .B(core_mi_32_), .Y(_abc_19068_n934_1) );
  AND2X2 AND2X2_410 ( .A(_abc_19068_n1620_bF_buf9), .B(word3_reg_1_), .Y(_abc_19068_n1625) );
  AND2X2 AND2X2_4100 ( .A(core__abc_21380_n7059), .B(core__abc_21380_n7116), .Y(core__abc_21380_n7117) );
  AND2X2 AND2X2_4101 ( .A(core__abc_21380_n7115), .B(core__abc_21380_n7066), .Y(core__abc_21380_n7118) );
  AND2X2 AND2X2_4102 ( .A(core__abc_21380_n7122), .B(core__abc_21380_n7123), .Y(core__abc_21380_n7124) );
  AND2X2 AND2X2_4103 ( .A(core__abc_21380_n7125), .B(core__abc_21380_n5436), .Y(core__abc_21380_n7126) );
  AND2X2 AND2X2_4104 ( .A(core__abc_21380_n7124), .B(core__abc_21380_n5435), .Y(core__abc_21380_n7127) );
  AND2X2 AND2X2_4105 ( .A(core__abc_21380_n7121), .B(core__abc_21380_n7128), .Y(core__abc_21380_n7129) );
  AND2X2 AND2X2_4106 ( .A(core__abc_21380_n7120), .B(core__abc_21380_n7130), .Y(core__abc_21380_n7131) );
  AND2X2 AND2X2_4107 ( .A(core__abc_21380_n7133), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n7134) );
  AND2X2 AND2X2_4108 ( .A(core__abc_21380_n3313_bF_buf10), .B(core_key_2_), .Y(core__abc_21380_n7135) );
  AND2X2 AND2X2_4109 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core__abc_21380_n1306), .Y(core__abc_21380_n7136) );
  AND2X2 AND2X2_411 ( .A(_abc_19068_n1626), .B(reset_n_bF_buf83), .Y(word3_reg_1__FF_INPUT) );
  AND2X2 AND2X2_4110 ( .A(core__abc_21380_n7140), .B(reset_n_bF_buf83), .Y(core__abc_21380_n7141) );
  AND2X2 AND2X2_4111 ( .A(core__abc_21380_n7139), .B(core__abc_21380_n7141), .Y(core_v2_reg_2__FF_INPUT) );
  AND2X2 AND2X2_4112 ( .A(core__abc_21380_n3463), .B(core__abc_21380_n1665), .Y(core__abc_21380_n7145) );
  AND2X2 AND2X2_4113 ( .A(core__abc_21380_n3477), .B(core_v1_reg_22_), .Y(core__abc_21380_n7146) );
  AND2X2 AND2X2_4114 ( .A(core__abc_21380_n7148), .B(core__abc_21380_n5479), .Y(core__abc_21380_n7149) );
  AND2X2 AND2X2_4115 ( .A(core__abc_21380_n7147), .B(core__abc_21380_n5480), .Y(core__abc_21380_n7151) );
  AND2X2 AND2X2_4116 ( .A(core__abc_21380_n7150), .B(core__abc_21380_n7152), .Y(core__abc_21380_n7153) );
  AND2X2 AND2X2_4117 ( .A(core__abc_21380_n7144), .B(core__abc_21380_n7154), .Y(core__abc_21380_n7155) );
  AND2X2 AND2X2_4118 ( .A(core__abc_21380_n7143), .B(core__abc_21380_n7153), .Y(core__abc_21380_n7156) );
  AND2X2 AND2X2_4119 ( .A(core__abc_21380_n7158), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n7159) );
  AND2X2 AND2X2_412 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_98_), .Y(_abc_19068_n1628) );
  AND2X2 AND2X2_4120 ( .A(core__abc_21380_n3313_bF_buf9), .B(core_key_3_), .Y(core__abc_21380_n7160) );
  AND2X2 AND2X2_4121 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core__abc_21380_n1324), .Y(core__abc_21380_n7161) );
  AND2X2 AND2X2_4122 ( .A(core__abc_21380_n7165), .B(reset_n_bF_buf82), .Y(core__abc_21380_n7166) );
  AND2X2 AND2X2_4123 ( .A(core__abc_21380_n7164), .B(core__abc_21380_n7166), .Y(core_v2_reg_3__FF_INPUT) );
  AND2X2 AND2X2_4124 ( .A(core__abc_21380_n7152), .B(core__abc_21380_n7126), .Y(core__abc_21380_n7168) );
  AND2X2 AND2X2_4125 ( .A(core__abc_21380_n7153), .B(core__abc_21380_n7130), .Y(core__abc_21380_n7170) );
  AND2X2 AND2X2_4126 ( .A(core__abc_21380_n7170), .B(core__abc_21380_n7119), .Y(core__abc_21380_n7171) );
  AND2X2 AND2X2_4127 ( .A(core__abc_21380_n7170), .B(core__abc_21380_n7116), .Y(core__abc_21380_n7173) );
  AND2X2 AND2X2_4128 ( .A(core__abc_21380_n7059), .B(core__abc_21380_n7173), .Y(core__abc_21380_n7174) );
  AND2X2 AND2X2_4129 ( .A(core__abc_21380_n7176), .B(core__abc_21380_n7177), .Y(core__abc_21380_n7178) );
  AND2X2 AND2X2_413 ( .A(_abc_19068_n1620_bF_buf8), .B(word3_reg_2_), .Y(_abc_19068_n1629) );
  AND2X2 AND2X2_4130 ( .A(core__abc_21380_n7179), .B(core__abc_21380_n5531), .Y(core__abc_21380_n7180) );
  AND2X2 AND2X2_4131 ( .A(core__abc_21380_n7178), .B(core__abc_21380_n5530), .Y(core__abc_21380_n7181) );
  AND2X2 AND2X2_4132 ( .A(core__abc_21380_n7175), .B(core__abc_21380_n7183), .Y(core__abc_21380_n7184) );
  AND2X2 AND2X2_4133 ( .A(core__abc_21380_n7185), .B(core__abc_21380_n7186), .Y(core__abc_21380_n7187) );
  AND2X2 AND2X2_4134 ( .A(core__abc_21380_n7187), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n7188) );
  AND2X2 AND2X2_4135 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_4_), .Y(core__abc_21380_n7189) );
  AND2X2 AND2X2_4136 ( .A(core__abc_21380_n7190), .B(core__abc_21380_n7191), .Y(core__abc_21380_n7192) );
  AND2X2 AND2X2_4137 ( .A(core__abc_21380_n3163_1_bF_buf1), .B(core__abc_21380_n7192), .Y(core__abc_21380_n7193) );
  AND2X2 AND2X2_4138 ( .A(core__abc_21380_n7197), .B(reset_n_bF_buf81), .Y(core__abc_21380_n7198) );
  AND2X2 AND2X2_4139 ( .A(core__abc_21380_n7196), .B(core__abc_21380_n7198), .Y(core_v2_reg_4__FF_INPUT) );
  AND2X2 AND2X2_414 ( .A(_abc_19068_n1630), .B(reset_n_bF_buf82), .Y(word3_reg_2__FF_INPUT) );
  AND2X2 AND2X2_4140 ( .A(core__abc_21380_n7185), .B(core__abc_21380_n7200), .Y(core__abc_21380_n7201) );
  AND2X2 AND2X2_4141 ( .A(core__abc_21380_n3603), .B(core__abc_21380_n1703), .Y(core__abc_21380_n7204) );
  AND2X2 AND2X2_4142 ( .A(core__abc_21380_n3604_1), .B(core_v1_reg_24_), .Y(core__abc_21380_n7205) );
  AND2X2 AND2X2_4143 ( .A(core__abc_21380_n7207), .B(core__abc_21380_n7203), .Y(core__abc_21380_n7208) );
  AND2X2 AND2X2_4144 ( .A(core__abc_21380_n7206), .B(core__abc_21380_n5572), .Y(core__abc_21380_n7210) );
  AND2X2 AND2X2_4145 ( .A(core__abc_21380_n7209), .B(core__abc_21380_n7211), .Y(core__abc_21380_n7212) );
  AND2X2 AND2X2_4146 ( .A(core__abc_21380_n7202), .B(core__abc_21380_n7213), .Y(core__abc_21380_n7214) );
  AND2X2 AND2X2_4147 ( .A(core__abc_21380_n7201), .B(core__abc_21380_n7212), .Y(core__abc_21380_n7215) );
  AND2X2 AND2X2_4148 ( .A(core__abc_21380_n7216), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n7217) );
  AND2X2 AND2X2_4149 ( .A(core__abc_21380_n3313_bF_buf7), .B(core__abc_21380_n7218), .Y(core__abc_21380_n7219) );
  AND2X2 AND2X2_415 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_99_), .Y(_abc_19068_n1632) );
  AND2X2 AND2X2_4150 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core__abc_21380_n1361), .Y(core__abc_21380_n7220) );
  AND2X2 AND2X2_4151 ( .A(core__abc_21380_n7224), .B(reset_n_bF_buf80), .Y(core__abc_21380_n7225) );
  AND2X2 AND2X2_4152 ( .A(core__abc_21380_n7223), .B(core__abc_21380_n7225), .Y(core_v2_reg_5__FF_INPUT) );
  AND2X2 AND2X2_4153 ( .A(core__abc_21380_n7228), .B(core__abc_21380_n7229), .Y(core__abc_21380_n7230) );
  AND2X2 AND2X2_4154 ( .A(core__abc_21380_n7231), .B(core__abc_21380_n5624), .Y(core__abc_21380_n7232) );
  AND2X2 AND2X2_4155 ( .A(core__abc_21380_n7230), .B(core__abc_21380_n5623), .Y(core__abc_21380_n7233) );
  AND2X2 AND2X2_4156 ( .A(core__abc_21380_n7209), .B(core__abc_21380_n7200), .Y(core__abc_21380_n7235) );
  AND2X2 AND2X2_4157 ( .A(core__abc_21380_n7185), .B(core__abc_21380_n7235), .Y(core__abc_21380_n7236) );
  AND2X2 AND2X2_4158 ( .A(core__abc_21380_n7237), .B(core__abc_21380_n7234), .Y(core__abc_21380_n7238) );
  AND2X2 AND2X2_4159 ( .A(core__abc_21380_n7242), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n7243) );
  AND2X2 AND2X2_416 ( .A(_abc_19068_n1620_bF_buf7), .B(word3_reg_3_), .Y(_abc_19068_n1633) );
  AND2X2 AND2X2_4160 ( .A(core__abc_21380_n3313_bF_buf6), .B(core__abc_21380_n7244), .Y(core__abc_21380_n7245) );
  AND2X2 AND2X2_4161 ( .A(core__abc_21380_n3163_1_bF_buf6), .B(core__abc_21380_n1381), .Y(core__abc_21380_n7246) );
  AND2X2 AND2X2_4162 ( .A(core__abc_21380_n7250), .B(reset_n_bF_buf79), .Y(core__abc_21380_n7251) );
  AND2X2 AND2X2_4163 ( .A(core__abc_21380_n7249), .B(core__abc_21380_n7251), .Y(core_v2_reg_6__FF_INPUT) );
  AND2X2 AND2X2_4164 ( .A(core__abc_21380_n7239), .B(core__abc_21380_n7253), .Y(core__abc_21380_n7254) );
  AND2X2 AND2X2_4165 ( .A(core__abc_21380_n3746), .B(core__abc_21380_n7256), .Y(core__abc_21380_n7257) );
  AND2X2 AND2X2_4166 ( .A(core__abc_21380_n3760), .B(core_v1_reg_26_), .Y(core__abc_21380_n7258) );
  AND2X2 AND2X2_4167 ( .A(core__abc_21380_n7255), .B(core__abc_21380_n7260), .Y(core__abc_21380_n7261) );
  AND2X2 AND2X2_4168 ( .A(core__abc_21380_n5668), .B(core__abc_21380_n7259), .Y(core__abc_21380_n7262) );
  AND2X2 AND2X2_4169 ( .A(core__abc_21380_n7254), .B(core__abc_21380_n7263), .Y(core__abc_21380_n7264) );
  AND2X2 AND2X2_417 ( .A(_abc_19068_n1634), .B(reset_n_bF_buf81), .Y(word3_reg_3__FF_INPUT) );
  AND2X2 AND2X2_4170 ( .A(core__abc_21380_n7265), .B(core__abc_21380_n7266), .Y(core__abc_21380_n7267) );
  AND2X2 AND2X2_4171 ( .A(core__abc_21380_n7267), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n7268) );
  AND2X2 AND2X2_4172 ( .A(core__abc_21380_n3313_bF_buf5), .B(core_key_7_), .Y(core__abc_21380_n7269) );
  AND2X2 AND2X2_4173 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core__abc_21380_n1400), .Y(core__abc_21380_n7270) );
  AND2X2 AND2X2_4174 ( .A(core__abc_21380_n7274), .B(reset_n_bF_buf78), .Y(core__abc_21380_n7275) );
  AND2X2 AND2X2_4175 ( .A(core__abc_21380_n7273), .B(core__abc_21380_n7275), .Y(core_v2_reg_7__FF_INPUT) );
  AND2X2 AND2X2_4176 ( .A(core__abc_21380_n7212), .B(core__abc_21380_n7183), .Y(core__abc_21380_n7277) );
  AND2X2 AND2X2_4177 ( .A(core__abc_21380_n7279), .B(core__abc_21380_n7277), .Y(core__abc_21380_n7280) );
  AND2X2 AND2X2_4178 ( .A(core__abc_21380_n7280), .B(core__abc_21380_n7173), .Y(core__abc_21380_n7281) );
  AND2X2 AND2X2_4179 ( .A(core__abc_21380_n7059), .B(core__abc_21380_n7281), .Y(core__abc_21380_n7282) );
  AND2X2 AND2X2_418 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_100_), .Y(_abc_19068_n1636) );
  AND2X2 AND2X2_4180 ( .A(core__abc_21380_n7280), .B(core__abc_21380_n7172), .Y(core__abc_21380_n7283) );
  AND2X2 AND2X2_4181 ( .A(core__abc_21380_n7287), .B(core__abc_21380_n7232), .Y(core__abc_21380_n7288) );
  AND2X2 AND2X2_4182 ( .A(core__abc_21380_n7286), .B(core__abc_21380_n7290), .Y(core__abc_21380_n7291) );
  AND2X2 AND2X2_4183 ( .A(core__abc_21380_n7284), .B(core__abc_21380_n7291), .Y(core__abc_21380_n7292) );
  AND2X2 AND2X2_4184 ( .A(core__abc_21380_n7295), .B(core__abc_21380_n7296), .Y(core__abc_21380_n7297) );
  AND2X2 AND2X2_4185 ( .A(core__abc_21380_n7298), .B(core__abc_21380_n5722), .Y(core__abc_21380_n7299) );
  AND2X2 AND2X2_4186 ( .A(core__abc_21380_n7297), .B(core__abc_21380_n5721), .Y(core__abc_21380_n7300) );
  AND2X2 AND2X2_4187 ( .A(core__abc_21380_n7294), .B(core__abc_21380_n7302), .Y(core__abc_21380_n7303) );
  AND2X2 AND2X2_4188 ( .A(core__abc_21380_n7304), .B(core__abc_21380_n7301), .Y(core__abc_21380_n7305) );
  AND2X2 AND2X2_4189 ( .A(core__abc_21380_n7307), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n7308) );
  AND2X2 AND2X2_419 ( .A(_abc_19068_n1620_bF_buf6), .B(word3_reg_4_), .Y(_abc_19068_n1637) );
  AND2X2 AND2X2_4190 ( .A(core__abc_21380_n3313_bF_buf4), .B(core_key_8_), .Y(core__abc_21380_n7309) );
  AND2X2 AND2X2_4191 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core_v2_reg_8_), .Y(core__abc_21380_n7310) );
  AND2X2 AND2X2_4192 ( .A(core__abc_21380_n7314), .B(reset_n_bF_buf77), .Y(core__abc_21380_n7315) );
  AND2X2 AND2X2_4193 ( .A(core__abc_21380_n7313), .B(core__abc_21380_n7315), .Y(core_v2_reg_8__FF_INPUT) );
  AND2X2 AND2X2_4194 ( .A(core__abc_21380_n7318), .B(core__abc_21380_n7317), .Y(core__abc_21380_n7319) );
  AND2X2 AND2X2_4195 ( .A(core__abc_21380_n3890), .B(core__abc_21380_n1778), .Y(core__abc_21380_n7320) );
  AND2X2 AND2X2_4196 ( .A(core__abc_21380_n7321), .B(core__abc_21380_n7322), .Y(core__abc_21380_n7323) );
  AND2X2 AND2X2_4197 ( .A(core__abc_21380_n7323), .B(core__abc_21380_n5768), .Y(core__abc_21380_n7324) );
  AND2X2 AND2X2_4198 ( .A(core__abc_21380_n7326), .B(core__abc_21380_n5766), .Y(core__abc_21380_n7327) );
  AND2X2 AND2X2_4199 ( .A(core__abc_21380_n7328), .B(core__abc_21380_n7325), .Y(core__abc_21380_n7329) );
  AND2X2 AND2X2_42 ( .A(_abc_19068_n897_1_bF_buf3), .B(word0_reg_0_), .Y(_abc_19068_n935) );
  AND2X2 AND2X2_420 ( .A(_abc_19068_n1638), .B(reset_n_bF_buf80), .Y(word3_reg_4__FF_INPUT) );
  AND2X2 AND2X2_4200 ( .A(core__abc_21380_n7319), .B(core__abc_21380_n7330), .Y(core__abc_21380_n7331) );
  AND2X2 AND2X2_4201 ( .A(core__abc_21380_n7332), .B(core__abc_21380_n7333), .Y(core__abc_21380_n7334) );
  AND2X2 AND2X2_4202 ( .A(core__abc_21380_n7334), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n7335) );
  AND2X2 AND2X2_4203 ( .A(core__abc_21380_n3313_bF_buf3), .B(core__abc_21380_n7336), .Y(core__abc_21380_n7337) );
  AND2X2 AND2X2_4204 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core_v2_reg_9_), .Y(core__abc_21380_n7338) );
  AND2X2 AND2X2_4205 ( .A(core__abc_21380_n7342), .B(reset_n_bF_buf76), .Y(core__abc_21380_n7343) );
  AND2X2 AND2X2_4206 ( .A(core__abc_21380_n7341), .B(core__abc_21380_n7343), .Y(core_v2_reg_9__FF_INPUT) );
  AND2X2 AND2X2_4207 ( .A(core__abc_21380_n7345), .B(core__abc_21380_n7325), .Y(core__abc_21380_n7346) );
  AND2X2 AND2X2_4208 ( .A(core__abc_21380_n7329), .B(core__abc_21380_n7302), .Y(core__abc_21380_n7348) );
  AND2X2 AND2X2_4209 ( .A(core__abc_21380_n7294), .B(core__abc_21380_n7348), .Y(core__abc_21380_n7349) );
  AND2X2 AND2X2_421 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_101_), .Y(_abc_19068_n1640) );
  AND2X2 AND2X2_4210 ( .A(core__abc_21380_n7352), .B(core__abc_21380_n7353), .Y(core__abc_21380_n7354) );
  AND2X2 AND2X2_4211 ( .A(core__abc_21380_n7355), .B(core__abc_21380_n5807), .Y(core__abc_21380_n7356) );
  AND2X2 AND2X2_4212 ( .A(core__abc_21380_n7354), .B(core__abc_21380_n5809), .Y(core__abc_21380_n7357) );
  AND2X2 AND2X2_4213 ( .A(core__abc_21380_n7351), .B(core__abc_21380_n7358), .Y(core__abc_21380_n7359) );
  AND2X2 AND2X2_4214 ( .A(core__abc_21380_n7350), .B(core__abc_21380_n7360), .Y(core__abc_21380_n7361) );
  AND2X2 AND2X2_4215 ( .A(core__abc_21380_n7363), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n7364) );
  AND2X2 AND2X2_4216 ( .A(core__abc_21380_n3313_bF_buf2), .B(core_key_10_), .Y(core__abc_21380_n7365) );
  AND2X2 AND2X2_4217 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core_v2_reg_10_), .Y(core__abc_21380_n7366) );
  AND2X2 AND2X2_4218 ( .A(core__abc_21380_n7370), .B(reset_n_bF_buf75), .Y(core__abc_21380_n7371) );
  AND2X2 AND2X2_4219 ( .A(core__abc_21380_n7369), .B(core__abc_21380_n7371), .Y(core_v2_reg_10__FF_INPUT) );
  AND2X2 AND2X2_422 ( .A(_abc_19068_n1620_bF_buf5), .B(word3_reg_5_), .Y(_abc_19068_n1641) );
  AND2X2 AND2X2_4220 ( .A(core__abc_21380_n4011), .B(core_v1_reg_30_), .Y(core__abc_21380_n7375) );
  AND2X2 AND2X2_4221 ( .A(core__abc_21380_n4072_1), .B(core__abc_21380_n1816_1), .Y(core__abc_21380_n7376) );
  AND2X2 AND2X2_4222 ( .A(core__abc_21380_n7377), .B(core__abc_21380_n3154), .Y(core__abc_21380_n7378) );
  AND2X2 AND2X2_4223 ( .A(core__abc_21380_n7379), .B(core__abc_21380_n3157), .Y(core__abc_21380_n7380) );
  AND2X2 AND2X2_4224 ( .A(core__abc_21380_n7374), .B(core__abc_21380_n7381), .Y(core__abc_21380_n7382) );
  AND2X2 AND2X2_4225 ( .A(core__abc_21380_n7373), .B(core__abc_21380_n7383), .Y(core__abc_21380_n7384) );
  AND2X2 AND2X2_4226 ( .A(core__abc_21380_n7386), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n7387) );
  AND2X2 AND2X2_4227 ( .A(core__abc_21380_n3313_bF_buf1), .B(core_key_11_), .Y(core__abc_21380_n7388) );
  AND2X2 AND2X2_4228 ( .A(core__abc_21380_n3163_1_bF_buf1), .B(core_v2_reg_11_), .Y(core__abc_21380_n7389) );
  AND2X2 AND2X2_4229 ( .A(core__abc_21380_n7393), .B(reset_n_bF_buf74), .Y(core__abc_21380_n7394) );
  AND2X2 AND2X2_423 ( .A(_abc_19068_n1642), .B(reset_n_bF_buf79), .Y(word3_reg_5__FF_INPUT) );
  AND2X2 AND2X2_4230 ( .A(core__abc_21380_n7392), .B(core__abc_21380_n7394), .Y(core_v2_reg_11__FF_INPUT) );
  AND2X2 AND2X2_4231 ( .A(core__abc_21380_n7383), .B(core__abc_21380_n7360), .Y(core__abc_21380_n7396) );
  AND2X2 AND2X2_4232 ( .A(core__abc_21380_n7396), .B(core__abc_21380_n7347), .Y(core__abc_21380_n7397) );
  AND2X2 AND2X2_4233 ( .A(core__abc_21380_n7383), .B(core__abc_21380_n7356), .Y(core__abc_21380_n7398) );
  AND2X2 AND2X2_4234 ( .A(core__abc_21380_n7396), .B(core__abc_21380_n7348), .Y(core__abc_21380_n7401) );
  AND2X2 AND2X2_4235 ( .A(core__abc_21380_n7294), .B(core__abc_21380_n7401), .Y(core__abc_21380_n7402) );
  AND2X2 AND2X2_4236 ( .A(core__abc_21380_n7405), .B(core__abc_21380_n7406), .Y(core__abc_21380_n7407) );
  AND2X2 AND2X2_4237 ( .A(core__abc_21380_n7408), .B(core__abc_21380_n3380), .Y(core__abc_21380_n7409) );
  AND2X2 AND2X2_4238 ( .A(core__abc_21380_n7407), .B(core__abc_21380_n3379), .Y(core__abc_21380_n7410) );
  AND2X2 AND2X2_4239 ( .A(core__abc_21380_n7404), .B(core__abc_21380_n7411), .Y(core__abc_21380_n7412) );
  AND2X2 AND2X2_424 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_102_), .Y(_abc_19068_n1644) );
  AND2X2 AND2X2_4240 ( .A(core__abc_21380_n7403), .B(core__abc_21380_n7413), .Y(core__abc_21380_n7414) );
  AND2X2 AND2X2_4241 ( .A(core__abc_21380_n7416), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n7417) );
  AND2X2 AND2X2_4242 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n7418), .Y(core__abc_21380_n7419) );
  AND2X2 AND2X2_4243 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core_v2_reg_12_), .Y(core__abc_21380_n7420) );
  AND2X2 AND2X2_4244 ( .A(core__abc_21380_n7424), .B(reset_n_bF_buf73), .Y(core__abc_21380_n7425) );
  AND2X2 AND2X2_4245 ( .A(core__abc_21380_n7423), .B(core__abc_21380_n7425), .Y(core_v2_reg_12__FF_INPUT) );
  AND2X2 AND2X2_4246 ( .A(core__abc_21380_n4174), .B(core__abc_21380_n1854), .Y(core__abc_21380_n7427) );
  AND2X2 AND2X2_4247 ( .A(core__abc_21380_n4160), .B(core_v1_reg_32_), .Y(core__abc_21380_n7428) );
  AND2X2 AND2X2_4248 ( .A(core__abc_21380_n7429), .B(core__abc_21380_n3434), .Y(core__abc_21380_n7431) );
  AND2X2 AND2X2_4249 ( .A(core__abc_21380_n7432), .B(core__abc_21380_n7430), .Y(core__abc_21380_n7433) );
  AND2X2 AND2X2_425 ( .A(_abc_19068_n1620_bF_buf4), .B(word3_reg_6_), .Y(_abc_19068_n1645) );
  AND2X2 AND2X2_4250 ( .A(core__abc_21380_n7436), .B(core__abc_21380_n7435), .Y(core__abc_21380_n7437) );
  AND2X2 AND2X2_4251 ( .A(core__abc_21380_n7437), .B(core__abc_21380_n7434), .Y(core__abc_21380_n7438) );
  AND2X2 AND2X2_4252 ( .A(core__abc_21380_n7442), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf2), .Y(core__abc_21380_n7443) );
  AND2X2 AND2X2_4253 ( .A(core__abc_21380_n3313_bF_buf12), .B(core__abc_21380_n7444), .Y(core__abc_21380_n7445) );
  AND2X2 AND2X2_4254 ( .A(core__abc_21380_n3163_1_bF_buf6), .B(core_v2_reg_13_), .Y(core__abc_21380_n7446) );
  AND2X2 AND2X2_4255 ( .A(core__abc_21380_n7450), .B(reset_n_bF_buf72), .Y(core__abc_21380_n7451) );
  AND2X2 AND2X2_4256 ( .A(core__abc_21380_n7449), .B(core__abc_21380_n7451), .Y(core_v2_reg_13__FF_INPUT) );
  AND2X2 AND2X2_4257 ( .A(core__abc_21380_n7433), .B(core__abc_21380_n7413), .Y(core__abc_21380_n7453) );
  AND2X2 AND2X2_4258 ( .A(core__abc_21380_n7403), .B(core__abc_21380_n7453), .Y(core__abc_21380_n7454) );
  AND2X2 AND2X2_4259 ( .A(core__abc_21380_n7432), .B(core__abc_21380_n7409), .Y(core__abc_21380_n7456) );
  AND2X2 AND2X2_426 ( .A(_abc_19068_n1646), .B(reset_n_bF_buf78), .Y(word3_reg_6__FF_INPUT) );
  AND2X2 AND2X2_4260 ( .A(core__abc_21380_n7460), .B(core__abc_21380_n7461), .Y(core__abc_21380_n7462) );
  AND2X2 AND2X2_4261 ( .A(core__abc_21380_n7463), .B(core__abc_21380_n3500), .Y(core__abc_21380_n7464) );
  AND2X2 AND2X2_4262 ( .A(core__abc_21380_n7462), .B(core__abc_21380_n3501_1), .Y(core__abc_21380_n7465) );
  AND2X2 AND2X2_4263 ( .A(core__abc_21380_n7459), .B(core__abc_21380_n7466), .Y(core__abc_21380_n7467) );
  AND2X2 AND2X2_4264 ( .A(core__abc_21380_n7458), .B(core__abc_21380_n7468), .Y(core__abc_21380_n7469) );
  AND2X2 AND2X2_4265 ( .A(core__abc_21380_n7471), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf2), .Y(core__abc_21380_n7472) );
  AND2X2 AND2X2_4266 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n7473), .Y(core__abc_21380_n7474) );
  AND2X2 AND2X2_4267 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core_v2_reg_14_), .Y(core__abc_21380_n7475) );
  AND2X2 AND2X2_4268 ( .A(core__abc_21380_n7479), .B(reset_n_bF_buf71), .Y(core__abc_21380_n7480) );
  AND2X2 AND2X2_4269 ( .A(core__abc_21380_n7478), .B(core__abc_21380_n7480), .Y(core_v2_reg_14__FF_INPUT) );
  AND2X2 AND2X2_427 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_103_), .Y(_abc_19068_n1648) );
  AND2X2 AND2X2_4270 ( .A(core__abc_21380_n4300), .B(core__abc_21380_n1890), .Y(core__abc_21380_n7484) );
  AND2X2 AND2X2_4271 ( .A(core__abc_21380_n4315), .B(core_v1_reg_34_), .Y(core__abc_21380_n7485) );
  AND2X2 AND2X2_4272 ( .A(core__abc_21380_n7487), .B(core__abc_21380_n3574), .Y(core__abc_21380_n7488) );
  AND2X2 AND2X2_4273 ( .A(core__abc_21380_n7486), .B(core__abc_21380_n3569_1), .Y(core__abc_21380_n7489) );
  AND2X2 AND2X2_4274 ( .A(core__abc_21380_n7483), .B(core__abc_21380_n7490), .Y(core__abc_21380_n7491) );
  AND2X2 AND2X2_4275 ( .A(core__abc_21380_n7482), .B(core__abc_21380_n7492), .Y(core__abc_21380_n7493) );
  AND2X2 AND2X2_4276 ( .A(core__abc_21380_n7495), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n7496) );
  AND2X2 AND2X2_4277 ( .A(core__abc_21380_n3313_bF_buf10), .B(core_key_15_), .Y(core__abc_21380_n7497) );
  AND2X2 AND2X2_4278 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core_v2_reg_15_), .Y(core__abc_21380_n7498) );
  AND2X2 AND2X2_4279 ( .A(core__abc_21380_n7502), .B(reset_n_bF_buf70), .Y(core__abc_21380_n7503) );
  AND2X2 AND2X2_428 ( .A(_abc_19068_n1620_bF_buf3), .B(word3_reg_7_), .Y(_abc_19068_n1649) );
  AND2X2 AND2X2_4280 ( .A(core__abc_21380_n7501), .B(core__abc_21380_n7503), .Y(core_v2_reg_15__FF_INPUT) );
  AND2X2 AND2X2_4281 ( .A(core__abc_21380_n7492), .B(core__abc_21380_n7468), .Y(core__abc_21380_n7505) );
  AND2X2 AND2X2_4282 ( .A(core__abc_21380_n7505), .B(core__abc_21380_n7453), .Y(core__abc_21380_n7506) );
  AND2X2 AND2X2_4283 ( .A(core__abc_21380_n7506), .B(core__abc_21380_n7400), .Y(core__abc_21380_n7507) );
  AND2X2 AND2X2_4284 ( .A(core__abc_21380_n7505), .B(core__abc_21380_n7457), .Y(core__abc_21380_n7508) );
  AND2X2 AND2X2_4285 ( .A(core__abc_21380_n7509), .B(core__abc_21380_n7465), .Y(core__abc_21380_n7510) );
  AND2X2 AND2X2_4286 ( .A(core__abc_21380_n7506), .B(core__abc_21380_n7401), .Y(core__abc_21380_n7514) );
  AND2X2 AND2X2_4287 ( .A(core__abc_21380_n7294), .B(core__abc_21380_n7514), .Y(core__abc_21380_n7515) );
  AND2X2 AND2X2_4288 ( .A(core__abc_21380_n7517), .B(core__abc_21380_n7518), .Y(core__abc_21380_n7519) );
  AND2X2 AND2X2_4289 ( .A(core__abc_21380_n3643), .B(core__abc_21380_n7519), .Y(core__abc_21380_n7520) );
  AND2X2 AND2X2_429 ( .A(_abc_19068_n1650), .B(reset_n_bF_buf77), .Y(word3_reg_7__FF_INPUT) );
  AND2X2 AND2X2_4290 ( .A(core__abc_21380_n3644), .B(core__abc_21380_n7521), .Y(core__abc_21380_n7522) );
  AND2X2 AND2X2_4291 ( .A(core__abc_21380_n7516), .B(core__abc_21380_n7524), .Y(core__abc_21380_n7525) );
  AND2X2 AND2X2_4292 ( .A(core__abc_21380_n7526), .B(core__abc_21380_n7528), .Y(core__abc_21380_n7529) );
  AND2X2 AND2X2_4293 ( .A(core__abc_21380_n7514), .B(core__abc_21380_n7281), .Y(core__abc_21380_n7530) );
  AND2X2 AND2X2_4294 ( .A(core__abc_21380_n7530), .B(core__abc_21380_n7059), .Y(core__abc_21380_n7531) );
  AND2X2 AND2X2_4295 ( .A(core__abc_21380_n7529), .B(core__abc_21380_n7532), .Y(core__abc_21380_n7533) );
  AND2X2 AND2X2_4296 ( .A(core__abc_21380_n7533), .B(core__abc_21380_n7523), .Y(core__abc_21380_n7534) );
  AND2X2 AND2X2_4297 ( .A(core__abc_21380_n7536), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n7537) );
  AND2X2 AND2X2_4298 ( .A(core__abc_21380_n3313_bF_buf9), .B(core__abc_21380_n7538), .Y(core__abc_21380_n7539) );
  AND2X2 AND2X2_4299 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core_v2_reg_16_), .Y(core__abc_21380_n7540) );
  AND2X2 AND2X2_43 ( .A(_abc_19068_n912_1), .B(_abc_19068_n901_1), .Y(_abc_19068_n939_1) );
  AND2X2 AND2X2_430 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_104_), .Y(_abc_19068_n1652) );
  AND2X2 AND2X2_4300 ( .A(core__abc_21380_n7544), .B(reset_n_bF_buf69), .Y(core__abc_21380_n7545) );
  AND2X2 AND2X2_4301 ( .A(core__abc_21380_n7543), .B(core__abc_21380_n7545), .Y(core_v2_reg_16__FF_INPUT) );
  AND2X2 AND2X2_4302 ( .A(core__abc_21380_n7548), .B(core__abc_21380_n7547), .Y(core__abc_21380_n7549) );
  AND2X2 AND2X2_4303 ( .A(core__abc_21380_n4474_1), .B(core__abc_21380_n1929), .Y(core__abc_21380_n7551) );
  AND2X2 AND2X2_4304 ( .A(core__abc_21380_n4461), .B(core_v1_reg_36_), .Y(core__abc_21380_n7552) );
  AND2X2 AND2X2_4305 ( .A(core__abc_21380_n3717), .B(core__abc_21380_n7554), .Y(core__abc_21380_n7555) );
  AND2X2 AND2X2_4306 ( .A(core__abc_21380_n3715), .B(core__abc_21380_n7553), .Y(core__abc_21380_n7557) );
  AND2X2 AND2X2_4307 ( .A(core__abc_21380_n7556), .B(core__abc_21380_n7558), .Y(core__abc_21380_n7559) );
  AND2X2 AND2X2_4308 ( .A(core__abc_21380_n7560), .B(core__abc_21380_n7562), .Y(core__abc_21380_n7563) );
  AND2X2 AND2X2_4309 ( .A(core__abc_21380_n7563), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n7564) );
  AND2X2 AND2X2_431 ( .A(_abc_19068_n1620_bF_buf2), .B(word3_reg_8_), .Y(_abc_19068_n1653) );
  AND2X2 AND2X2_4310 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_17_), .Y(core__abc_21380_n7565) );
  AND2X2 AND2X2_4311 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core_v2_reg_17_), .Y(core__abc_21380_n7566) );
  AND2X2 AND2X2_4312 ( .A(core__abc_21380_n7570), .B(reset_n_bF_buf68), .Y(core__abc_21380_n7571) );
  AND2X2 AND2X2_4313 ( .A(core__abc_21380_n7569), .B(core__abc_21380_n7571), .Y(core_v2_reg_17__FF_INPUT) );
  AND2X2 AND2X2_4314 ( .A(core__abc_21380_n7573), .B(core__abc_21380_n7558), .Y(core__abc_21380_n7574) );
  AND2X2 AND2X2_4315 ( .A(core__abc_21380_n7559), .B(core__abc_21380_n7524), .Y(core__abc_21380_n7575) );
  AND2X2 AND2X2_4316 ( .A(core__abc_21380_n7516), .B(core__abc_21380_n7575), .Y(core__abc_21380_n7576) );
  AND2X2 AND2X2_4317 ( .A(core__abc_21380_n7579), .B(core__abc_21380_n7580), .Y(core__abc_21380_n7581) );
  AND2X2 AND2X2_4318 ( .A(core__abc_21380_n3777), .B(core__abc_21380_n7581), .Y(core__abc_21380_n7582) );
  AND2X2 AND2X2_4319 ( .A(core__abc_21380_n3775), .B(core__abc_21380_n7583), .Y(core__abc_21380_n7584) );
  AND2X2 AND2X2_432 ( .A(_abc_19068_n1654), .B(reset_n_bF_buf76), .Y(word3_reg_8__FF_INPUT) );
  AND2X2 AND2X2_4320 ( .A(core__abc_21380_n7578), .B(core__abc_21380_n7585), .Y(core__abc_21380_n7586) );
  AND2X2 AND2X2_4321 ( .A(core__abc_21380_n7577), .B(core__abc_21380_n7587), .Y(core__abc_21380_n7588) );
  AND2X2 AND2X2_4322 ( .A(core__abc_21380_n7590), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n7591) );
  AND2X2 AND2X2_4323 ( .A(core__abc_21380_n3313_bF_buf7), .B(core__abc_21380_n7592), .Y(core__abc_21380_n7593) );
  AND2X2 AND2X2_4324 ( .A(core__abc_21380_n3163_1_bF_buf1), .B(core_v2_reg_18_), .Y(core__abc_21380_n7594) );
  AND2X2 AND2X2_4325 ( .A(core__abc_21380_n7598), .B(reset_n_bF_buf67), .Y(core__abc_21380_n7599) );
  AND2X2 AND2X2_4326 ( .A(core__abc_21380_n7597), .B(core__abc_21380_n7599), .Y(core_v2_reg_18__FF_INPUT) );
  AND2X2 AND2X2_4327 ( .A(core__abc_21380_n4606), .B(core__abc_21380_n1966), .Y(core__abc_21380_n7602) );
  AND2X2 AND2X2_4328 ( .A(core__abc_21380_n4594), .B(core_v1_reg_38_), .Y(core__abc_21380_n7603) );
  AND2X2 AND2X2_4329 ( .A(core__abc_21380_n3855), .B(core__abc_21380_n7605), .Y(core__abc_21380_n7606) );
  AND2X2 AND2X2_433 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_105_), .Y(_abc_19068_n1656) );
  AND2X2 AND2X2_4330 ( .A(core__abc_21380_n7607), .B(core__abc_21380_n7608), .Y(core__abc_21380_n7609) );
  AND2X2 AND2X2_4331 ( .A(core__abc_21380_n7613), .B(core__abc_21380_n7610), .Y(core__abc_21380_n7614) );
  AND2X2 AND2X2_4332 ( .A(core__abc_21380_n7614), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n7615) );
  AND2X2 AND2X2_4333 ( .A(core__abc_21380_n3313_bF_buf6), .B(core_key_19_), .Y(core__abc_21380_n7616) );
  AND2X2 AND2X2_4334 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core_v2_reg_19_), .Y(core__abc_21380_n7617) );
  AND2X2 AND2X2_4335 ( .A(core__abc_21380_n7621), .B(reset_n_bF_buf66), .Y(core__abc_21380_n7622) );
  AND2X2 AND2X2_4336 ( .A(core__abc_21380_n7620), .B(core__abc_21380_n7622), .Y(core_v2_reg_19__FF_INPUT) );
  AND2X2 AND2X2_4337 ( .A(core__abc_21380_n7609), .B(core__abc_21380_n7587), .Y(core__abc_21380_n7624) );
  AND2X2 AND2X2_4338 ( .A(core__abc_21380_n7624), .B(core__abc_21380_n7574), .Y(core__abc_21380_n7625) );
  AND2X2 AND2X2_4339 ( .A(core__abc_21380_n7626), .B(core__abc_21380_n7608), .Y(core__abc_21380_n7627) );
  AND2X2 AND2X2_434 ( .A(_abc_19068_n1620_bF_buf1), .B(word3_reg_9_), .Y(_abc_19068_n1657) );
  AND2X2 AND2X2_4340 ( .A(core__abc_21380_n7624), .B(core__abc_21380_n7575), .Y(core__abc_21380_n7630) );
  AND2X2 AND2X2_4341 ( .A(core__abc_21380_n7632), .B(core__abc_21380_n7629), .Y(core__abc_21380_n7633) );
  AND2X2 AND2X2_4342 ( .A(core__abc_21380_n7634), .B(core__abc_21380_n7635), .Y(core__abc_21380_n7636) );
  AND2X2 AND2X2_4343 ( .A(core__abc_21380_n3924), .B(core__abc_21380_n7637), .Y(core__abc_21380_n7638) );
  AND2X2 AND2X2_4344 ( .A(core__abc_21380_n3923), .B(core__abc_21380_n7636), .Y(core__abc_21380_n7639) );
  AND2X2 AND2X2_4345 ( .A(core__abc_21380_n7633), .B(core__abc_21380_n7640), .Y(core__abc_21380_n7641) );
  AND2X2 AND2X2_4346 ( .A(core__abc_21380_n7645), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n7646) );
  AND2X2 AND2X2_4347 ( .A(core__abc_21380_n3313_bF_buf5), .B(core_key_20_), .Y(core__abc_21380_n7647) );
  AND2X2 AND2X2_4348 ( .A(core__abc_21380_n3163_1_bF_buf6), .B(core_v2_reg_20_), .Y(core__abc_21380_n7648) );
  AND2X2 AND2X2_4349 ( .A(core__abc_21380_n7652), .B(reset_n_bF_buf65), .Y(core__abc_21380_n7653) );
  AND2X2 AND2X2_435 ( .A(_abc_19068_n1658), .B(reset_n_bF_buf75), .Y(word3_reg_9__FF_INPUT) );
  AND2X2 AND2X2_4350 ( .A(core__abc_21380_n7651), .B(core__abc_21380_n7653), .Y(core_v2_reg_20__FF_INPUT) );
  AND2X2 AND2X2_4351 ( .A(core__abc_21380_n4710), .B(core__abc_21380_n2005), .Y(core__abc_21380_n7655) );
  AND2X2 AND2X2_4352 ( .A(core__abc_21380_n4711), .B(core_v1_reg_40_), .Y(core__abc_21380_n7656) );
  AND2X2 AND2X2_4353 ( .A(core__abc_21380_n3985), .B(core__abc_21380_n7658), .Y(core__abc_21380_n7659) );
  AND2X2 AND2X2_4354 ( .A(core__abc_21380_n3983), .B(core__abc_21380_n7657), .Y(core__abc_21380_n7660) );
  AND2X2 AND2X2_4355 ( .A(core__abc_21380_n7642), .B(core__abc_21380_n7662), .Y(core__abc_21380_n7663) );
  AND2X2 AND2X2_4356 ( .A(core__abc_21380_n7663), .B(core__abc_21380_n7661), .Y(core__abc_21380_n7664) );
  AND2X2 AND2X2_4357 ( .A(core__abc_21380_n7665), .B(core__abc_21380_n7666), .Y(core__abc_21380_n7667) );
  AND2X2 AND2X2_4358 ( .A(core__abc_21380_n7667), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n7668) );
  AND2X2 AND2X2_4359 ( .A(core__abc_21380_n3313_bF_buf4), .B(core__abc_21380_n7669), .Y(core__abc_21380_n7670) );
  AND2X2 AND2X2_436 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_106_), .Y(_abc_19068_n1660) );
  AND2X2 AND2X2_4360 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core_v2_reg_21_), .Y(core__abc_21380_n7671) );
  AND2X2 AND2X2_4361 ( .A(core__abc_21380_n7675), .B(reset_n_bF_buf64), .Y(core__abc_21380_n7676) );
  AND2X2 AND2X2_4362 ( .A(core__abc_21380_n7674), .B(core__abc_21380_n7676), .Y(core_v2_reg_21__FF_INPUT) );
  AND2X2 AND2X2_4363 ( .A(core__abc_21380_n7643), .B(core__abc_21380_n7678), .Y(core__abc_21380_n7679) );
  AND2X2 AND2X2_4364 ( .A(core__abc_21380_n7678), .B(core__abc_21380_n7638), .Y(core__abc_21380_n7680) );
  AND2X2 AND2X2_4365 ( .A(core__abc_21380_n7684), .B(core__abc_21380_n7685), .Y(core__abc_21380_n7686) );
  AND2X2 AND2X2_4366 ( .A(core__abc_21380_n4042), .B(core__abc_21380_n7687), .Y(core__abc_21380_n7688) );
  AND2X2 AND2X2_4367 ( .A(core__abc_21380_n4041), .B(core__abc_21380_n7686), .Y(core__abc_21380_n7689) );
  AND2X2 AND2X2_4368 ( .A(core__abc_21380_n7683), .B(core__abc_21380_n7690), .Y(core__abc_21380_n7691) );
  AND2X2 AND2X2_4369 ( .A(core__abc_21380_n7682), .B(core__abc_21380_n7692), .Y(core__abc_21380_n7693) );
  AND2X2 AND2X2_437 ( .A(_abc_19068_n1620_bF_buf0), .B(word3_reg_10_), .Y(_abc_19068_n1661) );
  AND2X2 AND2X2_4370 ( .A(core__abc_21380_n7695), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n7696) );
  AND2X2 AND2X2_4371 ( .A(core__abc_21380_n3313_bF_buf3), .B(core__abc_21380_n7697), .Y(core__abc_21380_n7698) );
  AND2X2 AND2X2_4372 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core_v2_reg_22_), .Y(core__abc_21380_n7699) );
  AND2X2 AND2X2_4373 ( .A(core__abc_21380_n7703), .B(reset_n_bF_buf63), .Y(core__abc_21380_n7704) );
  AND2X2 AND2X2_4374 ( .A(core__abc_21380_n7702), .B(core__abc_21380_n7704), .Y(core_v2_reg_22__FF_INPUT) );
  AND2X2 AND2X2_4375 ( .A(core__abc_21380_n4809), .B(core__abc_21380_n2040), .Y(core__abc_21380_n7707) );
  AND2X2 AND2X2_4376 ( .A(core__abc_21380_n4822), .B(core_v1_reg_42_), .Y(core__abc_21380_n7708) );
  AND2X2 AND2X2_4377 ( .A(core__abc_21380_n4130), .B(core__abc_21380_n7710), .Y(core__abc_21380_n7711) );
  AND2X2 AND2X2_4378 ( .A(core__abc_21380_n4125), .B(core__abc_21380_n7709), .Y(core__abc_21380_n7713) );
  AND2X2 AND2X2_4379 ( .A(core__abc_21380_n7714), .B(core__abc_21380_n7712), .Y(core__abc_21380_n7715) );
  AND2X2 AND2X2_438 ( .A(_abc_19068_n1662), .B(reset_n_bF_buf74), .Y(word3_reg_10__FF_INPUT) );
  AND2X2 AND2X2_4380 ( .A(core__abc_21380_n7719), .B(core__abc_21380_n7717), .Y(core__abc_21380_n7720) );
  AND2X2 AND2X2_4381 ( .A(core__abc_21380_n7721), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n7722) );
  AND2X2 AND2X2_4382 ( .A(core__abc_21380_n3313_bF_buf2), .B(core_key_23_), .Y(core__abc_21380_n7723) );
  AND2X2 AND2X2_4383 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core_v2_reg_23_), .Y(core__abc_21380_n7724) );
  AND2X2 AND2X2_4384 ( .A(core__abc_21380_n7728), .B(reset_n_bF_buf62), .Y(core__abc_21380_n7729) );
  AND2X2 AND2X2_4385 ( .A(core__abc_21380_n7727), .B(core__abc_21380_n7729), .Y(core_v2_reg_23__FF_INPUT) );
  AND2X2 AND2X2_4386 ( .A(core__abc_21380_n7715), .B(core__abc_21380_n7692), .Y(core__abc_21380_n7732) );
  AND2X2 AND2X2_4387 ( .A(core__abc_21380_n7735), .B(core__abc_21380_n7630), .Y(core__abc_21380_n7736) );
  AND2X2 AND2X2_4388 ( .A(core__abc_21380_n7735), .B(core__abc_21380_n7628), .Y(core__abc_21380_n7739) );
  AND2X2 AND2X2_4389 ( .A(core__abc_21380_n7681), .B(core__abc_21380_n7732), .Y(core__abc_21380_n7740) );
  AND2X2 AND2X2_439 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_107_), .Y(_abc_19068_n1664) );
  AND2X2 AND2X2_4390 ( .A(core__abc_21380_n7714), .B(core__abc_21380_n7688), .Y(core__abc_21380_n7741) );
  AND2X2 AND2X2_4391 ( .A(core__abc_21380_n7738), .B(core__abc_21380_n7745), .Y(core__abc_21380_n7746) );
  AND2X2 AND2X2_4392 ( .A(core__abc_21380_n7747), .B(core__abc_21380_n7748), .Y(core__abc_21380_n7749) );
  AND2X2 AND2X2_4393 ( .A(core__abc_21380_n4198_1), .B(core__abc_21380_n7749), .Y(core__abc_21380_n7750) );
  AND2X2 AND2X2_4394 ( .A(core__abc_21380_n4199), .B(core__abc_21380_n7751), .Y(core__abc_21380_n7752) );
  AND2X2 AND2X2_4395 ( .A(core__abc_21380_n7746), .B(core__abc_21380_n7753), .Y(core__abc_21380_n7754) );
  AND2X2 AND2X2_4396 ( .A(core__abc_21380_n7758), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n7759) );
  AND2X2 AND2X2_4397 ( .A(core__abc_21380_n3313_bF_buf1), .B(core_key_24_), .Y(core__abc_21380_n7760) );
  AND2X2 AND2X2_4398 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core_v2_reg_24_), .Y(core__abc_21380_n7761) );
  AND2X2 AND2X2_4399 ( .A(core__abc_21380_n7765), .B(reset_n_bF_buf61), .Y(core__abc_21380_n7766) );
  AND2X2 AND2X2_44 ( .A(_abc_19068_n939_1_bF_buf4), .B(core_key_64_), .Y(_abc_19068_n940_1) );
  AND2X2 AND2X2_440 ( .A(_abc_19068_n1620_bF_buf10), .B(word3_reg_11_), .Y(_abc_19068_n1665) );
  AND2X2 AND2X2_4400 ( .A(core__abc_21380_n7764), .B(core__abc_21380_n7766), .Y(core_v2_reg_24__FF_INPUT) );
  AND2X2 AND2X2_4401 ( .A(core__abc_21380_n7755), .B(core__abc_21380_n7768), .Y(core__abc_21380_n7769) );
  AND2X2 AND2X2_4402 ( .A(core__abc_21380_n4936), .B(core__abc_21380_n2079), .Y(core__abc_21380_n7770) );
  AND2X2 AND2X2_4403 ( .A(core__abc_21380_n7771), .B(core__abc_21380_n7772), .Y(core__abc_21380_n7773) );
  AND2X2 AND2X2_4404 ( .A(core__abc_21380_n4270), .B(core__abc_21380_n7773), .Y(core__abc_21380_n7774) );
  AND2X2 AND2X2_4405 ( .A(core__abc_21380_n4268), .B(core__abc_21380_n7776), .Y(core__abc_21380_n7777) );
  AND2X2 AND2X2_4406 ( .A(core__abc_21380_n7775), .B(core__abc_21380_n7778), .Y(core__abc_21380_n7779) );
  AND2X2 AND2X2_4407 ( .A(core__abc_21380_n7783), .B(core__abc_21380_n7780), .Y(core__abc_21380_n7784) );
  AND2X2 AND2X2_4408 ( .A(core__abc_21380_n7785), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n7786) );
  AND2X2 AND2X2_4409 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n7787), .Y(core__abc_21380_n7788) );
  AND2X2 AND2X2_441 ( .A(_abc_19068_n1666), .B(reset_n_bF_buf73), .Y(word3_reg_11__FF_INPUT) );
  AND2X2 AND2X2_4410 ( .A(core__abc_21380_n3163_1_bF_buf1), .B(core_v2_reg_25_), .Y(core__abc_21380_n7789) );
  AND2X2 AND2X2_4411 ( .A(core__abc_21380_n7793), .B(reset_n_bF_buf60), .Y(core__abc_21380_n7794) );
  AND2X2 AND2X2_4412 ( .A(core__abc_21380_n7792), .B(core__abc_21380_n7794), .Y(core_v2_reg_25__FF_INPUT) );
  AND2X2 AND2X2_4413 ( .A(core__abc_21380_n7796), .B(core__abc_21380_n7797), .Y(core__abc_21380_n7798) );
  AND2X2 AND2X2_4414 ( .A(core__abc_21380_n4331), .B(core__abc_21380_n7798), .Y(core__abc_21380_n7799) );
  AND2X2 AND2X2_4415 ( .A(core__abc_21380_n4328), .B(core__abc_21380_n7800), .Y(core__abc_21380_n7801) );
  AND2X2 AND2X2_4416 ( .A(core__abc_21380_n7775), .B(core__abc_21380_n7768), .Y(core__abc_21380_n7805) );
  AND2X2 AND2X2_4417 ( .A(core__abc_21380_n7804), .B(core__abc_21380_n7806), .Y(core__abc_21380_n7807) );
  AND2X2 AND2X2_4418 ( .A(core__abc_21380_n7807), .B(core__abc_21380_n7802), .Y(core__abc_21380_n7808) );
  AND2X2 AND2X2_4419 ( .A(core__abc_21380_n7812), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n7813) );
  AND2X2 AND2X2_442 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_108_), .Y(_abc_19068_n1668) );
  AND2X2 AND2X2_4420 ( .A(core__abc_21380_n3313_bF_buf12), .B(core__abc_21380_n7814), .Y(core__abc_21380_n7815) );
  AND2X2 AND2X2_4421 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core_v2_reg_26_), .Y(core__abc_21380_n7816) );
  AND2X2 AND2X2_4422 ( .A(core__abc_21380_n7820), .B(reset_n_bF_buf59), .Y(core__abc_21380_n7821) );
  AND2X2 AND2X2_4423 ( .A(core__abc_21380_n7819), .B(core__abc_21380_n7821), .Y(core_v2_reg_26__FF_INPUT) );
  AND2X2 AND2X2_4424 ( .A(core__abc_21380_n7809), .B(core__abc_21380_n7823), .Y(core__abc_21380_n7824) );
  AND2X2 AND2X2_4425 ( .A(core__abc_21380_n5043), .B(core__abc_21380_n2117), .Y(core__abc_21380_n7825) );
  AND2X2 AND2X2_4426 ( .A(core__abc_21380_n5031), .B(core_v1_reg_46_), .Y(core__abc_21380_n7826) );
  AND2X2 AND2X2_4427 ( .A(core__abc_21380_n4422_1), .B(core__abc_21380_n7828), .Y(core__abc_21380_n7829) );
  AND2X2 AND2X2_4428 ( .A(core__abc_21380_n7831), .B(core__abc_21380_n7827), .Y(core__abc_21380_n7832) );
  AND2X2 AND2X2_4429 ( .A(core__abc_21380_n7833), .B(core__abc_21380_n7830), .Y(core__abc_21380_n7834) );
  AND2X2 AND2X2_443 ( .A(_abc_19068_n1620_bF_buf9), .B(word3_reg_12_), .Y(_abc_19068_n1669) );
  AND2X2 AND2X2_4430 ( .A(core__abc_21380_n7824), .B(core__abc_21380_n7835), .Y(core__abc_21380_n7836) );
  AND2X2 AND2X2_4431 ( .A(core__abc_21380_n7837), .B(core__abc_21380_n7834), .Y(core__abc_21380_n7838) );
  AND2X2 AND2X2_4432 ( .A(core__abc_21380_n7840), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n7841) );
  AND2X2 AND2X2_4433 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n7842), .Y(core__abc_21380_n7843) );
  AND2X2 AND2X2_4434 ( .A(core__abc_21380_n3163_1_bF_buf6), .B(core_v2_reg_27_), .Y(core__abc_21380_n7844) );
  AND2X2 AND2X2_4435 ( .A(core__abc_21380_n7848), .B(reset_n_bF_buf58), .Y(core__abc_21380_n7849) );
  AND2X2 AND2X2_4436 ( .A(core__abc_21380_n7847), .B(core__abc_21380_n7849), .Y(core_v2_reg_27__FF_INPUT) );
  AND2X2 AND2X2_4437 ( .A(core__abc_21380_n7516), .B(core__abc_21380_n7736), .Y(core__abc_21380_n7851) );
  AND2X2 AND2X2_4438 ( .A(core__abc_21380_n7852), .B(core__abc_21380_n7855), .Y(core__abc_21380_n7856) );
  AND2X2 AND2X2_4439 ( .A(core__abc_21380_n7833), .B(core__abc_21380_n7801), .Y(core__abc_21380_n7858) );
  AND2X2 AND2X2_444 ( .A(_abc_19068_n1670), .B(reset_n_bF_buf72), .Y(word3_reg_12__FF_INPUT) );
  AND2X2 AND2X2_4440 ( .A(core__abc_21380_n7857), .B(core__abc_21380_n7860), .Y(core__abc_21380_n7861) );
  AND2X2 AND2X2_4441 ( .A(core__abc_21380_n7864), .B(core__abc_21380_n7865), .Y(core__abc_21380_n7866) );
  AND2X2 AND2X2_4442 ( .A(core__abc_21380_n4490), .B(core__abc_21380_n7866), .Y(core__abc_21380_n7867) );
  AND2X2 AND2X2_4443 ( .A(core__abc_21380_n4491_1), .B(core__abc_21380_n7868), .Y(core__abc_21380_n7869) );
  AND2X2 AND2X2_4444 ( .A(core__abc_21380_n7863), .B(core__abc_21380_n7871), .Y(core__abc_21380_n7872) );
  AND2X2 AND2X2_4445 ( .A(core__abc_21380_n7873), .B(core__abc_21380_n7861), .Y(core__abc_21380_n7874) );
  AND2X2 AND2X2_4446 ( .A(core__abc_21380_n7874), .B(core__abc_21380_n7870), .Y(core__abc_21380_n7875) );
  AND2X2 AND2X2_4447 ( .A(core__abc_21380_n7877), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n7878) );
  AND2X2 AND2X2_4448 ( .A(core__abc_21380_n3313_bF_buf10), .B(core_key_28_), .Y(core__abc_21380_n7879) );
  AND2X2 AND2X2_4449 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core_v2_reg_28_), .Y(core__abc_21380_n7880) );
  AND2X2 AND2X2_445 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_109_), .Y(_abc_19068_n1672) );
  AND2X2 AND2X2_4450 ( .A(core__abc_21380_n7884), .B(reset_n_bF_buf57), .Y(core__abc_21380_n7885) );
  AND2X2 AND2X2_4451 ( .A(core__abc_21380_n7883), .B(core__abc_21380_n7885), .Y(core_v2_reg_28__FF_INPUT) );
  AND2X2 AND2X2_4452 ( .A(core__abc_21380_n5149), .B(core_v1_reg_48_), .Y(core__abc_21380_n7889) );
  AND2X2 AND2X2_4453 ( .A(core__abc_21380_n5148), .B(core__abc_21380_n2154), .Y(core__abc_21380_n7890) );
  AND2X2 AND2X2_4454 ( .A(core__abc_21380_n7888), .B(core__abc_21380_n7891), .Y(core__abc_21380_n7892) );
  AND2X2 AND2X2_4455 ( .A(core__abc_21380_n4550), .B(core__abc_21380_n7893), .Y(core__abc_21380_n7894) );
  AND2X2 AND2X2_4456 ( .A(core__abc_21380_n7899), .B(core__abc_21380_n7896), .Y(core__abc_21380_n7900) );
  AND2X2 AND2X2_4457 ( .A(core__abc_21380_n7901), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf1), .Y(core__abc_21380_n7902) );
  AND2X2 AND2X2_4458 ( .A(core__abc_21380_n3313_bF_buf9), .B(core__abc_21380_n7903), .Y(core__abc_21380_n7904) );
  AND2X2 AND2X2_4459 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core_v2_reg_29_), .Y(core__abc_21380_n7905) );
  AND2X2 AND2X2_446 ( .A(_abc_19068_n1620_bF_buf8), .B(word3_reg_13_), .Y(_abc_19068_n1673) );
  AND2X2 AND2X2_4460 ( .A(core__abc_21380_n7909), .B(reset_n_bF_buf56), .Y(core__abc_21380_n7910) );
  AND2X2 AND2X2_4461 ( .A(core__abc_21380_n7908), .B(core__abc_21380_n7910), .Y(core_v2_reg_29__FF_INPUT) );
  AND2X2 AND2X2_4462 ( .A(core__abc_21380_n7898), .B(core__abc_21380_n7871), .Y(core__abc_21380_n7912) );
  AND2X2 AND2X2_4463 ( .A(core__abc_21380_n7898), .B(core__abc_21380_n7869), .Y(core__abc_21380_n7915) );
  AND2X2 AND2X2_4464 ( .A(core__abc_21380_n7914), .B(core__abc_21380_n7917), .Y(core__abc_21380_n7918) );
  AND2X2 AND2X2_4465 ( .A(core__abc_21380_n7919), .B(core__abc_21380_n7920), .Y(core__abc_21380_n7921) );
  AND2X2 AND2X2_4466 ( .A(core__abc_21380_n4583), .B(core__abc_21380_n7922), .Y(core__abc_21380_n7923) );
  AND2X2 AND2X2_4467 ( .A(core__abc_21380_n4581), .B(core__abc_21380_n7921), .Y(core__abc_21380_n7924) );
  AND2X2 AND2X2_4468 ( .A(core__abc_21380_n7918), .B(core__abc_21380_n7925), .Y(core__abc_21380_n7926) );
  AND2X2 AND2X2_4469 ( .A(core__abc_21380_n7863), .B(core__abc_21380_n7912), .Y(core__abc_21380_n7927) );
  AND2X2 AND2X2_447 ( .A(_abc_19068_n1674), .B(reset_n_bF_buf71), .Y(word3_reg_13__FF_INPUT) );
  AND2X2 AND2X2_4470 ( .A(core__abc_21380_n7928), .B(core__abc_21380_n7929), .Y(core__abc_21380_n7930) );
  AND2X2 AND2X2_4471 ( .A(core__abc_21380_n7932), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf1), .Y(core__abc_21380_n7933) );
  AND2X2 AND2X2_4472 ( .A(core__abc_21380_n3313_bF_buf8), .B(core__abc_21380_n7934), .Y(core__abc_21380_n7935) );
  AND2X2 AND2X2_4473 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core_v2_reg_30_), .Y(core__abc_21380_n7936) );
  AND2X2 AND2X2_4474 ( .A(core__abc_21380_n7940), .B(reset_n_bF_buf55), .Y(core__abc_21380_n7941) );
  AND2X2 AND2X2_4475 ( .A(core__abc_21380_n7939), .B(core__abc_21380_n7941), .Y(core_v2_reg_30__FF_INPUT) );
  AND2X2 AND2X2_4476 ( .A(core__abc_21380_n7944), .B(core__abc_21380_n7943), .Y(core__abc_21380_n7945) );
  AND2X2 AND2X2_4477 ( .A(core__abc_21380_n5255), .B(core__abc_21380_n2191), .Y(core__abc_21380_n7946) );
  AND2X2 AND2X2_4478 ( .A(core__abc_21380_n5270), .B(core_v1_reg_50_), .Y(core__abc_21380_n7947) );
  AND2X2 AND2X2_4479 ( .A(core__abc_21380_n7950), .B(core__abc_21380_n7951), .Y(core__abc_21380_n7952) );
  AND2X2 AND2X2_448 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_110_), .Y(_abc_19068_n1676) );
  AND2X2 AND2X2_4480 ( .A(core__abc_21380_n7945), .B(core__abc_21380_n7953), .Y(core__abc_21380_n7954) );
  AND2X2 AND2X2_4481 ( .A(core__abc_21380_n7955), .B(core__abc_21380_n7956), .Y(core__abc_21380_n7957) );
  AND2X2 AND2X2_4482 ( .A(core__abc_21380_n7957), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n7958) );
  AND2X2 AND2X2_4483 ( .A(core__abc_21380_n3313_bF_buf7), .B(core_key_31_), .Y(core__abc_21380_n7959) );
  AND2X2 AND2X2_4484 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core_v2_reg_31_), .Y(core__abc_21380_n7960) );
  AND2X2 AND2X2_4485 ( .A(core__abc_21380_n7964), .B(reset_n_bF_buf54), .Y(core__abc_21380_n7965) );
  AND2X2 AND2X2_4486 ( .A(core__abc_21380_n7963), .B(core__abc_21380_n7965), .Y(core_v2_reg_31__FF_INPUT) );
  AND2X2 AND2X2_4487 ( .A(core__abc_21380_n3313_bF_buf6), .B(core__abc_21380_n7967), .Y(core__abc_21380_n7968) );
  AND2X2 AND2X2_4488 ( .A(core__abc_21380_n7969), .B(core__abc_21380_n1267), .Y(core__abc_21380_n7970) );
  AND2X2 AND2X2_4489 ( .A(core__abc_21380_n3167_1_bF_buf12), .B(core__abc_21380_n7972), .Y(core__abc_21380_n7973) );
  AND2X2 AND2X2_449 ( .A(_abc_19068_n1620_bF_buf7), .B(word3_reg_14_), .Y(_abc_19068_n1677) );
  AND2X2 AND2X2_4490 ( .A(core__abc_21380_n7087_bF_buf7), .B(core__abc_21380_n7974), .Y(core__abc_21380_n7975) );
  AND2X2 AND2X2_4491 ( .A(core__abc_21380_n7976), .B(core_v2_reg_32_), .Y(core__abc_21380_n7977) );
  AND2X2 AND2X2_4492 ( .A(core__abc_21380_n7978), .B(reset_n_bF_buf53), .Y(core_v2_reg_32__FF_INPUT) );
  AND2X2 AND2X2_4493 ( .A(core__abc_21380_n7980), .B(core__abc_21380_n7981), .Y(core__abc_21380_n7982) );
  AND2X2 AND2X2_4494 ( .A(core__abc_21380_n7982), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n7983) );
  AND2X2 AND2X2_4495 ( .A(core__abc_21380_n3313_bF_buf5), .B(core_key_33_), .Y(core__abc_21380_n7984) );
  AND2X2 AND2X2_4496 ( .A(core__abc_21380_n7985), .B(core__abc_21380_n7087_bF_buf6), .Y(core__abc_21380_n7986) );
  AND2X2 AND2X2_4497 ( .A(core__abc_21380_n7976), .B(core_v2_reg_33_), .Y(core__abc_21380_n7987) );
  AND2X2 AND2X2_4498 ( .A(core__abc_21380_n7988), .B(reset_n_bF_buf52), .Y(core_v2_reg_33__FF_INPUT) );
  AND2X2 AND2X2_4499 ( .A(core__abc_21380_n7976), .B(core_v2_reg_34_), .Y(core__abc_21380_n7990) );
  AND2X2 AND2X2_45 ( .A(_abc_19068_n912_1), .B(_abc_19068_n898_1), .Y(_abc_19068_n941) );
  AND2X2 AND2X2_450 ( .A(_abc_19068_n1678), .B(reset_n_bF_buf70), .Y(word3_reg_14__FF_INPUT) );
  AND2X2 AND2X2_4500 ( .A(core__abc_21380_n7991), .B(core__abc_21380_n7992), .Y(core__abc_21380_n7993) );
  AND2X2 AND2X2_4501 ( .A(core__abc_21380_n7993), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n7994) );
  AND2X2 AND2X2_4502 ( .A(core__abc_21380_n3313_bF_buf4), .B(core__abc_21380_n7995), .Y(core__abc_21380_n7996) );
  AND2X2 AND2X2_4503 ( .A(core__abc_21380_n7997), .B(core__abc_21380_n7087_bF_buf5), .Y(core__abc_21380_n7998) );
  AND2X2 AND2X2_4504 ( .A(core__abc_21380_n7999), .B(reset_n_bF_buf51), .Y(core_v2_reg_34__FF_INPUT) );
  AND2X2 AND2X2_4505 ( .A(core__abc_21380_n8001), .B(core__abc_21380_n8002), .Y(core__abc_21380_n8003) );
  AND2X2 AND2X2_4506 ( .A(core__abc_21380_n8003), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n8004) );
  AND2X2 AND2X2_4507 ( .A(core__abc_21380_n3313_bF_buf3), .B(core_key_35_), .Y(core__abc_21380_n8005) );
  AND2X2 AND2X2_4508 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core_v2_reg_35_), .Y(core__abc_21380_n8006) );
  AND2X2 AND2X2_4509 ( .A(core__abc_21380_n8010), .B(reset_n_bF_buf50), .Y(core__abc_21380_n8011) );
  AND2X2 AND2X2_451 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_111_), .Y(_abc_19068_n1680) );
  AND2X2 AND2X2_4510 ( .A(core__abc_21380_n8009), .B(core__abc_21380_n8011), .Y(core_v2_reg_35__FF_INPUT) );
  AND2X2 AND2X2_4511 ( .A(core__abc_21380_n8013), .B(core__abc_21380_n8014), .Y(core__abc_21380_n8015) );
  AND2X2 AND2X2_4512 ( .A(core__abc_21380_n8015), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n8016) );
  AND2X2 AND2X2_4513 ( .A(core__abc_21380_n3313_bF_buf2), .B(core_key_36_), .Y(core__abc_21380_n8017) );
  AND2X2 AND2X2_4514 ( .A(core__abc_21380_n3163_1_bF_buf6), .B(core_v2_reg_36_), .Y(core__abc_21380_n8018) );
  AND2X2 AND2X2_4515 ( .A(core__abc_21380_n8022), .B(reset_n_bF_buf49), .Y(core__abc_21380_n8023) );
  AND2X2 AND2X2_4516 ( .A(core__abc_21380_n8021), .B(core__abc_21380_n8023), .Y(core_v2_reg_36__FF_INPUT) );
  AND2X2 AND2X2_4517 ( .A(core__abc_21380_n8025), .B(core__abc_21380_n8026), .Y(core__abc_21380_n8027) );
  AND2X2 AND2X2_4518 ( .A(core__abc_21380_n8027), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n8028) );
  AND2X2 AND2X2_4519 ( .A(core__abc_21380_n3313_bF_buf1), .B(core__abc_21380_n8029), .Y(core__abc_21380_n8030) );
  AND2X2 AND2X2_452 ( .A(_abc_19068_n1620_bF_buf6), .B(word3_reg_15_), .Y(_abc_19068_n1681) );
  AND2X2 AND2X2_4520 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core_v2_reg_37_), .Y(core__abc_21380_n8031) );
  AND2X2 AND2X2_4521 ( .A(core__abc_21380_n8035), .B(reset_n_bF_buf48), .Y(core__abc_21380_n8036) );
  AND2X2 AND2X2_4522 ( .A(core__abc_21380_n8034), .B(core__abc_21380_n8036), .Y(core_v2_reg_37__FF_INPUT) );
  AND2X2 AND2X2_4523 ( .A(core__abc_21380_n7034), .B(core__abc_21380_n6976), .Y(core__abc_21380_n8038) );
  AND2X2 AND2X2_4524 ( .A(core__abc_21380_n8039), .B(core__abc_21380_n8040), .Y(core__abc_21380_n8041) );
  AND2X2 AND2X2_4525 ( .A(core__abc_21380_n8041), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n8042) );
  AND2X2 AND2X2_4526 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n8043), .Y(core__abc_21380_n8044) );
  AND2X2 AND2X2_4527 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core_v2_reg_38_), .Y(core__abc_21380_n8045) );
  AND2X2 AND2X2_4528 ( .A(core__abc_21380_n8049), .B(reset_n_bF_buf47), .Y(core__abc_21380_n8050) );
  AND2X2 AND2X2_4529 ( .A(core__abc_21380_n8048), .B(core__abc_21380_n8050), .Y(core_v2_reg_38__FF_INPUT) );
  AND2X2 AND2X2_453 ( .A(_abc_19068_n1682), .B(reset_n_bF_buf69), .Y(word3_reg_15__FF_INPUT) );
  AND2X2 AND2X2_4530 ( .A(core__abc_21380_n8056), .B(core__abc_21380_n8053), .Y(core__abc_21380_n8057) );
  AND2X2 AND2X2_4531 ( .A(core__abc_21380_n8057), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n8058) );
  AND2X2 AND2X2_4532 ( .A(core__abc_21380_n3313_bF_buf12), .B(core_key_39_), .Y(core__abc_21380_n8059) );
  AND2X2 AND2X2_4533 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core_v2_reg_39_), .Y(core__abc_21380_n8060) );
  AND2X2 AND2X2_4534 ( .A(core__abc_21380_n8064), .B(reset_n_bF_buf46), .Y(core__abc_21380_n8065) );
  AND2X2 AND2X2_4535 ( .A(core__abc_21380_n8063), .B(core__abc_21380_n8065), .Y(core_v2_reg_39__FF_INPUT) );
  AND2X2 AND2X2_4536 ( .A(core__abc_21380_n8067), .B(core__abc_21380_n7040), .Y(core__abc_21380_n8068) );
  AND2X2 AND2X2_4537 ( .A(core__abc_21380_n7036), .B(core__abc_21380_n7041), .Y(core__abc_21380_n8069) );
  AND2X2 AND2X2_4538 ( .A(core__abc_21380_n8071), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n8072) );
  AND2X2 AND2X2_4539 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n8073), .Y(core__abc_21380_n8074) );
  AND2X2 AND2X2_454 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_112_), .Y(_abc_19068_n1684) );
  AND2X2 AND2X2_4540 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core_v2_reg_40_), .Y(core__abc_21380_n8075) );
  AND2X2 AND2X2_4541 ( .A(core__abc_21380_n8079), .B(reset_n_bF_buf45), .Y(core__abc_21380_n8080) );
  AND2X2 AND2X2_4542 ( .A(core__abc_21380_n8078), .B(core__abc_21380_n8080), .Y(core_v2_reg_40__FF_INPUT) );
  AND2X2 AND2X2_4543 ( .A(core__abc_21380_n8084), .B(core__abc_21380_n8082), .Y(core__abc_21380_n8085) );
  AND2X2 AND2X2_4544 ( .A(core__abc_21380_n8083), .B(core__abc_21380_n7038), .Y(core__abc_21380_n8086) );
  AND2X2 AND2X2_4545 ( .A(core__abc_21380_n8088), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n8089) );
  AND2X2 AND2X2_4546 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n8090), .Y(core__abc_21380_n8091) );
  AND2X2 AND2X2_4547 ( .A(core__abc_21380_n3163_1_bF_buf1), .B(core_v2_reg_41_), .Y(core__abc_21380_n8092) );
  AND2X2 AND2X2_4548 ( .A(core__abc_21380_n8096), .B(reset_n_bF_buf44), .Y(core__abc_21380_n8097) );
  AND2X2 AND2X2_4549 ( .A(core__abc_21380_n8095), .B(core__abc_21380_n8097), .Y(core_v2_reg_41__FF_INPUT) );
  AND2X2 AND2X2_455 ( .A(_abc_19068_n1620_bF_buf5), .B(word3_reg_16_), .Y(_abc_19068_n1685) );
  AND2X2 AND2X2_4550 ( .A(core__abc_21380_n7036), .B(core__abc_21380_n7042), .Y(core__abc_21380_n8099) );
  AND2X2 AND2X2_4551 ( .A(core__abc_21380_n8100), .B(core__abc_21380_n6954), .Y(core__abc_21380_n8101) );
  AND2X2 AND2X2_4552 ( .A(core__abc_21380_n8102), .B(core__abc_21380_n8103), .Y(core__abc_21380_n8104) );
  AND2X2 AND2X2_4553 ( .A(core__abc_21380_n8104), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n8105) );
  AND2X2 AND2X2_4554 ( .A(core__abc_21380_n3313_bF_buf9), .B(core__abc_21380_n8106), .Y(core__abc_21380_n8107) );
  AND2X2 AND2X2_4555 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core_v2_reg_42_), .Y(core__abc_21380_n8108) );
  AND2X2 AND2X2_4556 ( .A(core__abc_21380_n8112), .B(reset_n_bF_buf43), .Y(core__abc_21380_n8113) );
  AND2X2 AND2X2_4557 ( .A(core__abc_21380_n8111), .B(core__abc_21380_n8113), .Y(core_v2_reg_42__FF_INPUT) );
  AND2X2 AND2X2_4558 ( .A(core__abc_21380_n8102), .B(core__abc_21380_n6929), .Y(core__abc_21380_n8116) );
  AND2X2 AND2X2_4559 ( .A(core__abc_21380_n8116), .B(core__abc_21380_n8115), .Y(core__abc_21380_n8117) );
  AND2X2 AND2X2_456 ( .A(_abc_19068_n1686), .B(reset_n_bF_buf68), .Y(word3_reg_16__FF_INPUT) );
  AND2X2 AND2X2_4560 ( .A(core__abc_21380_n8118), .B(core__abc_21380_n8119), .Y(core__abc_21380_n8120) );
  AND2X2 AND2X2_4561 ( .A(core__abc_21380_n8120), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n8121) );
  AND2X2 AND2X2_4562 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_43_), .Y(core__abc_21380_n8122) );
  AND2X2 AND2X2_4563 ( .A(core__abc_21380_n3163_1_bF_buf6), .B(core_v2_reg_43_), .Y(core__abc_21380_n8123) );
  AND2X2 AND2X2_4564 ( .A(core__abc_21380_n8127), .B(reset_n_bF_buf42), .Y(core__abc_21380_n8128) );
  AND2X2 AND2X2_4565 ( .A(core__abc_21380_n8126), .B(core__abc_21380_n8128), .Y(core_v2_reg_43__FF_INPUT) );
  AND2X2 AND2X2_4566 ( .A(core__abc_21380_n7045), .B(core__abc_21380_n6916), .Y(core__abc_21380_n8130) );
  AND2X2 AND2X2_4567 ( .A(core__abc_21380_n8131), .B(core__abc_21380_n6915), .Y(core__abc_21380_n8132) );
  AND2X2 AND2X2_4568 ( .A(core__abc_21380_n8134), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n8135) );
  AND2X2 AND2X2_4569 ( .A(core__abc_21380_n3313_bF_buf7), .B(core_key_44_), .Y(core__abc_21380_n8136) );
  AND2X2 AND2X2_457 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_113_), .Y(_abc_19068_n1688) );
  AND2X2 AND2X2_4570 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core_v2_reg_44_), .Y(core__abc_21380_n8137) );
  AND2X2 AND2X2_4571 ( .A(core__abc_21380_n8141), .B(reset_n_bF_buf41), .Y(core__abc_21380_n8142) );
  AND2X2 AND2X2_4572 ( .A(core__abc_21380_n8140), .B(core__abc_21380_n8142), .Y(core_v2_reg_44__FF_INPUT) );
  AND2X2 AND2X2_4573 ( .A(core__abc_21380_n8145), .B(core__abc_21380_n8144), .Y(core__abc_21380_n8146) );
  AND2X2 AND2X2_4574 ( .A(core__abc_21380_n8147), .B(core__abc_21380_n8148), .Y(core__abc_21380_n8149) );
  AND2X2 AND2X2_4575 ( .A(core__abc_21380_n8150), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf0), .Y(core__abc_21380_n8151) );
  AND2X2 AND2X2_4576 ( .A(core__abc_21380_n3313_bF_buf6), .B(core__abc_21380_n8152), .Y(core__abc_21380_n8153) );
  AND2X2 AND2X2_4577 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core_v2_reg_45_), .Y(core__abc_21380_n8154) );
  AND2X2 AND2X2_4578 ( .A(core__abc_21380_n8158), .B(reset_n_bF_buf40), .Y(core__abc_21380_n8159) );
  AND2X2 AND2X2_4579 ( .A(core__abc_21380_n8157), .B(core__abc_21380_n8159), .Y(core_v2_reg_45__FF_INPUT) );
  AND2X2 AND2X2_458 ( .A(_abc_19068_n1620_bF_buf4), .B(word3_reg_17_), .Y(_abc_19068_n1689) );
  AND2X2 AND2X2_4580 ( .A(core__abc_21380_n7045), .B(core__abc_21380_n6917), .Y(core__abc_21380_n8161) );
  AND2X2 AND2X2_4581 ( .A(core__abc_21380_n8162), .B(core__abc_21380_n6889), .Y(core__abc_21380_n8163) );
  AND2X2 AND2X2_4582 ( .A(core__abc_21380_n8164), .B(core__abc_21380_n8165), .Y(core__abc_21380_n8166) );
  AND2X2 AND2X2_4583 ( .A(core__abc_21380_n8166), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf0), .Y(core__abc_21380_n8167) );
  AND2X2 AND2X2_4584 ( .A(core__abc_21380_n3313_bF_buf5), .B(core__abc_21380_n8168), .Y(core__abc_21380_n8169) );
  AND2X2 AND2X2_4585 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core_v2_reg_46_), .Y(core__abc_21380_n8170) );
  AND2X2 AND2X2_4586 ( .A(core__abc_21380_n8174), .B(reset_n_bF_buf39), .Y(core__abc_21380_n8175) );
  AND2X2 AND2X2_4587 ( .A(core__abc_21380_n8173), .B(core__abc_21380_n8175), .Y(core_v2_reg_46__FF_INPUT) );
  AND2X2 AND2X2_4588 ( .A(core__abc_21380_n8179), .B(core__abc_21380_n8177), .Y(core__abc_21380_n8180) );
  AND2X2 AND2X2_4589 ( .A(core__abc_21380_n8178), .B(core__abc_21380_n6881), .Y(core__abc_21380_n8181) );
  AND2X2 AND2X2_459 ( .A(_abc_19068_n1690), .B(reset_n_bF_buf67), .Y(word3_reg_17__FF_INPUT) );
  AND2X2 AND2X2_4590 ( .A(core__abc_21380_n8183), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n8184) );
  AND2X2 AND2X2_4591 ( .A(core__abc_21380_n3313_bF_buf4), .B(core_key_47_), .Y(core__abc_21380_n8185) );
  AND2X2 AND2X2_4592 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core_v2_reg_47_), .Y(core__abc_21380_n8186) );
  AND2X2 AND2X2_4593 ( .A(core__abc_21380_n8190), .B(reset_n_bF_buf38), .Y(core__abc_21380_n8191) );
  AND2X2 AND2X2_4594 ( .A(core__abc_21380_n8189), .B(core__abc_21380_n8191), .Y(core_v2_reg_47__FF_INPUT) );
  AND2X2 AND2X2_4595 ( .A(core__abc_21380_n8193), .B(core__abc_21380_n7051), .Y(core__abc_21380_n8194) );
  AND2X2 AND2X2_4596 ( .A(core__abc_21380_n7047), .B(core__abc_21380_n7052), .Y(core__abc_21380_n8195) );
  AND2X2 AND2X2_4597 ( .A(core__abc_21380_n8197), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n8198) );
  AND2X2 AND2X2_4598 ( .A(core__abc_21380_n3313_bF_buf3), .B(core__abc_21380_n8199), .Y(core__abc_21380_n8200) );
  AND2X2 AND2X2_4599 ( .A(core__abc_21380_n3163_1_bF_buf1), .B(core_v2_reg_48_), .Y(core__abc_21380_n8201) );
  AND2X2 AND2X2_46 ( .A(_abc_19068_n941_bF_buf4), .B(core_key_96_), .Y(_abc_19068_n942_1) );
  AND2X2 AND2X2_460 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_114_), .Y(_abc_19068_n1692) );
  AND2X2 AND2X2_4600 ( .A(core__abc_21380_n8205), .B(reset_n_bF_buf37), .Y(core__abc_21380_n8206) );
  AND2X2 AND2X2_4601 ( .A(core__abc_21380_n8204), .B(core__abc_21380_n8206), .Y(core_v2_reg_48__FF_INPUT) );
  AND2X2 AND2X2_4602 ( .A(core__abc_21380_n8209), .B(core__abc_21380_n8208), .Y(core__abc_21380_n8210) );
  AND2X2 AND2X2_4603 ( .A(core__abc_21380_n8211), .B(core__abc_21380_n7049), .Y(core__abc_21380_n8212) );
  AND2X2 AND2X2_4604 ( .A(core__abc_21380_n8213), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n8214) );
  AND2X2 AND2X2_4605 ( .A(core__abc_21380_n3313_bF_buf2), .B(core_key_49_), .Y(core__abc_21380_n8215) );
  AND2X2 AND2X2_4606 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core_v2_reg_49_), .Y(core__abc_21380_n8216) );
  AND2X2 AND2X2_4607 ( .A(core__abc_21380_n8220), .B(reset_n_bF_buf36), .Y(core__abc_21380_n8221) );
  AND2X2 AND2X2_4608 ( .A(core__abc_21380_n8219), .B(core__abc_21380_n8221), .Y(core_v2_reg_49__FF_INPUT) );
  AND2X2 AND2X2_4609 ( .A(core__abc_21380_n8211), .B(core__abc_21380_n7048), .Y(core__abc_21380_n8223) );
  AND2X2 AND2X2_461 ( .A(_abc_19068_n1620_bF_buf3), .B(word3_reg_18_), .Y(_abc_19068_n1693) );
  AND2X2 AND2X2_4610 ( .A(core__abc_21380_n8225), .B(core__abc_21380_n6838), .Y(core__abc_21380_n8226) );
  AND2X2 AND2X2_4611 ( .A(core__abc_21380_n8224), .B(core__abc_21380_n6837), .Y(core__abc_21380_n8227) );
  AND2X2 AND2X2_4612 ( .A(core__abc_21380_n8229), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n8230) );
  AND2X2 AND2X2_4613 ( .A(core__abc_21380_n3313_bF_buf1), .B(core_key_50_), .Y(core__abc_21380_n8231) );
  AND2X2 AND2X2_4614 ( .A(core__abc_21380_n3163_1_bF_buf6), .B(core_v2_reg_50_), .Y(core__abc_21380_n8232) );
  AND2X2 AND2X2_4615 ( .A(core__abc_21380_n8236), .B(reset_n_bF_buf35), .Y(core__abc_21380_n8237) );
  AND2X2 AND2X2_4616 ( .A(core__abc_21380_n8235), .B(core__abc_21380_n8237), .Y(core_v2_reg_50__FF_INPUT) );
  AND2X2 AND2X2_4617 ( .A(core__abc_21380_n8241), .B(core__abc_21380_n8239), .Y(core__abc_21380_n8242) );
  AND2X2 AND2X2_4618 ( .A(core__abc_21380_n8240), .B(core__abc_21380_n6830), .Y(core__abc_21380_n8243) );
  AND2X2 AND2X2_4619 ( .A(core__abc_21380_n8245), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n8246) );
  AND2X2 AND2X2_462 ( .A(_abc_19068_n1694), .B(reset_n_bF_buf66), .Y(word3_reg_18__FF_INPUT) );
  AND2X2 AND2X2_4620 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n8247), .Y(core__abc_21380_n8248) );
  AND2X2 AND2X2_4621 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core_v2_reg_51_), .Y(core__abc_21380_n8249) );
  AND2X2 AND2X2_4622 ( .A(core__abc_21380_n8253), .B(reset_n_bF_buf34), .Y(core__abc_21380_n8254) );
  AND2X2 AND2X2_4623 ( .A(core__abc_21380_n8252), .B(core__abc_21380_n8254), .Y(core_v2_reg_51__FF_INPUT) );
  AND2X2 AND2X2_4624 ( .A(core__abc_21380_n7047), .B(core__abc_21380_n7054), .Y(core__abc_21380_n8256) );
  AND2X2 AND2X2_4625 ( .A(core__abc_21380_n8257), .B(core__abc_21380_n6821), .Y(core__abc_21380_n8258) );
  AND2X2 AND2X2_4626 ( .A(core__abc_21380_n8259), .B(core__abc_21380_n8260), .Y(core__abc_21380_n8261) );
  AND2X2 AND2X2_4627 ( .A(core__abc_21380_n8261), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n8262) );
  AND2X2 AND2X2_4628 ( .A(core__abc_21380_n3313_bF_buf12), .B(core__abc_21380_n8263), .Y(core__abc_21380_n8264) );
  AND2X2 AND2X2_4629 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core_v2_reg_52_), .Y(core__abc_21380_n8265) );
  AND2X2 AND2X2_463 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_115_), .Y(_abc_19068_n1696) );
  AND2X2 AND2X2_4630 ( .A(core__abc_21380_n8269), .B(reset_n_bF_buf33), .Y(core__abc_21380_n8270) );
  AND2X2 AND2X2_4631 ( .A(core__abc_21380_n8268), .B(core__abc_21380_n8270), .Y(core_v2_reg_52__FF_INPUT) );
  AND2X2 AND2X2_4632 ( .A(core__abc_21380_n8259), .B(core__abc_21380_n6863), .Y(core__abc_21380_n8273) );
  AND2X2 AND2X2_4633 ( .A(core__abc_21380_n8274), .B(core__abc_21380_n8272), .Y(core__abc_21380_n8275) );
  AND2X2 AND2X2_4634 ( .A(core__abc_21380_n8273), .B(core__abc_21380_n6813), .Y(core__abc_21380_n8276) );
  AND2X2 AND2X2_4635 ( .A(core__abc_21380_n8277), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n8278) );
  AND2X2 AND2X2_4636 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n8279), .Y(core__abc_21380_n8280) );
  AND2X2 AND2X2_4637 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core_v2_reg_53_), .Y(core__abc_21380_n8281) );
  AND2X2 AND2X2_4638 ( .A(core__abc_21380_n8285), .B(reset_n_bF_buf32), .Y(core__abc_21380_n8286) );
  AND2X2 AND2X2_4639 ( .A(core__abc_21380_n8284), .B(core__abc_21380_n8286), .Y(core_v2_reg_53__FF_INPUT) );
  AND2X2 AND2X2_464 ( .A(_abc_19068_n1620_bF_buf2), .B(word3_reg_19_), .Y(_abc_19068_n1697) );
  AND2X2 AND2X2_4640 ( .A(core__abc_21380_n8259), .B(core__abc_21380_n6864), .Y(core__abc_21380_n8288) );
  AND2X2 AND2X2_4641 ( .A(core__abc_21380_n8289), .B(core__abc_21380_n6801), .Y(core__abc_21380_n8290) );
  AND2X2 AND2X2_4642 ( .A(core__abc_21380_n8294), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n8295) );
  AND2X2 AND2X2_4643 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n8296), .Y(core__abc_21380_n8297) );
  AND2X2 AND2X2_4644 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core_v2_reg_54_), .Y(core__abc_21380_n8298) );
  AND2X2 AND2X2_4645 ( .A(core__abc_21380_n8302), .B(reset_n_bF_buf31), .Y(core__abc_21380_n8303) );
  AND2X2 AND2X2_4646 ( .A(core__abc_21380_n8301), .B(core__abc_21380_n8303), .Y(core_v2_reg_54__FF_INPUT) );
  AND2X2 AND2X2_4647 ( .A(core__abc_21380_n8291), .B(core__abc_21380_n6869), .Y(core__abc_21380_n8306) );
  AND2X2 AND2X2_4648 ( .A(core__abc_21380_n8306), .B(core__abc_21380_n8305), .Y(core__abc_21380_n8307) );
  AND2X2 AND2X2_4649 ( .A(core__abc_21380_n8308), .B(core__abc_21380_n8309), .Y(core__abc_21380_n8310) );
  AND2X2 AND2X2_465 ( .A(_abc_19068_n1698), .B(reset_n_bF_buf65), .Y(word3_reg_19__FF_INPUT) );
  AND2X2 AND2X2_4650 ( .A(core__abc_21380_n8310), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n8311) );
  AND2X2 AND2X2_4651 ( .A(core__abc_21380_n3313_bF_buf9), .B(core_key_55_), .Y(core__abc_21380_n8312) );
  AND2X2 AND2X2_4652 ( .A(core__abc_21380_n3163_1_bF_buf1), .B(core_v2_reg_55_), .Y(core__abc_21380_n8313) );
  AND2X2 AND2X2_4653 ( .A(core__abc_21380_n8317), .B(reset_n_bF_buf30), .Y(core__abc_21380_n8318) );
  AND2X2 AND2X2_4654 ( .A(core__abc_21380_n8316), .B(core__abc_21380_n8318), .Y(core_v2_reg_55__FF_INPUT) );
  AND2X2 AND2X2_4655 ( .A(core__abc_21380_n7057), .B(core__abc_21380_n6780), .Y(core__abc_21380_n8320) );
  AND2X2 AND2X2_4656 ( .A(core__abc_21380_n8321), .B(core__abc_21380_n6779), .Y(core__abc_21380_n8322) );
  AND2X2 AND2X2_4657 ( .A(core__abc_21380_n8324), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n8325) );
  AND2X2 AND2X2_4658 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_56_), .Y(core__abc_21380_n8326) );
  AND2X2 AND2X2_4659 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core_v2_reg_56_), .Y(core__abc_21380_n8327) );
  AND2X2 AND2X2_466 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_116_), .Y(_abc_19068_n1700) );
  AND2X2 AND2X2_4660 ( .A(core__abc_21380_n8331), .B(reset_n_bF_buf29), .Y(core__abc_21380_n8332) );
  AND2X2 AND2X2_4661 ( .A(core__abc_21380_n8330), .B(core__abc_21380_n8332), .Y(core_v2_reg_56__FF_INPUT) );
  AND2X2 AND2X2_4662 ( .A(core__abc_21380_n8335), .B(core__abc_21380_n6754), .Y(core__abc_21380_n8336) );
  AND2X2 AND2X2_4663 ( .A(core__abc_21380_n8337), .B(core__abc_21380_n8334), .Y(core__abc_21380_n8338) );
  AND2X2 AND2X2_4664 ( .A(core__abc_21380_n8336), .B(core__abc_21380_n6777), .Y(core__abc_21380_n8339) );
  AND2X2 AND2X2_4665 ( .A(core__abc_21380_n8340), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n8341) );
  AND2X2 AND2X2_4666 ( .A(core__abc_21380_n3313_bF_buf7), .B(core_key_57_), .Y(core__abc_21380_n8342) );
  AND2X2 AND2X2_4667 ( .A(core__abc_21380_n3163_1_bF_buf6), .B(core_v2_reg_57_), .Y(core__abc_21380_n8343) );
  AND2X2 AND2X2_4668 ( .A(core__abc_21380_n8347), .B(reset_n_bF_buf28), .Y(core__abc_21380_n8348) );
  AND2X2 AND2X2_4669 ( .A(core__abc_21380_n8346), .B(core__abc_21380_n8348), .Y(core_v2_reg_57__FF_INPUT) );
  AND2X2 AND2X2_467 ( .A(_abc_19068_n1620_bF_buf1), .B(word3_reg_20_), .Y(_abc_19068_n1701) );
  AND2X2 AND2X2_4670 ( .A(core__abc_21380_n8335), .B(core__abc_21380_n6755), .Y(core__abc_21380_n8350) );
  AND2X2 AND2X2_4671 ( .A(core__abc_21380_n8351), .B(core__abc_21380_n6737), .Y(core__abc_21380_n8352) );
  AND2X2 AND2X2_4672 ( .A(core__abc_21380_n8356), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n8357) );
  AND2X2 AND2X2_4673 ( .A(core__abc_21380_n3313_bF_buf6), .B(core__abc_21380_n8358), .Y(core__abc_21380_n8359) );
  AND2X2 AND2X2_4674 ( .A(core__abc_21380_n3163_1_bF_buf5), .B(core_v2_reg_58_), .Y(core__abc_21380_n8360) );
  AND2X2 AND2X2_4675 ( .A(core__abc_21380_n8364), .B(reset_n_bF_buf27), .Y(core__abc_21380_n8365) );
  AND2X2 AND2X2_4676 ( .A(core__abc_21380_n8363), .B(core__abc_21380_n8365), .Y(core_v2_reg_58__FF_INPUT) );
  AND2X2 AND2X2_4677 ( .A(core__abc_21380_n8353), .B(core__abc_21380_n6759), .Y(core__abc_21380_n8368) );
  AND2X2 AND2X2_4678 ( .A(core__abc_21380_n8368), .B(core__abc_21380_n8367), .Y(core__abc_21380_n8369) );
  AND2X2 AND2X2_4679 ( .A(core__abc_21380_n8370), .B(core__abc_21380_n8371), .Y(core__abc_21380_n8372) );
  AND2X2 AND2X2_468 ( .A(_abc_19068_n1702), .B(reset_n_bF_buf64), .Y(word3_reg_20__FF_INPUT) );
  AND2X2 AND2X2_4680 ( .A(core__abc_21380_n8372), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n8373) );
  AND2X2 AND2X2_4681 ( .A(core__abc_21380_n3313_bF_buf5), .B(core__abc_21380_n8374), .Y(core__abc_21380_n8375) );
  AND2X2 AND2X2_4682 ( .A(core__abc_21380_n3163_1_bF_buf4), .B(core_v2_reg_59_), .Y(core__abc_21380_n8376) );
  AND2X2 AND2X2_4683 ( .A(core__abc_21380_n8380), .B(reset_n_bF_buf26), .Y(core__abc_21380_n8381) );
  AND2X2 AND2X2_4684 ( .A(core__abc_21380_n8379), .B(core__abc_21380_n8381), .Y(core_v2_reg_59__FF_INPUT) );
  AND2X2 AND2X2_4685 ( .A(core__abc_21380_n7057), .B(core__abc_21380_n6782), .Y(core__abc_21380_n8383) );
  AND2X2 AND2X2_4686 ( .A(core__abc_21380_n8385), .B(core__abc_21380_n6719), .Y(core__abc_21380_n8386) );
  AND2X2 AND2X2_4687 ( .A(core__abc_21380_n8384), .B(core__abc_21380_n6720), .Y(core__abc_21380_n8387) );
  AND2X2 AND2X2_4688 ( .A(core__abc_21380_n8389), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n8390) );
  AND2X2 AND2X2_4689 ( .A(core__abc_21380_n3313_bF_buf4), .B(core_key_60_), .Y(core__abc_21380_n8391) );
  AND2X2 AND2X2_469 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_117_), .Y(_abc_19068_n1704) );
  AND2X2 AND2X2_4690 ( .A(core__abc_21380_n3163_1_bF_buf3), .B(core_v2_reg_60_), .Y(core__abc_21380_n8392) );
  AND2X2 AND2X2_4691 ( .A(core__abc_21380_n8396), .B(reset_n_bF_buf25), .Y(core__abc_21380_n8397) );
  AND2X2 AND2X2_4692 ( .A(core__abc_21380_n8395), .B(core__abc_21380_n8397), .Y(core_v2_reg_60__FF_INPUT) );
  AND2X2 AND2X2_4693 ( .A(core__abc_21380_n8400), .B(core__abc_21380_n6765), .Y(core__abc_21380_n8401) );
  AND2X2 AND2X2_4694 ( .A(core__abc_21380_n8402), .B(core__abc_21380_n8399), .Y(core__abc_21380_n8403) );
  AND2X2 AND2X2_4695 ( .A(core__abc_21380_n8401), .B(core__abc_21380_n6712), .Y(core__abc_21380_n8404) );
  AND2X2 AND2X2_4696 ( .A(core__abc_21380_n8405), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf3), .Y(core__abc_21380_n8406) );
  AND2X2 AND2X2_4697 ( .A(core__abc_21380_n3313_bF_buf3), .B(core__abc_21380_n8407), .Y(core__abc_21380_n8408) );
  AND2X2 AND2X2_4698 ( .A(core__abc_21380_n3163_1_bF_buf2), .B(core_v2_reg_61_), .Y(core__abc_21380_n8409) );
  AND2X2 AND2X2_4699 ( .A(core__abc_21380_n8413), .B(reset_n_bF_buf24), .Y(core__abc_21380_n8414) );
  AND2X2 AND2X2_47 ( .A(_abc_19068_n889_1), .B(core_initalize), .Y(_abc_19068_n944) );
  AND2X2 AND2X2_470 ( .A(_abc_19068_n1620_bF_buf0), .B(word3_reg_21_), .Y(_abc_19068_n1705) );
  AND2X2 AND2X2_4700 ( .A(core__abc_21380_n8412), .B(core__abc_21380_n8414), .Y(core_v2_reg_61__FF_INPUT) );
  AND2X2 AND2X2_4701 ( .A(core__abc_21380_n8400), .B(core__abc_21380_n6766), .Y(core__abc_21380_n8416) );
  AND2X2 AND2X2_4702 ( .A(core__abc_21380_n8417), .B(core__abc_21380_n6700), .Y(core__abc_21380_n8418) );
  AND2X2 AND2X2_4703 ( .A(core__abc_21380_n8422), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf3), .Y(core__abc_21380_n8423) );
  AND2X2 AND2X2_4704 ( .A(core__abc_21380_n3313_bF_buf2), .B(core__abc_21380_n8424), .Y(core__abc_21380_n8425) );
  AND2X2 AND2X2_4705 ( .A(core__abc_21380_n3163_1_bF_buf1), .B(core_v2_reg_62_), .Y(core__abc_21380_n8426) );
  AND2X2 AND2X2_4706 ( .A(core__abc_21380_n8430), .B(reset_n_bF_buf23), .Y(core__abc_21380_n8431) );
  AND2X2 AND2X2_4707 ( .A(core__abc_21380_n8429), .B(core__abc_21380_n8431), .Y(core_v2_reg_62__FF_INPUT) );
  AND2X2 AND2X2_4708 ( .A(core__abc_21380_n8419), .B(core__abc_21380_n6771), .Y(core__abc_21380_n8434) );
  AND2X2 AND2X2_4709 ( .A(core__abc_21380_n8434), .B(core__abc_21380_n8433), .Y(core__abc_21380_n8435) );
  AND2X2 AND2X2_471 ( .A(_abc_19068_n1706), .B(reset_n_bF_buf63), .Y(word3_reg_21__FF_INPUT) );
  AND2X2 AND2X2_4710 ( .A(core__abc_21380_n8436), .B(core__abc_21380_n8437), .Y(core__abc_21380_n8438) );
  AND2X2 AND2X2_4711 ( .A(core__abc_21380_n8438), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n8439) );
  AND2X2 AND2X2_4712 ( .A(core__abc_21380_n3313_bF_buf1), .B(core_key_63_), .Y(core__abc_21380_n8440) );
  AND2X2 AND2X2_4713 ( .A(core__abc_21380_n3163_1_bF_buf0), .B(core_v2_reg_63_), .Y(core__abc_21380_n8441) );
  AND2X2 AND2X2_4714 ( .A(core__abc_21380_n8445), .B(reset_n_bF_buf22), .Y(core__abc_21380_n8446) );
  AND2X2 AND2X2_4715 ( .A(core__abc_21380_n8444), .B(core__abc_21380_n8446), .Y(core_v2_reg_63__FF_INPUT) );
  AND2X2 AND2X2_4716 ( .A(core__abc_21380_n3167_1_bF_buf12), .B(core__abc_21380_n7971), .Y(core__abc_21380_n8449) );
  AND2X2 AND2X2_4717 ( .A(core__abc_21380_n8448), .B(core__abc_21380_n8450), .Y(core__abc_21380_n8451) );
  AND2X2 AND2X2_4718 ( .A(core__abc_21380_n8453), .B(core__abc_21380_n8452), .Y(core__abc_21380_n8454) );
  AND2X2 AND2X2_4719 ( .A(core__abc_21380_n3166), .B(core__abc_21380_n3160), .Y(core__abc_21380_n8456) );
  AND2X2 AND2X2_472 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_118_), .Y(_abc_19068_n1708) );
  AND2X2 AND2X2_4720 ( .A(core__abc_21380_n8456_bF_buf7), .B(core__abc_21380_n6891), .Y(core__abc_21380_n8457) );
  AND2X2 AND2X2_4721 ( .A(core__abc_21380_n8461), .B(reset_n_bF_buf21), .Y(core__abc_21380_n8462) );
  AND2X2 AND2X2_4722 ( .A(core__abc_21380_n8460), .B(core__abc_21380_n8462), .Y(core_v1_reg_0__FF_INPUT) );
  AND2X2 AND2X2_4723 ( .A(core__abc_21380_n8466), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n8467) );
  AND2X2 AND2X2_4724 ( .A(core__abc_21380_n8467), .B(core__abc_21380_n8464), .Y(core__abc_21380_n8468) );
  AND2X2 AND2X2_4725 ( .A(core__abc_21380_n8456_bF_buf6), .B(core_v1_reg_1_), .Y(core__abc_21380_n8469) );
  AND2X2 AND2X2_4726 ( .A(core__abc_21380_n3389), .B(core_long), .Y(core__abc_21380_n8470) );
  AND2X2 AND2X2_4727 ( .A(core__abc_21380_n7079), .B(core_key_65_), .Y(core__abc_21380_n8471) );
  AND2X2 AND2X2_4728 ( .A(core__abc_21380_n3313_bF_buf12), .B(core__abc_21380_n8472), .Y(core__abc_21380_n8473) );
  AND2X2 AND2X2_4729 ( .A(core__abc_21380_n8477), .B(reset_n_bF_buf20), .Y(core__abc_21380_n8478) );
  AND2X2 AND2X2_473 ( .A(_abc_19068_n1620_bF_buf10), .B(word3_reg_22_), .Y(_abc_19068_n1709) );
  AND2X2 AND2X2_4730 ( .A(core__abc_21380_n8476), .B(core__abc_21380_n8478), .Y(core_v1_reg_1__FF_INPUT) );
  AND2X2 AND2X2_4731 ( .A(core__abc_21380_n8480), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n8481) );
  AND2X2 AND2X2_4732 ( .A(core__abc_21380_n8483), .B(core__abc_21380_n8482), .Y(core__abc_21380_n8484) );
  AND2X2 AND2X2_4733 ( .A(core__abc_21380_n8456_bF_buf5), .B(core__abc_21380_n1299), .Y(core__abc_21380_n8485) );
  AND2X2 AND2X2_4734 ( .A(core__abc_21380_n8486), .B(core__abc_21380_n8488), .Y(core__abc_21380_n8489) );
  AND2X2 AND2X2_4735 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n8489), .Y(core__abc_21380_n8490) );
  AND2X2 AND2X2_4736 ( .A(core__abc_21380_n8494), .B(reset_n_bF_buf19), .Y(core__abc_21380_n8495) );
  AND2X2 AND2X2_4737 ( .A(core__abc_21380_n8493), .B(core__abc_21380_n8495), .Y(core_v1_reg_2__FF_INPUT) );
  AND2X2 AND2X2_4738 ( .A(core__abc_21380_n8499), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n8500) );
  AND2X2 AND2X2_4739 ( .A(core__abc_21380_n8500), .B(core__abc_21380_n8497), .Y(core__abc_21380_n8501) );
  AND2X2 AND2X2_474 ( .A(_abc_19068_n1710), .B(reset_n_bF_buf62), .Y(word3_reg_22__FF_INPUT) );
  AND2X2 AND2X2_4740 ( .A(core__abc_21380_n8456_bF_buf4), .B(core__abc_21380_n1319), .Y(core__abc_21380_n8502) );
  AND2X2 AND2X2_4741 ( .A(core__abc_21380_n8503), .B(core__abc_21380_n8505), .Y(core__abc_21380_n8506) );
  AND2X2 AND2X2_4742 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n8506), .Y(core__abc_21380_n8507) );
  AND2X2 AND2X2_4743 ( .A(core__abc_21380_n8511), .B(reset_n_bF_buf18), .Y(core__abc_21380_n8512) );
  AND2X2 AND2X2_4744 ( .A(core__abc_21380_n8510), .B(core__abc_21380_n8512), .Y(core_v1_reg_3__FF_INPUT) );
  AND2X2 AND2X2_4745 ( .A(core__abc_21380_n8514), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n8515) );
  AND2X2 AND2X2_4746 ( .A(core__abc_21380_n8517), .B(core__abc_21380_n8516), .Y(core__abc_21380_n8518) );
  AND2X2 AND2X2_4747 ( .A(core__abc_21380_n8456_bF_buf3), .B(core__abc_21380_n6840), .Y(core__abc_21380_n8519) );
  AND2X2 AND2X2_4748 ( .A(core__abc_21380_n3313_bF_buf9), .B(core_key_68_), .Y(core__abc_21380_n8520) );
  AND2X2 AND2X2_4749 ( .A(core__abc_21380_n8524), .B(reset_n_bF_buf17), .Y(core__abc_21380_n8525) );
  AND2X2 AND2X2_475 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_119_), .Y(_abc_19068_n1712) );
  AND2X2 AND2X2_4750 ( .A(core__abc_21380_n8523), .B(core__abc_21380_n8525), .Y(core_v1_reg_4__FF_INPUT) );
  AND2X2 AND2X2_4751 ( .A(core__abc_21380_n8529), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n8530) );
  AND2X2 AND2X2_4752 ( .A(core__abc_21380_n8530), .B(core__abc_21380_n8527), .Y(core__abc_21380_n8531) );
  AND2X2 AND2X2_4753 ( .A(core__abc_21380_n8456_bF_buf2), .B(core_v1_reg_5_), .Y(core__abc_21380_n8532) );
  AND2X2 AND2X2_4754 ( .A(core__abc_21380_n8533), .B(core__abc_21380_n8534), .Y(core__abc_21380_n8535) );
  AND2X2 AND2X2_4755 ( .A(core__abc_21380_n3313_bF_buf8), .B(core__abc_21380_n8535), .Y(core__abc_21380_n8536) );
  AND2X2 AND2X2_4756 ( .A(core__abc_21380_n8540), .B(reset_n_bF_buf16), .Y(core__abc_21380_n8541) );
  AND2X2 AND2X2_4757 ( .A(core__abc_21380_n8539), .B(core__abc_21380_n8541), .Y(core_v1_reg_5__FF_INPUT) );
  AND2X2 AND2X2_4758 ( .A(core__abc_21380_n8543), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n8544) );
  AND2X2 AND2X2_4759 ( .A(core__abc_21380_n8546), .B(core__abc_21380_n8545), .Y(core__abc_21380_n8547) );
  AND2X2 AND2X2_476 ( .A(_abc_19068_n1620_bF_buf9), .B(word3_reg_23_), .Y(_abc_19068_n1713) );
  AND2X2 AND2X2_4760 ( .A(core__abc_21380_n8456_bF_buf1), .B(core__abc_21380_n1374), .Y(core__abc_21380_n8548) );
  AND2X2 AND2X2_4761 ( .A(core__abc_21380_n3725), .B(core__abc_21380_n7079), .Y(core__abc_21380_n8549) );
  AND2X2 AND2X2_4762 ( .A(core_key_70_), .B(core_long), .Y(core__abc_21380_n8550) );
  AND2X2 AND2X2_4763 ( .A(core__abc_21380_n3313_bF_buf7), .B(core__abc_21380_n8551), .Y(core__abc_21380_n8552) );
  AND2X2 AND2X2_4764 ( .A(core__abc_21380_n8556), .B(reset_n_bF_buf15), .Y(core__abc_21380_n8557) );
  AND2X2 AND2X2_4765 ( .A(core__abc_21380_n8555), .B(core__abc_21380_n8557), .Y(core_v1_reg_6__FF_INPUT) );
  AND2X2 AND2X2_4766 ( .A(core__abc_21380_n8561), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n8562) );
  AND2X2 AND2X2_4767 ( .A(core__abc_21380_n8562), .B(core__abc_21380_n8559), .Y(core__abc_21380_n8563) );
  AND2X2 AND2X2_4768 ( .A(core__abc_21380_n8456_bF_buf0), .B(core__abc_21380_n1393), .Y(core__abc_21380_n8564) );
  AND2X2 AND2X2_4769 ( .A(core_key_71_), .B(core_long), .Y(core__abc_21380_n8565) );
  AND2X2 AND2X2_477 ( .A(_abc_19068_n1714), .B(reset_n_bF_buf61), .Y(word3_reg_23__FF_INPUT) );
  AND2X2 AND2X2_4770 ( .A(core__abc_21380_n8566), .B(core__abc_21380_n8567), .Y(core__abc_21380_n8568) );
  AND2X2 AND2X2_4771 ( .A(core__abc_21380_n3313_bF_buf6), .B(core__abc_21380_n8568), .Y(core__abc_21380_n8569) );
  AND2X2 AND2X2_4772 ( .A(core__abc_21380_n8573), .B(reset_n_bF_buf14), .Y(core__abc_21380_n8574) );
  AND2X2 AND2X2_4773 ( .A(core__abc_21380_n8572), .B(core__abc_21380_n8574), .Y(core_v1_reg_7__FF_INPUT) );
  AND2X2 AND2X2_4774 ( .A(core__abc_21380_n8070), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n8576) );
  AND2X2 AND2X2_4775 ( .A(core__abc_21380_n8578), .B(core__abc_21380_n8577), .Y(core__abc_21380_n8579) );
  AND2X2 AND2X2_4776 ( .A(core__abc_21380_n8456_bF_buf7), .B(core_v1_reg_8_), .Y(core__abc_21380_n8580) );
  AND2X2 AND2X2_4777 ( .A(core__abc_21380_n8584), .B(reset_n_bF_buf13), .Y(core__abc_21380_n8585) );
  AND2X2 AND2X2_4778 ( .A(core__abc_21380_n8583), .B(core__abc_21380_n8585), .Y(core_v1_reg_8__FF_INPUT) );
  AND2X2 AND2X2_4779 ( .A(core__abc_21380_n8588), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n8589) );
  AND2X2 AND2X2_478 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_120_), .Y(_abc_19068_n1716) );
  AND2X2 AND2X2_4780 ( .A(core__abc_21380_n8589), .B(core__abc_21380_n8587), .Y(core__abc_21380_n8590) );
  AND2X2 AND2X2_4781 ( .A(core__abc_21380_n8456_bF_buf6), .B(core_v1_reg_9_), .Y(core__abc_21380_n8591) );
  AND2X2 AND2X2_4782 ( .A(core__abc_21380_n3313_bF_buf5), .B(core__abc_21380_n8592), .Y(core__abc_21380_n8593) );
  AND2X2 AND2X2_4783 ( .A(core__abc_21380_n8597), .B(reset_n_bF_buf12), .Y(core__abc_21380_n8598) );
  AND2X2 AND2X2_4784 ( .A(core__abc_21380_n8596), .B(core__abc_21380_n8598), .Y(core_v1_reg_9__FF_INPUT) );
  AND2X2 AND2X2_4785 ( .A(core__abc_21380_n8602), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n8603) );
  AND2X2 AND2X2_4786 ( .A(core__abc_21380_n8603), .B(core__abc_21380_n8601), .Y(core__abc_21380_n8604) );
  AND2X2 AND2X2_4787 ( .A(core__abc_21380_n8456_bF_buf5), .B(core_v1_reg_10_), .Y(core__abc_21380_n8605) );
  AND2X2 AND2X2_4788 ( .A(core__abc_21380_n8609), .B(reset_n_bF_buf11), .Y(core__abc_21380_n8610) );
  AND2X2 AND2X2_4789 ( .A(core__abc_21380_n8608), .B(core__abc_21380_n8610), .Y(core_v1_reg_10__FF_INPUT) );
  AND2X2 AND2X2_479 ( .A(_abc_19068_n1620_bF_buf8), .B(word3_reg_24_), .Y(_abc_19068_n1717) );
  AND2X2 AND2X2_4790 ( .A(core__abc_21380_n8614), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n8615) );
  AND2X2 AND2X2_4791 ( .A(core__abc_21380_n8615), .B(core__abc_21380_n8612), .Y(core__abc_21380_n8616) );
  AND2X2 AND2X2_4792 ( .A(core__abc_21380_n8456_bF_buf4), .B(core_v1_reg_11_), .Y(core__abc_21380_n8617) );
  AND2X2 AND2X2_4793 ( .A(core__abc_21380_n3313_bF_buf4), .B(core__abc_21380_n8618), .Y(core__abc_21380_n8619) );
  AND2X2 AND2X2_4794 ( .A(core__abc_21380_n8623), .B(reset_n_bF_buf10), .Y(core__abc_21380_n8624) );
  AND2X2 AND2X2_4795 ( .A(core__abc_21380_n8622), .B(core__abc_21380_n8624), .Y(core_v1_reg_11__FF_INPUT) );
  AND2X2 AND2X2_4796 ( .A(core__abc_21380_n8627), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n8628) );
  AND2X2 AND2X2_4797 ( .A(core__abc_21380_n8628), .B(core__abc_21380_n8626), .Y(core__abc_21380_n8629) );
  AND2X2 AND2X2_4798 ( .A(core__abc_21380_n8456_bF_buf3), .B(core_v1_reg_12_), .Y(core__abc_21380_n8630) );
  AND2X2 AND2X2_4799 ( .A(core__abc_21380_n8634), .B(reset_n_bF_buf9), .Y(core__abc_21380_n8635) );
  AND2X2 AND2X2_48 ( .A(_abc_19068_n912_1), .B(_abc_19068_n888_1), .Y(_abc_19068_n945_1) );
  AND2X2 AND2X2_480 ( .A(_abc_19068_n1718), .B(reset_n_bF_buf60), .Y(word3_reg_24__FF_INPUT) );
  AND2X2 AND2X2_4800 ( .A(core__abc_21380_n8633), .B(core__abc_21380_n8635), .Y(core_v1_reg_12__FF_INPUT) );
  AND2X2 AND2X2_4801 ( .A(core__abc_21380_n8638), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf2), .Y(core__abc_21380_n8639) );
  AND2X2 AND2X2_4802 ( .A(core__abc_21380_n8639), .B(core__abc_21380_n8637), .Y(core__abc_21380_n8640) );
  AND2X2 AND2X2_4803 ( .A(core__abc_21380_n8456_bF_buf2), .B(core_v1_reg_13_), .Y(core__abc_21380_n8641) );
  AND2X2 AND2X2_4804 ( .A(core__abc_21380_n8645), .B(reset_n_bF_buf8), .Y(core__abc_21380_n8646) );
  AND2X2 AND2X2_4805 ( .A(core__abc_21380_n8644), .B(core__abc_21380_n8646), .Y(core_v1_reg_13__FF_INPUT) );
  AND2X2 AND2X2_4806 ( .A(core__abc_21380_n8650), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf2), .Y(core__abc_21380_n8651) );
  AND2X2 AND2X2_4807 ( .A(core__abc_21380_n8651), .B(core__abc_21380_n8649), .Y(core__abc_21380_n8652) );
  AND2X2 AND2X2_4808 ( .A(core__abc_21380_n8456_bF_buf1), .B(core_v1_reg_14_), .Y(core__abc_21380_n8653) );
  AND2X2 AND2X2_4809 ( .A(core__abc_21380_n8657), .B(reset_n_bF_buf7), .Y(core__abc_21380_n8658) );
  AND2X2 AND2X2_481 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_121_), .Y(_abc_19068_n1720) );
  AND2X2 AND2X2_4810 ( .A(core__abc_21380_n8656), .B(core__abc_21380_n8658), .Y(core_v1_reg_14__FF_INPUT) );
  AND2X2 AND2X2_4811 ( .A(core__abc_21380_n8661), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n8662) );
  AND2X2 AND2X2_4812 ( .A(core__abc_21380_n8662), .B(core__abc_21380_n8660), .Y(core__abc_21380_n8663) );
  AND2X2 AND2X2_4813 ( .A(core__abc_21380_n8456_bF_buf0), .B(core_v1_reg_15_), .Y(core__abc_21380_n8664) );
  AND2X2 AND2X2_4814 ( .A(core__abc_21380_n8668), .B(reset_n_bF_buf6), .Y(core__abc_21380_n8669) );
  AND2X2 AND2X2_4815 ( .A(core__abc_21380_n8667), .B(core__abc_21380_n8669), .Y(core_v1_reg_15__FF_INPUT) );
  AND2X2 AND2X2_4816 ( .A(core__abc_21380_n8672), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n8673) );
  AND2X2 AND2X2_4817 ( .A(core__abc_21380_n8673), .B(core__abc_21380_n8671), .Y(core__abc_21380_n8674) );
  AND2X2 AND2X2_4818 ( .A(core__abc_21380_n8456_bF_buf7), .B(core_v1_reg_16_), .Y(core__abc_21380_n8675) );
  AND2X2 AND2X2_4819 ( .A(core__abc_21380_n8679), .B(reset_n_bF_buf5), .Y(core__abc_21380_n8680) );
  AND2X2 AND2X2_482 ( .A(_abc_19068_n1620_bF_buf7), .B(word3_reg_25_), .Y(_abc_19068_n1721) );
  AND2X2 AND2X2_4820 ( .A(core__abc_21380_n8678), .B(core__abc_21380_n8680), .Y(core_v1_reg_16__FF_INPUT) );
  AND2X2 AND2X2_4821 ( .A(core__abc_21380_n8684), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n8685) );
  AND2X2 AND2X2_4822 ( .A(core__abc_21380_n8685), .B(core__abc_21380_n8682), .Y(core__abc_21380_n8686) );
  AND2X2 AND2X2_4823 ( .A(core__abc_21380_n8456_bF_buf6), .B(core_v1_reg_17_), .Y(core__abc_21380_n8687) );
  AND2X2 AND2X2_4824 ( .A(core__abc_21380_n8691), .B(reset_n_bF_buf4), .Y(core__abc_21380_n8692) );
  AND2X2 AND2X2_4825 ( .A(core__abc_21380_n8690), .B(core__abc_21380_n8692), .Y(core_v1_reg_17__FF_INPUT) );
  AND2X2 AND2X2_4826 ( .A(core__abc_21380_n8695), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n8696) );
  AND2X2 AND2X2_4827 ( .A(core__abc_21380_n8696), .B(core__abc_21380_n8694), .Y(core__abc_21380_n8697) );
  AND2X2 AND2X2_4828 ( .A(core__abc_21380_n8456_bF_buf5), .B(core_v1_reg_18_), .Y(core__abc_21380_n8698) );
  AND2X2 AND2X2_4829 ( .A(core__abc_21380_n8702), .B(reset_n_bF_buf3), .Y(core__abc_21380_n8703) );
  AND2X2 AND2X2_483 ( .A(_abc_19068_n1722), .B(reset_n_bF_buf59), .Y(word3_reg_25__FF_INPUT) );
  AND2X2 AND2X2_4830 ( .A(core__abc_21380_n8701), .B(core__abc_21380_n8703), .Y(core_v1_reg_18__FF_INPUT) );
  AND2X2 AND2X2_4831 ( .A(core__abc_21380_n8706), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n8707) );
  AND2X2 AND2X2_4832 ( .A(core__abc_21380_n8707), .B(core__abc_21380_n8705), .Y(core__abc_21380_n8708) );
  AND2X2 AND2X2_4833 ( .A(core__abc_21380_n8456_bF_buf4), .B(core_v1_reg_19_), .Y(core__abc_21380_n8709) );
  AND2X2 AND2X2_4834 ( .A(core__abc_21380_n8713), .B(reset_n_bF_buf2), .Y(core__abc_21380_n8714) );
  AND2X2 AND2X2_4835 ( .A(core__abc_21380_n8712), .B(core__abc_21380_n8714), .Y(core_v1_reg_19__FF_INPUT) );
  AND2X2 AND2X2_4836 ( .A(core__abc_21380_n8719), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n8720) );
  AND2X2 AND2X2_4837 ( .A(core__abc_21380_n8720), .B(core__abc_21380_n8717), .Y(core__abc_21380_n8721) );
  AND2X2 AND2X2_4838 ( .A(core__abc_21380_n8456_bF_buf3), .B(core_v1_reg_20_), .Y(core__abc_21380_n8722) );
  AND2X2 AND2X2_4839 ( .A(core__abc_21380_n3313_bF_buf3), .B(core_key_84_), .Y(core__abc_21380_n8723) );
  AND2X2 AND2X2_484 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_122_), .Y(_abc_19068_n1724) );
  AND2X2 AND2X2_4840 ( .A(core__abc_21380_n8727), .B(reset_n_bF_buf1), .Y(core__abc_21380_n8728) );
  AND2X2 AND2X2_4841 ( .A(core__abc_21380_n8726), .B(core__abc_21380_n8728), .Y(core_v1_reg_20__FF_INPUT) );
  AND2X2 AND2X2_4842 ( .A(core__abc_21380_n8732), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n8733) );
  AND2X2 AND2X2_4843 ( .A(core__abc_21380_n8733), .B(core__abc_21380_n8730), .Y(core__abc_21380_n8734) );
  AND2X2 AND2X2_4844 ( .A(core__abc_21380_n8456_bF_buf2), .B(core_v1_reg_21_), .Y(core__abc_21380_n8735) );
  AND2X2 AND2X2_4845 ( .A(core__abc_21380_n8739), .B(reset_n_bF_buf0), .Y(core__abc_21380_n8740) );
  AND2X2 AND2X2_4846 ( .A(core__abc_21380_n8738), .B(core__abc_21380_n8740), .Y(core_v1_reg_21__FF_INPUT) );
  AND2X2 AND2X2_4847 ( .A(core__abc_21380_n8743), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n8744) );
  AND2X2 AND2X2_4848 ( .A(core__abc_21380_n8744), .B(core__abc_21380_n8742), .Y(core__abc_21380_n8745) );
  AND2X2 AND2X2_4849 ( .A(core__abc_21380_n8456_bF_buf1), .B(core_v1_reg_22_), .Y(core__abc_21380_n8746) );
  AND2X2 AND2X2_485 ( .A(_abc_19068_n1620_bF_buf6), .B(word3_reg_26_), .Y(_abc_19068_n1725) );
  AND2X2 AND2X2_4850 ( .A(core__abc_21380_n8750), .B(reset_n_bF_buf84), .Y(core__abc_21380_n8751) );
  AND2X2 AND2X2_4851 ( .A(core__abc_21380_n8749), .B(core__abc_21380_n8751), .Y(core_v1_reg_22__FF_INPUT) );
  AND2X2 AND2X2_4852 ( .A(core__abc_21380_n8755), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n8756) );
  AND2X2 AND2X2_4853 ( .A(core__abc_21380_n8756), .B(core__abc_21380_n8753), .Y(core__abc_21380_n8757) );
  AND2X2 AND2X2_4854 ( .A(core__abc_21380_n8456_bF_buf0), .B(core_v1_reg_23_), .Y(core__abc_21380_n8758) );
  AND2X2 AND2X2_4855 ( .A(core__abc_21380_n8762), .B(reset_n_bF_buf83), .Y(core__abc_21380_n8763) );
  AND2X2 AND2X2_4856 ( .A(core__abc_21380_n8761), .B(core__abc_21380_n8763), .Y(core_v1_reg_23__FF_INPUT) );
  AND2X2 AND2X2_4857 ( .A(core__abc_21380_n8766), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n8767) );
  AND2X2 AND2X2_4858 ( .A(core__abc_21380_n8767), .B(core__abc_21380_n8765), .Y(core__abc_21380_n8768) );
  AND2X2 AND2X2_4859 ( .A(core__abc_21380_n8456_bF_buf7), .B(core_v1_reg_24_), .Y(core__abc_21380_n8769) );
  AND2X2 AND2X2_486 ( .A(_abc_19068_n1726), .B(reset_n_bF_buf58), .Y(word3_reg_26__FF_INPUT) );
  AND2X2 AND2X2_4860 ( .A(core__abc_21380_n3313_bF_buf2), .B(core_key_88_), .Y(core__abc_21380_n8770) );
  AND2X2 AND2X2_4861 ( .A(core__abc_21380_n8774), .B(reset_n_bF_buf82), .Y(core__abc_21380_n8775) );
  AND2X2 AND2X2_4862 ( .A(core__abc_21380_n8773), .B(core__abc_21380_n8775), .Y(core_v1_reg_24__FF_INPUT) );
  AND2X2 AND2X2_4863 ( .A(core__abc_21380_n8779), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n8780) );
  AND2X2 AND2X2_4864 ( .A(core__abc_21380_n8780), .B(core__abc_21380_n8777), .Y(core__abc_21380_n8781) );
  AND2X2 AND2X2_4865 ( .A(core__abc_21380_n8456_bF_buf6), .B(core_v1_reg_25_), .Y(core__abc_21380_n8782) );
  AND2X2 AND2X2_4866 ( .A(core__abc_21380_n3313_bF_buf1), .B(core__abc_21380_n8783), .Y(core__abc_21380_n8784) );
  AND2X2 AND2X2_4867 ( .A(core__abc_21380_n8788), .B(reset_n_bF_buf81), .Y(core__abc_21380_n8789) );
  AND2X2 AND2X2_4868 ( .A(core__abc_21380_n8787), .B(core__abc_21380_n8789), .Y(core_v1_reg_25__FF_INPUT) );
  AND2X2 AND2X2_4869 ( .A(core__abc_21380_n8792), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n8793) );
  AND2X2 AND2X2_487 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_123_), .Y(_abc_19068_n1728) );
  AND2X2 AND2X2_4870 ( .A(core__abc_21380_n8793), .B(core__abc_21380_n8791), .Y(core__abc_21380_n8794) );
  AND2X2 AND2X2_4871 ( .A(core__abc_21380_n8456_bF_buf5), .B(core_v1_reg_26_), .Y(core__abc_21380_n8795) );
  AND2X2 AND2X2_4872 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n8796), .Y(core__abc_21380_n8797) );
  AND2X2 AND2X2_4873 ( .A(core__abc_21380_n8801), .B(reset_n_bF_buf80), .Y(core__abc_21380_n8802) );
  AND2X2 AND2X2_4874 ( .A(core__abc_21380_n8800), .B(core__abc_21380_n8802), .Y(core_v1_reg_26__FF_INPUT) );
  AND2X2 AND2X2_4875 ( .A(core__abc_21380_n8806), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n8807) );
  AND2X2 AND2X2_4876 ( .A(core__abc_21380_n8807), .B(core__abc_21380_n8804), .Y(core__abc_21380_n8808) );
  AND2X2 AND2X2_4877 ( .A(core__abc_21380_n8456_bF_buf4), .B(core_v1_reg_27_), .Y(core__abc_21380_n8809) );
  AND2X2 AND2X2_4878 ( .A(core__abc_21380_n8813), .B(reset_n_bF_buf79), .Y(core__abc_21380_n8814) );
  AND2X2 AND2X2_4879 ( .A(core__abc_21380_n8812), .B(core__abc_21380_n8814), .Y(core_v1_reg_27__FF_INPUT) );
  AND2X2 AND2X2_488 ( .A(_abc_19068_n1620_bF_buf5), .B(word3_reg_27_), .Y(_abc_19068_n1729) );
  AND2X2 AND2X2_4880 ( .A(core__abc_21380_n8818), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n8819) );
  AND2X2 AND2X2_4881 ( .A(core__abc_21380_n8819), .B(core__abc_21380_n8817), .Y(core__abc_21380_n8820) );
  AND2X2 AND2X2_4882 ( .A(core__abc_21380_n8456_bF_buf3), .B(core_v1_reg_28_), .Y(core__abc_21380_n8821) );
  AND2X2 AND2X2_4883 ( .A(core__abc_21380_n3313_bF_buf12), .B(core_key_92_), .Y(core__abc_21380_n8822) );
  AND2X2 AND2X2_4884 ( .A(core__abc_21380_n8826), .B(reset_n_bF_buf78), .Y(core__abc_21380_n8827) );
  AND2X2 AND2X2_4885 ( .A(core__abc_21380_n8825), .B(core__abc_21380_n8827), .Y(core_v1_reg_28__FF_INPUT) );
  AND2X2 AND2X2_4886 ( .A(core__abc_21380_n8831), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf1), .Y(core__abc_21380_n8832) );
  AND2X2 AND2X2_4887 ( .A(core__abc_21380_n8832), .B(core__abc_21380_n8829), .Y(core__abc_21380_n8833) );
  AND2X2 AND2X2_4888 ( .A(core__abc_21380_n8456_bF_buf2), .B(core_v1_reg_29_), .Y(core__abc_21380_n8834) );
  AND2X2 AND2X2_4889 ( .A(core__abc_21380_n8838), .B(reset_n_bF_buf77), .Y(core__abc_21380_n8839) );
  AND2X2 AND2X2_489 ( .A(_abc_19068_n1730), .B(reset_n_bF_buf57), .Y(word3_reg_27__FF_INPUT) );
  AND2X2 AND2X2_4890 ( .A(core__abc_21380_n8837), .B(core__abc_21380_n8839), .Y(core_v1_reg_29__FF_INPUT) );
  AND2X2 AND2X2_4891 ( .A(core__abc_21380_n8842), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf1), .Y(core__abc_21380_n8843) );
  AND2X2 AND2X2_4892 ( .A(core__abc_21380_n8843), .B(core__abc_21380_n8841), .Y(core__abc_21380_n8844) );
  AND2X2 AND2X2_4893 ( .A(core__abc_21380_n8456_bF_buf1), .B(core_v1_reg_30_), .Y(core__abc_21380_n8845) );
  AND2X2 AND2X2_4894 ( .A(core__abc_21380_n8849), .B(reset_n_bF_buf76), .Y(core__abc_21380_n8850) );
  AND2X2 AND2X2_4895 ( .A(core__abc_21380_n8848), .B(core__abc_21380_n8850), .Y(core_v1_reg_30__FF_INPUT) );
  AND2X2 AND2X2_4896 ( .A(core__abc_21380_n8854), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n8855) );
  AND2X2 AND2X2_4897 ( .A(core__abc_21380_n8855), .B(core__abc_21380_n8852), .Y(core__abc_21380_n8856) );
  AND2X2 AND2X2_4898 ( .A(core__abc_21380_n8456_bF_buf0), .B(core_v1_reg_31_), .Y(core__abc_21380_n8857) );
  AND2X2 AND2X2_4899 ( .A(core__abc_21380_n8861), .B(reset_n_bF_buf75), .Y(core__abc_21380_n8862) );
  AND2X2 AND2X2_49 ( .A(_abc_19068_n945_1_bF_buf4), .B(core_mi_0_), .Y(_abc_19068_n946_1) );
  AND2X2 AND2X2_490 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_124_), .Y(_abc_19068_n1732) );
  AND2X2 AND2X2_4900 ( .A(core__abc_21380_n8860), .B(core__abc_21380_n8862), .Y(core_v1_reg_31__FF_INPUT) );
  AND2X2 AND2X2_4901 ( .A(core__abc_21380_n8866), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n8867) );
  AND2X2 AND2X2_4902 ( .A(core__abc_21380_n8867), .B(core__abc_21380_n8864), .Y(core__abc_21380_n8868) );
  AND2X2 AND2X2_4903 ( .A(core__abc_21380_n8456_bF_buf7), .B(core_v1_reg_32_), .Y(core__abc_21380_n8869) );
  AND2X2 AND2X2_4904 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n8870), .Y(core__abc_21380_n8871) );
  AND2X2 AND2X2_4905 ( .A(core__abc_21380_n8875), .B(reset_n_bF_buf74), .Y(core__abc_21380_n8876) );
  AND2X2 AND2X2_4906 ( .A(core__abc_21380_n8874), .B(core__abc_21380_n8876), .Y(core_v1_reg_32__FF_INPUT) );
  AND2X2 AND2X2_4907 ( .A(core__abc_21380_n8879), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n8880) );
  AND2X2 AND2X2_4908 ( .A(core__abc_21380_n8880), .B(core__abc_21380_n8878), .Y(core__abc_21380_n8881) );
  AND2X2 AND2X2_4909 ( .A(core__abc_21380_n8456_bF_buf6), .B(core_v1_reg_33_), .Y(core__abc_21380_n8882) );
  AND2X2 AND2X2_491 ( .A(_abc_19068_n1620_bF_buf4), .B(word3_reg_28_), .Y(_abc_19068_n1733) );
  AND2X2 AND2X2_4910 ( .A(core__abc_21380_n3313_bF_buf10), .B(core_key_97_), .Y(core__abc_21380_n8883) );
  AND2X2 AND2X2_4911 ( .A(core__abc_21380_n8887), .B(reset_n_bF_buf73), .Y(core__abc_21380_n8888) );
  AND2X2 AND2X2_4912 ( .A(core__abc_21380_n8886), .B(core__abc_21380_n8888), .Y(core_v1_reg_33__FF_INPUT) );
  AND2X2 AND2X2_4913 ( .A(core__abc_21380_n8891), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n8892) );
  AND2X2 AND2X2_4914 ( .A(core__abc_21380_n8892), .B(core__abc_21380_n8890), .Y(core__abc_21380_n8893) );
  AND2X2 AND2X2_4915 ( .A(core__abc_21380_n8456_bF_buf5), .B(core_v1_reg_34_), .Y(core__abc_21380_n8894) );
  AND2X2 AND2X2_4916 ( .A(core__abc_21380_n8898), .B(reset_n_bF_buf72), .Y(core__abc_21380_n8899) );
  AND2X2 AND2X2_4917 ( .A(core__abc_21380_n8897), .B(core__abc_21380_n8899), .Y(core_v1_reg_34__FF_INPUT) );
  AND2X2 AND2X2_4918 ( .A(core__abc_21380_n8902), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n8903) );
  AND2X2 AND2X2_4919 ( .A(core__abc_21380_n8903), .B(core__abc_21380_n8901), .Y(core__abc_21380_n8904) );
  AND2X2 AND2X2_492 ( .A(_abc_19068_n1734), .B(reset_n_bF_buf56), .Y(word3_reg_28__FF_INPUT) );
  AND2X2 AND2X2_4920 ( .A(core__abc_21380_n8456_bF_buf4), .B(core_v1_reg_35_), .Y(core__abc_21380_n8905) );
  AND2X2 AND2X2_4921 ( .A(core__abc_21380_n8909), .B(reset_n_bF_buf71), .Y(core__abc_21380_n8910) );
  AND2X2 AND2X2_4922 ( .A(core__abc_21380_n8908), .B(core__abc_21380_n8910), .Y(core_v1_reg_35__FF_INPUT) );
  AND2X2 AND2X2_4923 ( .A(core__abc_21380_n8915), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n8916) );
  AND2X2 AND2X2_4924 ( .A(core__abc_21380_n8916), .B(core__abc_21380_n8912), .Y(core__abc_21380_n8917) );
  AND2X2 AND2X2_4925 ( .A(core__abc_21380_n8456_bF_buf3), .B(core_v1_reg_36_), .Y(core__abc_21380_n8918) );
  AND2X2 AND2X2_4926 ( .A(core__abc_21380_n8922), .B(reset_n_bF_buf70), .Y(core__abc_21380_n8923) );
  AND2X2 AND2X2_4927 ( .A(core__abc_21380_n8921), .B(core__abc_21380_n8923), .Y(core_v1_reg_36__FF_INPUT) );
  AND2X2 AND2X2_4928 ( .A(core__abc_21380_n8927), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n8928) );
  AND2X2 AND2X2_4929 ( .A(core__abc_21380_n8928), .B(core__abc_21380_n8925), .Y(core__abc_21380_n8929) );
  AND2X2 AND2X2_493 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_125_), .Y(_abc_19068_n1736) );
  AND2X2 AND2X2_4930 ( .A(core__abc_21380_n8456_bF_buf2), .B(core_v1_reg_37_), .Y(core__abc_21380_n8930) );
  AND2X2 AND2X2_4931 ( .A(core__abc_21380_n8934), .B(reset_n_bF_buf69), .Y(core__abc_21380_n8935) );
  AND2X2 AND2X2_4932 ( .A(core__abc_21380_n8933), .B(core__abc_21380_n8935), .Y(core_v1_reg_37__FF_INPUT) );
  AND2X2 AND2X2_4933 ( .A(core__abc_21380_n8938), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n8939) );
  AND2X2 AND2X2_4934 ( .A(core__abc_21380_n8939), .B(core__abc_21380_n8937), .Y(core__abc_21380_n8940) );
  AND2X2 AND2X2_4935 ( .A(core__abc_21380_n8456_bF_buf1), .B(core_v1_reg_38_), .Y(core__abc_21380_n8941) );
  AND2X2 AND2X2_4936 ( .A(core__abc_21380_n8945), .B(reset_n_bF_buf68), .Y(core__abc_21380_n8946) );
  AND2X2 AND2X2_4937 ( .A(core__abc_21380_n8944), .B(core__abc_21380_n8946), .Y(core_v1_reg_38__FF_INPUT) );
  AND2X2 AND2X2_4938 ( .A(core__abc_21380_n8950), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n8951) );
  AND2X2 AND2X2_4939 ( .A(core__abc_21380_n8951), .B(core__abc_21380_n8948), .Y(core__abc_21380_n8952) );
  AND2X2 AND2X2_494 ( .A(_abc_19068_n1620_bF_buf3), .B(word3_reg_29_), .Y(_abc_19068_n1737) );
  AND2X2 AND2X2_4940 ( .A(core__abc_21380_n8456_bF_buf0), .B(core_v1_reg_39_), .Y(core__abc_21380_n8953) );
  AND2X2 AND2X2_4941 ( .A(core__abc_21380_n8957), .B(reset_n_bF_buf67), .Y(core__abc_21380_n8958) );
  AND2X2 AND2X2_4942 ( .A(core__abc_21380_n8956), .B(core__abc_21380_n8958), .Y(core_v1_reg_39__FF_INPUT) );
  AND2X2 AND2X2_4943 ( .A(core__abc_21380_n8961), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n8962) );
  AND2X2 AND2X2_4944 ( .A(core__abc_21380_n8962), .B(core__abc_21380_n8960), .Y(core__abc_21380_n8963) );
  AND2X2 AND2X2_4945 ( .A(core__abc_21380_n8456_bF_buf7), .B(core_v1_reg_40_), .Y(core__abc_21380_n8964) );
  AND2X2 AND2X2_4946 ( .A(core__abc_21380_n8968), .B(reset_n_bF_buf66), .Y(core__abc_21380_n8969) );
  AND2X2 AND2X2_4947 ( .A(core__abc_21380_n8967), .B(core__abc_21380_n8969), .Y(core_v1_reg_40__FF_INPUT) );
  AND2X2 AND2X2_4948 ( .A(core__abc_21380_n8973), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n8974) );
  AND2X2 AND2X2_4949 ( .A(core__abc_21380_n8974), .B(core__abc_21380_n8971), .Y(core__abc_21380_n8975) );
  AND2X2 AND2X2_495 ( .A(_abc_19068_n1738), .B(reset_n_bF_buf55), .Y(word3_reg_29__FF_INPUT) );
  AND2X2 AND2X2_4950 ( .A(core__abc_21380_n8456_bF_buf6), .B(core_v1_reg_41_), .Y(core__abc_21380_n8976) );
  AND2X2 AND2X2_4951 ( .A(core__abc_21380_n3313_bF_buf9), .B(core__abc_21380_n8977), .Y(core__abc_21380_n8978) );
  AND2X2 AND2X2_4952 ( .A(core__abc_21380_n8982), .B(reset_n_bF_buf65), .Y(core__abc_21380_n8983) );
  AND2X2 AND2X2_4953 ( .A(core__abc_21380_n8981), .B(core__abc_21380_n8983), .Y(core_v1_reg_41__FF_INPUT) );
  AND2X2 AND2X2_4954 ( .A(core__abc_21380_n8986), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n8987) );
  AND2X2 AND2X2_4955 ( .A(core__abc_21380_n8987), .B(core__abc_21380_n8985), .Y(core__abc_21380_n8988) );
  AND2X2 AND2X2_4956 ( .A(core__abc_21380_n8456_bF_buf5), .B(core_v1_reg_42_), .Y(core__abc_21380_n8989) );
  AND2X2 AND2X2_4957 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_106_), .Y(core__abc_21380_n8990) );
  AND2X2 AND2X2_4958 ( .A(core__abc_21380_n8994), .B(reset_n_bF_buf64), .Y(core__abc_21380_n8995) );
  AND2X2 AND2X2_4959 ( .A(core__abc_21380_n8993), .B(core__abc_21380_n8995), .Y(core_v1_reg_42__FF_INPUT) );
  AND2X2 AND2X2_496 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_126_), .Y(_abc_19068_n1740) );
  AND2X2 AND2X2_4960 ( .A(core__abc_21380_n8998), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n8999) );
  AND2X2 AND2X2_4961 ( .A(core__abc_21380_n8999), .B(core__abc_21380_n8997), .Y(core__abc_21380_n9000) );
  AND2X2 AND2X2_4962 ( .A(core__abc_21380_n8456_bF_buf4), .B(core_v1_reg_43_), .Y(core__abc_21380_n9001) );
  AND2X2 AND2X2_4963 ( .A(core__abc_21380_n9005), .B(reset_n_bF_buf63), .Y(core__abc_21380_n9006) );
  AND2X2 AND2X2_4964 ( .A(core__abc_21380_n9004), .B(core__abc_21380_n9006), .Y(core_v1_reg_43__FF_INPUT) );
  AND2X2 AND2X2_4965 ( .A(core__abc_21380_n9011), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n9012) );
  AND2X2 AND2X2_4966 ( .A(core__abc_21380_n9012), .B(core__abc_21380_n9010), .Y(core__abc_21380_n9013) );
  AND2X2 AND2X2_4967 ( .A(core__abc_21380_n8456_bF_buf3), .B(core_v1_reg_44_), .Y(core__abc_21380_n9014) );
  AND2X2 AND2X2_4968 ( .A(core__abc_21380_n3313_bF_buf7), .B(core__abc_21380_n9015), .Y(core__abc_21380_n9016) );
  AND2X2 AND2X2_4969 ( .A(core__abc_21380_n9020), .B(reset_n_bF_buf62), .Y(core__abc_21380_n9021) );
  AND2X2 AND2X2_497 ( .A(_abc_19068_n1620_bF_buf2), .B(word3_reg_30_), .Y(_abc_19068_n1741) );
  AND2X2 AND2X2_4970 ( .A(core__abc_21380_n9019), .B(core__abc_21380_n9021), .Y(core_v1_reg_44__FF_INPUT) );
  AND2X2 AND2X2_4971 ( .A(core__abc_21380_n9024), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf0), .Y(core__abc_21380_n9025) );
  AND2X2 AND2X2_4972 ( .A(core__abc_21380_n9025), .B(core__abc_21380_n9023), .Y(core__abc_21380_n9026) );
  AND2X2 AND2X2_4973 ( .A(core__abc_21380_n8456_bF_buf2), .B(core_v1_reg_45_), .Y(core__abc_21380_n9027) );
  AND2X2 AND2X2_4974 ( .A(core__abc_21380_n9031), .B(reset_n_bF_buf61), .Y(core__abc_21380_n9032) );
  AND2X2 AND2X2_4975 ( .A(core__abc_21380_n9030), .B(core__abc_21380_n9032), .Y(core_v1_reg_45__FF_INPUT) );
  AND2X2 AND2X2_4976 ( .A(core__abc_21380_n9035), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf0), .Y(core__abc_21380_n9036) );
  AND2X2 AND2X2_4977 ( .A(core__abc_21380_n9036), .B(core__abc_21380_n9034), .Y(core__abc_21380_n9037) );
  AND2X2 AND2X2_4978 ( .A(core__abc_21380_n8456_bF_buf1), .B(core_v1_reg_46_), .Y(core__abc_21380_n9038) );
  AND2X2 AND2X2_4979 ( .A(core__abc_21380_n9042), .B(reset_n_bF_buf60), .Y(core__abc_21380_n9043) );
  AND2X2 AND2X2_498 ( .A(_abc_19068_n1742), .B(reset_n_bF_buf54), .Y(word3_reg_30__FF_INPUT) );
  AND2X2 AND2X2_4980 ( .A(core__abc_21380_n9041), .B(core__abc_21380_n9043), .Y(core_v1_reg_46__FF_INPUT) );
  AND2X2 AND2X2_4981 ( .A(core__abc_21380_n9046), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n9047) );
  AND2X2 AND2X2_4982 ( .A(core__abc_21380_n9047), .B(core__abc_21380_n9045), .Y(core__abc_21380_n9048) );
  AND2X2 AND2X2_4983 ( .A(core__abc_21380_n8456_bF_buf0), .B(core_v1_reg_47_), .Y(core__abc_21380_n9049) );
  AND2X2 AND2X2_4984 ( .A(core__abc_21380_n9053), .B(reset_n_bF_buf59), .Y(core__abc_21380_n9054) );
  AND2X2 AND2X2_4985 ( .A(core__abc_21380_n9052), .B(core__abc_21380_n9054), .Y(core_v1_reg_47__FF_INPUT) );
  AND2X2 AND2X2_4986 ( .A(core__abc_21380_n9057), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n9058) );
  AND2X2 AND2X2_4987 ( .A(core__abc_21380_n9058), .B(core__abc_21380_n9056), .Y(core__abc_21380_n9059) );
  AND2X2 AND2X2_4988 ( .A(core__abc_21380_n8456_bF_buf7), .B(core_v1_reg_48_), .Y(core__abc_21380_n9060) );
  AND2X2 AND2X2_4989 ( .A(core__abc_21380_n9064), .B(reset_n_bF_buf58), .Y(core__abc_21380_n9065) );
  AND2X2 AND2X2_499 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_127_), .Y(_abc_19068_n1744) );
  AND2X2 AND2X2_4990 ( .A(core__abc_21380_n9063), .B(core__abc_21380_n9065), .Y(core_v1_reg_48__FF_INPUT) );
  AND2X2 AND2X2_4991 ( .A(core__abc_21380_n9069), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n9070) );
  AND2X2 AND2X2_4992 ( .A(core__abc_21380_n9070), .B(core__abc_21380_n9067), .Y(core__abc_21380_n9071) );
  AND2X2 AND2X2_4993 ( .A(core__abc_21380_n8456_bF_buf6), .B(core_v1_reg_49_), .Y(core__abc_21380_n9072) );
  AND2X2 AND2X2_4994 ( .A(core__abc_21380_n3313_bF_buf6), .B(core__abc_21380_n9073), .Y(core__abc_21380_n9074) );
  AND2X2 AND2X2_4995 ( .A(core__abc_21380_n9078), .B(reset_n_bF_buf57), .Y(core__abc_21380_n9079) );
  AND2X2 AND2X2_4996 ( .A(core__abc_21380_n9077), .B(core__abc_21380_n9079), .Y(core_v1_reg_49__FF_INPUT) );
  AND2X2 AND2X2_4997 ( .A(core__abc_21380_n9082), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n9083) );
  AND2X2 AND2X2_4998 ( .A(core__abc_21380_n9083), .B(core__abc_21380_n9081), .Y(core__abc_21380_n9084) );
  AND2X2 AND2X2_4999 ( .A(core__abc_21380_n8456_bF_buf5), .B(core_v1_reg_50_), .Y(core__abc_21380_n9085) );
  AND2X2 AND2X2_5 ( .A(_abc_19068_n878), .B(_abc_19068_n879_1), .Y(_abc_19068_n880_1) );
  AND2X2 AND2X2_50 ( .A(_abc_19068_n899_bF_buf3), .B(word3_reg_0_), .Y(_abc_19068_n948_1) );
  AND2X2 AND2X2_500 ( .A(_abc_19068_n1620_bF_buf1), .B(word3_reg_31_), .Y(_abc_19068_n1745) );
  AND2X2 AND2X2_5000 ( .A(core__abc_21380_n9089), .B(reset_n_bF_buf56), .Y(core__abc_21380_n9090) );
  AND2X2 AND2X2_5001 ( .A(core__abc_21380_n9088), .B(core__abc_21380_n9090), .Y(core_v1_reg_50__FF_INPUT) );
  AND2X2 AND2X2_5002 ( .A(core__abc_21380_n9094), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n9095) );
  AND2X2 AND2X2_5003 ( .A(core__abc_21380_n9095), .B(core__abc_21380_n9092), .Y(core__abc_21380_n9096) );
  AND2X2 AND2X2_5004 ( .A(core__abc_21380_n8456_bF_buf4), .B(core_v1_reg_51_), .Y(core__abc_21380_n9097) );
  AND2X2 AND2X2_5005 ( .A(core__abc_21380_n3313_bF_buf5), .B(core__abc_21380_n9098), .Y(core__abc_21380_n9099) );
  AND2X2 AND2X2_5006 ( .A(core__abc_21380_n9103), .B(reset_n_bF_buf55), .Y(core__abc_21380_n9104) );
  AND2X2 AND2X2_5007 ( .A(core__abc_21380_n9102), .B(core__abc_21380_n9104), .Y(core_v1_reg_51__FF_INPUT) );
  AND2X2 AND2X2_5008 ( .A(core__abc_21380_n9107), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n9108) );
  AND2X2 AND2X2_5009 ( .A(core__abc_21380_n9108), .B(core__abc_21380_n9106), .Y(core__abc_21380_n9109) );
  AND2X2 AND2X2_501 ( .A(_abc_19068_n1746), .B(reset_n_bF_buf53), .Y(word3_reg_31__FF_INPUT) );
  AND2X2 AND2X2_5010 ( .A(core__abc_21380_n8456_bF_buf3), .B(core_v1_reg_52_), .Y(core__abc_21380_n9110) );
  AND2X2 AND2X2_5011 ( .A(core__abc_21380_n9114), .B(reset_n_bF_buf54), .Y(core__abc_21380_n9115) );
  AND2X2 AND2X2_5012 ( .A(core__abc_21380_n9113), .B(core__abc_21380_n9115), .Y(core_v1_reg_52__FF_INPUT) );
  AND2X2 AND2X2_5013 ( .A(core__abc_21380_n9119), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n9120) );
  AND2X2 AND2X2_5014 ( .A(core__abc_21380_n9120), .B(core__abc_21380_n9117), .Y(core__abc_21380_n9121) );
  AND2X2 AND2X2_5015 ( .A(core__abc_21380_n8456_bF_buf2), .B(core_v1_reg_53_), .Y(core__abc_21380_n9122) );
  AND2X2 AND2X2_5016 ( .A(core__abc_21380_n9126), .B(reset_n_bF_buf53), .Y(core__abc_21380_n9127) );
  AND2X2 AND2X2_5017 ( .A(core__abc_21380_n9125), .B(core__abc_21380_n9127), .Y(core_v1_reg_53__FF_INPUT) );
  AND2X2 AND2X2_5018 ( .A(core__abc_21380_n9130), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n9131) );
  AND2X2 AND2X2_5019 ( .A(core__abc_21380_n9131), .B(core__abc_21380_n9129), .Y(core__abc_21380_n9132) );
  AND2X2 AND2X2_502 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_64_), .Y(_abc_19068_n1748) );
  AND2X2 AND2X2_5020 ( .A(core__abc_21380_n8456_bF_buf1), .B(core_v1_reg_54_), .Y(core__abc_21380_n9133) );
  AND2X2 AND2X2_5021 ( .A(core__abc_21380_n9137), .B(reset_n_bF_buf52), .Y(core__abc_21380_n9138) );
  AND2X2 AND2X2_5022 ( .A(core__abc_21380_n9136), .B(core__abc_21380_n9138), .Y(core_v1_reg_54__FF_INPUT) );
  AND2X2 AND2X2_5023 ( .A(core__abc_21380_n9141), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n9142) );
  AND2X2 AND2X2_5024 ( .A(core__abc_21380_n9142), .B(core__abc_21380_n9140), .Y(core__abc_21380_n9143) );
  AND2X2 AND2X2_5025 ( .A(core__abc_21380_n8456_bF_buf0), .B(core_v1_reg_55_), .Y(core__abc_21380_n9144) );
  AND2X2 AND2X2_5026 ( .A(core__abc_21380_n9148), .B(reset_n_bF_buf51), .Y(core__abc_21380_n9149) );
  AND2X2 AND2X2_5027 ( .A(core__abc_21380_n9147), .B(core__abc_21380_n9149), .Y(core_v1_reg_55__FF_INPUT) );
  AND2X2 AND2X2_5028 ( .A(core__abc_21380_n9152), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n9153) );
  AND2X2 AND2X2_5029 ( .A(core__abc_21380_n9153), .B(core__abc_21380_n9151), .Y(core__abc_21380_n9154) );
  AND2X2 AND2X2_503 ( .A(_abc_19068_n1620_bF_buf0), .B(word2_reg_0_), .Y(_abc_19068_n1749) );
  AND2X2 AND2X2_5030 ( .A(core__abc_21380_n8456_bF_buf7), .B(core_v1_reg_56_), .Y(core__abc_21380_n9155) );
  AND2X2 AND2X2_5031 ( .A(core__abc_21380_n9159), .B(reset_n_bF_buf50), .Y(core__abc_21380_n9160) );
  AND2X2 AND2X2_5032 ( .A(core__abc_21380_n9158), .B(core__abc_21380_n9160), .Y(core_v1_reg_56__FF_INPUT) );
  AND2X2 AND2X2_5033 ( .A(core__abc_21380_n9163), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n9164) );
  AND2X2 AND2X2_5034 ( .A(core__abc_21380_n9164), .B(core__abc_21380_n9162), .Y(core__abc_21380_n9165) );
  AND2X2 AND2X2_5035 ( .A(core__abc_21380_n8456_bF_buf6), .B(core_v1_reg_57_), .Y(core__abc_21380_n9166) );
  AND2X2 AND2X2_5036 ( .A(core__abc_21380_n9170), .B(reset_n_bF_buf49), .Y(core__abc_21380_n9171) );
  AND2X2 AND2X2_5037 ( .A(core__abc_21380_n9169), .B(core__abc_21380_n9171), .Y(core_v1_reg_57__FF_INPUT) );
  AND2X2 AND2X2_5038 ( .A(core__abc_21380_n9174), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n9175) );
  AND2X2 AND2X2_5039 ( .A(core__abc_21380_n9175), .B(core__abc_21380_n9173), .Y(core__abc_21380_n9176) );
  AND2X2 AND2X2_504 ( .A(_abc_19068_n1750), .B(reset_n_bF_buf52), .Y(word2_reg_0__FF_INPUT) );
  AND2X2 AND2X2_5040 ( .A(core__abc_21380_n8456_bF_buf5), .B(core_v1_reg_58_), .Y(core__abc_21380_n9177) );
  AND2X2 AND2X2_5041 ( .A(core__abc_21380_n9181), .B(reset_n_bF_buf48), .Y(core__abc_21380_n9182) );
  AND2X2 AND2X2_5042 ( .A(core__abc_21380_n9180), .B(core__abc_21380_n9182), .Y(core_v1_reg_58__FF_INPUT) );
  AND2X2 AND2X2_5043 ( .A(core__abc_21380_n9185), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n9186) );
  AND2X2 AND2X2_5044 ( .A(core__abc_21380_n9186), .B(core__abc_21380_n9184), .Y(core__abc_21380_n9187) );
  AND2X2 AND2X2_5045 ( .A(core__abc_21380_n8456_bF_buf4), .B(core_v1_reg_59_), .Y(core__abc_21380_n9188) );
  AND2X2 AND2X2_5046 ( .A(core__abc_21380_n9192), .B(reset_n_bF_buf47), .Y(core__abc_21380_n9193) );
  AND2X2 AND2X2_5047 ( .A(core__abc_21380_n9191), .B(core__abc_21380_n9193), .Y(core_v1_reg_59__FF_INPUT) );
  AND2X2 AND2X2_5048 ( .A(core__abc_21380_n9196), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n9197) );
  AND2X2 AND2X2_5049 ( .A(core__abc_21380_n9197), .B(core__abc_21380_n9195), .Y(core__abc_21380_n9198) );
  AND2X2 AND2X2_505 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_65_), .Y(_abc_19068_n1752) );
  AND2X2 AND2X2_5050 ( .A(core__abc_21380_n8456_bF_buf3), .B(core_v1_reg_60_), .Y(core__abc_21380_n9199) );
  AND2X2 AND2X2_5051 ( .A(core__abc_21380_n3313_bF_buf4), .B(core_key_124_), .Y(core__abc_21380_n9200) );
  AND2X2 AND2X2_5052 ( .A(core__abc_21380_n9204), .B(reset_n_bF_buf46), .Y(core__abc_21380_n9205) );
  AND2X2 AND2X2_5053 ( .A(core__abc_21380_n9203), .B(core__abc_21380_n9205), .Y(core_v1_reg_60__FF_INPUT) );
  AND2X2 AND2X2_5054 ( .A(core__abc_21380_n9208), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf3), .Y(core__abc_21380_n9209) );
  AND2X2 AND2X2_5055 ( .A(core__abc_21380_n9209), .B(core__abc_21380_n9207), .Y(core__abc_21380_n9210) );
  AND2X2 AND2X2_5056 ( .A(core__abc_21380_n8456_bF_buf2), .B(core_v1_reg_61_), .Y(core__abc_21380_n9211) );
  AND2X2 AND2X2_5057 ( .A(core__abc_21380_n9215), .B(reset_n_bF_buf45), .Y(core__abc_21380_n9216) );
  AND2X2 AND2X2_5058 ( .A(core__abc_21380_n9214), .B(core__abc_21380_n9216), .Y(core_v1_reg_61__FF_INPUT) );
  AND2X2 AND2X2_5059 ( .A(core__abc_21380_n9220), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf3), .Y(core__abc_21380_n9221) );
  AND2X2 AND2X2_506 ( .A(_abc_19068_n1620_bF_buf10), .B(word2_reg_1_), .Y(_abc_19068_n1753) );
  AND2X2 AND2X2_5060 ( .A(core__abc_21380_n9221), .B(core__abc_21380_n9218), .Y(core__abc_21380_n9222) );
  AND2X2 AND2X2_5061 ( .A(core__abc_21380_n8456_bF_buf1), .B(core_v1_reg_62_), .Y(core__abc_21380_n9223) );
  AND2X2 AND2X2_5062 ( .A(core__abc_21380_n9227), .B(reset_n_bF_buf44), .Y(core__abc_21380_n9228) );
  AND2X2 AND2X2_5063 ( .A(core__abc_21380_n9226), .B(core__abc_21380_n9228), .Y(core_v1_reg_62__FF_INPUT) );
  AND2X2 AND2X2_5064 ( .A(core__abc_21380_n7957), .B(core__abc_21380_n7463), .Y(core__abc_21380_n9230) );
  AND2X2 AND2X2_5065 ( .A(core__abc_21380_n9231), .B(core__abc_21380_n7952), .Y(core__abc_21380_n9232) );
  AND2X2 AND2X2_5066 ( .A(core__abc_21380_n9233), .B(core__abc_21380_n7462), .Y(core__abc_21380_n9234) );
  AND2X2 AND2X2_5067 ( .A(core__abc_21380_n9235), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n9236) );
  AND2X2 AND2X2_5068 ( .A(core__abc_21380_n8456_bF_buf0), .B(core_v1_reg_63_), .Y(core__abc_21380_n9237) );
  AND2X2 AND2X2_5069 ( .A(core__abc_21380_n9241), .B(reset_n_bF_buf43), .Y(core__abc_21380_n9242) );
  AND2X2 AND2X2_507 ( .A(_abc_19068_n1754), .B(reset_n_bF_buf51), .Y(word2_reg_1__FF_INPUT) );
  AND2X2 AND2X2_5070 ( .A(core__abc_21380_n9240), .B(core__abc_21380_n9242), .Y(core_v1_reg_63__FF_INPUT) );
  AND2X2 AND2X2_5071 ( .A(core__abc_21380_n9244), .B(core__abc_21380_n8452), .Y(core__abc_21380_n9245) );
  AND2X2 AND2X2_5072 ( .A(core__abc_21380_n9247), .B(core__abc_21380_n3312), .Y(core__abc_21380_n9248) );
  AND2X2 AND2X2_5073 ( .A(core_v0_reg_0_), .B(core_mi_reg_0_), .Y(core__abc_21380_n9249) );
  AND2X2 AND2X2_5074 ( .A(core__abc_21380_n9250), .B(core__abc_21380_n9251), .Y(core__abc_21380_n9252) );
  AND2X2 AND2X2_5075 ( .A(core__abc_21380_n9248_bF_buf7), .B(core__abc_21380_n9252), .Y(core__abc_21380_n9253) );
  AND2X2 AND2X2_5076 ( .A(core__abc_21380_n9257), .B(reset_n_bF_buf42), .Y(core__abc_21380_n9258) );
  AND2X2 AND2X2_5077 ( .A(core__abc_21380_n9256), .B(core__abc_21380_n9258), .Y(core_v0_reg_0__FF_INPUT) );
  AND2X2 AND2X2_5078 ( .A(core__abc_21380_n3364), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n9260) );
  AND2X2 AND2X2_5079 ( .A(core__abc_21380_n9261), .B(core_v0_reg_1_), .Y(core__abc_21380_n9262) );
  AND2X2 AND2X2_508 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_66_), .Y(_abc_19068_n1756) );
  AND2X2 AND2X2_5080 ( .A(core__abc_21380_n1288_1), .B(core_mi_reg_1_), .Y(core__abc_21380_n9263) );
  AND2X2 AND2X2_5081 ( .A(core__abc_21380_n9248_bF_buf6), .B(core__abc_21380_n9264), .Y(core__abc_21380_n9265) );
  AND2X2 AND2X2_5082 ( .A(core__abc_21380_n9269), .B(reset_n_bF_buf41), .Y(core__abc_21380_n9270) );
  AND2X2 AND2X2_5083 ( .A(core__abc_21380_n9268), .B(core__abc_21380_n9270), .Y(core_v0_reg_1__FF_INPUT) );
  AND2X2 AND2X2_5084 ( .A(core__abc_21380_n3440), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n9272) );
  AND2X2 AND2X2_5085 ( .A(core__abc_21380_n3313_bF_buf3), .B(core__abc_21380_n9273), .Y(core__abc_21380_n9274) );
  AND2X2 AND2X2_5086 ( .A(core__abc_21380_n9275), .B(core_v0_reg_2_), .Y(core__abc_21380_n9276) );
  AND2X2 AND2X2_5087 ( .A(core__abc_21380_n1298), .B(core_mi_reg_2_), .Y(core__abc_21380_n9277) );
  AND2X2 AND2X2_5088 ( .A(core__abc_21380_n9248_bF_buf5), .B(core__abc_21380_n9278), .Y(core__abc_21380_n9279) );
  AND2X2 AND2X2_5089 ( .A(core__abc_21380_n9283), .B(reset_n_bF_buf40), .Y(core__abc_21380_n9284) );
  AND2X2 AND2X2_509 ( .A(_abc_19068_n1620_bF_buf9), .B(word2_reg_2_), .Y(_abc_19068_n1757) );
  AND2X2 AND2X2_5090 ( .A(core__abc_21380_n9282), .B(core__abc_21380_n9284), .Y(core_v0_reg_2__FF_INPUT) );
  AND2X2 AND2X2_5091 ( .A(core__abc_21380_n3489), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n9286) );
  AND2X2 AND2X2_5092 ( .A(core__abc_21380_n9287), .B(core_v0_reg_3_), .Y(core__abc_21380_n9288) );
  AND2X2 AND2X2_5093 ( .A(core__abc_21380_n1318), .B(core_mi_reg_3_), .Y(core__abc_21380_n9289) );
  AND2X2 AND2X2_5094 ( .A(core__abc_21380_n9248_bF_buf4), .B(core__abc_21380_n9290), .Y(core__abc_21380_n9291) );
  AND2X2 AND2X2_5095 ( .A(core__abc_21380_n9295), .B(reset_n_bF_buf39), .Y(core__abc_21380_n9296) );
  AND2X2 AND2X2_5096 ( .A(core__abc_21380_n9294), .B(core__abc_21380_n9296), .Y(core_v0_reg_3__FF_INPUT) );
  AND2X2 AND2X2_5097 ( .A(core__abc_21380_n3563), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n9298) );
  AND2X2 AND2X2_5098 ( .A(core__abc_21380_n3313_bF_buf2), .B(core__abc_21380_n9299), .Y(core__abc_21380_n9300) );
  AND2X2 AND2X2_5099 ( .A(core_v0_reg_4_), .B(core_mi_reg_4_), .Y(core__abc_21380_n9301) );
  AND2X2 AND2X2_51 ( .A(_abc_19068_n916_1_bF_buf3), .B(word1_reg_0_), .Y(_abc_19068_n949_1) );
  AND2X2 AND2X2_510 ( .A(_abc_19068_n1758), .B(reset_n_bF_buf50), .Y(word2_reg_2__FF_INPUT) );
  AND2X2 AND2X2_5100 ( .A(core__abc_21380_n9302), .B(core__abc_21380_n9303), .Y(core__abc_21380_n9304) );
  AND2X2 AND2X2_5101 ( .A(core__abc_21380_n9248_bF_buf3), .B(core__abc_21380_n9304), .Y(core__abc_21380_n9305) );
  AND2X2 AND2X2_5102 ( .A(core__abc_21380_n9309), .B(reset_n_bF_buf38), .Y(core__abc_21380_n9310) );
  AND2X2 AND2X2_5103 ( .A(core__abc_21380_n9308), .B(core__abc_21380_n9310), .Y(core_v0_reg_4__FF_INPUT) );
  AND2X2 AND2X2_5104 ( .A(core__abc_21380_n3623_1), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n9312) );
  AND2X2 AND2X2_5105 ( .A(core__abc_21380_n9313), .B(core_v0_reg_5_), .Y(core__abc_21380_n9314) );
  AND2X2 AND2X2_5106 ( .A(core__abc_21380_n1355), .B(core_mi_reg_5_), .Y(core__abc_21380_n9315) );
  AND2X2 AND2X2_5107 ( .A(core__abc_21380_n9248_bF_buf2), .B(core__abc_21380_n9316), .Y(core__abc_21380_n9317) );
  AND2X2 AND2X2_5108 ( .A(core__abc_21380_n9321), .B(reset_n_bF_buf37), .Y(core__abc_21380_n9322) );
  AND2X2 AND2X2_5109 ( .A(core__abc_21380_n9320), .B(core__abc_21380_n9322), .Y(core_v0_reg_5__FF_INPUT) );
  AND2X2 AND2X2_511 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_67_), .Y(_abc_19068_n1760) );
  AND2X2 AND2X2_5110 ( .A(core__abc_21380_n3706), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n9324) );
  AND2X2 AND2X2_5111 ( .A(core__abc_21380_n9325), .B(core_v0_reg_6_), .Y(core__abc_21380_n9326) );
  AND2X2 AND2X2_5112 ( .A(core__abc_21380_n1373), .B(core_mi_reg_6_), .Y(core__abc_21380_n9327) );
  AND2X2 AND2X2_5113 ( .A(core__abc_21380_n9248_bF_buf1), .B(core__abc_21380_n9328), .Y(core__abc_21380_n9329) );
  AND2X2 AND2X2_5114 ( .A(core__abc_21380_n9333), .B(reset_n_bF_buf36), .Y(core__abc_21380_n9334) );
  AND2X2 AND2X2_5115 ( .A(core__abc_21380_n9332), .B(core__abc_21380_n9334), .Y(core_v0_reg_6__FF_INPUT) );
  AND2X2 AND2X2_5116 ( .A(core__abc_21380_n3768), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n9336) );
  AND2X2 AND2X2_5117 ( .A(core__abc_21380_n9337), .B(core_v0_reg_7_), .Y(core__abc_21380_n9338) );
  AND2X2 AND2X2_5118 ( .A(core__abc_21380_n1392), .B(core_mi_reg_7_), .Y(core__abc_21380_n9339) );
  AND2X2 AND2X2_5119 ( .A(core__abc_21380_n9248_bF_buf0), .B(core__abc_21380_n9340), .Y(core__abc_21380_n9341) );
  AND2X2 AND2X2_512 ( .A(_abc_19068_n1620_bF_buf8), .B(word2_reg_3_), .Y(_abc_19068_n1761) );
  AND2X2 AND2X2_5120 ( .A(core__abc_21380_n9345), .B(reset_n_bF_buf35), .Y(core__abc_21380_n9346) );
  AND2X2 AND2X2_5121 ( .A(core__abc_21380_n9344), .B(core__abc_21380_n9346), .Y(core_v0_reg_7__FF_INPUT) );
  AND2X2 AND2X2_5122 ( .A(core__abc_21380_n3849), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n9348) );
  AND2X2 AND2X2_5123 ( .A(core__abc_21380_n3313_bF_buf1), .B(core__abc_21380_n9349), .Y(core__abc_21380_n9350) );
  AND2X2 AND2X2_5124 ( .A(core_v0_reg_8_), .B(core_mi_reg_8_), .Y(core__abc_21380_n9351) );
  AND2X2 AND2X2_5125 ( .A(core__abc_21380_n9352), .B(core__abc_21380_n9353), .Y(core__abc_21380_n9354) );
  AND2X2 AND2X2_5126 ( .A(core__abc_21380_n9248_bF_buf7), .B(core__abc_21380_n9354), .Y(core__abc_21380_n9355) );
  AND2X2 AND2X2_5127 ( .A(core__abc_21380_n9359), .B(reset_n_bF_buf34), .Y(core__abc_21380_n9360) );
  AND2X2 AND2X2_5128 ( .A(core__abc_21380_n9358), .B(core__abc_21380_n9360), .Y(core_v0_reg_8__FF_INPUT) );
  AND2X2 AND2X2_5129 ( .A(core__abc_21380_n3908), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n9362) );
  AND2X2 AND2X2_513 ( .A(_abc_19068_n1762), .B(reset_n_bF_buf49), .Y(word2_reg_3__FF_INPUT) );
  AND2X2 AND2X2_5130 ( .A(core__abc_21380_n3313_bF_buf0), .B(core_key_9_), .Y(core__abc_21380_n9363) );
  AND2X2 AND2X2_5131 ( .A(core__abc_21380_n9364), .B(core_v0_reg_9_), .Y(core__abc_21380_n9365) );
  AND2X2 AND2X2_5132 ( .A(core__abc_21380_n1430), .B(core_mi_reg_9_), .Y(core__abc_21380_n9366) );
  AND2X2 AND2X2_5133 ( .A(core__abc_21380_n9248_bF_buf6), .B(core__abc_21380_n9367), .Y(core__abc_21380_n9368) );
  AND2X2 AND2X2_5134 ( .A(core__abc_21380_n9372), .B(reset_n_bF_buf33), .Y(core__abc_21380_n9373) );
  AND2X2 AND2X2_5135 ( .A(core__abc_21380_n9371), .B(core__abc_21380_n9373), .Y(core_v0_reg_9__FF_INPUT) );
  AND2X2 AND2X2_5136 ( .A(core__abc_21380_n3977), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n9375) );
  AND2X2 AND2X2_5137 ( .A(core__abc_21380_n3313_bF_buf12), .B(core__abc_21380_n9376), .Y(core__abc_21380_n9377) );
  AND2X2 AND2X2_5138 ( .A(core_v0_reg_10_), .B(core_mi_reg_10_), .Y(core__abc_21380_n9378) );
  AND2X2 AND2X2_5139 ( .A(core__abc_21380_n9379), .B(core__abc_21380_n9380), .Y(core__abc_21380_n9381) );
  AND2X2 AND2X2_514 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_68_), .Y(_abc_19068_n1764) );
  AND2X2 AND2X2_5140 ( .A(core__abc_21380_n9248_bF_buf5), .B(core__abc_21380_n9381), .Y(core__abc_21380_n9382) );
  AND2X2 AND2X2_5141 ( .A(core__abc_21380_n9386), .B(reset_n_bF_buf32), .Y(core__abc_21380_n9387) );
  AND2X2 AND2X2_5142 ( .A(core__abc_21380_n9385), .B(core__abc_21380_n9387), .Y(core_v0_reg_10__FF_INPUT) );
  AND2X2 AND2X2_5143 ( .A(core__abc_21380_n4029), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n9389) );
  AND2X2 AND2X2_5144 ( .A(core__abc_21380_n9390), .B(core_v0_reg_11_), .Y(core__abc_21380_n9391) );
  AND2X2 AND2X2_5145 ( .A(core__abc_21380_n9392), .B(core_mi_reg_11_), .Y(core__abc_21380_n9393) );
  AND2X2 AND2X2_5146 ( .A(core__abc_21380_n9248_bF_buf4), .B(core__abc_21380_n9394), .Y(core__abc_21380_n9395) );
  AND2X2 AND2X2_5147 ( .A(core__abc_21380_n9399), .B(reset_n_bF_buf31), .Y(core__abc_21380_n9400) );
  AND2X2 AND2X2_5148 ( .A(core__abc_21380_n9398), .B(core__abc_21380_n9400), .Y(core_v0_reg_11__FF_INPUT) );
  AND2X2 AND2X2_5149 ( .A(core__abc_21380_n4119), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n9402) );
  AND2X2 AND2X2_515 ( .A(_abc_19068_n1620_bF_buf7), .B(word2_reg_4_), .Y(_abc_19068_n1765) );
  AND2X2 AND2X2_5150 ( .A(core__abc_21380_n3313_bF_buf11), .B(core_key_12_), .Y(core__abc_21380_n9403) );
  AND2X2 AND2X2_5151 ( .A(core__abc_21380_n9404), .B(core_v0_reg_12_), .Y(core__abc_21380_n9405) );
  AND2X2 AND2X2_5152 ( .A(core__abc_21380_n1483), .B(core_mi_reg_12_), .Y(core__abc_21380_n9406) );
  AND2X2 AND2X2_5153 ( .A(core__abc_21380_n9248_bF_buf3), .B(core__abc_21380_n9407), .Y(core__abc_21380_n9408) );
  AND2X2 AND2X2_5154 ( .A(core__abc_21380_n9412), .B(reset_n_bF_buf30), .Y(core__abc_21380_n9413) );
  AND2X2 AND2X2_5155 ( .A(core__abc_21380_n9411), .B(core__abc_21380_n9413), .Y(core_v0_reg_12__FF_INPUT) );
  AND2X2 AND2X2_5156 ( .A(core__abc_21380_n4181), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf2), .Y(core__abc_21380_n9415) );
  AND2X2 AND2X2_5157 ( .A(core__abc_21380_n9416), .B(core_v0_reg_13_), .Y(core__abc_21380_n9417) );
  AND2X2 AND2X2_5158 ( .A(core__abc_21380_n1500), .B(core_mi_reg_13_), .Y(core__abc_21380_n9418) );
  AND2X2 AND2X2_5159 ( .A(core__abc_21380_n9248_bF_buf2), .B(core__abc_21380_n9419), .Y(core__abc_21380_n9420) );
  AND2X2 AND2X2_516 ( .A(_abc_19068_n1766), .B(reset_n_bF_buf48), .Y(word2_reg_4__FF_INPUT) );
  AND2X2 AND2X2_5160 ( .A(core__abc_21380_n9424), .B(reset_n_bF_buf29), .Y(core__abc_21380_n9425) );
  AND2X2 AND2X2_5161 ( .A(core__abc_21380_n9423), .B(core__abc_21380_n9425), .Y(core_v0_reg_13__FF_INPUT) );
  AND2X2 AND2X2_5162 ( .A(core__abc_21380_n4274), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf2), .Y(core__abc_21380_n9427) );
  AND2X2 AND2X2_5163 ( .A(core__abc_21380_n9428), .B(core_v0_reg_14_), .Y(core__abc_21380_n9429) );
  AND2X2 AND2X2_5164 ( .A(core__abc_21380_n1518), .B(core_mi_reg_14_), .Y(core__abc_21380_n9430) );
  AND2X2 AND2X2_5165 ( .A(core__abc_21380_n9248_bF_buf1), .B(core__abc_21380_n9431), .Y(core__abc_21380_n9432) );
  AND2X2 AND2X2_5166 ( .A(core__abc_21380_n9436), .B(reset_n_bF_buf28), .Y(core__abc_21380_n9437) );
  AND2X2 AND2X2_5167 ( .A(core__abc_21380_n9435), .B(core__abc_21380_n9437), .Y(core_v0_reg_14__FF_INPUT) );
  AND2X2 AND2X2_5168 ( .A(core__abc_21380_n4321), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n9439) );
  AND2X2 AND2X2_5169 ( .A(core__abc_21380_n9440), .B(core_v0_reg_15_), .Y(core__abc_21380_n9441) );
  AND2X2 AND2X2_517 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_69_), .Y(_abc_19068_n1768) );
  AND2X2 AND2X2_5170 ( .A(core__abc_21380_n1536), .B(core_mi_reg_15_), .Y(core__abc_21380_n9442) );
  AND2X2 AND2X2_5171 ( .A(core__abc_21380_n9248_bF_buf0), .B(core__abc_21380_n9443), .Y(core__abc_21380_n9444) );
  AND2X2 AND2X2_5172 ( .A(core__abc_21380_n9448), .B(reset_n_bF_buf27), .Y(core__abc_21380_n9449) );
  AND2X2 AND2X2_5173 ( .A(core__abc_21380_n9447), .B(core__abc_21380_n9449), .Y(core_v0_reg_15__FF_INPUT) );
  AND2X2 AND2X2_5174 ( .A(core__abc_21380_n4428), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n9451) );
  AND2X2 AND2X2_5175 ( .A(core__abc_21380_n9452), .B(core_v0_reg_16_), .Y(core__abc_21380_n9453) );
  AND2X2 AND2X2_5176 ( .A(core__abc_21380_n1557), .B(core_mi_reg_16_), .Y(core__abc_21380_n9454) );
  AND2X2 AND2X2_5177 ( .A(core__abc_21380_n9248_bF_buf7), .B(core__abc_21380_n9455), .Y(core__abc_21380_n9456) );
  AND2X2 AND2X2_5178 ( .A(core__abc_21380_n9460), .B(reset_n_bF_buf26), .Y(core__abc_21380_n9461) );
  AND2X2 AND2X2_5179 ( .A(core__abc_21380_n9459), .B(core__abc_21380_n9461), .Y(core_v0_reg_16__FF_INPUT) );
  AND2X2 AND2X2_518 ( .A(_abc_19068_n1620_bF_buf6), .B(word2_reg_5_), .Y(_abc_19068_n1769) );
  AND2X2 AND2X2_5180 ( .A(core__abc_21380_n4481), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n9463) );
  AND2X2 AND2X2_5181 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n9464), .Y(core__abc_21380_n9465) );
  AND2X2 AND2X2_5182 ( .A(core__abc_21380_n9466), .B(core_v0_reg_17_), .Y(core__abc_21380_n9467) );
  AND2X2 AND2X2_5183 ( .A(core__abc_21380_n1576), .B(core_mi_reg_17_), .Y(core__abc_21380_n9468) );
  AND2X2 AND2X2_5184 ( .A(core__abc_21380_n9248_bF_buf6), .B(core__abc_21380_n9469), .Y(core__abc_21380_n9470) );
  AND2X2 AND2X2_5185 ( .A(core__abc_21380_n9474), .B(reset_n_bF_buf25), .Y(core__abc_21380_n9475) );
  AND2X2 AND2X2_5186 ( .A(core__abc_21380_n9473), .B(core__abc_21380_n9475), .Y(core_v0_reg_17__FF_INPUT) );
  AND2X2 AND2X2_5187 ( .A(core__abc_21380_n4557), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n9477) );
  AND2X2 AND2X2_5188 ( .A(core__abc_21380_n3313_bF_buf9), .B(core_key_18_), .Y(core__abc_21380_n9478) );
  AND2X2 AND2X2_5189 ( .A(core__abc_21380_n9479), .B(core_v0_reg_18_), .Y(core__abc_21380_n9480) );
  AND2X2 AND2X2_519 ( .A(_abc_19068_n1770), .B(reset_n_bF_buf47), .Y(word2_reg_5__FF_INPUT) );
  AND2X2 AND2X2_5190 ( .A(core__abc_21380_n9481), .B(core_mi_reg_18_), .Y(core__abc_21380_n9482) );
  AND2X2 AND2X2_5191 ( .A(core__abc_21380_n9248_bF_buf5), .B(core__abc_21380_n9483), .Y(core__abc_21380_n9484) );
  AND2X2 AND2X2_5192 ( .A(core__abc_21380_n9488), .B(reset_n_bF_buf24), .Y(core__abc_21380_n9489) );
  AND2X2 AND2X2_5193 ( .A(core__abc_21380_n9487), .B(core__abc_21380_n9489), .Y(core_v0_reg_18__FF_INPUT) );
  AND2X2 AND2X2_5194 ( .A(core__abc_21380_n9491), .B(core_v0_reg_19_), .Y(core__abc_21380_n9492) );
  AND2X2 AND2X2_5195 ( .A(core__abc_21380_n9493), .B(core_mi_reg_19_), .Y(core__abc_21380_n9494) );
  AND2X2 AND2X2_5196 ( .A(core__abc_21380_n9248_bF_buf4), .B(core__abc_21380_n9495), .Y(core__abc_21380_n9496) );
  AND2X2 AND2X2_5197 ( .A(core__abc_21380_n9500), .B(reset_n_bF_buf23), .Y(core__abc_21380_n9501) );
  AND2X2 AND2X2_5198 ( .A(core__abc_21380_n9499), .B(core__abc_21380_n9501), .Y(core_v0_reg_19__FF_INPUT) );
  AND2X2 AND2X2_5199 ( .A(core__abc_21380_n4686_1), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n9503) );
  AND2X2 AND2X2_52 ( .A(_abc_19068_n953), .B(_abc_19068_n923_bF_buf4), .Y(_auto_iopadmap_cc_313_execute_30317_0_) );
  AND2X2 AND2X2_520 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_70_), .Y(_abc_19068_n1772) );
  AND2X2 AND2X2_5200 ( .A(core__abc_21380_n3313_bF_buf8), .B(core__abc_21380_n9504), .Y(core__abc_21380_n9505) );
  AND2X2 AND2X2_5201 ( .A(core__abc_21380_n9506), .B(core_v0_reg_20_), .Y(core__abc_21380_n9507) );
  AND2X2 AND2X2_5202 ( .A(core__abc_21380_n1628), .B(core_mi_reg_20_), .Y(core__abc_21380_n9508) );
  AND2X2 AND2X2_5203 ( .A(core__abc_21380_n9248_bF_buf3), .B(core__abc_21380_n9509), .Y(core__abc_21380_n9510) );
  AND2X2 AND2X2_5204 ( .A(core__abc_21380_n9514), .B(reset_n_bF_buf22), .Y(core__abc_21380_n9515) );
  AND2X2 AND2X2_5205 ( .A(core__abc_21380_n9513), .B(core__abc_21380_n9515), .Y(core_v0_reg_20__FF_INPUT) );
  AND2X2 AND2X2_5206 ( .A(core__abc_21380_n4731), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n9517) );
  AND2X2 AND2X2_5207 ( .A(core__abc_21380_n9518), .B(core_v0_reg_21_), .Y(core__abc_21380_n9519) );
  AND2X2 AND2X2_5208 ( .A(core__abc_21380_n1646), .B(core_mi_reg_21_), .Y(core__abc_21380_n9520) );
  AND2X2 AND2X2_5209 ( .A(core__abc_21380_n9248_bF_buf2), .B(core__abc_21380_n9521), .Y(core__abc_21380_n9522) );
  AND2X2 AND2X2_521 ( .A(_abc_19068_n1620_bF_buf5), .B(word2_reg_6_), .Y(_abc_19068_n1773) );
  AND2X2 AND2X2_5210 ( .A(core__abc_21380_n9526), .B(reset_n_bF_buf21), .Y(core__abc_21380_n9527) );
  AND2X2 AND2X2_5211 ( .A(core__abc_21380_n9525), .B(core__abc_21380_n9527), .Y(core_v0_reg_21__FF_INPUT) );
  AND2X2 AND2X2_5212 ( .A(core__abc_21380_n4784), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n9529) );
  AND2X2 AND2X2_5213 ( .A(core__abc_21380_n9530), .B(core_v0_reg_22_), .Y(core__abc_21380_n9531) );
  AND2X2 AND2X2_5214 ( .A(core__abc_21380_n1664), .B(core_mi_reg_22_), .Y(core__abc_21380_n9532) );
  AND2X2 AND2X2_5215 ( .A(core__abc_21380_n9248_bF_buf1), .B(core__abc_21380_n9533), .Y(core__abc_21380_n9534) );
  AND2X2 AND2X2_5216 ( .A(core__abc_21380_n9538), .B(reset_n_bF_buf20), .Y(core__abc_21380_n9539) );
  AND2X2 AND2X2_5217 ( .A(core__abc_21380_n9537), .B(core__abc_21380_n9539), .Y(core_v0_reg_22__FF_INPUT) );
  AND2X2 AND2X2_5218 ( .A(core__abc_21380_n4832), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n9541) );
  AND2X2 AND2X2_5219 ( .A(core__abc_21380_n9542), .B(core_v0_reg_23_), .Y(core__abc_21380_n9543) );
  AND2X2 AND2X2_522 ( .A(_abc_19068_n1774), .B(reset_n_bF_buf46), .Y(word2_reg_6__FF_INPUT) );
  AND2X2 AND2X2_5220 ( .A(core__abc_21380_n1682), .B(core_mi_reg_23_), .Y(core__abc_21380_n9544) );
  AND2X2 AND2X2_5221 ( .A(core__abc_21380_n9248_bF_buf0), .B(core__abc_21380_n9545), .Y(core__abc_21380_n9546) );
  AND2X2 AND2X2_5222 ( .A(core__abc_21380_n9550), .B(reset_n_bF_buf19), .Y(core__abc_21380_n9551) );
  AND2X2 AND2X2_5223 ( .A(core__abc_21380_n9549), .B(core__abc_21380_n9551), .Y(core_v0_reg_23__FF_INPUT) );
  AND2X2 AND2X2_5224 ( .A(core__abc_21380_n4908), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n9553) );
  AND2X2 AND2X2_5225 ( .A(core__abc_21380_n9554), .B(core_v0_reg_24_), .Y(core__abc_21380_n9555) );
  AND2X2 AND2X2_5226 ( .A(core__abc_21380_n1702), .B(core_mi_reg_24_), .Y(core__abc_21380_n9556) );
  AND2X2 AND2X2_5227 ( .A(core__abc_21380_n9248_bF_buf7), .B(core__abc_21380_n9557), .Y(core__abc_21380_n9558) );
  AND2X2 AND2X2_5228 ( .A(core__abc_21380_n9562), .B(reset_n_bF_buf18), .Y(core__abc_21380_n9563) );
  AND2X2 AND2X2_5229 ( .A(core__abc_21380_n9561), .B(core__abc_21380_n9563), .Y(core_v0_reg_24__FF_INPUT) );
  AND2X2 AND2X2_523 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_71_), .Y(_abc_19068_n1776) );
  AND2X2 AND2X2_5230 ( .A(core__abc_21380_n4956), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n9565) );
  AND2X2 AND2X2_5231 ( .A(core__abc_21380_n3313_bF_buf7), .B(core_key_25_), .Y(core__abc_21380_n9566) );
  AND2X2 AND2X2_5232 ( .A(core__abc_21380_n9567), .B(core_v0_reg_25_), .Y(core__abc_21380_n9568) );
  AND2X2 AND2X2_5233 ( .A(core__abc_21380_n1720), .B(core_mi_reg_25_), .Y(core__abc_21380_n9569) );
  AND2X2 AND2X2_5234 ( .A(core__abc_21380_n9248_bF_buf6), .B(core__abc_21380_n9570), .Y(core__abc_21380_n9571) );
  AND2X2 AND2X2_5235 ( .A(core__abc_21380_n9575), .B(reset_n_bF_buf17), .Y(core__abc_21380_n9576) );
  AND2X2 AND2X2_5236 ( .A(core__abc_21380_n9574), .B(core__abc_21380_n9576), .Y(core_v0_reg_25__FF_INPUT) );
  AND2X2 AND2X2_5237 ( .A(core__abc_21380_n5006), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n9578) );
  AND2X2 AND2X2_5238 ( .A(core__abc_21380_n3313_bF_buf6), .B(core_key_26_), .Y(core__abc_21380_n9579) );
  AND2X2 AND2X2_5239 ( .A(core_v0_reg_26_), .B(core_mi_reg_26_), .Y(core__abc_21380_n9580) );
  AND2X2 AND2X2_524 ( .A(_abc_19068_n1620_bF_buf4), .B(word2_reg_7_), .Y(_abc_19068_n1777) );
  AND2X2 AND2X2_5240 ( .A(core__abc_21380_n9581), .B(core__abc_21380_n9582), .Y(core__abc_21380_n9583) );
  AND2X2 AND2X2_5241 ( .A(core__abc_21380_n9248_bF_buf5), .B(core__abc_21380_n9583), .Y(core__abc_21380_n9584) );
  AND2X2 AND2X2_5242 ( .A(core__abc_21380_n9588), .B(reset_n_bF_buf16), .Y(core__abc_21380_n9589) );
  AND2X2 AND2X2_5243 ( .A(core__abc_21380_n9587), .B(core__abc_21380_n9589), .Y(core_v0_reg_26__FF_INPUT) );
  AND2X2 AND2X2_5244 ( .A(core__abc_21380_n5054), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n9591) );
  AND2X2 AND2X2_5245 ( .A(core__abc_21380_n3313_bF_buf5), .B(core_key_27_), .Y(core__abc_21380_n9592) );
  AND2X2 AND2X2_5246 ( .A(core__abc_21380_n9593), .B(core_v0_reg_27_), .Y(core__abc_21380_n9594) );
  AND2X2 AND2X2_5247 ( .A(core__abc_21380_n1757), .B(core_mi_reg_27_), .Y(core__abc_21380_n9595) );
  AND2X2 AND2X2_5248 ( .A(core__abc_21380_n9248_bF_buf4), .B(core__abc_21380_n9596), .Y(core__abc_21380_n9597) );
  AND2X2 AND2X2_5249 ( .A(core__abc_21380_n9601), .B(reset_n_bF_buf15), .Y(core__abc_21380_n9602) );
  AND2X2 AND2X2_525 ( .A(_abc_19068_n1778), .B(reset_n_bF_buf45), .Y(word2_reg_7__FF_INPUT) );
  AND2X2 AND2X2_5250 ( .A(core__abc_21380_n9600), .B(core__abc_21380_n9602), .Y(core_v0_reg_27__FF_INPUT) );
  AND2X2 AND2X2_5251 ( .A(core__abc_21380_n5122), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n9604) );
  AND2X2 AND2X2_5252 ( .A(core__abc_21380_n3313_bF_buf4), .B(core__abc_21380_n9605), .Y(core__abc_21380_n9606) );
  AND2X2 AND2X2_5253 ( .A(core__abc_21380_n9607), .B(core_v0_reg_28_), .Y(core__abc_21380_n9608) );
  AND2X2 AND2X2_5254 ( .A(core__abc_21380_n1777), .B(core_mi_reg_28_), .Y(core__abc_21380_n9609) );
  AND2X2 AND2X2_5255 ( .A(core__abc_21380_n9248_bF_buf3), .B(core__abc_21380_n9610), .Y(core__abc_21380_n9611) );
  AND2X2 AND2X2_5256 ( .A(core__abc_21380_n9615), .B(reset_n_bF_buf14), .Y(core__abc_21380_n9616) );
  AND2X2 AND2X2_5257 ( .A(core__abc_21380_n9614), .B(core__abc_21380_n9616), .Y(core_v0_reg_28__FF_INPUT) );
  AND2X2 AND2X2_5258 ( .A(core__abc_21380_n5176), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n9618) );
  AND2X2 AND2X2_5259 ( .A(core__abc_21380_n9619), .B(core_v0_reg_29_), .Y(core__abc_21380_n9620) );
  AND2X2 AND2X2_526 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_72_), .Y(_abc_19068_n1780) );
  AND2X2 AND2X2_5260 ( .A(core__abc_21380_n1795), .B(core_mi_reg_29_), .Y(core__abc_21380_n9621) );
  AND2X2 AND2X2_5261 ( .A(core__abc_21380_n9248_bF_buf2), .B(core__abc_21380_n9622), .Y(core__abc_21380_n9623) );
  AND2X2 AND2X2_5262 ( .A(core__abc_21380_n9627), .B(reset_n_bF_buf13), .Y(core__abc_21380_n9628) );
  AND2X2 AND2X2_5263 ( .A(core__abc_21380_n9626), .B(core__abc_21380_n9628), .Y(core_v0_reg_29__FF_INPUT) );
  AND2X2 AND2X2_5264 ( .A(core__abc_21380_n5228), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf1), .Y(core__abc_21380_n9630) );
  AND2X2 AND2X2_5265 ( .A(core__abc_21380_n9631), .B(core_v0_reg_30_), .Y(core__abc_21380_n9632) );
  AND2X2 AND2X2_5266 ( .A(core__abc_21380_n1815), .B(core_mi_reg_30_), .Y(core__abc_21380_n9633) );
  AND2X2 AND2X2_5267 ( .A(core__abc_21380_n9248_bF_buf1), .B(core__abc_21380_n9634), .Y(core__abc_21380_n9635) );
  AND2X2 AND2X2_5268 ( .A(core__abc_21380_n9639), .B(reset_n_bF_buf12), .Y(core__abc_21380_n9640) );
  AND2X2 AND2X2_5269 ( .A(core__abc_21380_n9638), .B(core__abc_21380_n9640), .Y(core_v0_reg_30__FF_INPUT) );
  AND2X2 AND2X2_527 ( .A(_abc_19068_n1620_bF_buf3), .B(word2_reg_8_), .Y(_abc_19068_n1781) );
  AND2X2 AND2X2_5270 ( .A(core__abc_21380_n5281), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf1), .Y(core__abc_21380_n9642) );
  AND2X2 AND2X2_5271 ( .A(core__abc_21380_n9643), .B(core_v0_reg_31_), .Y(core__abc_21380_n9644) );
  AND2X2 AND2X2_5272 ( .A(core__abc_21380_n1833), .B(core_mi_reg_31_), .Y(core__abc_21380_n9645) );
  AND2X2 AND2X2_5273 ( .A(core__abc_21380_n9248_bF_buf0), .B(core__abc_21380_n9646), .Y(core__abc_21380_n9647) );
  AND2X2 AND2X2_5274 ( .A(core__abc_21380_n9651), .B(reset_n_bF_buf11), .Y(core__abc_21380_n9652) );
  AND2X2 AND2X2_5275 ( .A(core__abc_21380_n9650), .B(core__abc_21380_n9652), .Y(core_v0_reg_31__FF_INPUT) );
  AND2X2 AND2X2_5276 ( .A(core__abc_21380_n5358), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n9654) );
  AND2X2 AND2X2_5277 ( .A(core__abc_21380_n9655), .B(core_v0_reg_32_), .Y(core__abc_21380_n9656) );
  AND2X2 AND2X2_5278 ( .A(core__abc_21380_n1853), .B(core_mi_reg_32_), .Y(core__abc_21380_n9657) );
  AND2X2 AND2X2_5279 ( .A(core__abc_21380_n9248_bF_buf7), .B(core__abc_21380_n9658), .Y(core__abc_21380_n9659) );
  AND2X2 AND2X2_528 ( .A(_abc_19068_n1782), .B(reset_n_bF_buf44), .Y(word2_reg_8__FF_INPUT) );
  AND2X2 AND2X2_5280 ( .A(core__abc_21380_n9663), .B(reset_n_bF_buf10), .Y(core__abc_21380_n9664) );
  AND2X2 AND2X2_5281 ( .A(core__abc_21380_n9662), .B(core__abc_21380_n9664), .Y(core_v0_reg_32__FF_INPUT) );
  AND2X2 AND2X2_5282 ( .A(core__abc_21380_n5398), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n9666) );
  AND2X2 AND2X2_5283 ( .A(core__abc_21380_n9667), .B(core_v0_reg_33_), .Y(core__abc_21380_n9668) );
  AND2X2 AND2X2_5284 ( .A(core__abc_21380_n1871), .B(core_mi_reg_33_), .Y(core__abc_21380_n9669) );
  AND2X2 AND2X2_5285 ( .A(core__abc_21380_n9248_bF_buf6), .B(core__abc_21380_n9670), .Y(core__abc_21380_n9671) );
  AND2X2 AND2X2_5286 ( .A(core__abc_21380_n9675), .B(reset_n_bF_buf9), .Y(core__abc_21380_n9676) );
  AND2X2 AND2X2_5287 ( .A(core__abc_21380_n9674), .B(core__abc_21380_n9676), .Y(core_v0_reg_33__FF_INPUT) );
  AND2X2 AND2X2_5288 ( .A(core__abc_21380_n5449), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n9678) );
  AND2X2 AND2X2_5289 ( .A(core__abc_21380_n9679), .B(core_v0_reg_34_), .Y(core__abc_21380_n9680) );
  AND2X2 AND2X2_529 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_73_), .Y(_abc_19068_n1784) );
  AND2X2 AND2X2_5290 ( .A(core__abc_21380_n1889), .B(core_mi_reg_34_), .Y(core__abc_21380_n9681) );
  AND2X2 AND2X2_5291 ( .A(core__abc_21380_n9248_bF_buf5), .B(core__abc_21380_n9682), .Y(core__abc_21380_n9683) );
  AND2X2 AND2X2_5292 ( .A(core__abc_21380_n9687), .B(reset_n_bF_buf8), .Y(core__abc_21380_n9688) );
  AND2X2 AND2X2_5293 ( .A(core__abc_21380_n9686), .B(core__abc_21380_n9688), .Y(core_v0_reg_34__FF_INPUT) );
  AND2X2 AND2X2_5294 ( .A(core__abc_21380_n5491), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n9690) );
  AND2X2 AND2X2_5295 ( .A(core__abc_21380_n9691), .B(core_v0_reg_35_), .Y(core__abc_21380_n9692) );
  AND2X2 AND2X2_5296 ( .A(core__abc_21380_n1907), .B(core_mi_reg_35_), .Y(core__abc_21380_n9693) );
  AND2X2 AND2X2_5297 ( .A(core__abc_21380_n9248_bF_buf4), .B(core__abc_21380_n9694), .Y(core__abc_21380_n9695) );
  AND2X2 AND2X2_5298 ( .A(core__abc_21380_n9699), .B(reset_n_bF_buf7), .Y(core__abc_21380_n9700) );
  AND2X2 AND2X2_5299 ( .A(core__abc_21380_n9698), .B(core__abc_21380_n9700), .Y(core_v0_reg_35__FF_INPUT) );
  AND2X2 AND2X2_53 ( .A(_abc_19068_n924_1_bF_buf3), .B(core_key_33_), .Y(_abc_19068_n955_1) );
  AND2X2 AND2X2_530 ( .A(_abc_19068_n1620_bF_buf2), .B(word2_reg_9_), .Y(_abc_19068_n1785) );
  AND2X2 AND2X2_5300 ( .A(core__abc_21380_n5545), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n9702) );
  AND2X2 AND2X2_5301 ( .A(core__abc_21380_n9703), .B(core_v0_reg_36_), .Y(core__abc_21380_n9704) );
  AND2X2 AND2X2_5302 ( .A(core__abc_21380_n1928_1), .B(core_mi_reg_36_), .Y(core__abc_21380_n9705) );
  AND2X2 AND2X2_5303 ( .A(core__abc_21380_n9248_bF_buf3), .B(core__abc_21380_n9706), .Y(core__abc_21380_n9707) );
  AND2X2 AND2X2_5304 ( .A(core__abc_21380_n9711), .B(reset_n_bF_buf6), .Y(core__abc_21380_n9712) );
  AND2X2 AND2X2_5305 ( .A(core__abc_21380_n9710), .B(core__abc_21380_n9712), .Y(core_v0_reg_36__FF_INPUT) );
  AND2X2 AND2X2_5306 ( .A(core__abc_21380_n5587), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n9714) );
  AND2X2 AND2X2_5307 ( .A(core__abc_21380_n9715), .B(core_v0_reg_37_), .Y(core__abc_21380_n9716) );
  AND2X2 AND2X2_5308 ( .A(core__abc_21380_n1947), .B(core_mi_reg_37_), .Y(core__abc_21380_n9717) );
  AND2X2 AND2X2_5309 ( .A(core__abc_21380_n9248_bF_buf2), .B(core__abc_21380_n9718), .Y(core__abc_21380_n9719) );
  AND2X2 AND2X2_531 ( .A(_abc_19068_n1786), .B(reset_n_bF_buf43), .Y(word2_reg_9__FF_INPUT) );
  AND2X2 AND2X2_5310 ( .A(core__abc_21380_n9723), .B(reset_n_bF_buf5), .Y(core__abc_21380_n9724) );
  AND2X2 AND2X2_5311 ( .A(core__abc_21380_n9722), .B(core__abc_21380_n9724), .Y(core_v0_reg_37__FF_INPUT) );
  AND2X2 AND2X2_5312 ( .A(core__abc_21380_n5639), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n9726) );
  AND2X2 AND2X2_5313 ( .A(core__abc_21380_n9727), .B(core_v0_reg_38_), .Y(core__abc_21380_n9728) );
  AND2X2 AND2X2_5314 ( .A(core__abc_21380_n1965_1), .B(core_mi_reg_38_), .Y(core__abc_21380_n9729) );
  AND2X2 AND2X2_5315 ( .A(core__abc_21380_n9248_bF_buf1), .B(core__abc_21380_n9730), .Y(core__abc_21380_n9731) );
  AND2X2 AND2X2_5316 ( .A(core__abc_21380_n9735), .B(reset_n_bF_buf4), .Y(core__abc_21380_n9736) );
  AND2X2 AND2X2_5317 ( .A(core__abc_21380_n9734), .B(core__abc_21380_n9736), .Y(core_v0_reg_38__FF_INPUT) );
  AND2X2 AND2X2_5318 ( .A(core__abc_21380_n5685), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n9738) );
  AND2X2 AND2X2_5319 ( .A(core__abc_21380_n9739), .B(core_v0_reg_39_), .Y(core__abc_21380_n9740) );
  AND2X2 AND2X2_532 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_74_), .Y(_abc_19068_n1788) );
  AND2X2 AND2X2_5320 ( .A(core__abc_21380_n1983), .B(core_mi_reg_39_), .Y(core__abc_21380_n9741) );
  AND2X2 AND2X2_5321 ( .A(core__abc_21380_n9248_bF_buf0), .B(core__abc_21380_n9742), .Y(core__abc_21380_n9743) );
  AND2X2 AND2X2_5322 ( .A(core__abc_21380_n9747), .B(reset_n_bF_buf3), .Y(core__abc_21380_n9748) );
  AND2X2 AND2X2_5323 ( .A(core__abc_21380_n9746), .B(core__abc_21380_n9748), .Y(core_v0_reg_39__FF_INPUT) );
  AND2X2 AND2X2_5324 ( .A(core__abc_21380_n5735), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n9750) );
  AND2X2 AND2X2_5325 ( .A(core__abc_21380_n9751), .B(core_v0_reg_40_), .Y(core__abc_21380_n9752) );
  AND2X2 AND2X2_5326 ( .A(core__abc_21380_n2004), .B(core_mi_reg_40_), .Y(core__abc_21380_n9753) );
  AND2X2 AND2X2_5327 ( .A(core__abc_21380_n9248_bF_buf7), .B(core__abc_21380_n9754), .Y(core__abc_21380_n9755) );
  AND2X2 AND2X2_5328 ( .A(core__abc_21380_n9759), .B(reset_n_bF_buf2), .Y(core__abc_21380_n9760) );
  AND2X2 AND2X2_5329 ( .A(core__abc_21380_n9758), .B(core__abc_21380_n9760), .Y(core_v0_reg_40__FF_INPUT) );
  AND2X2 AND2X2_533 ( .A(_abc_19068_n1620_bF_buf1), .B(word2_reg_10_), .Y(_abc_19068_n1789) );
  AND2X2 AND2X2_5330 ( .A(core__abc_21380_n5782), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n9762) );
  AND2X2 AND2X2_5331 ( .A(core__abc_21380_n3313_bF_buf3), .B(core_key_41_), .Y(core__abc_21380_n9763) );
  AND2X2 AND2X2_5332 ( .A(core__abc_21380_n9764), .B(core_v0_reg_41_), .Y(core__abc_21380_n9765) );
  AND2X2 AND2X2_5333 ( .A(core__abc_21380_n2022), .B(core_mi_reg_41_), .Y(core__abc_21380_n9766) );
  AND2X2 AND2X2_5334 ( .A(core__abc_21380_n9248_bF_buf6), .B(core__abc_21380_n9767), .Y(core__abc_21380_n9768) );
  AND2X2 AND2X2_5335 ( .A(core__abc_21380_n9772), .B(reset_n_bF_buf1), .Y(core__abc_21380_n9773) );
  AND2X2 AND2X2_5336 ( .A(core__abc_21380_n9771), .B(core__abc_21380_n9773), .Y(core_v0_reg_41__FF_INPUT) );
  AND2X2 AND2X2_5337 ( .A(core__abc_21380_n5825), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n9775) );
  AND2X2 AND2X2_5338 ( .A(core__abc_21380_n9776), .B(core_v0_reg_42_), .Y(core__abc_21380_n9777) );
  AND2X2 AND2X2_5339 ( .A(core__abc_21380_n2039_1), .B(core_mi_reg_42_), .Y(core__abc_21380_n9778) );
  AND2X2 AND2X2_534 ( .A(_abc_19068_n1790), .B(reset_n_bF_buf42), .Y(word2_reg_10__FF_INPUT) );
  AND2X2 AND2X2_5340 ( .A(core__abc_21380_n9248_bF_buf5), .B(core__abc_21380_n9779), .Y(core__abc_21380_n9780) );
  AND2X2 AND2X2_5341 ( .A(core__abc_21380_n9784), .B(reset_n_bF_buf0), .Y(core__abc_21380_n9785) );
  AND2X2 AND2X2_5342 ( .A(core__abc_21380_n9783), .B(core__abc_21380_n9785), .Y(core_v0_reg_42__FF_INPUT) );
  AND2X2 AND2X2_5343 ( .A(core__abc_21380_n5858), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n9787) );
  AND2X2 AND2X2_5344 ( .A(core__abc_21380_n3313_bF_buf2), .B(core__abc_21380_n9788), .Y(core__abc_21380_n9789) );
  AND2X2 AND2X2_5345 ( .A(core__abc_21380_n9790), .B(core_v0_reg_43_), .Y(core__abc_21380_n9791) );
  AND2X2 AND2X2_5346 ( .A(core__abc_21380_n2057), .B(core_mi_reg_43_), .Y(core__abc_21380_n9792) );
  AND2X2 AND2X2_5347 ( .A(core__abc_21380_n9248_bF_buf4), .B(core__abc_21380_n9793), .Y(core__abc_21380_n9794) );
  AND2X2 AND2X2_5348 ( .A(core__abc_21380_n9798), .B(reset_n_bF_buf84), .Y(core__abc_21380_n9799) );
  AND2X2 AND2X2_5349 ( .A(core__abc_21380_n9797), .B(core__abc_21380_n9799), .Y(core_v0_reg_43__FF_INPUT) );
  AND2X2 AND2X2_535 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_75_), .Y(_abc_19068_n1792) );
  AND2X2 AND2X2_5350 ( .A(core__abc_21380_n5905), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n9801) );
  AND2X2 AND2X2_5351 ( .A(core__abc_21380_n9802), .B(core_v0_reg_44_), .Y(core__abc_21380_n9803) );
  AND2X2 AND2X2_5352 ( .A(core__abc_21380_n2078), .B(core_mi_reg_44_), .Y(core__abc_21380_n9804) );
  AND2X2 AND2X2_5353 ( .A(core__abc_21380_n9248_bF_buf3), .B(core__abc_21380_n9805), .Y(core__abc_21380_n9806) );
  AND2X2 AND2X2_5354 ( .A(core__abc_21380_n9810), .B(reset_n_bF_buf83), .Y(core__abc_21380_n9811) );
  AND2X2 AND2X2_5355 ( .A(core__abc_21380_n9809), .B(core__abc_21380_n9811), .Y(core_v0_reg_44__FF_INPUT) );
  AND2X2 AND2X2_5356 ( .A(core__abc_21380_n5938), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n9813) );
  AND2X2 AND2X2_5357 ( .A(core__abc_21380_n9814), .B(core_v0_reg_45_), .Y(core__abc_21380_n9815) );
  AND2X2 AND2X2_5358 ( .A(core__abc_21380_n2095), .B(core_mi_reg_45_), .Y(core__abc_21380_n9816) );
  AND2X2 AND2X2_5359 ( .A(core__abc_21380_n9248_bF_buf2), .B(core__abc_21380_n9817), .Y(core__abc_21380_n9818) );
  AND2X2 AND2X2_536 ( .A(_abc_19068_n1620_bF_buf0), .B(word2_reg_11_), .Y(_abc_19068_n1793) );
  AND2X2 AND2X2_5360 ( .A(core__abc_21380_n9822), .B(reset_n_bF_buf82), .Y(core__abc_21380_n9823) );
  AND2X2 AND2X2_5361 ( .A(core__abc_21380_n9821), .B(core__abc_21380_n9823), .Y(core_v0_reg_45__FF_INPUT) );
  AND2X2 AND2X2_5362 ( .A(core__abc_21380_n5979), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf0), .Y(core__abc_21380_n9825) );
  AND2X2 AND2X2_5363 ( .A(core__abc_21380_n9826), .B(core_v0_reg_46_), .Y(core__abc_21380_n9827) );
  AND2X2 AND2X2_5364 ( .A(core__abc_21380_n2116), .B(core_mi_reg_46_), .Y(core__abc_21380_n9828) );
  AND2X2 AND2X2_5365 ( .A(core__abc_21380_n9248_bF_buf1), .B(core__abc_21380_n9829), .Y(core__abc_21380_n9830) );
  AND2X2 AND2X2_5366 ( .A(core__abc_21380_n9834), .B(reset_n_bF_buf81), .Y(core__abc_21380_n9835) );
  AND2X2 AND2X2_5367 ( .A(core__abc_21380_n9833), .B(core__abc_21380_n9835), .Y(core_v0_reg_46__FF_INPUT) );
  AND2X2 AND2X2_5368 ( .A(core__abc_21380_n6013), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf0), .Y(core__abc_21380_n9837) );
  AND2X2 AND2X2_5369 ( .A(core__abc_21380_n9838), .B(core_v0_reg_47_), .Y(core__abc_21380_n9839) );
  AND2X2 AND2X2_537 ( .A(_abc_19068_n1794), .B(reset_n_bF_buf41), .Y(word2_reg_11__FF_INPUT) );
  AND2X2 AND2X2_5370 ( .A(core__abc_21380_n2135), .B(core_mi_reg_47_), .Y(core__abc_21380_n9840) );
  AND2X2 AND2X2_5371 ( .A(core__abc_21380_n9248_bF_buf0), .B(core__abc_21380_n9841), .Y(core__abc_21380_n9842) );
  AND2X2 AND2X2_5372 ( .A(core__abc_21380_n9846), .B(reset_n_bF_buf80), .Y(core__abc_21380_n9847) );
  AND2X2 AND2X2_5373 ( .A(core__abc_21380_n9845), .B(core__abc_21380_n9847), .Y(core_v0_reg_47__FF_INPUT) );
  AND2X2 AND2X2_5374 ( .A(core__abc_21380_n6076), .B(core__abc_21380_n3167_1_bF_buf13), .Y(core__abc_21380_n9849) );
  AND2X2 AND2X2_5375 ( .A(core__abc_21380_n9850), .B(core_v0_reg_48_), .Y(core__abc_21380_n9851) );
  AND2X2 AND2X2_5376 ( .A(core__abc_21380_n2153), .B(core_mi_reg_48_), .Y(core__abc_21380_n9852) );
  AND2X2 AND2X2_5377 ( .A(core__abc_21380_n9248_bF_buf7), .B(core__abc_21380_n9853), .Y(core__abc_21380_n9854) );
  AND2X2 AND2X2_5378 ( .A(core__abc_21380_n9858), .B(reset_n_bF_buf79), .Y(core__abc_21380_n9859) );
  AND2X2 AND2X2_5379 ( .A(core__abc_21380_n9857), .B(core__abc_21380_n9859), .Y(core_v0_reg_48__FF_INPUT) );
  AND2X2 AND2X2_538 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_76_), .Y(_abc_19068_n1796) );
  AND2X2 AND2X2_5380 ( .A(core__abc_21380_n6112), .B(core__abc_21380_n3167_1_bF_buf12), .Y(core__abc_21380_n9861) );
  AND2X2 AND2X2_5381 ( .A(core__abc_21380_n3313_bF_buf1), .B(core__abc_21380_n9862), .Y(core__abc_21380_n9863) );
  AND2X2 AND2X2_5382 ( .A(core__abc_21380_n9864), .B(core_v0_reg_49_), .Y(core__abc_21380_n9865) );
  AND2X2 AND2X2_5383 ( .A(core__abc_21380_n2172), .B(core_mi_reg_49_), .Y(core__abc_21380_n9866) );
  AND2X2 AND2X2_5384 ( .A(core__abc_21380_n9248_bF_buf6), .B(core__abc_21380_n9867), .Y(core__abc_21380_n9868) );
  AND2X2 AND2X2_5385 ( .A(core__abc_21380_n9872), .B(reset_n_bF_buf78), .Y(core__abc_21380_n9873) );
  AND2X2 AND2X2_5386 ( .A(core__abc_21380_n9871), .B(core__abc_21380_n9873), .Y(core_v0_reg_49__FF_INPUT) );
  AND2X2 AND2X2_5387 ( .A(core__abc_21380_n6152), .B(core__abc_21380_n3167_1_bF_buf11), .Y(core__abc_21380_n9875) );
  AND2X2 AND2X2_5388 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n9876), .Y(core__abc_21380_n9877) );
  AND2X2 AND2X2_5389 ( .A(core__abc_21380_n9878), .B(core_v0_reg_50_), .Y(core__abc_21380_n9879) );
  AND2X2 AND2X2_539 ( .A(_abc_19068_n1620_bF_buf10), .B(word2_reg_12_), .Y(_abc_19068_n1797) );
  AND2X2 AND2X2_5390 ( .A(core__abc_21380_n2190), .B(core_mi_reg_50_), .Y(core__abc_21380_n9880) );
  AND2X2 AND2X2_5391 ( .A(core__abc_21380_n9248_bF_buf5), .B(core__abc_21380_n9881), .Y(core__abc_21380_n9882) );
  AND2X2 AND2X2_5392 ( .A(core__abc_21380_n9886), .B(reset_n_bF_buf77), .Y(core__abc_21380_n9887) );
  AND2X2 AND2X2_5393 ( .A(core__abc_21380_n9885), .B(core__abc_21380_n9887), .Y(core_v0_reg_50__FF_INPUT) );
  AND2X2 AND2X2_5394 ( .A(core__abc_21380_n6185), .B(core__abc_21380_n3167_1_bF_buf10), .Y(core__abc_21380_n9889) );
  AND2X2 AND2X2_5395 ( .A(core__abc_21380_n9890), .B(core_v0_reg_51_), .Y(core__abc_21380_n9891) );
  AND2X2 AND2X2_5396 ( .A(core__abc_21380_n2209), .B(core_mi_reg_51_), .Y(core__abc_21380_n9892) );
  AND2X2 AND2X2_5397 ( .A(core__abc_21380_n9248_bF_buf4), .B(core__abc_21380_n9893), .Y(core__abc_21380_n9894) );
  AND2X2 AND2X2_5398 ( .A(core__abc_21380_n9898), .B(reset_n_bF_buf76), .Y(core__abc_21380_n9899) );
  AND2X2 AND2X2_5399 ( .A(core__abc_21380_n9897), .B(core__abc_21380_n9899), .Y(core_v0_reg_51__FF_INPUT) );
  AND2X2 AND2X2_54 ( .A(_abc_19068_n926_bF_buf3), .B(core_key_1_), .Y(_abc_19068_n956) );
  AND2X2 AND2X2_540 ( .A(_abc_19068_n1798), .B(reset_n_bF_buf40), .Y(word2_reg_12__FF_INPUT) );
  AND2X2 AND2X2_5400 ( .A(core__abc_21380_n6227), .B(core__abc_21380_n3167_1_bF_buf9), .Y(core__abc_21380_n9901) );
  AND2X2 AND2X2_5401 ( .A(core__abc_21380_n3313_bF_buf12), .B(core_key_52_), .Y(core__abc_21380_n9902) );
  AND2X2 AND2X2_5402 ( .A(core_v0_reg_52_), .B(core_mi_reg_52_), .Y(core__abc_21380_n9903) );
  AND2X2 AND2X2_5403 ( .A(core__abc_21380_n9904), .B(core__abc_21380_n9905), .Y(core__abc_21380_n9906) );
  AND2X2 AND2X2_5404 ( .A(core__abc_21380_n9248_bF_buf3), .B(core__abc_21380_n9906), .Y(core__abc_21380_n9907) );
  AND2X2 AND2X2_5405 ( .A(core__abc_21380_n9911), .B(reset_n_bF_buf75), .Y(core__abc_21380_n9912) );
  AND2X2 AND2X2_5406 ( .A(core__abc_21380_n9910), .B(core__abc_21380_n9912), .Y(core_v0_reg_52__FF_INPUT) );
  AND2X2 AND2X2_5407 ( .A(core__abc_21380_n6257), .B(core__abc_21380_n3167_1_bF_buf8), .Y(core__abc_21380_n9914) );
  AND2X2 AND2X2_5408 ( .A(core__abc_21380_n9915), .B(core_v0_reg_53_), .Y(core__abc_21380_n9916) );
  AND2X2 AND2X2_5409 ( .A(core__abc_21380_n2246), .B(core_mi_reg_53_), .Y(core__abc_21380_n9917) );
  AND2X2 AND2X2_541 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_77_), .Y(_abc_19068_n1800) );
  AND2X2 AND2X2_5410 ( .A(core__abc_21380_n9248_bF_buf2), .B(core__abc_21380_n9918), .Y(core__abc_21380_n9919) );
  AND2X2 AND2X2_5411 ( .A(core__abc_21380_n9923), .B(reset_n_bF_buf74), .Y(core__abc_21380_n9924) );
  AND2X2 AND2X2_5412 ( .A(core__abc_21380_n9922), .B(core__abc_21380_n9924), .Y(core_v0_reg_53__FF_INPUT) );
  AND2X2 AND2X2_5413 ( .A(core__abc_21380_n6301), .B(core__abc_21380_n3167_1_bF_buf7), .Y(core__abc_21380_n9926) );
  AND2X2 AND2X2_5414 ( .A(core__abc_21380_n9927), .B(core_v0_reg_54_), .Y(core__abc_21380_n9928) );
  AND2X2 AND2X2_5415 ( .A(core__abc_21380_n2264), .B(core_mi_reg_54_), .Y(core__abc_21380_n9929) );
  AND2X2 AND2X2_5416 ( .A(core__abc_21380_n9248_bF_buf1), .B(core__abc_21380_n9930), .Y(core__abc_21380_n9931) );
  AND2X2 AND2X2_5417 ( .A(core__abc_21380_n9935), .B(reset_n_bF_buf73), .Y(core__abc_21380_n9936) );
  AND2X2 AND2X2_5418 ( .A(core__abc_21380_n9934), .B(core__abc_21380_n9936), .Y(core_v0_reg_54__FF_INPUT) );
  AND2X2 AND2X2_5419 ( .A(core__abc_21380_n6335), .B(core__abc_21380_n3167_1_bF_buf6), .Y(core__abc_21380_n9938) );
  AND2X2 AND2X2_542 ( .A(_abc_19068_n1620_bF_buf9), .B(word2_reg_13_), .Y(_abc_19068_n1801) );
  AND2X2 AND2X2_5420 ( .A(core__abc_21380_n9939), .B(core_v0_reg_55_), .Y(core__abc_21380_n9940) );
  AND2X2 AND2X2_5421 ( .A(core__abc_21380_n2282), .B(core_mi_reg_55_), .Y(core__abc_21380_n9941) );
  AND2X2 AND2X2_5422 ( .A(core__abc_21380_n9248_bF_buf0), .B(core__abc_21380_n9942), .Y(core__abc_21380_n9943) );
  AND2X2 AND2X2_5423 ( .A(core__abc_21380_n9947), .B(reset_n_bF_buf72), .Y(core__abc_21380_n9948) );
  AND2X2 AND2X2_5424 ( .A(core__abc_21380_n9946), .B(core__abc_21380_n9948), .Y(core_v0_reg_55__FF_INPUT) );
  AND2X2 AND2X2_5425 ( .A(core__abc_21380_n6395), .B(core__abc_21380_n3167_1_bF_buf5), .Y(core__abc_21380_n9950) );
  AND2X2 AND2X2_5426 ( .A(core__abc_21380_n9951), .B(core_v0_reg_56_), .Y(core__abc_21380_n9952) );
  AND2X2 AND2X2_5427 ( .A(core__abc_21380_n2302), .B(core_mi_reg_56_), .Y(core__abc_21380_n9953) );
  AND2X2 AND2X2_5428 ( .A(core__abc_21380_n9248_bF_buf7), .B(core__abc_21380_n9954), .Y(core__abc_21380_n9955) );
  AND2X2 AND2X2_5429 ( .A(core__abc_21380_n3313_bF_buf11), .B(core__abc_21380_n9956), .Y(core__abc_21380_n9957) );
  AND2X2 AND2X2_543 ( .A(_abc_19068_n1802), .B(reset_n_bF_buf39), .Y(word2_reg_13__FF_INPUT) );
  AND2X2 AND2X2_5430 ( .A(core__abc_21380_n9961), .B(reset_n_bF_buf71), .Y(core__abc_21380_n9962) );
  AND2X2 AND2X2_5431 ( .A(core__abc_21380_n9960), .B(core__abc_21380_n9962), .Y(core_v0_reg_56__FF_INPUT) );
  AND2X2 AND2X2_5432 ( .A(core__abc_21380_n6430), .B(core__abc_21380_n3167_1_bF_buf4), .Y(core__abc_21380_n9964) );
  AND2X2 AND2X2_5433 ( .A(core__abc_21380_n3313_bF_buf10), .B(core__abc_21380_n9965), .Y(core__abc_21380_n9966) );
  AND2X2 AND2X2_5434 ( .A(core__abc_21380_n9967), .B(core_v0_reg_57_), .Y(core__abc_21380_n9968) );
  AND2X2 AND2X2_5435 ( .A(core__abc_21380_n2320), .B(core_mi_reg_57_), .Y(core__abc_21380_n9969) );
  AND2X2 AND2X2_5436 ( .A(core__abc_21380_n9248_bF_buf6), .B(core__abc_21380_n9970), .Y(core__abc_21380_n9971) );
  AND2X2 AND2X2_5437 ( .A(core__abc_21380_n9975), .B(reset_n_bF_buf70), .Y(core__abc_21380_n9976) );
  AND2X2 AND2X2_5438 ( .A(core__abc_21380_n9974), .B(core__abc_21380_n9976), .Y(core_v0_reg_57__FF_INPUT) );
  AND2X2 AND2X2_5439 ( .A(core__abc_21380_n6470), .B(core__abc_21380_n3167_1_bF_buf3), .Y(core__abc_21380_n9978) );
  AND2X2 AND2X2_544 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_78_), .Y(_abc_19068_n1804) );
  AND2X2 AND2X2_5440 ( .A(core__abc_21380_n3313_bF_buf9), .B(core_key_58_), .Y(core__abc_21380_n9979) );
  AND2X2 AND2X2_5441 ( .A(core__abc_21380_n9980), .B(core_v0_reg_58_), .Y(core__abc_21380_n9981) );
  AND2X2 AND2X2_5442 ( .A(core__abc_21380_n2338), .B(core_mi_reg_58_), .Y(core__abc_21380_n9982) );
  AND2X2 AND2X2_5443 ( .A(core__abc_21380_n9248_bF_buf5), .B(core__abc_21380_n9983), .Y(core__abc_21380_n9984) );
  AND2X2 AND2X2_5444 ( .A(core__abc_21380_n9988), .B(reset_n_bF_buf69), .Y(core__abc_21380_n9989) );
  AND2X2 AND2X2_5445 ( .A(core__abc_21380_n9987), .B(core__abc_21380_n9989), .Y(core_v0_reg_58__FF_INPUT) );
  AND2X2 AND2X2_5446 ( .A(core__abc_21380_n6504), .B(core__abc_21380_n3167_1_bF_buf2), .Y(core__abc_21380_n9991) );
  AND2X2 AND2X2_5447 ( .A(core__abc_21380_n3313_bF_buf8), .B(core_key_59_), .Y(core__abc_21380_n9992) );
  AND2X2 AND2X2_5448 ( .A(core__abc_21380_n9993), .B(core_v0_reg_59_), .Y(core__abc_21380_n9994) );
  AND2X2 AND2X2_5449 ( .A(core__abc_21380_n2356), .B(core_mi_reg_59_), .Y(core__abc_21380_n9995) );
  AND2X2 AND2X2_545 ( .A(_abc_19068_n1620_bF_buf8), .B(word2_reg_14_), .Y(_abc_19068_n1805) );
  AND2X2 AND2X2_5450 ( .A(core__abc_21380_n9248_bF_buf4), .B(core__abc_21380_n9996), .Y(core__abc_21380_n9997) );
  AND2X2 AND2X2_5451 ( .A(core__abc_21380_n10001), .B(reset_n_bF_buf68), .Y(core__abc_21380_n10002) );
  AND2X2 AND2X2_5452 ( .A(core__abc_21380_n10000), .B(core__abc_21380_n10002), .Y(core_v0_reg_59__FF_INPUT) );
  AND2X2 AND2X2_5453 ( .A(core__abc_21380_n6553), .B(core__abc_21380_n3167_1_bF_buf1), .Y(core__abc_21380_n10004) );
  AND2X2 AND2X2_5454 ( .A(core__abc_21380_n3313_bF_buf7), .B(core__abc_21380_n10005), .Y(core__abc_21380_n10006) );
  AND2X2 AND2X2_5455 ( .A(core__abc_21380_n10007), .B(core_v0_reg_60_), .Y(core__abc_21380_n10008) );
  AND2X2 AND2X2_5456 ( .A(core__abc_21380_n2376), .B(core_mi_reg_60_), .Y(core__abc_21380_n10009) );
  AND2X2 AND2X2_5457 ( .A(core__abc_21380_n9248_bF_buf3), .B(core__abc_21380_n10010), .Y(core__abc_21380_n10011) );
  AND2X2 AND2X2_5458 ( .A(core__abc_21380_n10015), .B(reset_n_bF_buf67), .Y(core__abc_21380_n10016) );
  AND2X2 AND2X2_5459 ( .A(core__abc_21380_n10014), .B(core__abc_21380_n10016), .Y(core_v0_reg_60__FF_INPUT) );
  AND2X2 AND2X2_546 ( .A(_abc_19068_n1806), .B(reset_n_bF_buf38), .Y(word2_reg_14__FF_INPUT) );
  AND2X2 AND2X2_5460 ( .A(core__abc_21380_n6588), .B(core__abc_21380_n3167_1_bF_buf0), .Y(core__abc_21380_n10018) );
  AND2X2 AND2X2_5461 ( .A(core__abc_21380_n10019), .B(core_v0_reg_61_), .Y(core__abc_21380_n10020) );
  AND2X2 AND2X2_5462 ( .A(core__abc_21380_n2394), .B(core_mi_reg_61_), .Y(core__abc_21380_n10021) );
  AND2X2 AND2X2_5463 ( .A(core__abc_21380_n9248_bF_buf2), .B(core__abc_21380_n10022), .Y(core__abc_21380_n10023) );
  AND2X2 AND2X2_5464 ( .A(core__abc_21380_n10027), .B(reset_n_bF_buf66), .Y(core__abc_21380_n10028) );
  AND2X2 AND2X2_5465 ( .A(core__abc_21380_n10026), .B(core__abc_21380_n10028), .Y(core_v0_reg_61__FF_INPUT) );
  AND2X2 AND2X2_5466 ( .A(core__abc_21380_n6629), .B(core__abc_21380_n3167_1_bF_buf15_bF_buf3), .Y(core__abc_21380_n10030) );
  AND2X2 AND2X2_5467 ( .A(core__abc_21380_n10031), .B(core_v0_reg_62_), .Y(core__abc_21380_n10032) );
  AND2X2 AND2X2_5468 ( .A(core__abc_21380_n2412), .B(core_mi_reg_62_), .Y(core__abc_21380_n10033) );
  AND2X2 AND2X2_5469 ( .A(core__abc_21380_n9248_bF_buf1), .B(core__abc_21380_n10034), .Y(core__abc_21380_n10035) );
  AND2X2 AND2X2_547 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_79_), .Y(_abc_19068_n1808) );
  AND2X2 AND2X2_5470 ( .A(core__abc_21380_n10039), .B(reset_n_bF_buf65), .Y(core__abc_21380_n10040) );
  AND2X2 AND2X2_5471 ( .A(core__abc_21380_n10038), .B(core__abc_21380_n10040), .Y(core_v0_reg_62__FF_INPUT) );
  AND2X2 AND2X2_5472 ( .A(core__abc_21380_n6667), .B(core__abc_21380_n3167_1_bF_buf14_bF_buf3), .Y(core__abc_21380_n10042) );
  AND2X2 AND2X2_5473 ( .A(core__abc_21380_n10043), .B(core_v0_reg_63_), .Y(core__abc_21380_n10044) );
  AND2X2 AND2X2_5474 ( .A(core__abc_21380_n2430_1), .B(core_mi_reg_63_), .Y(core__abc_21380_n10045) );
  AND2X2 AND2X2_5475 ( .A(core__abc_21380_n9248_bF_buf0), .B(core__abc_21380_n10046), .Y(core__abc_21380_n10047) );
  AND2X2 AND2X2_5476 ( .A(core__abc_21380_n10051), .B(reset_n_bF_buf64), .Y(core__abc_21380_n10052) );
  AND2X2 AND2X2_5477 ( .A(core__abc_21380_n10050), .B(core__abc_21380_n10052), .Y(core_v0_reg_63__FF_INPUT) );
  AND2X2 AND2X2_5478 ( .A(core__abc_21380_n1225_1), .B(core__abc_21380_n1220_1), .Y(core__abc_21380_n10054) );
  AND2X2 AND2X2_5479 ( .A(core_siphash_ctrl_reg_6_), .B(reset_n_bF_buf63), .Y(core__abc_21380_n10055) );
  AND2X2 AND2X2_548 ( .A(_abc_19068_n1620_bF_buf7), .B(word2_reg_15_), .Y(_abc_19068_n1809) );
  AND2X2 AND2X2_5480 ( .A(core__abc_21380_n10054), .B(core__abc_21380_n10055), .Y(core__abc_21380_n10056) );
  AND2X2 AND2X2_5481 ( .A(core__abc_21380_n10056), .B(core__abc_21380_n7079), .Y(core__abc_14829_n6021) );
  AND2X2 AND2X2_5482 ( .A(core__abc_21380_n1226_1), .B(core__abc_21380_n1185_1), .Y(core__abc_14829_n6022) );
  AND2X2 AND2X2_5483 ( .A(core__abc_21380_n10056), .B(core_long), .Y(core__abc_14829_n6023) );
  AND2X2 AND2X2_5484 ( .A(core__abc_21380_n10054), .B(core__abc_21380_n1249_1), .Y(core__abc_14829_n6024) );
  AND2X2 AND2X2_5485 ( .A(core__abc_21380_n10062), .B(core_siphash_valid_reg_bF_buf1), .Y(core__abc_21380_n10063) );
  AND2X2 AND2X2_5486 ( .A(core__abc_21380_n10064), .B(reset_n_bF_buf62), .Y(core_siphash_valid_reg_FF_INPUT) );
  AND2X2 AND2X2_549 ( .A(_abc_19068_n1810), .B(reset_n_bF_buf37), .Y(word2_reg_15__FF_INPUT) );
  AND2X2 AND2X2_55 ( .A(_abc_19068_n882_1), .B(core_siphash_valid_reg_bF_buf10), .Y(_abc_19068_n958_1) );
  AND2X2 AND2X2_550 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_80_), .Y(_abc_19068_n1812) );
  AND2X2 AND2X2_551 ( .A(_abc_19068_n1620_bF_buf6), .B(word2_reg_16_), .Y(_abc_19068_n1813) );
  AND2X2 AND2X2_552 ( .A(_abc_19068_n1814), .B(reset_n_bF_buf36), .Y(word2_reg_16__FF_INPUT) );
  AND2X2 AND2X2_553 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_81_), .Y(_abc_19068_n1816) );
  AND2X2 AND2X2_554 ( .A(_abc_19068_n1620_bF_buf5), .B(word2_reg_17_), .Y(_abc_19068_n1817) );
  AND2X2 AND2X2_555 ( .A(_abc_19068_n1818), .B(reset_n_bF_buf35), .Y(word2_reg_17__FF_INPUT) );
  AND2X2 AND2X2_556 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_82_), .Y(_abc_19068_n1820) );
  AND2X2 AND2X2_557 ( .A(_abc_19068_n1620_bF_buf4), .B(word2_reg_18_), .Y(_abc_19068_n1821) );
  AND2X2 AND2X2_558 ( .A(_abc_19068_n1822), .B(reset_n_bF_buf34), .Y(word2_reg_18__FF_INPUT) );
  AND2X2 AND2X2_559 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_83_), .Y(_abc_19068_n1824) );
  AND2X2 AND2X2_56 ( .A(_abc_19068_n885_1), .B(core_compression_rounds_1_), .Y(_abc_19068_n959) );
  AND2X2 AND2X2_560 ( .A(_abc_19068_n1620_bF_buf3), .B(word2_reg_19_), .Y(_abc_19068_n1825) );
  AND2X2 AND2X2_561 ( .A(_abc_19068_n1826), .B(reset_n_bF_buf33), .Y(word2_reg_19__FF_INPUT) );
  AND2X2 AND2X2_562 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_84_), .Y(_abc_19068_n1828) );
  AND2X2 AND2X2_563 ( .A(_abc_19068_n1620_bF_buf2), .B(word2_reg_20_), .Y(_abc_19068_n1829) );
  AND2X2 AND2X2_564 ( .A(_abc_19068_n1830), .B(reset_n_bF_buf32), .Y(word2_reg_20__FF_INPUT) );
  AND2X2 AND2X2_565 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_85_), .Y(_abc_19068_n1832) );
  AND2X2 AND2X2_566 ( .A(_abc_19068_n1620_bF_buf1), .B(word2_reg_21_), .Y(_abc_19068_n1833) );
  AND2X2 AND2X2_567 ( .A(_abc_19068_n1834), .B(reset_n_bF_buf31), .Y(word2_reg_21__FF_INPUT) );
  AND2X2 AND2X2_568 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_86_), .Y(_abc_19068_n1836) );
  AND2X2 AND2X2_569 ( .A(_abc_19068_n1620_bF_buf0), .B(word2_reg_22_), .Y(_abc_19068_n1837) );
  AND2X2 AND2X2_57 ( .A(_abc_19068_n902_bF_buf2), .B(word2_reg_1_), .Y(_abc_19068_n962) );
  AND2X2 AND2X2_570 ( .A(_abc_19068_n1838), .B(reset_n_bF_buf30), .Y(word2_reg_22__FF_INPUT) );
  AND2X2 AND2X2_571 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_87_), .Y(_abc_19068_n1840) );
  AND2X2 AND2X2_572 ( .A(_abc_19068_n1620_bF_buf10), .B(word2_reg_23_), .Y(_abc_19068_n1841) );
  AND2X2 AND2X2_573 ( .A(_abc_19068_n1842), .B(reset_n_bF_buf29), .Y(word2_reg_23__FF_INPUT) );
  AND2X2 AND2X2_574 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_88_), .Y(_abc_19068_n1844) );
  AND2X2 AND2X2_575 ( .A(_abc_19068_n1620_bF_buf9), .B(word2_reg_24_), .Y(_abc_19068_n1845) );
  AND2X2 AND2X2_576 ( .A(_abc_19068_n1846), .B(reset_n_bF_buf28), .Y(word2_reg_24__FF_INPUT) );
  AND2X2 AND2X2_577 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_89_), .Y(_abc_19068_n1848) );
  AND2X2 AND2X2_578 ( .A(_abc_19068_n1620_bF_buf8), .B(word2_reg_25_), .Y(_abc_19068_n1849) );
  AND2X2 AND2X2_579 ( .A(_abc_19068_n1850), .B(reset_n_bF_buf27), .Y(word2_reg_25__FF_INPUT) );
  AND2X2 AND2X2_58 ( .A(_abc_19068_n915_1_bF_buf2), .B(core_mi_33_), .Y(_abc_19068_n963_1) );
  AND2X2 AND2X2_580 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_90_), .Y(_abc_19068_n1852) );
  AND2X2 AND2X2_581 ( .A(_abc_19068_n1620_bF_buf7), .B(word2_reg_26_), .Y(_abc_19068_n1853) );
  AND2X2 AND2X2_582 ( .A(_abc_19068_n1854), .B(reset_n_bF_buf26), .Y(word2_reg_26__FF_INPUT) );
  AND2X2 AND2X2_583 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_91_), .Y(_abc_19068_n1856) );
  AND2X2 AND2X2_584 ( .A(_abc_19068_n1620_bF_buf6), .B(word2_reg_27_), .Y(_abc_19068_n1857) );
  AND2X2 AND2X2_585 ( .A(_abc_19068_n1858), .B(reset_n_bF_buf25), .Y(word2_reg_27__FF_INPUT) );
  AND2X2 AND2X2_586 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_92_), .Y(_abc_19068_n1860) );
  AND2X2 AND2X2_587 ( .A(_abc_19068_n1620_bF_buf5), .B(word2_reg_28_), .Y(_abc_19068_n1861) );
  AND2X2 AND2X2_588 ( .A(_abc_19068_n1862), .B(reset_n_bF_buf24), .Y(word2_reg_28__FF_INPUT) );
  AND2X2 AND2X2_589 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_93_), .Y(_abc_19068_n1864) );
  AND2X2 AND2X2_59 ( .A(_abc_19068_n897_1_bF_buf2), .B(word0_reg_1_), .Y(_abc_19068_n964_1) );
  AND2X2 AND2X2_590 ( .A(_abc_19068_n1620_bF_buf4), .B(word2_reg_29_), .Y(_abc_19068_n1865) );
  AND2X2 AND2X2_591 ( .A(_abc_19068_n1866), .B(reset_n_bF_buf23), .Y(word2_reg_29__FF_INPUT) );
  AND2X2 AND2X2_592 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_94_), .Y(_abc_19068_n1868) );
  AND2X2 AND2X2_593 ( .A(_abc_19068_n1620_bF_buf3), .B(word2_reg_30_), .Y(_abc_19068_n1869) );
  AND2X2 AND2X2_594 ( .A(_abc_19068_n1870), .B(reset_n_bF_buf22), .Y(word2_reg_30__FF_INPUT) );
  AND2X2 AND2X2_595 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_95_), .Y(_abc_19068_n1872) );
  AND2X2 AND2X2_596 ( .A(_abc_19068_n1620_bF_buf2), .B(word2_reg_31_), .Y(_abc_19068_n1873) );
  AND2X2 AND2X2_597 ( .A(_abc_19068_n1874), .B(reset_n_bF_buf21), .Y(word2_reg_31__FF_INPUT) );
  AND2X2 AND2X2_598 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_32_), .Y(_abc_19068_n1876) );
  AND2X2 AND2X2_599 ( .A(_abc_19068_n1620_bF_buf1), .B(word1_reg_0_), .Y(_abc_19068_n1877) );
  AND2X2 AND2X2_6 ( .A(_abc_19068_n877_1), .B(_abc_19068_n880_1), .Y(_abc_19068_n881) );
  AND2X2 AND2X2_60 ( .A(_abc_19068_n939_1_bF_buf3), .B(core_key_65_), .Y(_abc_19068_n968) );
  AND2X2 AND2X2_600 ( .A(_abc_19068_n1878), .B(reset_n_bF_buf20), .Y(word1_reg_0__FF_INPUT) );
  AND2X2 AND2X2_601 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_33_), .Y(_abc_19068_n1880) );
  AND2X2 AND2X2_602 ( .A(_abc_19068_n1620_bF_buf0), .B(word1_reg_1_), .Y(_abc_19068_n1881) );
  AND2X2 AND2X2_603 ( .A(_abc_19068_n1882), .B(reset_n_bF_buf19), .Y(word1_reg_1__FF_INPUT) );
  AND2X2 AND2X2_604 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_34_), .Y(_abc_19068_n1884) );
  AND2X2 AND2X2_605 ( .A(_abc_19068_n1620_bF_buf10), .B(word1_reg_2_), .Y(_abc_19068_n1885) );
  AND2X2 AND2X2_606 ( .A(_abc_19068_n1886), .B(reset_n_bF_buf18), .Y(word1_reg_2__FF_INPUT) );
  AND2X2 AND2X2_607 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_35_), .Y(_abc_19068_n1888) );
  AND2X2 AND2X2_608 ( .A(_abc_19068_n1620_bF_buf9), .B(word1_reg_3_), .Y(_abc_19068_n1889) );
  AND2X2 AND2X2_609 ( .A(_abc_19068_n1890), .B(reset_n_bF_buf17), .Y(word1_reg_3__FF_INPUT) );
  AND2X2 AND2X2_61 ( .A(_abc_19068_n941_bF_buf3), .B(core_key_97_), .Y(_abc_19068_n969_1) );
  AND2X2 AND2X2_610 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_36_), .Y(_abc_19068_n1892) );
  AND2X2 AND2X2_611 ( .A(_abc_19068_n1620_bF_buf8), .B(word1_reg_4_), .Y(_abc_19068_n1893) );
  AND2X2 AND2X2_612 ( .A(_abc_19068_n1894), .B(reset_n_bF_buf16), .Y(word1_reg_4__FF_INPUT) );
  AND2X2 AND2X2_613 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_37_), .Y(_abc_19068_n1896) );
  AND2X2 AND2X2_614 ( .A(_abc_19068_n1620_bF_buf7), .B(word1_reg_5_), .Y(_abc_19068_n1897) );
  AND2X2 AND2X2_615 ( .A(_abc_19068_n1898), .B(reset_n_bF_buf15), .Y(word1_reg_5__FF_INPUT) );
  AND2X2 AND2X2_616 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_38_), .Y(_abc_19068_n1900) );
  AND2X2 AND2X2_617 ( .A(_abc_19068_n1620_bF_buf6), .B(word1_reg_6_), .Y(_abc_19068_n1901) );
  AND2X2 AND2X2_618 ( .A(_abc_19068_n1902), .B(reset_n_bF_buf14), .Y(word1_reg_6__FF_INPUT) );
  AND2X2 AND2X2_619 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_39_), .Y(_abc_19068_n1904) );
  AND2X2 AND2X2_62 ( .A(_abc_19068_n889_1), .B(core_compress), .Y(_abc_19068_n971) );
  AND2X2 AND2X2_620 ( .A(_abc_19068_n1620_bF_buf5), .B(word1_reg_7_), .Y(_abc_19068_n1905) );
  AND2X2 AND2X2_621 ( .A(_abc_19068_n1906), .B(reset_n_bF_buf13), .Y(word1_reg_7__FF_INPUT) );
  AND2X2 AND2X2_622 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_40_), .Y(_abc_19068_n1908) );
  AND2X2 AND2X2_623 ( .A(_abc_19068_n1620_bF_buf4), .B(word1_reg_8_), .Y(_abc_19068_n1909) );
  AND2X2 AND2X2_624 ( .A(_abc_19068_n1910), .B(reset_n_bF_buf12), .Y(word1_reg_8__FF_INPUT) );
  AND2X2 AND2X2_625 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_41_), .Y(_abc_19068_n1912) );
  AND2X2 AND2X2_626 ( .A(_abc_19068_n1620_bF_buf3), .B(word1_reg_9_), .Y(_abc_19068_n1913) );
  AND2X2 AND2X2_627 ( .A(_abc_19068_n1914), .B(reset_n_bF_buf11), .Y(word1_reg_9__FF_INPUT) );
  AND2X2 AND2X2_628 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_42_), .Y(_abc_19068_n1916) );
  AND2X2 AND2X2_629 ( .A(_abc_19068_n1620_bF_buf2), .B(word1_reg_10_), .Y(_abc_19068_n1917) );
  AND2X2 AND2X2_63 ( .A(_abc_19068_n945_1_bF_buf3), .B(core_mi_1_), .Y(_abc_19068_n972_1) );
  AND2X2 AND2X2_630 ( .A(_abc_19068_n1918), .B(reset_n_bF_buf10), .Y(word1_reg_10__FF_INPUT) );
  AND2X2 AND2X2_631 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_43_), .Y(_abc_19068_n1920) );
  AND2X2 AND2X2_632 ( .A(_abc_19068_n1620_bF_buf1), .B(word1_reg_11_), .Y(_abc_19068_n1921) );
  AND2X2 AND2X2_633 ( .A(_abc_19068_n1922), .B(reset_n_bF_buf9), .Y(word1_reg_11__FF_INPUT) );
  AND2X2 AND2X2_634 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_44_), .Y(_abc_19068_n1924) );
  AND2X2 AND2X2_635 ( .A(_abc_19068_n1620_bF_buf0), .B(word1_reg_12_), .Y(_abc_19068_n1925) );
  AND2X2 AND2X2_636 ( .A(_abc_19068_n1926), .B(reset_n_bF_buf8), .Y(word1_reg_12__FF_INPUT) );
  AND2X2 AND2X2_637 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_45_), .Y(_abc_19068_n1928) );
  AND2X2 AND2X2_638 ( .A(_abc_19068_n1620_bF_buf10), .B(word1_reg_13_), .Y(_abc_19068_n1929) );
  AND2X2 AND2X2_639 ( .A(_abc_19068_n1930), .B(reset_n_bF_buf7), .Y(word1_reg_13__FF_INPUT) );
  AND2X2 AND2X2_64 ( .A(_abc_19068_n899_bF_buf2), .B(word3_reg_1_), .Y(_abc_19068_n974) );
  AND2X2 AND2X2_640 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_46_), .Y(_abc_19068_n1932) );
  AND2X2 AND2X2_641 ( .A(_abc_19068_n1620_bF_buf9), .B(word1_reg_14_), .Y(_abc_19068_n1933) );
  AND2X2 AND2X2_642 ( .A(_abc_19068_n1934), .B(reset_n_bF_buf6), .Y(word1_reg_14__FF_INPUT) );
  AND2X2 AND2X2_643 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_47_), .Y(_abc_19068_n1936) );
  AND2X2 AND2X2_644 ( .A(_abc_19068_n1620_bF_buf8), .B(word1_reg_15_), .Y(_abc_19068_n1937) );
  AND2X2 AND2X2_645 ( .A(_abc_19068_n1938), .B(reset_n_bF_buf5), .Y(word1_reg_15__FF_INPUT) );
  AND2X2 AND2X2_646 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_48_), .Y(_abc_19068_n1940) );
  AND2X2 AND2X2_647 ( .A(_abc_19068_n1620_bF_buf7), .B(word1_reg_16_), .Y(_abc_19068_n1941) );
  AND2X2 AND2X2_648 ( .A(_abc_19068_n1942), .B(reset_n_bF_buf4), .Y(word1_reg_16__FF_INPUT) );
  AND2X2 AND2X2_649 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_49_), .Y(_abc_19068_n1944) );
  AND2X2 AND2X2_65 ( .A(_abc_19068_n916_1_bF_buf2), .B(word1_reg_1_), .Y(_abc_19068_n975_1) );
  AND2X2 AND2X2_650 ( .A(_abc_19068_n1620_bF_buf6), .B(word1_reg_17_), .Y(_abc_19068_n1945) );
  AND2X2 AND2X2_651 ( .A(_abc_19068_n1946), .B(reset_n_bF_buf3), .Y(word1_reg_17__FF_INPUT) );
  AND2X2 AND2X2_652 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_50_), .Y(_abc_19068_n1948) );
  AND2X2 AND2X2_653 ( .A(_abc_19068_n1620_bF_buf5), .B(word1_reg_18_), .Y(_abc_19068_n1949) );
  AND2X2 AND2X2_654 ( .A(_abc_19068_n1950), .B(reset_n_bF_buf2), .Y(word1_reg_18__FF_INPUT) );
  AND2X2 AND2X2_655 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_51_), .Y(_abc_19068_n1952) );
  AND2X2 AND2X2_656 ( .A(_abc_19068_n1620_bF_buf4), .B(word1_reg_19_), .Y(_abc_19068_n1953) );
  AND2X2 AND2X2_657 ( .A(_abc_19068_n1954), .B(reset_n_bF_buf1), .Y(word1_reg_19__FF_INPUT) );
  AND2X2 AND2X2_658 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_52_), .Y(_abc_19068_n1956) );
  AND2X2 AND2X2_659 ( .A(_abc_19068_n1620_bF_buf3), .B(word1_reg_20_), .Y(_abc_19068_n1957) );
  AND2X2 AND2X2_66 ( .A(_abc_19068_n979_1), .B(_abc_19068_n923_bF_buf3), .Y(_auto_iopadmap_cc_313_execute_30317_1_) );
  AND2X2 AND2X2_660 ( .A(_abc_19068_n1958), .B(reset_n_bF_buf0), .Y(word1_reg_20__FF_INPUT) );
  AND2X2 AND2X2_661 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_53_), .Y(_abc_19068_n1960) );
  AND2X2 AND2X2_662 ( .A(_abc_19068_n1620_bF_buf2), .B(word1_reg_21_), .Y(_abc_19068_n1961) );
  AND2X2 AND2X2_663 ( .A(_abc_19068_n1962), .B(reset_n_bF_buf84), .Y(word1_reg_21__FF_INPUT) );
  AND2X2 AND2X2_664 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_54_), .Y(_abc_19068_n1964) );
  AND2X2 AND2X2_665 ( .A(_abc_19068_n1620_bF_buf1), .B(word1_reg_22_), .Y(_abc_19068_n1965) );
  AND2X2 AND2X2_666 ( .A(_abc_19068_n1966), .B(reset_n_bF_buf83), .Y(word1_reg_22__FF_INPUT) );
  AND2X2 AND2X2_667 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_55_), .Y(_abc_19068_n1968) );
  AND2X2 AND2X2_668 ( .A(_abc_19068_n1620_bF_buf0), .B(word1_reg_23_), .Y(_abc_19068_n1969) );
  AND2X2 AND2X2_669 ( .A(_abc_19068_n1970), .B(reset_n_bF_buf82), .Y(word1_reg_23__FF_INPUT) );
  AND2X2 AND2X2_67 ( .A(_abc_19068_n926_bF_buf2), .B(core_key_2_), .Y(_abc_19068_n981_1) );
  AND2X2 AND2X2_670 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_56_), .Y(_abc_19068_n1972) );
  AND2X2 AND2X2_671 ( .A(_abc_19068_n1620_bF_buf10), .B(word1_reg_24_), .Y(_abc_19068_n1973) );
  AND2X2 AND2X2_672 ( .A(_abc_19068_n1974), .B(reset_n_bF_buf81), .Y(word1_reg_24__FF_INPUT) );
  AND2X2 AND2X2_673 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_57_), .Y(_abc_19068_n1976) );
  AND2X2 AND2X2_674 ( .A(_abc_19068_n1620_bF_buf9), .B(word1_reg_25_), .Y(_abc_19068_n1977) );
  AND2X2 AND2X2_675 ( .A(_abc_19068_n1978), .B(reset_n_bF_buf80), .Y(word1_reg_25__FF_INPUT) );
  AND2X2 AND2X2_676 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_58_), .Y(_abc_19068_n1980) );
  AND2X2 AND2X2_677 ( .A(_abc_19068_n1620_bF_buf8), .B(word1_reg_26_), .Y(_abc_19068_n1981) );
  AND2X2 AND2X2_678 ( .A(_abc_19068_n1982), .B(reset_n_bF_buf79), .Y(word1_reg_26__FF_INPUT) );
  AND2X2 AND2X2_679 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_59_), .Y(_abc_19068_n1984) );
  AND2X2 AND2X2_68 ( .A(_abc_19068_n939_1_bF_buf2), .B(core_key_66_), .Y(_abc_19068_n982_1) );
  AND2X2 AND2X2_680 ( .A(_abc_19068_n1620_bF_buf7), .B(word1_reg_27_), .Y(_abc_19068_n1985) );
  AND2X2 AND2X2_681 ( .A(_abc_19068_n1986), .B(reset_n_bF_buf78), .Y(word1_reg_27__FF_INPUT) );
  AND2X2 AND2X2_682 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_60_), .Y(_abc_19068_n1988) );
  AND2X2 AND2X2_683 ( .A(_abc_19068_n1620_bF_buf6), .B(word1_reg_28_), .Y(_abc_19068_n1989) );
  AND2X2 AND2X2_684 ( .A(_abc_19068_n1990), .B(reset_n_bF_buf77), .Y(word1_reg_28__FF_INPUT) );
  AND2X2 AND2X2_685 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_61_), .Y(_abc_19068_n1992) );
  AND2X2 AND2X2_686 ( .A(_abc_19068_n1620_bF_buf5), .B(word1_reg_29_), .Y(_abc_19068_n1993) );
  AND2X2 AND2X2_687 ( .A(_abc_19068_n1994), .B(reset_n_bF_buf76), .Y(word1_reg_29__FF_INPUT) );
  AND2X2 AND2X2_688 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_62_), .Y(_abc_19068_n1996) );
  AND2X2 AND2X2_689 ( .A(_abc_19068_n1620_bF_buf4), .B(word1_reg_30_), .Y(_abc_19068_n1997) );
  AND2X2 AND2X2_69 ( .A(_abc_19068_n941_bF_buf2), .B(core_key_98_), .Y(_abc_19068_n983) );
  AND2X2 AND2X2_690 ( .A(_abc_19068_n1998), .B(reset_n_bF_buf75), .Y(word1_reg_30__FF_INPUT) );
  AND2X2 AND2X2_691 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_63_), .Y(_abc_19068_n2000) );
  AND2X2 AND2X2_692 ( .A(_abc_19068_n1620_bF_buf3), .B(word1_reg_31_), .Y(_abc_19068_n2001) );
  AND2X2 AND2X2_693 ( .A(_abc_19068_n2002), .B(reset_n_bF_buf74), .Y(word1_reg_31__FF_INPUT) );
  AND2X2 AND2X2_694 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_0_), .Y(_abc_19068_n2004) );
  AND2X2 AND2X2_695 ( .A(_abc_19068_n1620_bF_buf2), .B(word0_reg_0_), .Y(_abc_19068_n2005) );
  AND2X2 AND2X2_696 ( .A(_abc_19068_n2006), .B(reset_n_bF_buf73), .Y(word0_reg_0__FF_INPUT) );
  AND2X2 AND2X2_697 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_1_), .Y(_abc_19068_n2008) );
  AND2X2 AND2X2_698 ( .A(_abc_19068_n1620_bF_buf1), .B(word0_reg_1_), .Y(_abc_19068_n2009) );
  AND2X2 AND2X2_699 ( .A(_abc_19068_n2010), .B(reset_n_bF_buf72), .Y(word0_reg_1__FF_INPUT) );
  AND2X2 AND2X2_7 ( .A(_abc_19068_n881), .B(_abc_19068_n874_1), .Y(_abc_19068_n882_1) );
  AND2X2 AND2X2_70 ( .A(_abc_19068_n899_bF_buf1), .B(word3_reg_2_), .Y(_abc_19068_n985_1) );
  AND2X2 AND2X2_700 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_2_), .Y(_abc_19068_n2012) );
  AND2X2 AND2X2_701 ( .A(_abc_19068_n1620_bF_buf0), .B(word0_reg_2_), .Y(_abc_19068_n2013) );
  AND2X2 AND2X2_702 ( .A(_abc_19068_n2014), .B(reset_n_bF_buf71), .Y(word0_reg_2__FF_INPUT) );
  AND2X2 AND2X2_703 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_3_), .Y(_abc_19068_n2016) );
  AND2X2 AND2X2_704 ( .A(_abc_19068_n1620_bF_buf10), .B(word0_reg_3_), .Y(_abc_19068_n2017) );
  AND2X2 AND2X2_705 ( .A(_abc_19068_n2018), .B(reset_n_bF_buf70), .Y(word0_reg_3__FF_INPUT) );
  AND2X2 AND2X2_706 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_4_), .Y(_abc_19068_n2020) );
  AND2X2 AND2X2_707 ( .A(_abc_19068_n1620_bF_buf9), .B(word0_reg_4_), .Y(_abc_19068_n2021) );
  AND2X2 AND2X2_708 ( .A(_abc_19068_n2022), .B(reset_n_bF_buf69), .Y(word0_reg_4__FF_INPUT) );
  AND2X2 AND2X2_709 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_5_), .Y(_abc_19068_n2024) );
  AND2X2 AND2X2_71 ( .A(_abc_19068_n902_bF_buf1), .B(word2_reg_2_), .Y(_abc_19068_n986) );
  AND2X2 AND2X2_710 ( .A(_abc_19068_n1620_bF_buf8), .B(word0_reg_5_), .Y(_abc_19068_n2025) );
  AND2X2 AND2X2_711 ( .A(_abc_19068_n2026), .B(reset_n_bF_buf68), .Y(word0_reg_5__FF_INPUT) );
  AND2X2 AND2X2_712 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_6_), .Y(_abc_19068_n2028) );
  AND2X2 AND2X2_713 ( .A(_abc_19068_n1620_bF_buf7), .B(word0_reg_6_), .Y(_abc_19068_n2029) );
  AND2X2 AND2X2_714 ( .A(_abc_19068_n2030), .B(reset_n_bF_buf67), .Y(word0_reg_6__FF_INPUT) );
  AND2X2 AND2X2_715 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_7_), .Y(_abc_19068_n2032) );
  AND2X2 AND2X2_716 ( .A(_abc_19068_n1620_bF_buf6), .B(word0_reg_7_), .Y(_abc_19068_n2033) );
  AND2X2 AND2X2_717 ( .A(_abc_19068_n2034), .B(reset_n_bF_buf66), .Y(word0_reg_7__FF_INPUT) );
  AND2X2 AND2X2_718 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_8_), .Y(_abc_19068_n2036) );
  AND2X2 AND2X2_719 ( .A(_abc_19068_n1620_bF_buf5), .B(word0_reg_8_), .Y(_abc_19068_n2037) );
  AND2X2 AND2X2_72 ( .A(_abc_19068_n924_1_bF_buf2), .B(core_key_34_), .Y(_abc_19068_n990_1) );
  AND2X2 AND2X2_720 ( .A(_abc_19068_n2038), .B(reset_n_bF_buf65), .Y(word0_reg_8__FF_INPUT) );
  AND2X2 AND2X2_721 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_9_), .Y(_abc_19068_n2040) );
  AND2X2 AND2X2_722 ( .A(_abc_19068_n1620_bF_buf4), .B(word0_reg_9_), .Y(_abc_19068_n2041) );
  AND2X2 AND2X2_723 ( .A(_abc_19068_n2042), .B(reset_n_bF_buf64), .Y(word0_reg_9__FF_INPUT) );
  AND2X2 AND2X2_724 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_10_), .Y(_abc_19068_n2044) );
  AND2X2 AND2X2_725 ( .A(_abc_19068_n1620_bF_buf3), .B(word0_reg_10_), .Y(_abc_19068_n2045) );
  AND2X2 AND2X2_726 ( .A(_abc_19068_n2046), .B(reset_n_bF_buf63), .Y(word0_reg_10__FF_INPUT) );
  AND2X2 AND2X2_727 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_11_), .Y(_abc_19068_n2048) );
  AND2X2 AND2X2_728 ( .A(_abc_19068_n1620_bF_buf2), .B(word0_reg_11_), .Y(_abc_19068_n2049) );
  AND2X2 AND2X2_729 ( .A(_abc_19068_n2050), .B(reset_n_bF_buf62), .Y(word0_reg_11__FF_INPUT) );
  AND2X2 AND2X2_73 ( .A(_abc_19068_n885_1), .B(core_compression_rounds_2_), .Y(_abc_19068_n991_1) );
  AND2X2 AND2X2_730 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_12_), .Y(_abc_19068_n2052) );
  AND2X2 AND2X2_731 ( .A(_abc_19068_n1620_bF_buf1), .B(word0_reg_12_), .Y(_abc_19068_n2053) );
  AND2X2 AND2X2_732 ( .A(_abc_19068_n2054), .B(reset_n_bF_buf61), .Y(word0_reg_12__FF_INPUT) );
  AND2X2 AND2X2_733 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_13_), .Y(_abc_19068_n2056) );
  AND2X2 AND2X2_734 ( .A(_abc_19068_n1620_bF_buf0), .B(word0_reg_13_), .Y(_abc_19068_n2057) );
  AND2X2 AND2X2_735 ( .A(_abc_19068_n2058), .B(reset_n_bF_buf60), .Y(word0_reg_13__FF_INPUT) );
  AND2X2 AND2X2_736 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_14_), .Y(_abc_19068_n2060) );
  AND2X2 AND2X2_737 ( .A(_abc_19068_n1620_bF_buf10), .B(word0_reg_14_), .Y(_abc_19068_n2061) );
  AND2X2 AND2X2_738 ( .A(_abc_19068_n2062), .B(reset_n_bF_buf59), .Y(word0_reg_14__FF_INPUT) );
  AND2X2 AND2X2_739 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_15_), .Y(_abc_19068_n2064) );
  AND2X2 AND2X2_74 ( .A(_abc_19068_n889_1), .B(core_finalize), .Y(_abc_19068_n992) );
  AND2X2 AND2X2_740 ( .A(_abc_19068_n1620_bF_buf9), .B(word0_reg_15_), .Y(_abc_19068_n2065) );
  AND2X2 AND2X2_741 ( .A(_abc_19068_n2066), .B(reset_n_bF_buf58), .Y(word0_reg_15__FF_INPUT) );
  AND2X2 AND2X2_742 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_16_), .Y(_abc_19068_n2068) );
  AND2X2 AND2X2_743 ( .A(_abc_19068_n1620_bF_buf8), .B(word0_reg_16_), .Y(_abc_19068_n2069) );
  AND2X2 AND2X2_744 ( .A(_abc_19068_n2070), .B(reset_n_bF_buf57), .Y(word0_reg_16__FF_INPUT) );
  AND2X2 AND2X2_745 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_17_), .Y(_abc_19068_n2072) );
  AND2X2 AND2X2_746 ( .A(_abc_19068_n1620_bF_buf7), .B(word0_reg_17_), .Y(_abc_19068_n2073) );
  AND2X2 AND2X2_747 ( .A(_abc_19068_n2074), .B(reset_n_bF_buf56), .Y(word0_reg_17__FF_INPUT) );
  AND2X2 AND2X2_748 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_18_), .Y(_abc_19068_n2076) );
  AND2X2 AND2X2_749 ( .A(_abc_19068_n1620_bF_buf6), .B(word0_reg_18_), .Y(_abc_19068_n2077) );
  AND2X2 AND2X2_75 ( .A(_abc_19068_n897_1_bF_buf1), .B(word0_reg_2_), .Y(_abc_19068_n995) );
  AND2X2 AND2X2_750 ( .A(_abc_19068_n2078), .B(reset_n_bF_buf55), .Y(word0_reg_18__FF_INPUT) );
  AND2X2 AND2X2_751 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_19_), .Y(_abc_19068_n2080) );
  AND2X2 AND2X2_752 ( .A(_abc_19068_n1620_bF_buf5), .B(word0_reg_19_), .Y(_abc_19068_n2081) );
  AND2X2 AND2X2_753 ( .A(_abc_19068_n2082), .B(reset_n_bF_buf54), .Y(word0_reg_19__FF_INPUT) );
  AND2X2 AND2X2_754 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_20_), .Y(_abc_19068_n2084) );
  AND2X2 AND2X2_755 ( .A(_abc_19068_n1620_bF_buf4), .B(word0_reg_20_), .Y(_abc_19068_n2085) );
  AND2X2 AND2X2_756 ( .A(_abc_19068_n2086), .B(reset_n_bF_buf53), .Y(word0_reg_20__FF_INPUT) );
  AND2X2 AND2X2_757 ( .A(core_siphash_valid_reg_bF_buf1), .B(core_siphash_word_21_), .Y(_abc_19068_n2088) );
  AND2X2 AND2X2_758 ( .A(_abc_19068_n1620_bF_buf3), .B(word0_reg_21_), .Y(_abc_19068_n2089) );
  AND2X2 AND2X2_759 ( .A(_abc_19068_n2090), .B(reset_n_bF_buf52), .Y(word0_reg_21__FF_INPUT) );
  AND2X2 AND2X2_76 ( .A(_abc_19068_n916_1_bF_buf1), .B(word1_reg_2_), .Y(_abc_19068_n996_1) );
  AND2X2 AND2X2_760 ( .A(core_siphash_valid_reg_bF_buf0), .B(core_siphash_word_22_), .Y(_abc_19068_n2092) );
  AND2X2 AND2X2_761 ( .A(_abc_19068_n1620_bF_buf2), .B(word0_reg_22_), .Y(_abc_19068_n2093) );
  AND2X2 AND2X2_762 ( .A(_abc_19068_n2094), .B(reset_n_bF_buf51), .Y(word0_reg_22__FF_INPUT) );
  AND2X2 AND2X2_763 ( .A(core_siphash_valid_reg_bF_buf10), .B(core_siphash_word_23_), .Y(_abc_19068_n2096) );
  AND2X2 AND2X2_764 ( .A(_abc_19068_n1620_bF_buf1), .B(word0_reg_23_), .Y(_abc_19068_n2097) );
  AND2X2 AND2X2_765 ( .A(_abc_19068_n2098), .B(reset_n_bF_buf50), .Y(word0_reg_23__FF_INPUT) );
  AND2X2 AND2X2_766 ( .A(core_siphash_valid_reg_bF_buf9), .B(core_siphash_word_24_), .Y(_abc_19068_n2100) );
  AND2X2 AND2X2_767 ( .A(_abc_19068_n1620_bF_buf0), .B(word0_reg_24_), .Y(_abc_19068_n2101) );
  AND2X2 AND2X2_768 ( .A(_abc_19068_n2102), .B(reset_n_bF_buf49), .Y(word0_reg_24__FF_INPUT) );
  AND2X2 AND2X2_769 ( .A(core_siphash_valid_reg_bF_buf8), .B(core_siphash_word_25_), .Y(_abc_19068_n2104) );
  AND2X2 AND2X2_77 ( .A(_abc_19068_n915_1_bF_buf1), .B(core_mi_34_), .Y(_abc_19068_n998) );
  AND2X2 AND2X2_770 ( .A(_abc_19068_n1620_bF_buf10), .B(word0_reg_25_), .Y(_abc_19068_n2105) );
  AND2X2 AND2X2_771 ( .A(_abc_19068_n2106), .B(reset_n_bF_buf48), .Y(word0_reg_25__FF_INPUT) );
  AND2X2 AND2X2_772 ( .A(core_siphash_valid_reg_bF_buf7), .B(core_siphash_word_26_), .Y(_abc_19068_n2108) );
  AND2X2 AND2X2_773 ( .A(_abc_19068_n1620_bF_buf9), .B(word0_reg_26_), .Y(_abc_19068_n2109) );
  AND2X2 AND2X2_774 ( .A(_abc_19068_n2110), .B(reset_n_bF_buf47), .Y(word0_reg_26__FF_INPUT) );
  AND2X2 AND2X2_775 ( .A(core_siphash_valid_reg_bF_buf6), .B(core_siphash_word_27_), .Y(_abc_19068_n2112) );
  AND2X2 AND2X2_776 ( .A(_abc_19068_n1620_bF_buf8), .B(word0_reg_27_), .Y(_abc_19068_n2113) );
  AND2X2 AND2X2_777 ( .A(_abc_19068_n2114), .B(reset_n_bF_buf46), .Y(word0_reg_27__FF_INPUT) );
  AND2X2 AND2X2_778 ( .A(core_siphash_valid_reg_bF_buf5), .B(core_siphash_word_28_), .Y(_abc_19068_n2116) );
  AND2X2 AND2X2_779 ( .A(_abc_19068_n1620_bF_buf7), .B(word0_reg_28_), .Y(_abc_19068_n2117) );
  AND2X2 AND2X2_78 ( .A(_abc_19068_n945_1_bF_buf2), .B(core_mi_2_), .Y(_abc_19068_n999_1) );
  AND2X2 AND2X2_780 ( .A(_abc_19068_n2118), .B(reset_n_bF_buf45), .Y(word0_reg_28__FF_INPUT) );
  AND2X2 AND2X2_781 ( .A(core_siphash_valid_reg_bF_buf4), .B(core_siphash_word_29_), .Y(_abc_19068_n2120) );
  AND2X2 AND2X2_782 ( .A(_abc_19068_n1620_bF_buf6), .B(word0_reg_29_), .Y(_abc_19068_n2121) );
  AND2X2 AND2X2_783 ( .A(_abc_19068_n2122), .B(reset_n_bF_buf44), .Y(word0_reg_29__FF_INPUT) );
  AND2X2 AND2X2_784 ( .A(core_siphash_valid_reg_bF_buf3), .B(core_siphash_word_30_), .Y(_abc_19068_n2124) );
  AND2X2 AND2X2_785 ( .A(_abc_19068_n1620_bF_buf5), .B(word0_reg_30_), .Y(_abc_19068_n2125) );
  AND2X2 AND2X2_786 ( .A(_abc_19068_n2126), .B(reset_n_bF_buf43), .Y(word0_reg_30__FF_INPUT) );
  AND2X2 AND2X2_787 ( .A(core_siphash_valid_reg_bF_buf2), .B(core_siphash_word_31_), .Y(_abc_19068_n2128) );
  AND2X2 AND2X2_788 ( .A(_abc_19068_n1620_bF_buf4), .B(word0_reg_31_), .Y(_abc_19068_n2129) );
  AND2X2 AND2X2_789 ( .A(_abc_19068_n2130), .B(reset_n_bF_buf42), .Y(word0_reg_31__FF_INPUT) );
  AND2X2 AND2X2_79 ( .A(_abc_19068_n1003_1), .B(_abc_19068_n923_bF_buf2), .Y(_auto_iopadmap_cc_313_execute_30317_2_) );
  AND2X2 AND2X2_790 ( .A(we), .B(cs), .Y(_abc_19068_n2132) );
  AND2X2 AND2X2_791 ( .A(_abc_19068_n915_1_bF_buf1), .B(_abc_19068_n2132), .Y(_abc_19068_n2133) );
  AND2X2 AND2X2_792 ( .A(_abc_19068_n2133_bF_buf6), .B(_abc_19068_n2135), .Y(_abc_19068_n2136) );
  AND2X2 AND2X2_793 ( .A(_abc_19068_n2137), .B(reset_n_bF_buf41), .Y(_abc_19068_n2138) );
  AND2X2 AND2X2_794 ( .A(_abc_19068_n2138), .B(_abc_19068_n2134), .Y(mi1_reg_0__FF_INPUT) );
  AND2X2 AND2X2_795 ( .A(_abc_19068_n2133_bF_buf4), .B(_abc_19068_n2141), .Y(_abc_19068_n2142) );
  AND2X2 AND2X2_796 ( .A(_abc_19068_n2143), .B(reset_n_bF_buf40), .Y(_abc_19068_n2144) );
  AND2X2 AND2X2_797 ( .A(_abc_19068_n2144), .B(_abc_19068_n2140), .Y(mi1_reg_1__FF_INPUT) );
  AND2X2 AND2X2_798 ( .A(_abc_19068_n2133_bF_buf2), .B(_abc_19068_n2147), .Y(_abc_19068_n2148) );
  AND2X2 AND2X2_799 ( .A(_abc_19068_n2149), .B(reset_n_bF_buf39), .Y(_abc_19068_n2150) );
  AND2X2 AND2X2_8 ( .A(\addr[0] ), .B(\addr[1] ), .Y(_abc_19068_n883_1) );
  AND2X2 AND2X2_80 ( .A(_abc_19068_n897_1_bF_buf0), .B(word0_reg_3_), .Y(_abc_19068_n1005_1) );
  AND2X2 AND2X2_800 ( .A(_abc_19068_n2150), .B(_abc_19068_n2146), .Y(mi1_reg_2__FF_INPUT) );
  AND2X2 AND2X2_801 ( .A(_abc_19068_n2133_bF_buf0), .B(_abc_19068_n2153), .Y(_abc_19068_n2154) );
  AND2X2 AND2X2_802 ( .A(_abc_19068_n2155), .B(reset_n_bF_buf38), .Y(_abc_19068_n2156) );
  AND2X2 AND2X2_803 ( .A(_abc_19068_n2156), .B(_abc_19068_n2152), .Y(mi1_reg_3__FF_INPUT) );
  AND2X2 AND2X2_804 ( .A(_abc_19068_n2133_bF_buf6), .B(_abc_19068_n2159), .Y(_abc_19068_n2160) );
  AND2X2 AND2X2_805 ( .A(_abc_19068_n2161), .B(reset_n_bF_buf37), .Y(_abc_19068_n2162) );
  AND2X2 AND2X2_806 ( .A(_abc_19068_n2162), .B(_abc_19068_n2158), .Y(mi1_reg_4__FF_INPUT) );
  AND2X2 AND2X2_807 ( .A(_abc_19068_n2133_bF_buf4), .B(_abc_19068_n2165), .Y(_abc_19068_n2166) );
  AND2X2 AND2X2_808 ( .A(_abc_19068_n2167), .B(reset_n_bF_buf36), .Y(_abc_19068_n2168) );
  AND2X2 AND2X2_809 ( .A(_abc_19068_n2168), .B(_abc_19068_n2164), .Y(mi1_reg_5__FF_INPUT) );
  AND2X2 AND2X2_81 ( .A(_abc_19068_n915_1_bF_buf0), .B(core_mi_35_), .Y(_abc_19068_n1006_1) );
  AND2X2 AND2X2_810 ( .A(_abc_19068_n2133_bF_buf2), .B(_abc_19068_n2171), .Y(_abc_19068_n2172) );
  AND2X2 AND2X2_811 ( .A(_abc_19068_n2173), .B(reset_n_bF_buf35), .Y(_abc_19068_n2174) );
  AND2X2 AND2X2_812 ( .A(_abc_19068_n2174), .B(_abc_19068_n2170), .Y(mi1_reg_6__FF_INPUT) );
  AND2X2 AND2X2_813 ( .A(_abc_19068_n2133_bF_buf0), .B(_abc_19068_n2177), .Y(_abc_19068_n2178) );
  AND2X2 AND2X2_814 ( .A(_abc_19068_n2179), .B(reset_n_bF_buf34), .Y(_abc_19068_n2180) );
  AND2X2 AND2X2_815 ( .A(_abc_19068_n2180), .B(_abc_19068_n2176), .Y(mi1_reg_7__FF_INPUT) );
  AND2X2 AND2X2_816 ( .A(_abc_19068_n2133_bF_buf6), .B(_abc_19068_n2183), .Y(_abc_19068_n2184) );
  AND2X2 AND2X2_817 ( .A(_abc_19068_n2185), .B(reset_n_bF_buf33), .Y(_abc_19068_n2186) );
  AND2X2 AND2X2_818 ( .A(_abc_19068_n2186), .B(_abc_19068_n2182), .Y(mi1_reg_8__FF_INPUT) );
  AND2X2 AND2X2_819 ( .A(_abc_19068_n2133_bF_buf4), .B(_abc_19068_n2189), .Y(_abc_19068_n2190) );
  AND2X2 AND2X2_82 ( .A(_abc_19068_n945_1_bF_buf1), .B(core_mi_3_), .Y(_abc_19068_n1008_1) );
  AND2X2 AND2X2_820 ( .A(_abc_19068_n2191), .B(reset_n_bF_buf32), .Y(_abc_19068_n2192) );
  AND2X2 AND2X2_821 ( .A(_abc_19068_n2192), .B(_abc_19068_n2188), .Y(mi1_reg_9__FF_INPUT) );
  AND2X2 AND2X2_822 ( .A(_abc_19068_n2133_bF_buf2), .B(_abc_19068_n2195), .Y(_abc_19068_n2196) );
  AND2X2 AND2X2_823 ( .A(_abc_19068_n2197), .B(reset_n_bF_buf31), .Y(_abc_19068_n2198) );
  AND2X2 AND2X2_824 ( .A(_abc_19068_n2198), .B(_abc_19068_n2194), .Y(mi1_reg_10__FF_INPUT) );
  AND2X2 AND2X2_825 ( .A(_abc_19068_n2133_bF_buf0), .B(_abc_19068_n2201), .Y(_abc_19068_n2202) );
  AND2X2 AND2X2_826 ( .A(_abc_19068_n2203), .B(reset_n_bF_buf30), .Y(_abc_19068_n2204) );
  AND2X2 AND2X2_827 ( .A(_abc_19068_n2204), .B(_abc_19068_n2200), .Y(mi1_reg_11__FF_INPUT) );
  AND2X2 AND2X2_828 ( .A(_abc_19068_n2133_bF_buf6), .B(_abc_19068_n2207), .Y(_abc_19068_n2208) );
  AND2X2 AND2X2_829 ( .A(_abc_19068_n2209), .B(reset_n_bF_buf29), .Y(_abc_19068_n2210) );
  AND2X2 AND2X2_83 ( .A(_abc_19068_n941_bF_buf1), .B(core_key_99_), .Y(_abc_19068_n1009_1) );
  AND2X2 AND2X2_830 ( .A(_abc_19068_n2210), .B(_abc_19068_n2206), .Y(mi1_reg_12__FF_INPUT) );
  AND2X2 AND2X2_831 ( .A(_abc_19068_n2133_bF_buf4), .B(_abc_19068_n2213), .Y(_abc_19068_n2214) );
  AND2X2 AND2X2_832 ( .A(_abc_19068_n2215), .B(reset_n_bF_buf28), .Y(_abc_19068_n2216) );
  AND2X2 AND2X2_833 ( .A(_abc_19068_n2216), .B(_abc_19068_n2212), .Y(mi1_reg_13__FF_INPUT) );
  AND2X2 AND2X2_834 ( .A(_abc_19068_n2133_bF_buf2), .B(_abc_19068_n2219), .Y(_abc_19068_n2220) );
  AND2X2 AND2X2_835 ( .A(_abc_19068_n2221), .B(reset_n_bF_buf27), .Y(_abc_19068_n2222) );
  AND2X2 AND2X2_836 ( .A(_abc_19068_n2222), .B(_abc_19068_n2218), .Y(mi1_reg_14__FF_INPUT) );
  AND2X2 AND2X2_837 ( .A(_abc_19068_n2133_bF_buf0), .B(_abc_19068_n2225), .Y(_abc_19068_n2226) );
  AND2X2 AND2X2_838 ( .A(_abc_19068_n2227), .B(reset_n_bF_buf26), .Y(_abc_19068_n2228) );
  AND2X2 AND2X2_839 ( .A(_abc_19068_n2228), .B(_abc_19068_n2224), .Y(mi1_reg_15__FF_INPUT) );
  AND2X2 AND2X2_84 ( .A(_abc_19068_n916_1_bF_buf0), .B(word1_reg_3_), .Y(_abc_19068_n1012_1) );
  AND2X2 AND2X2_840 ( .A(_abc_19068_n2133_bF_buf6), .B(_abc_19068_n2231), .Y(_abc_19068_n2232) );
  AND2X2 AND2X2_841 ( .A(_abc_19068_n2233), .B(reset_n_bF_buf25), .Y(_abc_19068_n2234) );
  AND2X2 AND2X2_842 ( .A(_abc_19068_n2234), .B(_abc_19068_n2230), .Y(mi1_reg_16__FF_INPUT) );
  AND2X2 AND2X2_843 ( .A(_abc_19068_n2133_bF_buf4), .B(_abc_19068_n2237), .Y(_abc_19068_n2238) );
  AND2X2 AND2X2_844 ( .A(_abc_19068_n2239), .B(reset_n_bF_buf24), .Y(_abc_19068_n2240) );
  AND2X2 AND2X2_845 ( .A(_abc_19068_n2240), .B(_abc_19068_n2236), .Y(mi1_reg_17__FF_INPUT) );
  AND2X2 AND2X2_846 ( .A(_abc_19068_n2133_bF_buf2), .B(_abc_19068_n2243), .Y(_abc_19068_n2244) );
  AND2X2 AND2X2_847 ( .A(_abc_19068_n2245), .B(reset_n_bF_buf23), .Y(_abc_19068_n2246) );
  AND2X2 AND2X2_848 ( .A(_abc_19068_n2246), .B(_abc_19068_n2242), .Y(mi1_reg_18__FF_INPUT) );
  AND2X2 AND2X2_849 ( .A(_abc_19068_n2133_bF_buf0), .B(_abc_19068_n2249), .Y(_abc_19068_n2250) );
  AND2X2 AND2X2_85 ( .A(_abc_19068_n902_bF_buf0), .B(word2_reg_3_), .Y(_abc_19068_n1013) );
  AND2X2 AND2X2_850 ( .A(_abc_19068_n2251), .B(reset_n_bF_buf22), .Y(_abc_19068_n2252) );
  AND2X2 AND2X2_851 ( .A(_abc_19068_n2252), .B(_abc_19068_n2248), .Y(mi1_reg_19__FF_INPUT) );
  AND2X2 AND2X2_852 ( .A(_abc_19068_n2133_bF_buf6), .B(_abc_19068_n2255), .Y(_abc_19068_n2256) );
  AND2X2 AND2X2_853 ( .A(_abc_19068_n2257), .B(reset_n_bF_buf21), .Y(_abc_19068_n2258) );
  AND2X2 AND2X2_854 ( .A(_abc_19068_n2258), .B(_abc_19068_n2254), .Y(mi1_reg_20__FF_INPUT) );
  AND2X2 AND2X2_855 ( .A(_abc_19068_n2133_bF_buf4), .B(_abc_19068_n2261), .Y(_abc_19068_n2262) );
  AND2X2 AND2X2_856 ( .A(_abc_19068_n2263), .B(reset_n_bF_buf20), .Y(_abc_19068_n2264) );
  AND2X2 AND2X2_857 ( .A(_abc_19068_n2264), .B(_abc_19068_n2260), .Y(mi1_reg_21__FF_INPUT) );
  AND2X2 AND2X2_858 ( .A(_abc_19068_n2133_bF_buf2), .B(_abc_19068_n2267), .Y(_abc_19068_n2268) );
  AND2X2 AND2X2_859 ( .A(_abc_19068_n2269), .B(reset_n_bF_buf19), .Y(_abc_19068_n2270) );
  AND2X2 AND2X2_86 ( .A(_abc_19068_n899_bF_buf0), .B(word3_reg_3_), .Y(_abc_19068_n1015_1) );
  AND2X2 AND2X2_860 ( .A(_abc_19068_n2270), .B(_abc_19068_n2266), .Y(mi1_reg_22__FF_INPUT) );
  AND2X2 AND2X2_861 ( .A(_abc_19068_n2133_bF_buf0), .B(_abc_19068_n2273), .Y(_abc_19068_n2274) );
  AND2X2 AND2X2_862 ( .A(_abc_19068_n2275), .B(reset_n_bF_buf18), .Y(_abc_19068_n2276) );
  AND2X2 AND2X2_863 ( .A(_abc_19068_n2276), .B(_abc_19068_n2272), .Y(mi1_reg_23__FF_INPUT) );
  AND2X2 AND2X2_864 ( .A(_abc_19068_n2133_bF_buf6), .B(_abc_19068_n2279), .Y(_abc_19068_n2280) );
  AND2X2 AND2X2_865 ( .A(_abc_19068_n2281), .B(reset_n_bF_buf17), .Y(_abc_19068_n2282) );
  AND2X2 AND2X2_866 ( .A(_abc_19068_n2282), .B(_abc_19068_n2278), .Y(mi1_reg_24__FF_INPUT) );
  AND2X2 AND2X2_867 ( .A(_abc_19068_n2133_bF_buf4), .B(_abc_19068_n2285), .Y(_abc_19068_n2286) );
  AND2X2 AND2X2_868 ( .A(_abc_19068_n2287), .B(reset_n_bF_buf16), .Y(_abc_19068_n2288) );
  AND2X2 AND2X2_869 ( .A(_abc_19068_n2288), .B(_abc_19068_n2284), .Y(mi1_reg_25__FF_INPUT) );
  AND2X2 AND2X2_87 ( .A(_abc_19068_n885_1), .B(core_compression_rounds_3_), .Y(_abc_19068_n1019) );
  AND2X2 AND2X2_870 ( .A(_abc_19068_n2133_bF_buf2), .B(_abc_19068_n2291), .Y(_abc_19068_n2292) );
  AND2X2 AND2X2_871 ( .A(_abc_19068_n2293), .B(reset_n_bF_buf15), .Y(_abc_19068_n2294) );
  AND2X2 AND2X2_872 ( .A(_abc_19068_n2294), .B(_abc_19068_n2290), .Y(mi1_reg_26__FF_INPUT) );
  AND2X2 AND2X2_873 ( .A(_abc_19068_n2133_bF_buf0), .B(_abc_19068_n2297), .Y(_abc_19068_n2298) );
  AND2X2 AND2X2_874 ( .A(_abc_19068_n2299), .B(reset_n_bF_buf14), .Y(_abc_19068_n2300) );
  AND2X2 AND2X2_875 ( .A(_abc_19068_n2300), .B(_abc_19068_n2296), .Y(mi1_reg_27__FF_INPUT) );
  AND2X2 AND2X2_876 ( .A(_abc_19068_n2133_bF_buf6), .B(_abc_19068_n2303), .Y(_abc_19068_n2304) );
  AND2X2 AND2X2_877 ( .A(_abc_19068_n2305), .B(reset_n_bF_buf13), .Y(_abc_19068_n2306) );
  AND2X2 AND2X2_878 ( .A(_abc_19068_n2306), .B(_abc_19068_n2302), .Y(mi1_reg_28__FF_INPUT) );
  AND2X2 AND2X2_879 ( .A(_abc_19068_n2133_bF_buf4), .B(_abc_19068_n2309), .Y(_abc_19068_n2310) );
  AND2X2 AND2X2_88 ( .A(_abc_19068_n926_bF_buf1), .B(core_key_3_), .Y(_abc_19068_n1020_1) );
  AND2X2 AND2X2_880 ( .A(_abc_19068_n2311), .B(reset_n_bF_buf12), .Y(_abc_19068_n2312) );
  AND2X2 AND2X2_881 ( .A(_abc_19068_n2312), .B(_abc_19068_n2308), .Y(mi1_reg_29__FF_INPUT) );
  AND2X2 AND2X2_882 ( .A(_abc_19068_n2133_bF_buf2), .B(_abc_19068_n2315), .Y(_abc_19068_n2316) );
  AND2X2 AND2X2_883 ( .A(_abc_19068_n2317), .B(reset_n_bF_buf11), .Y(_abc_19068_n2318) );
  AND2X2 AND2X2_884 ( .A(_abc_19068_n2318), .B(_abc_19068_n2314), .Y(mi1_reg_30__FF_INPUT) );
  AND2X2 AND2X2_885 ( .A(_abc_19068_n2133_bF_buf0), .B(_abc_19068_n2321), .Y(_abc_19068_n2322) );
  AND2X2 AND2X2_886 ( .A(_abc_19068_n2323), .B(reset_n_bF_buf10), .Y(_abc_19068_n2324) );
  AND2X2 AND2X2_887 ( .A(_abc_19068_n2324), .B(_abc_19068_n2320), .Y(mi1_reg_31__FF_INPUT) );
  AND2X2 AND2X2_888 ( .A(_abc_19068_n945_1_bF_buf2), .B(_abc_19068_n2132), .Y(_abc_19068_n2326) );
  AND2X2 AND2X2_889 ( .A(_abc_19068_n2326_bF_buf6), .B(_abc_19068_n2135), .Y(_abc_19068_n2328) );
  AND2X2 AND2X2_89 ( .A(_abc_19068_n924_1_bF_buf1), .B(core_key_35_), .Y(_abc_19068_n1022) );
  AND2X2 AND2X2_890 ( .A(_abc_19068_n2329), .B(reset_n_bF_buf9), .Y(_abc_19068_n2330) );
  AND2X2 AND2X2_891 ( .A(_abc_19068_n2330), .B(_abc_19068_n2327), .Y(mi0_reg_0__FF_INPUT) );
  AND2X2 AND2X2_892 ( .A(_abc_19068_n2326_bF_buf4), .B(_abc_19068_n2141), .Y(_abc_19068_n2333) );
  AND2X2 AND2X2_893 ( .A(_abc_19068_n2334), .B(reset_n_bF_buf8), .Y(_abc_19068_n2335) );
  AND2X2 AND2X2_894 ( .A(_abc_19068_n2335), .B(_abc_19068_n2332), .Y(mi0_reg_1__FF_INPUT) );
  AND2X2 AND2X2_895 ( .A(_abc_19068_n2326_bF_buf2), .B(_abc_19068_n2147), .Y(_abc_19068_n2338) );
  AND2X2 AND2X2_896 ( .A(_abc_19068_n2339), .B(reset_n_bF_buf7), .Y(_abc_19068_n2340) );
  AND2X2 AND2X2_897 ( .A(_abc_19068_n2340), .B(_abc_19068_n2337), .Y(mi0_reg_2__FF_INPUT) );
  AND2X2 AND2X2_898 ( .A(_abc_19068_n2326_bF_buf0), .B(_abc_19068_n2153), .Y(_abc_19068_n2343) );
  AND2X2 AND2X2_899 ( .A(_abc_19068_n2344), .B(reset_n_bF_buf6), .Y(_abc_19068_n2345) );
  AND2X2 AND2X2_9 ( .A(_abc_19068_n871_1), .B(_abc_19068_n883_1), .Y(_abc_19068_n884) );
  AND2X2 AND2X2_90 ( .A(_abc_19068_n939_1_bF_buf1), .B(core_key_67_), .Y(_abc_19068_n1023_1) );
  AND2X2 AND2X2_900 ( .A(_abc_19068_n2345), .B(_abc_19068_n2342), .Y(mi0_reg_3__FF_INPUT) );
  AND2X2 AND2X2_901 ( .A(_abc_19068_n2326_bF_buf6), .B(_abc_19068_n2159), .Y(_abc_19068_n2348) );
  AND2X2 AND2X2_902 ( .A(_abc_19068_n2349), .B(reset_n_bF_buf5), .Y(_abc_19068_n2350) );
  AND2X2 AND2X2_903 ( .A(_abc_19068_n2350), .B(_abc_19068_n2347), .Y(mi0_reg_4__FF_INPUT) );
  AND2X2 AND2X2_904 ( .A(_abc_19068_n2326_bF_buf4), .B(_abc_19068_n2165), .Y(_abc_19068_n2353) );
  AND2X2 AND2X2_905 ( .A(_abc_19068_n2354), .B(reset_n_bF_buf4), .Y(_abc_19068_n2355) );
  AND2X2 AND2X2_906 ( .A(_abc_19068_n2355), .B(_abc_19068_n2352), .Y(mi0_reg_5__FF_INPUT) );
  AND2X2 AND2X2_907 ( .A(_abc_19068_n2326_bF_buf2), .B(_abc_19068_n2171), .Y(_abc_19068_n2358) );
  AND2X2 AND2X2_908 ( .A(_abc_19068_n2359), .B(reset_n_bF_buf3), .Y(_abc_19068_n2360) );
  AND2X2 AND2X2_909 ( .A(_abc_19068_n2360), .B(_abc_19068_n2357), .Y(mi0_reg_6__FF_INPUT) );
  AND2X2 AND2X2_91 ( .A(_abc_19068_n923_bF_buf1), .B(_abc_19068_n1026_1), .Y(_auto_iopadmap_cc_313_execute_30317_3_) );
  AND2X2 AND2X2_910 ( .A(_abc_19068_n2326_bF_buf0), .B(_abc_19068_n2177), .Y(_abc_19068_n2363) );
  AND2X2 AND2X2_911 ( .A(_abc_19068_n2364), .B(reset_n_bF_buf2), .Y(_abc_19068_n2365) );
  AND2X2 AND2X2_912 ( .A(_abc_19068_n2365), .B(_abc_19068_n2362), .Y(mi0_reg_7__FF_INPUT) );
  AND2X2 AND2X2_913 ( .A(_abc_19068_n2326_bF_buf6), .B(_abc_19068_n2183), .Y(_abc_19068_n2368) );
  AND2X2 AND2X2_914 ( .A(_abc_19068_n2369), .B(reset_n_bF_buf1), .Y(_abc_19068_n2370) );
  AND2X2 AND2X2_915 ( .A(_abc_19068_n2370), .B(_abc_19068_n2367), .Y(mi0_reg_8__FF_INPUT) );
  AND2X2 AND2X2_916 ( .A(_abc_19068_n2326_bF_buf4), .B(_abc_19068_n2189), .Y(_abc_19068_n2373) );
  AND2X2 AND2X2_917 ( .A(_abc_19068_n2374), .B(reset_n_bF_buf0), .Y(_abc_19068_n2375) );
  AND2X2 AND2X2_918 ( .A(_abc_19068_n2375), .B(_abc_19068_n2372), .Y(mi0_reg_9__FF_INPUT) );
  AND2X2 AND2X2_919 ( .A(_abc_19068_n2326_bF_buf2), .B(_abc_19068_n2195), .Y(_abc_19068_n2378) );
  AND2X2 AND2X2_92 ( .A(_abc_19068_n897_1_bF_buf4), .B(word0_reg_4_), .Y(_abc_19068_n1028) );
  AND2X2 AND2X2_920 ( .A(_abc_19068_n2379), .B(reset_n_bF_buf84), .Y(_abc_19068_n2380) );
  AND2X2 AND2X2_921 ( .A(_abc_19068_n2380), .B(_abc_19068_n2377), .Y(mi0_reg_10__FF_INPUT) );
  AND2X2 AND2X2_922 ( .A(_abc_19068_n2326_bF_buf0), .B(_abc_19068_n2201), .Y(_abc_19068_n2383) );
  AND2X2 AND2X2_923 ( .A(_abc_19068_n2384), .B(reset_n_bF_buf83), .Y(_abc_19068_n2385) );
  AND2X2 AND2X2_924 ( .A(_abc_19068_n2385), .B(_abc_19068_n2382), .Y(mi0_reg_11__FF_INPUT) );
  AND2X2 AND2X2_925 ( .A(_abc_19068_n2326_bF_buf6), .B(_abc_19068_n2207), .Y(_abc_19068_n2388) );
  AND2X2 AND2X2_926 ( .A(_abc_19068_n2389), .B(reset_n_bF_buf82), .Y(_abc_19068_n2390) );
  AND2X2 AND2X2_927 ( .A(_abc_19068_n2390), .B(_abc_19068_n2387), .Y(mi0_reg_12__FF_INPUT) );
  AND2X2 AND2X2_928 ( .A(_abc_19068_n2326_bF_buf4), .B(_abc_19068_n2213), .Y(_abc_19068_n2393) );
  AND2X2 AND2X2_929 ( .A(_abc_19068_n2394), .B(reset_n_bF_buf81), .Y(_abc_19068_n2395) );
  AND2X2 AND2X2_93 ( .A(_abc_19068_n915_1_bF_buf4), .B(core_mi_36_), .Y(_abc_19068_n1029_1) );
  AND2X2 AND2X2_930 ( .A(_abc_19068_n2395), .B(_abc_19068_n2392), .Y(mi0_reg_13__FF_INPUT) );
  AND2X2 AND2X2_931 ( .A(_abc_19068_n2326_bF_buf2), .B(_abc_19068_n2219), .Y(_abc_19068_n2398) );
  AND2X2 AND2X2_932 ( .A(_abc_19068_n2399), .B(reset_n_bF_buf80), .Y(_abc_19068_n2400) );
  AND2X2 AND2X2_933 ( .A(_abc_19068_n2400), .B(_abc_19068_n2397), .Y(mi0_reg_14__FF_INPUT) );
  AND2X2 AND2X2_934 ( .A(_abc_19068_n2326_bF_buf0), .B(_abc_19068_n2225), .Y(_abc_19068_n2403) );
  AND2X2 AND2X2_935 ( .A(_abc_19068_n2404), .B(reset_n_bF_buf79), .Y(_abc_19068_n2405) );
  AND2X2 AND2X2_936 ( .A(_abc_19068_n2405), .B(_abc_19068_n2402), .Y(mi0_reg_15__FF_INPUT) );
  AND2X2 AND2X2_937 ( .A(_abc_19068_n2326_bF_buf6), .B(_abc_19068_n2231), .Y(_abc_19068_n2408) );
  AND2X2 AND2X2_938 ( .A(_abc_19068_n2409), .B(reset_n_bF_buf78), .Y(_abc_19068_n2410) );
  AND2X2 AND2X2_939 ( .A(_abc_19068_n2410), .B(_abc_19068_n2407), .Y(mi0_reg_16__FF_INPUT) );
  AND2X2 AND2X2_94 ( .A(_abc_19068_n945_1_bF_buf0), .B(core_mi_4_), .Y(_abc_19068_n1031) );
  AND2X2 AND2X2_940 ( .A(_abc_19068_n2326_bF_buf4), .B(_abc_19068_n2237), .Y(_abc_19068_n2413) );
  AND2X2 AND2X2_941 ( .A(_abc_19068_n2414), .B(reset_n_bF_buf77), .Y(_abc_19068_n2415) );
  AND2X2 AND2X2_942 ( .A(_abc_19068_n2415), .B(_abc_19068_n2412), .Y(mi0_reg_17__FF_INPUT) );
  AND2X2 AND2X2_943 ( .A(_abc_19068_n2326_bF_buf2), .B(_abc_19068_n2243), .Y(_abc_19068_n2418) );
  AND2X2 AND2X2_944 ( .A(_abc_19068_n2419), .B(reset_n_bF_buf76), .Y(_abc_19068_n2420) );
  AND2X2 AND2X2_945 ( .A(_abc_19068_n2420), .B(_abc_19068_n2417), .Y(mi0_reg_18__FF_INPUT) );
  AND2X2 AND2X2_946 ( .A(_abc_19068_n2326_bF_buf0), .B(_abc_19068_n2249), .Y(_abc_19068_n2423) );
  AND2X2 AND2X2_947 ( .A(_abc_19068_n2424), .B(reset_n_bF_buf75), .Y(_abc_19068_n2425) );
  AND2X2 AND2X2_948 ( .A(_abc_19068_n2425), .B(_abc_19068_n2422), .Y(mi0_reg_19__FF_INPUT) );
  AND2X2 AND2X2_949 ( .A(_abc_19068_n2326_bF_buf6), .B(_abc_19068_n2255), .Y(_abc_19068_n2428) );
  AND2X2 AND2X2_95 ( .A(_abc_19068_n941_bF_buf0), .B(core_key_100_), .Y(_abc_19068_n1032_1) );
  AND2X2 AND2X2_950 ( .A(_abc_19068_n2429), .B(reset_n_bF_buf74), .Y(_abc_19068_n2430) );
  AND2X2 AND2X2_951 ( .A(_abc_19068_n2430), .B(_abc_19068_n2427), .Y(mi0_reg_20__FF_INPUT) );
  AND2X2 AND2X2_952 ( .A(_abc_19068_n2326_bF_buf4), .B(_abc_19068_n2261), .Y(_abc_19068_n2433) );
  AND2X2 AND2X2_953 ( .A(_abc_19068_n2434), .B(reset_n_bF_buf73), .Y(_abc_19068_n2435) );
  AND2X2 AND2X2_954 ( .A(_abc_19068_n2435), .B(_abc_19068_n2432), .Y(mi0_reg_21__FF_INPUT) );
  AND2X2 AND2X2_955 ( .A(_abc_19068_n2326_bF_buf2), .B(_abc_19068_n2267), .Y(_abc_19068_n2438) );
  AND2X2 AND2X2_956 ( .A(_abc_19068_n2439), .B(reset_n_bF_buf72), .Y(_abc_19068_n2440) );
  AND2X2 AND2X2_957 ( .A(_abc_19068_n2440), .B(_abc_19068_n2437), .Y(mi0_reg_22__FF_INPUT) );
  AND2X2 AND2X2_958 ( .A(_abc_19068_n2326_bF_buf0), .B(_abc_19068_n2273), .Y(_abc_19068_n2443) );
  AND2X2 AND2X2_959 ( .A(_abc_19068_n2444), .B(reset_n_bF_buf71), .Y(_abc_19068_n2445) );
  AND2X2 AND2X2_96 ( .A(_abc_19068_n916_1_bF_buf4), .B(word1_reg_4_), .Y(_abc_19068_n1035_1) );
  AND2X2 AND2X2_960 ( .A(_abc_19068_n2445), .B(_abc_19068_n2442), .Y(mi0_reg_23__FF_INPUT) );
  AND2X2 AND2X2_961 ( .A(_abc_19068_n2326_bF_buf6), .B(_abc_19068_n2279), .Y(_abc_19068_n2448) );
  AND2X2 AND2X2_962 ( .A(_abc_19068_n2449), .B(reset_n_bF_buf70), .Y(_abc_19068_n2450) );
  AND2X2 AND2X2_963 ( .A(_abc_19068_n2450), .B(_abc_19068_n2447), .Y(mi0_reg_24__FF_INPUT) );
  AND2X2 AND2X2_964 ( .A(_abc_19068_n2326_bF_buf4), .B(_abc_19068_n2285), .Y(_abc_19068_n2453) );
  AND2X2 AND2X2_965 ( .A(_abc_19068_n2454), .B(reset_n_bF_buf69), .Y(_abc_19068_n2455) );
  AND2X2 AND2X2_966 ( .A(_abc_19068_n2455), .B(_abc_19068_n2452), .Y(mi0_reg_25__FF_INPUT) );
  AND2X2 AND2X2_967 ( .A(_abc_19068_n2326_bF_buf2), .B(_abc_19068_n2291), .Y(_abc_19068_n2458) );
  AND2X2 AND2X2_968 ( .A(_abc_19068_n2459), .B(reset_n_bF_buf68), .Y(_abc_19068_n2460) );
  AND2X2 AND2X2_969 ( .A(_abc_19068_n2460), .B(_abc_19068_n2457), .Y(mi0_reg_26__FF_INPUT) );
  AND2X2 AND2X2_97 ( .A(_abc_19068_n902_bF_buf4), .B(word2_reg_4_), .Y(_abc_19068_n1036_1) );
  AND2X2 AND2X2_970 ( .A(_abc_19068_n2326_bF_buf0), .B(_abc_19068_n2297), .Y(_abc_19068_n2463) );
  AND2X2 AND2X2_971 ( .A(_abc_19068_n2464), .B(reset_n_bF_buf67), .Y(_abc_19068_n2465) );
  AND2X2 AND2X2_972 ( .A(_abc_19068_n2465), .B(_abc_19068_n2462), .Y(mi0_reg_27__FF_INPUT) );
  AND2X2 AND2X2_973 ( .A(_abc_19068_n2326_bF_buf6), .B(_abc_19068_n2303), .Y(_abc_19068_n2468) );
  AND2X2 AND2X2_974 ( .A(_abc_19068_n2469), .B(reset_n_bF_buf66), .Y(_abc_19068_n2470) );
  AND2X2 AND2X2_975 ( .A(_abc_19068_n2470), .B(_abc_19068_n2467), .Y(mi0_reg_28__FF_INPUT) );
  AND2X2 AND2X2_976 ( .A(_abc_19068_n2326_bF_buf4), .B(_abc_19068_n2309), .Y(_abc_19068_n2473) );
  AND2X2 AND2X2_977 ( .A(_abc_19068_n2474), .B(reset_n_bF_buf65), .Y(_abc_19068_n2475) );
  AND2X2 AND2X2_978 ( .A(_abc_19068_n2475), .B(_abc_19068_n2472), .Y(mi0_reg_29__FF_INPUT) );
  AND2X2 AND2X2_979 ( .A(_abc_19068_n2326_bF_buf2), .B(_abc_19068_n2315), .Y(_abc_19068_n2478) );
  AND2X2 AND2X2_98 ( .A(_abc_19068_n881), .B(_abc_19068_n901_1), .Y(_abc_19068_n1038_1) );
  AND2X2 AND2X2_980 ( .A(_abc_19068_n2479), .B(reset_n_bF_buf64), .Y(_abc_19068_n2480) );
  AND2X2 AND2X2_981 ( .A(_abc_19068_n2480), .B(_abc_19068_n2477), .Y(mi0_reg_30__FF_INPUT) );
  AND2X2 AND2X2_982 ( .A(_abc_19068_n2326_bF_buf0), .B(_abc_19068_n2321), .Y(_abc_19068_n2483) );
  AND2X2 AND2X2_983 ( .A(_abc_19068_n2484), .B(reset_n_bF_buf63), .Y(_abc_19068_n2485) );
  AND2X2 AND2X2_984 ( .A(_abc_19068_n2485), .B(_abc_19068_n2482), .Y(mi0_reg_31__FF_INPUT) );
  AND2X2 AND2X2_985 ( .A(_abc_19068_n941_bF_buf2), .B(_abc_19068_n2132), .Y(_abc_19068_n2487) );
  AND2X2 AND2X2_986 ( .A(_abc_19068_n2487_bF_buf6), .B(_abc_19068_n2135), .Y(_abc_19068_n2489) );
  AND2X2 AND2X2_987 ( .A(_abc_19068_n2490), .B(reset_n_bF_buf62), .Y(_abc_19068_n2491) );
  AND2X2 AND2X2_988 ( .A(_abc_19068_n2491), .B(_abc_19068_n2488), .Y(key3_reg_0__FF_INPUT) );
  AND2X2 AND2X2_989 ( .A(_abc_19068_n2487_bF_buf4), .B(_abc_19068_n2141), .Y(_abc_19068_n2494) );
  AND2X2 AND2X2_99 ( .A(_abc_19068_n899_bF_buf4), .B(word3_reg_4_), .Y(_abc_19068_n1039_1) );
  AND2X2 AND2X2_990 ( .A(_abc_19068_n2495), .B(reset_n_bF_buf61), .Y(_abc_19068_n2496) );
  AND2X2 AND2X2_991 ( .A(_abc_19068_n2496), .B(_abc_19068_n2493), .Y(key3_reg_1__FF_INPUT) );
  AND2X2 AND2X2_992 ( .A(_abc_19068_n2487_bF_buf2), .B(_abc_19068_n2147), .Y(_abc_19068_n2499) );
  AND2X2 AND2X2_993 ( .A(_abc_19068_n2500), .B(reset_n_bF_buf60), .Y(_abc_19068_n2501) );
  AND2X2 AND2X2_994 ( .A(_abc_19068_n2501), .B(_abc_19068_n2498), .Y(key3_reg_2__FF_INPUT) );
  AND2X2 AND2X2_995 ( .A(_abc_19068_n2487_bF_buf0), .B(_abc_19068_n2153), .Y(_abc_19068_n2504) );
  AND2X2 AND2X2_996 ( .A(_abc_19068_n2505), .B(reset_n_bF_buf59), .Y(_abc_19068_n2506) );
  AND2X2 AND2X2_997 ( .A(_abc_19068_n2506), .B(_abc_19068_n2503), .Y(key3_reg_3__FF_INPUT) );
  AND2X2 AND2X2_998 ( .A(_abc_19068_n2487_bF_buf6), .B(_abc_19068_n2159), .Y(_abc_19068_n2509) );
  AND2X2 AND2X2_999 ( .A(_abc_19068_n2510), .B(reset_n_bF_buf58), .Y(_abc_19068_n2511) );
  BUFX2 BUFX2_1 ( .A(clk), .Y(clk_hier0_bF_buf8) );
  BUFX2 BUFX2_10 ( .A(reset_n), .Y(reset_n_hier0_bF_buf8) );
  BUFX2 BUFX2_100 ( .A(core__abc_21380_n2451_1), .Y(core__abc_21380_n2451_1_bF_buf3) );
  BUFX2 BUFX2_101 ( .A(core__abc_21380_n2451_1), .Y(core__abc_21380_n2451_1_bF_buf2) );
  BUFX2 BUFX2_102 ( .A(core__abc_21380_n2451_1), .Y(core__abc_21380_n2451_1_bF_buf1) );
  BUFX2 BUFX2_103 ( .A(core__abc_21380_n2451_1), .Y(core__abc_21380_n2451_1_bF_buf0) );
  BUFX2 BUFX2_104 ( .A(core__abc_21380_n7076), .Y(core__abc_21380_n7076_bF_buf6) );
  BUFX2 BUFX2_105 ( .A(core__abc_21380_n7076), .Y(core__abc_21380_n7076_bF_buf5) );
  BUFX2 BUFX2_106 ( .A(core__abc_21380_n7076), .Y(core__abc_21380_n7076_bF_buf4) );
  BUFX2 BUFX2_107 ( .A(core__abc_21380_n7076), .Y(core__abc_21380_n7076_bF_buf3) );
  BUFX2 BUFX2_108 ( .A(core__abc_21380_n7076), .Y(core__abc_21380_n7076_bF_buf2) );
  BUFX2 BUFX2_109 ( .A(core__abc_21380_n7076), .Y(core__abc_21380_n7076_bF_buf1) );
  BUFX2 BUFX2_11 ( .A(reset_n), .Y(reset_n_hier0_bF_buf7) );
  BUFX2 BUFX2_110 ( .A(core__abc_21380_n7076), .Y(core__abc_21380_n7076_bF_buf0) );
  BUFX2 BUFX2_111 ( .A(core__abc_21380_n1134_1), .Y(core__abc_21380_n1134_1_bF_buf7) );
  BUFX2 BUFX2_112 ( .A(core__abc_21380_n1134_1), .Y(core__abc_21380_n1134_1_bF_buf6) );
  BUFX2 BUFX2_113 ( .A(core__abc_21380_n1134_1), .Y(core__abc_21380_n1134_1_bF_buf5) );
  BUFX2 BUFX2_114 ( .A(core__abc_21380_n1134_1), .Y(core__abc_21380_n1134_1_bF_buf4) );
  BUFX2 BUFX2_115 ( .A(core__abc_21380_n1134_1), .Y(core__abc_21380_n1134_1_bF_buf3) );
  BUFX2 BUFX2_116 ( .A(core__abc_21380_n1134_1), .Y(core__abc_21380_n1134_1_bF_buf2) );
  BUFX2 BUFX2_117 ( .A(core__abc_21380_n1134_1), .Y(core__abc_21380_n1134_1_bF_buf1) );
  BUFX2 BUFX2_118 ( .A(core__abc_21380_n1134_1), .Y(core__abc_21380_n1134_1_bF_buf0) );
  BUFX2 BUFX2_119 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf84) );
  BUFX2 BUFX2_12 ( .A(reset_n), .Y(reset_n_hier0_bF_buf6) );
  BUFX2 BUFX2_120 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf83) );
  BUFX2 BUFX2_121 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf82) );
  BUFX2 BUFX2_122 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf81) );
  BUFX2 BUFX2_123 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf80) );
  BUFX2 BUFX2_124 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf79) );
  BUFX2 BUFX2_125 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf78) );
  BUFX2 BUFX2_126 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf77) );
  BUFX2 BUFX2_127 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf76) );
  BUFX2 BUFX2_128 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf75) );
  BUFX2 BUFX2_129 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf74) );
  BUFX2 BUFX2_13 ( .A(reset_n), .Y(reset_n_hier0_bF_buf5) );
  BUFX2 BUFX2_130 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf73) );
  BUFX2 BUFX2_131 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf72) );
  BUFX2 BUFX2_132 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf71) );
  BUFX2 BUFX2_133 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf70) );
  BUFX2 BUFX2_134 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf69) );
  BUFX2 BUFX2_135 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf68) );
  BUFX2 BUFX2_136 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf67) );
  BUFX2 BUFX2_137 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf66) );
  BUFX2 BUFX2_138 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf65) );
  BUFX2 BUFX2_139 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf64) );
  BUFX2 BUFX2_14 ( .A(reset_n), .Y(reset_n_hier0_bF_buf4) );
  BUFX2 BUFX2_140 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf63) );
  BUFX2 BUFX2_141 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf62) );
  BUFX2 BUFX2_142 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf61) );
  BUFX2 BUFX2_143 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf60) );
  BUFX2 BUFX2_144 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf59) );
  BUFX2 BUFX2_145 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf58) );
  BUFX2 BUFX2_146 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf57) );
  BUFX2 BUFX2_147 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf56) );
  BUFX2 BUFX2_148 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf55) );
  BUFX2 BUFX2_149 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf54) );
  BUFX2 BUFX2_15 ( .A(reset_n), .Y(reset_n_hier0_bF_buf3) );
  BUFX2 BUFX2_150 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf53) );
  BUFX2 BUFX2_151 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf52) );
  BUFX2 BUFX2_152 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf51) );
  BUFX2 BUFX2_153 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf50) );
  BUFX2 BUFX2_154 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf49) );
  BUFX2 BUFX2_155 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf48) );
  BUFX2 BUFX2_156 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf47) );
  BUFX2 BUFX2_157 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf46) );
  BUFX2 BUFX2_158 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf45) );
  BUFX2 BUFX2_159 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf44) );
  BUFX2 BUFX2_16 ( .A(reset_n), .Y(reset_n_hier0_bF_buf2) );
  BUFX2 BUFX2_160 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf43) );
  BUFX2 BUFX2_161 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf42) );
  BUFX2 BUFX2_162 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf41) );
  BUFX2 BUFX2_163 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf40) );
  BUFX2 BUFX2_164 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf39) );
  BUFX2 BUFX2_165 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf38) );
  BUFX2 BUFX2_166 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf37) );
  BUFX2 BUFX2_167 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf36) );
  BUFX2 BUFX2_168 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf35) );
  BUFX2 BUFX2_169 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf34) );
  BUFX2 BUFX2_17 ( .A(reset_n), .Y(reset_n_hier0_bF_buf1) );
  BUFX2 BUFX2_170 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf33) );
  BUFX2 BUFX2_171 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf32) );
  BUFX2 BUFX2_172 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf31) );
  BUFX2 BUFX2_173 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf30) );
  BUFX2 BUFX2_174 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf29) );
  BUFX2 BUFX2_175 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf28) );
  BUFX2 BUFX2_176 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf27) );
  BUFX2 BUFX2_177 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf26) );
  BUFX2 BUFX2_178 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf25) );
  BUFX2 BUFX2_179 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf24) );
  BUFX2 BUFX2_18 ( .A(reset_n), .Y(reset_n_hier0_bF_buf0) );
  BUFX2 BUFX2_180 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf23) );
  BUFX2 BUFX2_181 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf22) );
  BUFX2 BUFX2_182 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf21) );
  BUFX2 BUFX2_183 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf20) );
  BUFX2 BUFX2_184 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf19) );
  BUFX2 BUFX2_185 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf18) );
  BUFX2 BUFX2_186 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf17) );
  BUFX2 BUFX2_187 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf16) );
  BUFX2 BUFX2_188 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf15) );
  BUFX2 BUFX2_189 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf14) );
  BUFX2 BUFX2_19 ( .A(core__abc_21380_n3167_1_bF_buf14), .Y(core__abc_21380_n3167_1_bF_buf14_bF_buf3) );
  BUFX2 BUFX2_190 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf13) );
  BUFX2 BUFX2_191 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf12) );
  BUFX2 BUFX2_192 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf11) );
  BUFX2 BUFX2_193 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf10) );
  BUFX2 BUFX2_194 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf9) );
  BUFX2 BUFX2_195 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf8) );
  BUFX2 BUFX2_196 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf7) );
  BUFX2 BUFX2_197 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf6) );
  BUFX2 BUFX2_198 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf5) );
  BUFX2 BUFX2_199 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf4) );
  BUFX2 BUFX2_2 ( .A(clk), .Y(clk_hier0_bF_buf7) );
  BUFX2 BUFX2_20 ( .A(core__abc_21380_n3167_1_bF_buf14), .Y(core__abc_21380_n3167_1_bF_buf14_bF_buf2) );
  BUFX2 BUFX2_200 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf3) );
  BUFX2 BUFX2_201 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf2) );
  BUFX2 BUFX2_202 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf1) );
  BUFX2 BUFX2_203 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf0) );
  BUFX2 BUFX2_204 ( .A(core__abc_21380_n9245), .Y(core__abc_21380_n9245_bF_buf7) );
  BUFX2 BUFX2_205 ( .A(core__abc_21380_n9245), .Y(core__abc_21380_n9245_bF_buf6) );
  BUFX2 BUFX2_206 ( .A(core__abc_21380_n9245), .Y(core__abc_21380_n9245_bF_buf5) );
  BUFX2 BUFX2_207 ( .A(core__abc_21380_n9245), .Y(core__abc_21380_n9245_bF_buf4) );
  BUFX2 BUFX2_208 ( .A(core__abc_21380_n9245), .Y(core__abc_21380_n9245_bF_buf3) );
  BUFX2 BUFX2_209 ( .A(core__abc_21380_n9245), .Y(core__abc_21380_n9245_bF_buf2) );
  BUFX2 BUFX2_21 ( .A(core__abc_21380_n3167_1_bF_buf14), .Y(core__abc_21380_n3167_1_bF_buf14_bF_buf1) );
  BUFX2 BUFX2_210 ( .A(core__abc_21380_n9245), .Y(core__abc_21380_n9245_bF_buf1) );
  BUFX2 BUFX2_211 ( .A(core__abc_21380_n9245), .Y(core__abc_21380_n9245_bF_buf0) );
  BUFX2 BUFX2_212 ( .A(core__abc_21380_n9246), .Y(core__abc_21380_n9246_bF_buf7) );
  BUFX2 BUFX2_213 ( .A(core__abc_21380_n9246), .Y(core__abc_21380_n9246_bF_buf6) );
  BUFX2 BUFX2_214 ( .A(core__abc_21380_n9246), .Y(core__abc_21380_n9246_bF_buf5) );
  BUFX2 BUFX2_215 ( .A(core__abc_21380_n9246), .Y(core__abc_21380_n9246_bF_buf4) );
  BUFX2 BUFX2_216 ( .A(core__abc_21380_n9246), .Y(core__abc_21380_n9246_bF_buf3) );
  BUFX2 BUFX2_217 ( .A(core__abc_21380_n9246), .Y(core__abc_21380_n9246_bF_buf2) );
  BUFX2 BUFX2_218 ( .A(core__abc_21380_n9246), .Y(core__abc_21380_n9246_bF_buf1) );
  BUFX2 BUFX2_219 ( .A(core__abc_21380_n9246), .Y(core__abc_21380_n9246_bF_buf0) );
  BUFX2 BUFX2_22 ( .A(core__abc_21380_n3167_1_bF_buf14), .Y(core__abc_21380_n3167_1_bF_buf14_bF_buf0) );
  BUFX2 BUFX2_220 ( .A(core__abc_21380_n9248), .Y(core__abc_21380_n9248_bF_buf7) );
  BUFX2 BUFX2_221 ( .A(core__abc_21380_n9248), .Y(core__abc_21380_n9248_bF_buf6) );
  BUFX2 BUFX2_222 ( .A(core__abc_21380_n9248), .Y(core__abc_21380_n9248_bF_buf5) );
  BUFX2 BUFX2_223 ( .A(core__abc_21380_n9248), .Y(core__abc_21380_n9248_bF_buf4) );
  BUFX2 BUFX2_224 ( .A(core__abc_21380_n9248), .Y(core__abc_21380_n9248_bF_buf3) );
  BUFX2 BUFX2_225 ( .A(core__abc_21380_n9248), .Y(core__abc_21380_n9248_bF_buf2) );
  BUFX2 BUFX2_226 ( .A(core__abc_21380_n9248), .Y(core__abc_21380_n9248_bF_buf1) );
  BUFX2 BUFX2_227 ( .A(core__abc_21380_n9248), .Y(core__abc_21380_n9248_bF_buf0) );
  BUFX2 BUFX2_228 ( .A(_abc_19068_n2326), .Y(_abc_19068_n2326_bF_buf7) );
  BUFX2 BUFX2_229 ( .A(_abc_19068_n2326), .Y(_abc_19068_n2326_bF_buf6) );
  BUFX2 BUFX2_23 ( .A(core__abc_21380_n3167_1_bF_buf15), .Y(core__abc_21380_n3167_1_bF_buf15_bF_buf3) );
  BUFX2 BUFX2_230 ( .A(_abc_19068_n2326), .Y(_abc_19068_n2326_bF_buf5) );
  BUFX2 BUFX2_231 ( .A(_abc_19068_n2326), .Y(_abc_19068_n2326_bF_buf4) );
  BUFX2 BUFX2_232 ( .A(_abc_19068_n2326), .Y(_abc_19068_n2326_bF_buf3) );
  BUFX2 BUFX2_233 ( .A(_abc_19068_n2326), .Y(_abc_19068_n2326_bF_buf2) );
  BUFX2 BUFX2_234 ( .A(_abc_19068_n2326), .Y(_abc_19068_n2326_bF_buf1) );
  BUFX2 BUFX2_235 ( .A(_abc_19068_n2326), .Y(_abc_19068_n2326_bF_buf0) );
  BUFX2 BUFX2_236 ( .A(_abc_19068_n902), .Y(_abc_19068_n902_bF_buf4) );
  BUFX2 BUFX2_237 ( .A(_abc_19068_n902), .Y(_abc_19068_n902_bF_buf3) );
  BUFX2 BUFX2_238 ( .A(_abc_19068_n902), .Y(_abc_19068_n902_bF_buf2) );
  BUFX2 BUFX2_239 ( .A(_abc_19068_n902), .Y(_abc_19068_n902_bF_buf1) );
  BUFX2 BUFX2_24 ( .A(core__abc_21380_n3167_1_bF_buf15), .Y(core__abc_21380_n3167_1_bF_buf15_bF_buf2) );
  BUFX2 BUFX2_240 ( .A(_abc_19068_n902), .Y(_abc_19068_n902_bF_buf0) );
  BUFX2 BUFX2_241 ( .A(_abc_19068_n2648), .Y(_abc_19068_n2648_bF_buf7) );
  BUFX2 BUFX2_242 ( .A(_abc_19068_n2648), .Y(_abc_19068_n2648_bF_buf6) );
  BUFX2 BUFX2_243 ( .A(_abc_19068_n2648), .Y(_abc_19068_n2648_bF_buf5) );
  BUFX2 BUFX2_244 ( .A(_abc_19068_n2648), .Y(_abc_19068_n2648_bF_buf4) );
  BUFX2 BUFX2_245 ( .A(_abc_19068_n2648), .Y(_abc_19068_n2648_bF_buf3) );
  BUFX2 BUFX2_246 ( .A(_abc_19068_n2648), .Y(_abc_19068_n2648_bF_buf2) );
  BUFX2 BUFX2_247 ( .A(_abc_19068_n2648), .Y(_abc_19068_n2648_bF_buf1) );
  BUFX2 BUFX2_248 ( .A(_abc_19068_n2648), .Y(_abc_19068_n2648_bF_buf0) );
  BUFX2 BUFX2_249 ( .A(_abc_19068_n945_1), .Y(_abc_19068_n945_1_bF_buf4) );
  BUFX2 BUFX2_25 ( .A(core__abc_21380_n3167_1_bF_buf15), .Y(core__abc_21380_n3167_1_bF_buf15_bF_buf1) );
  BUFX2 BUFX2_250 ( .A(_abc_19068_n945_1), .Y(_abc_19068_n945_1_bF_buf3) );
  BUFX2 BUFX2_251 ( .A(_abc_19068_n945_1), .Y(_abc_19068_n945_1_bF_buf2) );
  BUFX2 BUFX2_252 ( .A(_abc_19068_n945_1), .Y(_abc_19068_n945_1_bF_buf1) );
  BUFX2 BUFX2_253 ( .A(_abc_19068_n945_1), .Y(_abc_19068_n945_1_bF_buf0) );
  BUFX2 BUFX2_254 ( .A(core__abc_21380_n2452), .Y(core__abc_21380_n2452_bF_buf7) );
  BUFX2 BUFX2_255 ( .A(core__abc_21380_n2452), .Y(core__abc_21380_n2452_bF_buf6) );
  BUFX2 BUFX2_256 ( .A(core__abc_21380_n2452), .Y(core__abc_21380_n2452_bF_buf5) );
  BUFX2 BUFX2_257 ( .A(core__abc_21380_n2452), .Y(core__abc_21380_n2452_bF_buf4) );
  BUFX2 BUFX2_258 ( .A(core__abc_21380_n2452), .Y(core__abc_21380_n2452_bF_buf3) );
  BUFX2 BUFX2_259 ( .A(core__abc_21380_n2452), .Y(core__abc_21380_n2452_bF_buf2) );
  BUFX2 BUFX2_26 ( .A(core__abc_21380_n3167_1_bF_buf15), .Y(core__abc_21380_n3167_1_bF_buf15_bF_buf0) );
  BUFX2 BUFX2_260 ( .A(core__abc_21380_n2452), .Y(core__abc_21380_n2452_bF_buf1) );
  BUFX2 BUFX2_261 ( .A(core__abc_21380_n2452), .Y(core__abc_21380_n2452_bF_buf0) );
  BUFX2 BUFX2_262 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf10) );
  BUFX2 BUFX2_263 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf9) );
  BUFX2 BUFX2_264 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf8) );
  BUFX2 BUFX2_265 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf7) );
  BUFX2 BUFX2_266 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf6) );
  BUFX2 BUFX2_267 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf5) );
  BUFX2 BUFX2_268 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf4) );
  BUFX2 BUFX2_269 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf3) );
  BUFX2 BUFX2_27 ( .A(_abc_19068_n916_1), .Y(_abc_19068_n916_1_bF_buf4) );
  BUFX2 BUFX2_270 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf2) );
  BUFX2 BUFX2_271 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf1) );
  BUFX2 BUFX2_272 ( .A(core__abc_21380_n2749), .Y(core__abc_21380_n2749_bF_buf0) );
  BUFX2 BUFX2_273 ( .A(_abc_19068_n915_1), .Y(_abc_19068_n915_1_bF_buf4) );
  BUFX2 BUFX2_274 ( .A(_abc_19068_n915_1), .Y(_abc_19068_n915_1_bF_buf3) );
  BUFX2 BUFX2_275 ( .A(_abc_19068_n915_1), .Y(_abc_19068_n915_1_bF_buf2) );
  BUFX2 BUFX2_276 ( .A(_abc_19068_n915_1), .Y(_abc_19068_n915_1_bF_buf1) );
  BUFX2 BUFX2_277 ( .A(_abc_19068_n915_1), .Y(_abc_19068_n915_1_bF_buf0) );
  BUFX2 BUFX2_278 ( .A(_abc_19068_n897_1), .Y(_abc_19068_n897_1_bF_buf4) );
  BUFX2 BUFX2_279 ( .A(_abc_19068_n897_1), .Y(_abc_19068_n897_1_bF_buf3) );
  BUFX2 BUFX2_28 ( .A(_abc_19068_n916_1), .Y(_abc_19068_n916_1_bF_buf3) );
  BUFX2 BUFX2_280 ( .A(_abc_19068_n897_1), .Y(_abc_19068_n897_1_bF_buf2) );
  BUFX2 BUFX2_281 ( .A(_abc_19068_n897_1), .Y(_abc_19068_n897_1_bF_buf1) );
  BUFX2 BUFX2_282 ( .A(_abc_19068_n897_1), .Y(_abc_19068_n897_1_bF_buf0) );
  BUFX2 BUFX2_283 ( .A(core__abc_21380_n3163_1), .Y(core__abc_21380_n3163_1_bF_buf6) );
  BUFX2 BUFX2_284 ( .A(core__abc_21380_n3163_1), .Y(core__abc_21380_n3163_1_bF_buf5) );
  BUFX2 BUFX2_285 ( .A(core__abc_21380_n3163_1), .Y(core__abc_21380_n3163_1_bF_buf4) );
  BUFX2 BUFX2_286 ( .A(core__abc_21380_n3163_1), .Y(core__abc_21380_n3163_1_bF_buf3) );
  BUFX2 BUFX2_287 ( .A(core__abc_21380_n3163_1), .Y(core__abc_21380_n3163_1_bF_buf2) );
  BUFX2 BUFX2_288 ( .A(core__abc_21380_n3163_1), .Y(core__abc_21380_n3163_1_bF_buf1) );
  BUFX2 BUFX2_289 ( .A(core__abc_21380_n3163_1), .Y(core__abc_21380_n3163_1_bF_buf0) );
  BUFX2 BUFX2_29 ( .A(_abc_19068_n916_1), .Y(_abc_19068_n916_1_bF_buf2) );
  BUFX2 BUFX2_290 ( .A(_abc_19068_n923), .Y(_abc_19068_n923_bF_buf4) );
  BUFX2 BUFX2_291 ( .A(_abc_19068_n923), .Y(_abc_19068_n923_bF_buf3) );
  BUFX2 BUFX2_292 ( .A(_abc_19068_n923), .Y(_abc_19068_n923_bF_buf2) );
  BUFX2 BUFX2_293 ( .A(_abc_19068_n923), .Y(_abc_19068_n923_bF_buf1) );
  BUFX2 BUFX2_294 ( .A(_abc_19068_n923), .Y(_abc_19068_n923_bF_buf0) );
  BUFX2 BUFX2_295 ( .A(_abc_19068_n926), .Y(_abc_19068_n926_bF_buf4) );
  BUFX2 BUFX2_296 ( .A(_abc_19068_n926), .Y(_abc_19068_n926_bF_buf3) );
  BUFX2 BUFX2_297 ( .A(_abc_19068_n926), .Y(_abc_19068_n926_bF_buf2) );
  BUFX2 BUFX2_298 ( .A(_abc_19068_n926), .Y(_abc_19068_n926_bF_buf1) );
  BUFX2 BUFX2_299 ( .A(_abc_19068_n926), .Y(_abc_19068_n926_bF_buf0) );
  BUFX2 BUFX2_3 ( .A(clk), .Y(clk_hier0_bF_buf6) );
  BUFX2 BUFX2_30 ( .A(_abc_19068_n916_1), .Y(_abc_19068_n916_1_bF_buf1) );
  BUFX2 BUFX2_300 ( .A(_abc_19068_n899), .Y(_abc_19068_n899_bF_buf4) );
  BUFX2 BUFX2_301 ( .A(_abc_19068_n899), .Y(_abc_19068_n899_bF_buf3) );
  BUFX2 BUFX2_302 ( .A(_abc_19068_n899), .Y(_abc_19068_n899_bF_buf2) );
  BUFX2 BUFX2_303 ( .A(_abc_19068_n899), .Y(_abc_19068_n899_bF_buf1) );
  BUFX2 BUFX2_304 ( .A(_abc_19068_n899), .Y(_abc_19068_n899_bF_buf0) );
  BUFX2 BUFX2_305 ( .A(_abc_19068_n939_1), .Y(_abc_19068_n939_1_bF_buf4) );
  BUFX2 BUFX2_306 ( .A(_abc_19068_n939_1), .Y(_abc_19068_n939_1_bF_buf3) );
  BUFX2 BUFX2_307 ( .A(_abc_19068_n939_1), .Y(_abc_19068_n939_1_bF_buf2) );
  BUFX2 BUFX2_308 ( .A(_abc_19068_n939_1), .Y(_abc_19068_n939_1_bF_buf1) );
  BUFX2 BUFX2_309 ( .A(_abc_19068_n939_1), .Y(_abc_19068_n939_1_bF_buf0) );
  BUFX2 BUFX2_31 ( .A(_abc_19068_n916_1), .Y(_abc_19068_n916_1_bF_buf0) );
  BUFX2 BUFX2_310 ( .A(core__abc_21380_n3328), .Y(core__abc_21380_n3328_bF_buf7) );
  BUFX2 BUFX2_311 ( .A(core__abc_21380_n3328), .Y(core__abc_21380_n3328_bF_buf6) );
  BUFX2 BUFX2_312 ( .A(core__abc_21380_n3328), .Y(core__abc_21380_n3328_bF_buf5) );
  BUFX2 BUFX2_313 ( .A(core__abc_21380_n3328), .Y(core__abc_21380_n3328_bF_buf4) );
  BUFX2 BUFX2_314 ( .A(core__abc_21380_n3328), .Y(core__abc_21380_n3328_bF_buf3) );
  BUFX2 BUFX2_315 ( .A(core__abc_21380_n3328), .Y(core__abc_21380_n3328_bF_buf2) );
  BUFX2 BUFX2_316 ( .A(core__abc_21380_n3328), .Y(core__abc_21380_n3328_bF_buf1) );
  BUFX2 BUFX2_317 ( .A(core__abc_21380_n3328), .Y(core__abc_21380_n3328_bF_buf0) );
  BUFX2 BUFX2_318 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf7) );
  BUFX2 BUFX2_319 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf6) );
  BUFX2 BUFX2_32 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf10) );
  BUFX2 BUFX2_320 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf5) );
  BUFX2 BUFX2_321 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf4) );
  BUFX2 BUFX2_322 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf3) );
  BUFX2 BUFX2_323 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf2) );
  BUFX2 BUFX2_324 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf1) );
  BUFX2 BUFX2_325 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf0) );
  BUFX2 BUFX2_326 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf84) );
  BUFX2 BUFX2_327 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf83) );
  BUFX2 BUFX2_328 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf82) );
  BUFX2 BUFX2_329 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf81) );
  BUFX2 BUFX2_33 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf9) );
  BUFX2 BUFX2_330 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf80) );
  BUFX2 BUFX2_331 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf79) );
  BUFX2 BUFX2_332 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf78) );
  BUFX2 BUFX2_333 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf77) );
  BUFX2 BUFX2_334 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf76) );
  BUFX2 BUFX2_335 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf75) );
  BUFX2 BUFX2_336 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf74) );
  BUFX2 BUFX2_337 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf73) );
  BUFX2 BUFX2_338 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf72) );
  BUFX2 BUFX2_339 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf71) );
  BUFX2 BUFX2_34 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf8) );
  BUFX2 BUFX2_340 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf70) );
  BUFX2 BUFX2_341 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf69) );
  BUFX2 BUFX2_342 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf68) );
  BUFX2 BUFX2_343 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf67) );
  BUFX2 BUFX2_344 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf66) );
  BUFX2 BUFX2_345 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf65) );
  BUFX2 BUFX2_346 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf64) );
  BUFX2 BUFX2_347 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf63) );
  BUFX2 BUFX2_348 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf62) );
  BUFX2 BUFX2_349 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf61) );
  BUFX2 BUFX2_35 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf7) );
  BUFX2 BUFX2_350 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf60) );
  BUFX2 BUFX2_351 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf59) );
  BUFX2 BUFX2_352 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf58) );
  BUFX2 BUFX2_353 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf57) );
  BUFX2 BUFX2_354 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf56) );
  BUFX2 BUFX2_355 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf55) );
  BUFX2 BUFX2_356 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf54) );
  BUFX2 BUFX2_357 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf53) );
  BUFX2 BUFX2_358 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf52) );
  BUFX2 BUFX2_359 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf51) );
  BUFX2 BUFX2_36 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf6) );
  BUFX2 BUFX2_360 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf50) );
  BUFX2 BUFX2_361 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf49) );
  BUFX2 BUFX2_362 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf48) );
  BUFX2 BUFX2_363 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf47) );
  BUFX2 BUFX2_364 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf46) );
  BUFX2 BUFX2_365 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf45) );
  BUFX2 BUFX2_366 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf44) );
  BUFX2 BUFX2_367 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf43) );
  BUFX2 BUFX2_368 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf42) );
  BUFX2 BUFX2_369 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf41) );
  BUFX2 BUFX2_37 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf5) );
  BUFX2 BUFX2_370 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf40) );
  BUFX2 BUFX2_371 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf39) );
  BUFX2 BUFX2_372 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf38) );
  BUFX2 BUFX2_373 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf37) );
  BUFX2 BUFX2_374 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf36) );
  BUFX2 BUFX2_375 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf35) );
  BUFX2 BUFX2_376 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf34) );
  BUFX2 BUFX2_377 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf33) );
  BUFX2 BUFX2_378 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf32) );
  BUFX2 BUFX2_379 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf31) );
  BUFX2 BUFX2_38 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf4) );
  BUFX2 BUFX2_380 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf30) );
  BUFX2 BUFX2_381 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf29) );
  BUFX2 BUFX2_382 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf28) );
  BUFX2 BUFX2_383 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf27) );
  BUFX2 BUFX2_384 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf26) );
  BUFX2 BUFX2_385 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf25) );
  BUFX2 BUFX2_386 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf24) );
  BUFX2 BUFX2_387 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf23) );
  BUFX2 BUFX2_388 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf22) );
  BUFX2 BUFX2_389 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf21) );
  BUFX2 BUFX2_39 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf3) );
  BUFX2 BUFX2_390 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf20) );
  BUFX2 BUFX2_391 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf19) );
  BUFX2 BUFX2_392 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf18) );
  BUFX2 BUFX2_393 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf17) );
  BUFX2 BUFX2_394 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf16) );
  BUFX2 BUFX2_395 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf15) );
  BUFX2 BUFX2_396 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf14) );
  BUFX2 BUFX2_397 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf13) );
  BUFX2 BUFX2_398 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf12) );
  BUFX2 BUFX2_399 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf11) );
  BUFX2 BUFX2_4 ( .A(clk), .Y(clk_hier0_bF_buf5) );
  BUFX2 BUFX2_40 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf2) );
  BUFX2 BUFX2_400 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf10) );
  BUFX2 BUFX2_401 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf9) );
  BUFX2 BUFX2_402 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf8) );
  BUFX2 BUFX2_403 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf7) );
  BUFX2 BUFX2_404 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf6) );
  BUFX2 BUFX2_405 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf5) );
  BUFX2 BUFX2_406 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf4) );
  BUFX2 BUFX2_407 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf3) );
  BUFX2 BUFX2_408 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf2) );
  BUFX2 BUFX2_409 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf1) );
  BUFX2 BUFX2_41 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf1) );
  BUFX2 BUFX2_410 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf0) );
  BUFX2 BUFX2_411 ( .A(_abc_19068_n2133), .Y(_abc_19068_n2133_bF_buf7) );
  BUFX2 BUFX2_412 ( .A(_abc_19068_n2133), .Y(_abc_19068_n2133_bF_buf6) );
  BUFX2 BUFX2_413 ( .A(_abc_19068_n2133), .Y(_abc_19068_n2133_bF_buf5) );
  BUFX2 BUFX2_414 ( .A(_abc_19068_n2133), .Y(_abc_19068_n2133_bF_buf4) );
  BUFX2 BUFX2_415 ( .A(_abc_19068_n2133), .Y(_abc_19068_n2133_bF_buf3) );
  BUFX2 BUFX2_416 ( .A(_abc_19068_n2133), .Y(_abc_19068_n2133_bF_buf2) );
  BUFX2 BUFX2_417 ( .A(_abc_19068_n2133), .Y(_abc_19068_n2133_bF_buf1) );
  BUFX2 BUFX2_418 ( .A(_abc_19068_n2133), .Y(_abc_19068_n2133_bF_buf0) );
  BUFX2 BUFX2_419 ( .A(_abc_19068_n2487), .Y(_abc_19068_n2487_bF_buf7) );
  BUFX2 BUFX2_42 ( .A(_abc_19068_n1620), .Y(_abc_19068_n1620_bF_buf0) );
  BUFX2 BUFX2_420 ( .A(_abc_19068_n2487), .Y(_abc_19068_n2487_bF_buf6) );
  BUFX2 BUFX2_421 ( .A(_abc_19068_n2487), .Y(_abc_19068_n2487_bF_buf5) );
  BUFX2 BUFX2_422 ( .A(_abc_19068_n2487), .Y(_abc_19068_n2487_bF_buf4) );
  BUFX2 BUFX2_423 ( .A(_abc_19068_n2487), .Y(_abc_19068_n2487_bF_buf3) );
  BUFX2 BUFX2_424 ( .A(_abc_19068_n2487), .Y(_abc_19068_n2487_bF_buf2) );
  BUFX2 BUFX2_425 ( .A(_abc_19068_n2487), .Y(_abc_19068_n2487_bF_buf1) );
  BUFX2 BUFX2_426 ( .A(_abc_19068_n2487), .Y(_abc_19068_n2487_bF_buf0) );
  BUFX2 BUFX2_427 ( .A(core__abc_21380_n7087), .Y(core__abc_21380_n7087_bF_buf7) );
  BUFX2 BUFX2_428 ( .A(core__abc_21380_n7087), .Y(core__abc_21380_n7087_bF_buf6) );
  BUFX2 BUFX2_429 ( .A(core__abc_21380_n7087), .Y(core__abc_21380_n7087_bF_buf5) );
  BUFX2 BUFX2_43 ( .A(core__abc_21380_n2750), .Y(core__abc_21380_n2750_bF_buf7) );
  BUFX2 BUFX2_430 ( .A(core__abc_21380_n7087), .Y(core__abc_21380_n7087_bF_buf4) );
  BUFX2 BUFX2_431 ( .A(core__abc_21380_n7087), .Y(core__abc_21380_n7087_bF_buf3) );
  BUFX2 BUFX2_432 ( .A(core__abc_21380_n7087), .Y(core__abc_21380_n7087_bF_buf2) );
  BUFX2 BUFX2_433 ( .A(core__abc_21380_n7087), .Y(core__abc_21380_n7087_bF_buf1) );
  BUFX2 BUFX2_434 ( .A(core__abc_21380_n7087), .Y(core__abc_21380_n7087_bF_buf0) );
  BUFX2 BUFX2_435 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf15) );
  BUFX2 BUFX2_436 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf14) );
  BUFX2 BUFX2_437 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf13) );
  BUFX2 BUFX2_438 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf12) );
  BUFX2 BUFX2_439 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf11) );
  BUFX2 BUFX2_44 ( .A(core__abc_21380_n2750), .Y(core__abc_21380_n2750_bF_buf6) );
  BUFX2 BUFX2_440 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf10) );
  BUFX2 BUFX2_441 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf9) );
  BUFX2 BUFX2_442 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf8) );
  BUFX2 BUFX2_443 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf7) );
  BUFX2 BUFX2_444 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf6) );
  BUFX2 BUFX2_445 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf5) );
  BUFX2 BUFX2_446 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf4) );
  BUFX2 BUFX2_447 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf3) );
  BUFX2 BUFX2_448 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf2) );
  BUFX2 BUFX2_449 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf1) );
  BUFX2 BUFX2_45 ( .A(core__abc_21380_n2750), .Y(core__abc_21380_n2750_bF_buf5) );
  BUFX2 BUFX2_450 ( .A(core__abc_21380_n3167_1), .Y(core__abc_21380_n3167_1_bF_buf0) );
  BUFX2 BUFX2_451 ( .A(_abc_19068_n924_1), .Y(_abc_19068_n924_1_bF_buf4) );
  BUFX2 BUFX2_452 ( .A(_abc_19068_n924_1), .Y(_abc_19068_n924_1_bF_buf3) );
  BUFX2 BUFX2_453 ( .A(_abc_19068_n924_1), .Y(_abc_19068_n924_1_bF_buf2) );
  BUFX2 BUFX2_454 ( .A(_abc_19068_n924_1), .Y(_abc_19068_n924_1_bF_buf1) );
  BUFX2 BUFX2_455 ( .A(_abc_19068_n924_1), .Y(_abc_19068_n924_1_bF_buf0) );
  BUFX2 BUFX2_456 ( .A(_abc_19068_n2809), .Y(_abc_19068_n2809_bF_buf7) );
  BUFX2 BUFX2_457 ( .A(_abc_19068_n2809), .Y(_abc_19068_n2809_bF_buf6) );
  BUFX2 BUFX2_458 ( .A(_abc_19068_n2809), .Y(_abc_19068_n2809_bF_buf5) );
  BUFX2 BUFX2_459 ( .A(_abc_19068_n2809), .Y(_abc_19068_n2809_bF_buf4) );
  BUFX2 BUFX2_46 ( .A(core__abc_21380_n2750), .Y(core__abc_21380_n2750_bF_buf4) );
  BUFX2 BUFX2_460 ( .A(_abc_19068_n2809), .Y(_abc_19068_n2809_bF_buf3) );
  BUFX2 BUFX2_461 ( .A(_abc_19068_n2809), .Y(_abc_19068_n2809_bF_buf2) );
  BUFX2 BUFX2_462 ( .A(_abc_19068_n2809), .Y(_abc_19068_n2809_bF_buf1) );
  BUFX2 BUFX2_463 ( .A(_abc_19068_n2809), .Y(_abc_19068_n2809_bF_buf0) );
  BUFX2 BUFX2_464 ( .A(_abc_19068_n941), .Y(_abc_19068_n941_bF_buf4) );
  BUFX2 BUFX2_465 ( .A(_abc_19068_n941), .Y(_abc_19068_n941_bF_buf3) );
  BUFX2 BUFX2_466 ( .A(_abc_19068_n941), .Y(_abc_19068_n941_bF_buf2) );
  BUFX2 BUFX2_467 ( .A(_abc_19068_n941), .Y(_abc_19068_n941_bF_buf1) );
  BUFX2 BUFX2_468 ( .A(_abc_19068_n941), .Y(_abc_19068_n941_bF_buf0) );
  BUFX2 BUFX2_469 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf10) );
  BUFX2 BUFX2_47 ( .A(core__abc_21380_n2750), .Y(core__abc_21380_n2750_bF_buf3) );
  BUFX2 BUFX2_470 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf9) );
  BUFX2 BUFX2_471 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf8) );
  BUFX2 BUFX2_472 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf7) );
  BUFX2 BUFX2_473 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf6) );
  BUFX2 BUFX2_474 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf5) );
  BUFX2 BUFX2_475 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf4) );
  BUFX2 BUFX2_476 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf3) );
  BUFX2 BUFX2_477 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf2) );
  BUFX2 BUFX2_478 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf1) );
  BUFX2 BUFX2_479 ( .A(core_siphash_valid_reg), .Y(core_siphash_valid_reg_bF_buf0) );
  BUFX2 BUFX2_48 ( .A(core__abc_21380_n2750), .Y(core__abc_21380_n2750_bF_buf2) );
  BUFX2 BUFX2_480 ( .A(_abc_19068_n2970), .Y(_abc_19068_n2970_bF_buf7) );
  BUFX2 BUFX2_481 ( .A(_abc_19068_n2970), .Y(_abc_19068_n2970_bF_buf6) );
  BUFX2 BUFX2_482 ( .A(_abc_19068_n2970), .Y(_abc_19068_n2970_bF_buf5) );
  BUFX2 BUFX2_483 ( .A(_abc_19068_n2970), .Y(_abc_19068_n2970_bF_buf4) );
  BUFX2 BUFX2_484 ( .A(_abc_19068_n2970), .Y(_abc_19068_n2970_bF_buf3) );
  BUFX2 BUFX2_485 ( .A(_abc_19068_n2970), .Y(_abc_19068_n2970_bF_buf2) );
  BUFX2 BUFX2_486 ( .A(_abc_19068_n2970), .Y(_abc_19068_n2970_bF_buf1) );
  BUFX2 BUFX2_487 ( .A(_abc_19068_n2970), .Y(_abc_19068_n2970_bF_buf0) );
  BUFX2 BUFX2_488 ( .A(_auto_iopadmap_cc_313_execute_30317_0_), .Y(\read_data[0] ) );
  BUFX2 BUFX2_489 ( .A(_auto_iopadmap_cc_313_execute_30317_1_), .Y(\read_data[1] ) );
  BUFX2 BUFX2_49 ( .A(core__abc_21380_n2750), .Y(core__abc_21380_n2750_bF_buf1) );
  BUFX2 BUFX2_490 ( .A(_auto_iopadmap_cc_313_execute_30317_2_), .Y(\read_data[2] ) );
  BUFX2 BUFX2_491 ( .A(_auto_iopadmap_cc_313_execute_30317_3_), .Y(\read_data[3] ) );
  BUFX2 BUFX2_492 ( .A(_auto_iopadmap_cc_313_execute_30317_4_), .Y(\read_data[4] ) );
  BUFX2 BUFX2_493 ( .A(_auto_iopadmap_cc_313_execute_30317_5_), .Y(\read_data[5] ) );
  BUFX2 BUFX2_494 ( .A(_auto_iopadmap_cc_313_execute_30317_6_), .Y(\read_data[6] ) );
  BUFX2 BUFX2_495 ( .A(_auto_iopadmap_cc_313_execute_30317_7_), .Y(\read_data[7] ) );
  BUFX2 BUFX2_496 ( .A(_auto_iopadmap_cc_313_execute_30317_8_), .Y(\read_data[8] ) );
  BUFX2 BUFX2_497 ( .A(_auto_iopadmap_cc_313_execute_30317_9_), .Y(\read_data[9] ) );
  BUFX2 BUFX2_498 ( .A(_auto_iopadmap_cc_313_execute_30317_10_), .Y(\read_data[10] ) );
  BUFX2 BUFX2_499 ( .A(_auto_iopadmap_cc_313_execute_30317_11_), .Y(\read_data[11] ) );
  BUFX2 BUFX2_5 ( .A(clk), .Y(clk_hier0_bF_buf4) );
  BUFX2 BUFX2_50 ( .A(core__abc_21380_n2750), .Y(core__abc_21380_n2750_bF_buf0) );
  BUFX2 BUFX2_500 ( .A(_auto_iopadmap_cc_313_execute_30317_12_), .Y(\read_data[12] ) );
  BUFX2 BUFX2_501 ( .A(_auto_iopadmap_cc_313_execute_30317_13_), .Y(\read_data[13] ) );
  BUFX2 BUFX2_502 ( .A(_auto_iopadmap_cc_313_execute_30317_14_), .Y(\read_data[14] ) );
  BUFX2 BUFX2_503 ( .A(_auto_iopadmap_cc_313_execute_30317_15_), .Y(\read_data[15] ) );
  BUFX2 BUFX2_504 ( .A(_auto_iopadmap_cc_313_execute_30317_16_), .Y(\read_data[16] ) );
  BUFX2 BUFX2_505 ( .A(_auto_iopadmap_cc_313_execute_30317_17_), .Y(\read_data[17] ) );
  BUFX2 BUFX2_506 ( .A(_auto_iopadmap_cc_313_execute_30317_18_), .Y(\read_data[18] ) );
  BUFX2 BUFX2_507 ( .A(_auto_iopadmap_cc_313_execute_30317_19_), .Y(\read_data[19] ) );
  BUFX2 BUFX2_508 ( .A(_auto_iopadmap_cc_313_execute_30317_20_), .Y(\read_data[20] ) );
  BUFX2 BUFX2_509 ( .A(_auto_iopadmap_cc_313_execute_30317_21_), .Y(\read_data[21] ) );
  BUFX2 BUFX2_51 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf12) );
  BUFX2 BUFX2_510 ( .A(_auto_iopadmap_cc_313_execute_30317_22_), .Y(\read_data[22] ) );
  BUFX2 BUFX2_511 ( .A(_auto_iopadmap_cc_313_execute_30317_23_), .Y(\read_data[23] ) );
  BUFX2 BUFX2_512 ( .A(_auto_iopadmap_cc_313_execute_30317_24_), .Y(\read_data[24] ) );
  BUFX2 BUFX2_513 ( .A(_auto_iopadmap_cc_313_execute_30317_25_), .Y(\read_data[25] ) );
  BUFX2 BUFX2_514 ( .A(_auto_iopadmap_cc_313_execute_30317_26_), .Y(\read_data[26] ) );
  BUFX2 BUFX2_515 ( .A(_auto_iopadmap_cc_313_execute_30317_27_), .Y(\read_data[27] ) );
  BUFX2 BUFX2_516 ( .A(_auto_iopadmap_cc_313_execute_30317_28_), .Y(\read_data[28] ) );
  BUFX2 BUFX2_517 ( .A(_auto_iopadmap_cc_313_execute_30317_29_), .Y(\read_data[29] ) );
  BUFX2 BUFX2_518 ( .A(_auto_iopadmap_cc_313_execute_30317_30_), .Y(\read_data[30] ) );
  BUFX2 BUFX2_519 ( .A(_auto_iopadmap_cc_313_execute_30317_31_), .Y(\read_data[31] ) );
  BUFX2 BUFX2_52 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf11) );
  BUFX2 BUFX2_53 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf10) );
  BUFX2 BUFX2_54 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf9) );
  BUFX2 BUFX2_55 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf8) );
  BUFX2 BUFX2_56 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf7) );
  BUFX2 BUFX2_57 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf6) );
  BUFX2 BUFX2_58 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf5) );
  BUFX2 BUFX2_59 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf4) );
  BUFX2 BUFX2_6 ( .A(clk), .Y(clk_hier0_bF_buf3) );
  BUFX2 BUFX2_60 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf3) );
  BUFX2 BUFX2_61 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf2) );
  BUFX2 BUFX2_62 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf1) );
  BUFX2 BUFX2_63 ( .A(core__abc_21380_n3313), .Y(core__abc_21380_n3313_bF_buf0) );
  BUFX2 BUFX2_64 ( .A(core__abc_21380_n3317), .Y(core__abc_21380_n3317_bF_buf7) );
  BUFX2 BUFX2_65 ( .A(core__abc_21380_n3317), .Y(core__abc_21380_n3317_bF_buf6) );
  BUFX2 BUFX2_66 ( .A(core__abc_21380_n3317), .Y(core__abc_21380_n3317_bF_buf5) );
  BUFX2 BUFX2_67 ( .A(core__abc_21380_n3317), .Y(core__abc_21380_n3317_bF_buf4) );
  BUFX2 BUFX2_68 ( .A(core__abc_21380_n3317), .Y(core__abc_21380_n3317_bF_buf3) );
  BUFX2 BUFX2_69 ( .A(core__abc_21380_n3317), .Y(core__abc_21380_n3317_bF_buf2) );
  BUFX2 BUFX2_7 ( .A(clk), .Y(clk_hier0_bF_buf2) );
  BUFX2 BUFX2_70 ( .A(core__abc_21380_n3317), .Y(core__abc_21380_n3317_bF_buf1) );
  BUFX2 BUFX2_71 ( .A(core__abc_21380_n3317), .Y(core__abc_21380_n3317_bF_buf0) );
  BUFX2 BUFX2_72 ( .A(core__abc_21380_n8454), .Y(core__abc_21380_n8454_bF_buf7) );
  BUFX2 BUFX2_73 ( .A(core__abc_21380_n8454), .Y(core__abc_21380_n8454_bF_buf6) );
  BUFX2 BUFX2_74 ( .A(core__abc_21380_n8454), .Y(core__abc_21380_n8454_bF_buf5) );
  BUFX2 BUFX2_75 ( .A(core__abc_21380_n8454), .Y(core__abc_21380_n8454_bF_buf4) );
  BUFX2 BUFX2_76 ( .A(core__abc_21380_n8454), .Y(core__abc_21380_n8454_bF_buf3) );
  BUFX2 BUFX2_77 ( .A(core__abc_21380_n8454), .Y(core__abc_21380_n8454_bF_buf2) );
  BUFX2 BUFX2_78 ( .A(core__abc_21380_n8454), .Y(core__abc_21380_n8454_bF_buf1) );
  BUFX2 BUFX2_79 ( .A(core__abc_21380_n8454), .Y(core__abc_21380_n8454_bF_buf0) );
  BUFX2 BUFX2_8 ( .A(clk), .Y(clk_hier0_bF_buf1) );
  BUFX2 BUFX2_80 ( .A(core__abc_21380_n8455), .Y(core__abc_21380_n8455_bF_buf7) );
  BUFX2 BUFX2_81 ( .A(core__abc_21380_n8455), .Y(core__abc_21380_n8455_bF_buf6) );
  BUFX2 BUFX2_82 ( .A(core__abc_21380_n8455), .Y(core__abc_21380_n8455_bF_buf5) );
  BUFX2 BUFX2_83 ( .A(core__abc_21380_n8455), .Y(core__abc_21380_n8455_bF_buf4) );
  BUFX2 BUFX2_84 ( .A(core__abc_21380_n8455), .Y(core__abc_21380_n8455_bF_buf3) );
  BUFX2 BUFX2_85 ( .A(core__abc_21380_n8455), .Y(core__abc_21380_n8455_bF_buf2) );
  BUFX2 BUFX2_86 ( .A(core__abc_21380_n8455), .Y(core__abc_21380_n8455_bF_buf1) );
  BUFX2 BUFX2_87 ( .A(core__abc_21380_n8455), .Y(core__abc_21380_n8455_bF_buf0) );
  BUFX2 BUFX2_88 ( .A(core__abc_21380_n8456), .Y(core__abc_21380_n8456_bF_buf7) );
  BUFX2 BUFX2_89 ( .A(core__abc_21380_n8456), .Y(core__abc_21380_n8456_bF_buf6) );
  BUFX2 BUFX2_9 ( .A(clk), .Y(clk_hier0_bF_buf0) );
  BUFX2 BUFX2_90 ( .A(core__abc_21380_n8456), .Y(core__abc_21380_n8456_bF_buf5) );
  BUFX2 BUFX2_91 ( .A(core__abc_21380_n8456), .Y(core__abc_21380_n8456_bF_buf4) );
  BUFX2 BUFX2_92 ( .A(core__abc_21380_n8456), .Y(core__abc_21380_n8456_bF_buf3) );
  BUFX2 BUFX2_93 ( .A(core__abc_21380_n8456), .Y(core__abc_21380_n8456_bF_buf2) );
  BUFX2 BUFX2_94 ( .A(core__abc_21380_n8456), .Y(core__abc_21380_n8456_bF_buf1) );
  BUFX2 BUFX2_95 ( .A(core__abc_21380_n8456), .Y(core__abc_21380_n8456_bF_buf0) );
  BUFX2 BUFX2_96 ( .A(core__abc_21380_n2451_1), .Y(core__abc_21380_n2451_1_bF_buf7) );
  BUFX2 BUFX2_97 ( .A(core__abc_21380_n2451_1), .Y(core__abc_21380_n2451_1_bF_buf6) );
  BUFX2 BUFX2_98 ( .A(core__abc_21380_n2451_1), .Y(core__abc_21380_n2451_1_bF_buf5) );
  BUFX2 BUFX2_99 ( .A(core__abc_21380_n2451_1), .Y(core__abc_21380_n2451_1_bF_buf4) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf84), .D(ctrl_reg_0__FF_INPUT), .Q(core_initalize) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf75), .D(param_reg_5__FF_INPUT), .Q(core_final_rounds_1_) );
  DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf70), .D(key2_reg_23__FF_INPUT), .Q(core_key_87_) );
  DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf69), .D(key2_reg_24__FF_INPUT), .Q(core_key_88_) );
  DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf68), .D(key2_reg_25__FF_INPUT), .Q(core_key_89_) );
  DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf67), .D(key2_reg_26__FF_INPUT), .Q(core_key_90_) );
  DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf66), .D(key2_reg_27__FF_INPUT), .Q(core_key_91_) );
  DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf65), .D(key2_reg_28__FF_INPUT), .Q(core_key_92_) );
  DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf64), .D(key2_reg_29__FF_INPUT), .Q(core_key_93_) );
  DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf63), .D(key2_reg_30__FF_INPUT), .Q(core_key_94_) );
  DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf62), .D(key2_reg_31__FF_INPUT), .Q(core_key_95_) );
  DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf61), .D(key3_reg_0__FF_INPUT), .Q(core_key_96_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf74), .D(param_reg_6__FF_INPUT), .Q(core_final_rounds_2_) );
  DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf60), .D(key3_reg_1__FF_INPUT), .Q(core_key_97_) );
  DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf59), .D(key3_reg_2__FF_INPUT), .Q(core_key_98_) );
  DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf58), .D(key3_reg_3__FF_INPUT), .Q(core_key_99_) );
  DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf57), .D(key3_reg_4__FF_INPUT), .Q(core_key_100_) );
  DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf56), .D(key3_reg_5__FF_INPUT), .Q(core_key_101_) );
  DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf55), .D(key3_reg_6__FF_INPUT), .Q(core_key_102_) );
  DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf54), .D(key3_reg_7__FF_INPUT), .Q(core_key_103_) );
  DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf53), .D(key3_reg_8__FF_INPUT), .Q(core_key_104_) );
  DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf52), .D(key3_reg_9__FF_INPUT), .Q(core_key_105_) );
  DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf51), .D(key3_reg_10__FF_INPUT), .Q(core_key_106_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf73), .D(param_reg_7__FF_INPUT), .Q(core_final_rounds_3_) );
  DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf50), .D(key3_reg_11__FF_INPUT), .Q(core_key_107_) );
  DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf49), .D(key3_reg_12__FF_INPUT), .Q(core_key_108_) );
  DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf48), .D(key3_reg_13__FF_INPUT), .Q(core_key_109_) );
  DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf47), .D(key3_reg_14__FF_INPUT), .Q(core_key_110_) );
  DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf46), .D(key3_reg_15__FF_INPUT), .Q(core_key_111_) );
  DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf45), .D(key3_reg_16__FF_INPUT), .Q(core_key_112_) );
  DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf44), .D(key3_reg_17__FF_INPUT), .Q(core_key_113_) );
  DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf43), .D(key3_reg_18__FF_INPUT), .Q(core_key_114_) );
  DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf42), .D(key3_reg_19__FF_INPUT), .Q(core_key_115_) );
  DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf41), .D(key3_reg_20__FF_INPUT), .Q(core_key_116_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf72), .D(key0_reg_0__FF_INPUT), .Q(core_key_0_) );
  DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf40), .D(key3_reg_21__FF_INPUT), .Q(core_key_117_) );
  DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf39), .D(key3_reg_22__FF_INPUT), .Q(core_key_118_) );
  DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf38), .D(key3_reg_23__FF_INPUT), .Q(core_key_119_) );
  DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf37), .D(key3_reg_24__FF_INPUT), .Q(core_key_120_) );
  DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf36), .D(key3_reg_25__FF_INPUT), .Q(core_key_121_) );
  DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf35), .D(key3_reg_26__FF_INPUT), .Q(core_key_122_) );
  DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf34), .D(key3_reg_27__FF_INPUT), .Q(core_key_123_) );
  DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf33), .D(key3_reg_28__FF_INPUT), .Q(core_key_124_) );
  DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf32), .D(key3_reg_29__FF_INPUT), .Q(core_key_125_) );
  DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf31), .D(key3_reg_30__FF_INPUT), .Q(core_key_126_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf71), .D(key0_reg_1__FF_INPUT), .Q(core_key_1_) );
  DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf30), .D(key3_reg_31__FF_INPUT), .Q(core_key_127_) );
  DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf29), .D(mi0_reg_0__FF_INPUT), .Q(core_mi_0_) );
  DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf28), .D(mi0_reg_1__FF_INPUT), .Q(core_mi_1_) );
  DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf27), .D(mi0_reg_2__FF_INPUT), .Q(core_mi_2_) );
  DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf26), .D(mi0_reg_3__FF_INPUT), .Q(core_mi_3_) );
  DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf25), .D(mi0_reg_4__FF_INPUT), .Q(core_mi_4_) );
  DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf24), .D(mi0_reg_5__FF_INPUT), .Q(core_mi_5_) );
  DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf23), .D(mi0_reg_6__FF_INPUT), .Q(core_mi_6_) );
  DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf22), .D(mi0_reg_7__FF_INPUT), .Q(core_mi_7_) );
  DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf21), .D(mi0_reg_8__FF_INPUT), .Q(core_mi_8_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf70), .D(key0_reg_2__FF_INPUT), .Q(core_key_2_) );
  DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf20), .D(mi0_reg_9__FF_INPUT), .Q(core_mi_9_) );
  DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf19), .D(mi0_reg_10__FF_INPUT), .Q(core_mi_10_) );
  DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf18), .D(mi0_reg_11__FF_INPUT), .Q(core_mi_11_) );
  DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf17), .D(mi0_reg_12__FF_INPUT), .Q(core_mi_12_) );
  DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf16), .D(mi0_reg_13__FF_INPUT), .Q(core_mi_13_) );
  DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf15), .D(mi0_reg_14__FF_INPUT), .Q(core_mi_14_) );
  DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf14), .D(mi0_reg_15__FF_INPUT), .Q(core_mi_15_) );
  DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf13), .D(mi0_reg_16__FF_INPUT), .Q(core_mi_16_) );
  DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf12), .D(mi0_reg_17__FF_INPUT), .Q(core_mi_17_) );
  DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf11), .D(mi0_reg_18__FF_INPUT), .Q(core_mi_18_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf69), .D(key0_reg_3__FF_INPUT), .Q(core_key_3_) );
  DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf10), .D(mi0_reg_19__FF_INPUT), .Q(core_mi_19_) );
  DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf9), .D(mi0_reg_20__FF_INPUT), .Q(core_mi_20_) );
  DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf8), .D(mi0_reg_21__FF_INPUT), .Q(core_mi_21_) );
  DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf7), .D(mi0_reg_22__FF_INPUT), .Q(core_mi_22_) );
  DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf6), .D(mi0_reg_23__FF_INPUT), .Q(core_mi_23_) );
  DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf5), .D(mi0_reg_24__FF_INPUT), .Q(core_mi_24_) );
  DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf4), .D(mi0_reg_25__FF_INPUT), .Q(core_mi_25_) );
  DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf3), .D(mi0_reg_26__FF_INPUT), .Q(core_mi_26_) );
  DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf2), .D(mi0_reg_27__FF_INPUT), .Q(core_mi_27_) );
  DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf1), .D(mi0_reg_28__FF_INPUT), .Q(core_mi_28_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf68), .D(key0_reg_4__FF_INPUT), .Q(core_key_4_) );
  DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf0), .D(mi0_reg_29__FF_INPUT), .Q(core_mi_29_) );
  DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf84), .D(mi0_reg_30__FF_INPUT), .Q(core_mi_30_) );
  DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf83), .D(mi0_reg_31__FF_INPUT), .Q(core_mi_31_) );
  DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf82), .D(mi1_reg_0__FF_INPUT), .Q(core_mi_32_) );
  DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf81), .D(mi1_reg_1__FF_INPUT), .Q(core_mi_33_) );
  DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf80), .D(mi1_reg_2__FF_INPUT), .Q(core_mi_34_) );
  DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf79), .D(mi1_reg_3__FF_INPUT), .Q(core_mi_35_) );
  DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf78), .D(mi1_reg_4__FF_INPUT), .Q(core_mi_36_) );
  DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf77), .D(mi1_reg_5__FF_INPUT), .Q(core_mi_37_) );
  DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf76), .D(mi1_reg_6__FF_INPUT), .Q(core_mi_38_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf67), .D(key0_reg_5__FF_INPUT), .Q(core_key_5_) );
  DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf75), .D(mi1_reg_7__FF_INPUT), .Q(core_mi_39_) );
  DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf74), .D(mi1_reg_8__FF_INPUT), .Q(core_mi_40_) );
  DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf73), .D(mi1_reg_9__FF_INPUT), .Q(core_mi_41_) );
  DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf72), .D(mi1_reg_10__FF_INPUT), .Q(core_mi_42_) );
  DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf71), .D(mi1_reg_11__FF_INPUT), .Q(core_mi_43_) );
  DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf70), .D(mi1_reg_12__FF_INPUT), .Q(core_mi_44_) );
  DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf69), .D(mi1_reg_13__FF_INPUT), .Q(core_mi_45_) );
  DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf68), .D(mi1_reg_14__FF_INPUT), .Q(core_mi_46_) );
  DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf67), .D(mi1_reg_15__FF_INPUT), .Q(core_mi_47_) );
  DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf66), .D(mi1_reg_16__FF_INPUT), .Q(core_mi_48_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf66), .D(key0_reg_6__FF_INPUT), .Q(core_key_6_) );
  DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf65), .D(mi1_reg_17__FF_INPUT), .Q(core_mi_49_) );
  DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf64), .D(mi1_reg_18__FF_INPUT), .Q(core_mi_50_) );
  DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf63), .D(mi1_reg_19__FF_INPUT), .Q(core_mi_51_) );
  DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf62), .D(mi1_reg_20__FF_INPUT), .Q(core_mi_52_) );
  DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf61), .D(mi1_reg_21__FF_INPUT), .Q(core_mi_53_) );
  DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf60), .D(mi1_reg_22__FF_INPUT), .Q(core_mi_54_) );
  DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf59), .D(mi1_reg_23__FF_INPUT), .Q(core_mi_55_) );
  DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf58), .D(mi1_reg_24__FF_INPUT), .Q(core_mi_56_) );
  DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf57), .D(mi1_reg_25__FF_INPUT), .Q(core_mi_57_) );
  DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf56), .D(mi1_reg_26__FF_INPUT), .Q(core_mi_58_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf83), .D(ctrl_reg_1__FF_INPUT), .Q(core_compress) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf65), .D(key0_reg_7__FF_INPUT), .Q(core_key_7_) );
  DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf55), .D(mi1_reg_27__FF_INPUT), .Q(core_mi_59_) );
  DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf54), .D(mi1_reg_28__FF_INPUT), .Q(core_mi_60_) );
  DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf53), .D(mi1_reg_29__FF_INPUT), .Q(core_mi_61_) );
  DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf52), .D(mi1_reg_30__FF_INPUT), .Q(core_mi_62_) );
  DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf51), .D(mi1_reg_31__FF_INPUT), .Q(core_mi_63_) );
  DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf50), .D(word0_reg_0__FF_INPUT), .Q(word0_reg_0_) );
  DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf49), .D(word0_reg_1__FF_INPUT), .Q(word0_reg_1_) );
  DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf48), .D(word0_reg_2__FF_INPUT), .Q(word0_reg_2_) );
  DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf47), .D(word0_reg_3__FF_INPUT), .Q(word0_reg_3_) );
  DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf46), .D(word0_reg_4__FF_INPUT), .Q(word0_reg_4_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf64), .D(key0_reg_8__FF_INPUT), .Q(core_key_8_) );
  DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf45), .D(word0_reg_5__FF_INPUT), .Q(word0_reg_5_) );
  DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf44), .D(word0_reg_6__FF_INPUT), .Q(word0_reg_6_) );
  DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf43), .D(word0_reg_7__FF_INPUT), .Q(word0_reg_7_) );
  DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf42), .D(word0_reg_8__FF_INPUT), .Q(word0_reg_8_) );
  DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf41), .D(word0_reg_9__FF_INPUT), .Q(word0_reg_9_) );
  DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf40), .D(word0_reg_10__FF_INPUT), .Q(word0_reg_10_) );
  DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf39), .D(word0_reg_11__FF_INPUT), .Q(word0_reg_11_) );
  DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf38), .D(word0_reg_12__FF_INPUT), .Q(word0_reg_12_) );
  DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf37), .D(word0_reg_13__FF_INPUT), .Q(word0_reg_13_) );
  DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf36), .D(word0_reg_14__FF_INPUT), .Q(word0_reg_14_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf63), .D(key0_reg_9__FF_INPUT), .Q(core_key_9_) );
  DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf35), .D(word0_reg_15__FF_INPUT), .Q(word0_reg_15_) );
  DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf34), .D(word0_reg_16__FF_INPUT), .Q(word0_reg_16_) );
  DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf33), .D(word0_reg_17__FF_INPUT), .Q(word0_reg_17_) );
  DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf32), .D(word0_reg_18__FF_INPUT), .Q(word0_reg_18_) );
  DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf31), .D(word0_reg_19__FF_INPUT), .Q(word0_reg_19_) );
  DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf30), .D(word0_reg_20__FF_INPUT), .Q(word0_reg_20_) );
  DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf29), .D(word0_reg_21__FF_INPUT), .Q(word0_reg_21_) );
  DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf28), .D(word0_reg_22__FF_INPUT), .Q(word0_reg_22_) );
  DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf27), .D(word0_reg_23__FF_INPUT), .Q(word0_reg_23_) );
  DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf26), .D(word0_reg_24__FF_INPUT), .Q(word0_reg_24_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf62), .D(key0_reg_10__FF_INPUT), .Q(core_key_10_) );
  DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf25), .D(word0_reg_25__FF_INPUT), .Q(word0_reg_25_) );
  DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf24), .D(word0_reg_26__FF_INPUT), .Q(word0_reg_26_) );
  DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf23), .D(word0_reg_27__FF_INPUT), .Q(word0_reg_27_) );
  DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf22), .D(word0_reg_28__FF_INPUT), .Q(word0_reg_28_) );
  DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf21), .D(word0_reg_29__FF_INPUT), .Q(word0_reg_29_) );
  DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf20), .D(word0_reg_30__FF_INPUT), .Q(word0_reg_30_) );
  DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf19), .D(word0_reg_31__FF_INPUT), .Q(word0_reg_31_) );
  DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf18), .D(word1_reg_0__FF_INPUT), .Q(word1_reg_0_) );
  DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf17), .D(word1_reg_1__FF_INPUT), .Q(word1_reg_1_) );
  DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf16), .D(word1_reg_2__FF_INPUT), .Q(word1_reg_2_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf61), .D(key0_reg_11__FF_INPUT), .Q(core_key_11_) );
  DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf15), .D(word1_reg_3__FF_INPUT), .Q(word1_reg_3_) );
  DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf14), .D(word1_reg_4__FF_INPUT), .Q(word1_reg_4_) );
  DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf13), .D(word1_reg_5__FF_INPUT), .Q(word1_reg_5_) );
  DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf12), .D(word1_reg_6__FF_INPUT), .Q(word1_reg_6_) );
  DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf11), .D(word1_reg_7__FF_INPUT), .Q(word1_reg_7_) );
  DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf10), .D(word1_reg_8__FF_INPUT), .Q(word1_reg_8_) );
  DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf9), .D(word1_reg_9__FF_INPUT), .Q(word1_reg_9_) );
  DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf8), .D(word1_reg_10__FF_INPUT), .Q(word1_reg_10_) );
  DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf7), .D(word1_reg_11__FF_INPUT), .Q(word1_reg_11_) );
  DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf6), .D(word1_reg_12__FF_INPUT), .Q(word1_reg_12_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf60), .D(key0_reg_12__FF_INPUT), .Q(core_key_12_) );
  DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf5), .D(word1_reg_13__FF_INPUT), .Q(word1_reg_13_) );
  DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf4), .D(word1_reg_14__FF_INPUT), .Q(word1_reg_14_) );
  DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf3), .D(word1_reg_15__FF_INPUT), .Q(word1_reg_15_) );
  DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf2), .D(word1_reg_16__FF_INPUT), .Q(word1_reg_16_) );
  DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf1), .D(word1_reg_17__FF_INPUT), .Q(word1_reg_17_) );
  DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf0), .D(word1_reg_18__FF_INPUT), .Q(word1_reg_18_) );
  DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf84), .D(word1_reg_19__FF_INPUT), .Q(word1_reg_19_) );
  DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf83), .D(word1_reg_20__FF_INPUT), .Q(word1_reg_20_) );
  DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf82), .D(word1_reg_21__FF_INPUT), .Q(word1_reg_21_) );
  DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf81), .D(word1_reg_22__FF_INPUT), .Q(word1_reg_22_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf59), .D(key0_reg_13__FF_INPUT), .Q(core_key_13_) );
  DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf80), .D(word1_reg_23__FF_INPUT), .Q(word1_reg_23_) );
  DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf79), .D(word1_reg_24__FF_INPUT), .Q(word1_reg_24_) );
  DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf78), .D(word1_reg_25__FF_INPUT), .Q(word1_reg_25_) );
  DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf77), .D(word1_reg_26__FF_INPUT), .Q(word1_reg_26_) );
  DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf76), .D(word1_reg_27__FF_INPUT), .Q(word1_reg_27_) );
  DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf75), .D(word1_reg_28__FF_INPUT), .Q(word1_reg_28_) );
  DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf74), .D(word1_reg_29__FF_INPUT), .Q(word1_reg_29_) );
  DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf73), .D(word1_reg_30__FF_INPUT), .Q(word1_reg_30_) );
  DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf72), .D(word1_reg_31__FF_INPUT), .Q(word1_reg_31_) );
  DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf71), .D(word2_reg_0__FF_INPUT), .Q(word2_reg_0_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf58), .D(key0_reg_14__FF_INPUT), .Q(core_key_14_) );
  DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf70), .D(word2_reg_1__FF_INPUT), .Q(word2_reg_1_) );
  DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf69), .D(word2_reg_2__FF_INPUT), .Q(word2_reg_2_) );
  DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf68), .D(word2_reg_3__FF_INPUT), .Q(word2_reg_3_) );
  DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf67), .D(word2_reg_4__FF_INPUT), .Q(word2_reg_4_) );
  DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf66), .D(word2_reg_5__FF_INPUT), .Q(word2_reg_5_) );
  DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf65), .D(word2_reg_6__FF_INPUT), .Q(word2_reg_6_) );
  DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf64), .D(word2_reg_7__FF_INPUT), .Q(word2_reg_7_) );
  DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf63), .D(word2_reg_8__FF_INPUT), .Q(word2_reg_8_) );
  DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf62), .D(word2_reg_9__FF_INPUT), .Q(word2_reg_9_) );
  DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf61), .D(word2_reg_10__FF_INPUT), .Q(word2_reg_10_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf57), .D(key0_reg_15__FF_INPUT), .Q(core_key_15_) );
  DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf60), .D(word2_reg_11__FF_INPUT), .Q(word2_reg_11_) );
  DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf59), .D(word2_reg_12__FF_INPUT), .Q(word2_reg_12_) );
  DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf58), .D(word2_reg_13__FF_INPUT), .Q(word2_reg_13_) );
  DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf57), .D(word2_reg_14__FF_INPUT), .Q(word2_reg_14_) );
  DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf56), .D(word2_reg_15__FF_INPUT), .Q(word2_reg_15_) );
  DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf55), .D(word2_reg_16__FF_INPUT), .Q(word2_reg_16_) );
  DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf54), .D(word2_reg_17__FF_INPUT), .Q(word2_reg_17_) );
  DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf53), .D(word2_reg_18__FF_INPUT), .Q(word2_reg_18_) );
  DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf52), .D(word2_reg_19__FF_INPUT), .Q(word2_reg_19_) );
  DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf51), .D(word2_reg_20__FF_INPUT), .Q(word2_reg_20_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf56), .D(key0_reg_16__FF_INPUT), .Q(core_key_16_) );
  DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf50), .D(word2_reg_21__FF_INPUT), .Q(word2_reg_21_) );
  DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf49), .D(word2_reg_22__FF_INPUT), .Q(word2_reg_22_) );
  DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf48), .D(word2_reg_23__FF_INPUT), .Q(word2_reg_23_) );
  DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf47), .D(word2_reg_24__FF_INPUT), .Q(word2_reg_24_) );
  DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf46), .D(word2_reg_25__FF_INPUT), .Q(word2_reg_25_) );
  DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf45), .D(word2_reg_26__FF_INPUT), .Q(word2_reg_26_) );
  DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf44), .D(word2_reg_27__FF_INPUT), .Q(word2_reg_27_) );
  DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf43), .D(word2_reg_28__FF_INPUT), .Q(word2_reg_28_) );
  DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf42), .D(word2_reg_29__FF_INPUT), .Q(word2_reg_29_) );
  DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf41), .D(word2_reg_30__FF_INPUT), .Q(word2_reg_30_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf82), .D(ctrl_reg_2__FF_INPUT), .Q(core_finalize) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf55), .D(key0_reg_17__FF_INPUT), .Q(core_key_17_) );
  DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf40), .D(word2_reg_31__FF_INPUT), .Q(word2_reg_31_) );
  DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf39), .D(word3_reg_0__FF_INPUT), .Q(word3_reg_0_) );
  DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf38), .D(word3_reg_1__FF_INPUT), .Q(word3_reg_1_) );
  DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf37), .D(word3_reg_2__FF_INPUT), .Q(word3_reg_2_) );
  DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf36), .D(word3_reg_3__FF_INPUT), .Q(word3_reg_3_) );
  DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf35), .D(word3_reg_4__FF_INPUT), .Q(word3_reg_4_) );
  DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf34), .D(word3_reg_5__FF_INPUT), .Q(word3_reg_5_) );
  DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf33), .D(word3_reg_6__FF_INPUT), .Q(word3_reg_6_) );
  DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf32), .D(word3_reg_7__FF_INPUT), .Q(word3_reg_7_) );
  DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf31), .D(word3_reg_8__FF_INPUT), .Q(word3_reg_8_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf54), .D(key0_reg_18__FF_INPUT), .Q(core_key_18_) );
  DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf30), .D(word3_reg_9__FF_INPUT), .Q(word3_reg_9_) );
  DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf29), .D(word3_reg_10__FF_INPUT), .Q(word3_reg_10_) );
  DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf28), .D(word3_reg_11__FF_INPUT), .Q(word3_reg_11_) );
  DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf27), .D(word3_reg_12__FF_INPUT), .Q(word3_reg_12_) );
  DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf26), .D(word3_reg_13__FF_INPUT), .Q(word3_reg_13_) );
  DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf25), .D(word3_reg_14__FF_INPUT), .Q(word3_reg_14_) );
  DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf24), .D(word3_reg_15__FF_INPUT), .Q(word3_reg_15_) );
  DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf23), .D(word3_reg_16__FF_INPUT), .Q(word3_reg_16_) );
  DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf22), .D(word3_reg_17__FF_INPUT), .Q(word3_reg_17_) );
  DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf21), .D(word3_reg_18__FF_INPUT), .Q(word3_reg_18_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf53), .D(key0_reg_19__FF_INPUT), .Q(core_key_19_) );
  DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf20), .D(word3_reg_19__FF_INPUT), .Q(word3_reg_19_) );
  DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf19), .D(word3_reg_20__FF_INPUT), .Q(word3_reg_20_) );
  DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf18), .D(word3_reg_21__FF_INPUT), .Q(word3_reg_21_) );
  DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf17), .D(word3_reg_22__FF_INPUT), .Q(word3_reg_22_) );
  DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf16), .D(word3_reg_23__FF_INPUT), .Q(word3_reg_23_) );
  DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf15), .D(word3_reg_24__FF_INPUT), .Q(word3_reg_24_) );
  DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf14), .D(word3_reg_25__FF_INPUT), .Q(word3_reg_25_) );
  DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf13), .D(word3_reg_26__FF_INPUT), .Q(word3_reg_26_) );
  DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf12), .D(word3_reg_27__FF_INPUT), .Q(word3_reg_27_) );
  DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf11), .D(word3_reg_28__FF_INPUT), .Q(word3_reg_28_) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf52), .D(key0_reg_20__FF_INPUT), .Q(core_key_20_) );
  DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf10), .D(word3_reg_29__FF_INPUT), .Q(word3_reg_29_) );
  DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf9), .D(word3_reg_30__FF_INPUT), .Q(word3_reg_30_) );
  DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf8), .D(word3_reg_31__FF_INPUT), .Q(word3_reg_31_) );
  DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf7), .D(core__abc_14829_n1285), .Q(core_siphash_ctrl_reg_0_) );
  DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf6), .D(core__abc_14829_n6021), .Q(core_siphash_ctrl_reg_1_) );
  DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf5), .D(core__abc_14829_n6022), .Q(core_siphash_ctrl_reg_2_) );
  DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf4), .D(core__abc_14829_n1310), .Q(core_siphash_ctrl_reg_3_) );
  DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf3), .D(core__abc_14829_n1316), .Q(core_siphash_ctrl_reg_4_) );
  DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf2), .D(core__abc_14829_n6023), .Q(core_siphash_ctrl_reg_5_) );
  DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf1), .D(core__abc_14829_n1330), .Q(core_siphash_ctrl_reg_6_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf51), .D(key0_reg_21__FF_INPUT), .Q(core_key_21_) );
  DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf0), .D(core__abc_14829_n6024), .Q(core_siphash_word1_we) );
  DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf84), .D(core_v0_reg_0__FF_INPUT), .Q(core_v0_reg_0_) );
  DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf83), .D(core_v0_reg_1__FF_INPUT), .Q(core_v0_reg_1_) );
  DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf82), .D(core_v0_reg_2__FF_INPUT), .Q(core_v0_reg_2_) );
  DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf81), .D(core_v0_reg_3__FF_INPUT), .Q(core_v0_reg_3_) );
  DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf80), .D(core_v0_reg_4__FF_INPUT), .Q(core_v0_reg_4_) );
  DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf79), .D(core_v0_reg_5__FF_INPUT), .Q(core_v0_reg_5_) );
  DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf78), .D(core_v0_reg_6__FF_INPUT), .Q(core_v0_reg_6_) );
  DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf77), .D(core_v0_reg_7__FF_INPUT), .Q(core_v0_reg_7_) );
  DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf76), .D(core_v0_reg_8__FF_INPUT), .Q(core_v0_reg_8_) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf50), .D(key0_reg_22__FF_INPUT), .Q(core_key_22_) );
  DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf75), .D(core_v0_reg_9__FF_INPUT), .Q(core_v0_reg_9_) );
  DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf74), .D(core_v0_reg_10__FF_INPUT), .Q(core_v0_reg_10_) );
  DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf73), .D(core_v0_reg_11__FF_INPUT), .Q(core_v0_reg_11_) );
  DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf72), .D(core_v0_reg_12__FF_INPUT), .Q(core_v0_reg_12_) );
  DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf71), .D(core_v0_reg_13__FF_INPUT), .Q(core_v0_reg_13_) );
  DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf70), .D(core_v0_reg_14__FF_INPUT), .Q(core_v0_reg_14_) );
  DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf69), .D(core_v0_reg_15__FF_INPUT), .Q(core_v0_reg_15_) );
  DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf68), .D(core_v0_reg_16__FF_INPUT), .Q(core_v0_reg_16_) );
  DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf67), .D(core_v0_reg_17__FF_INPUT), .Q(core_v0_reg_17_) );
  DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf66), .D(core_v0_reg_18__FF_INPUT), .Q(core_v0_reg_18_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf49), .D(key0_reg_23__FF_INPUT), .Q(core_key_23_) );
  DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf65), .D(core_v0_reg_19__FF_INPUT), .Q(core_v0_reg_19_) );
  DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf64), .D(core_v0_reg_20__FF_INPUT), .Q(core_v0_reg_20_) );
  DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf63), .D(core_v0_reg_21__FF_INPUT), .Q(core_v0_reg_21_) );
  DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf62), .D(core_v0_reg_22__FF_INPUT), .Q(core_v0_reg_22_) );
  DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf61), .D(core_v0_reg_23__FF_INPUT), .Q(core_v0_reg_23_) );
  DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf60), .D(core_v0_reg_24__FF_INPUT), .Q(core_v0_reg_24_) );
  DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf59), .D(core_v0_reg_25__FF_INPUT), .Q(core_v0_reg_25_) );
  DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf58), .D(core_v0_reg_26__FF_INPUT), .Q(core_v0_reg_26_) );
  DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf57), .D(core_v0_reg_27__FF_INPUT), .Q(core_v0_reg_27_) );
  DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf56), .D(core_v0_reg_28__FF_INPUT), .Q(core_v0_reg_28_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf48), .D(key0_reg_24__FF_INPUT), .Q(core_key_24_) );
  DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf55), .D(core_v0_reg_29__FF_INPUT), .Q(core_v0_reg_29_) );
  DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf54), .D(core_v0_reg_30__FF_INPUT), .Q(core_v0_reg_30_) );
  DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf53), .D(core_v0_reg_31__FF_INPUT), .Q(core_v0_reg_31_) );
  DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf52), .D(core_v0_reg_32__FF_INPUT), .Q(core_v0_reg_32_) );
  DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf51), .D(core_v0_reg_33__FF_INPUT), .Q(core_v0_reg_33_) );
  DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf50), .D(core_v0_reg_34__FF_INPUT), .Q(core_v0_reg_34_) );
  DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf49), .D(core_v0_reg_35__FF_INPUT), .Q(core_v0_reg_35_) );
  DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf48), .D(core_v0_reg_36__FF_INPUT), .Q(core_v0_reg_36_) );
  DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf47), .D(core_v0_reg_37__FF_INPUT), .Q(core_v0_reg_37_) );
  DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf46), .D(core_v0_reg_38__FF_INPUT), .Q(core_v0_reg_38_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf47), .D(key0_reg_25__FF_INPUT), .Q(core_key_25_) );
  DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf45), .D(core_v0_reg_39__FF_INPUT), .Q(core_v0_reg_39_) );
  DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf44), .D(core_v0_reg_40__FF_INPUT), .Q(core_v0_reg_40_) );
  DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf43), .D(core_v0_reg_41__FF_INPUT), .Q(core_v0_reg_41_) );
  DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf42), .D(core_v0_reg_42__FF_INPUT), .Q(core_v0_reg_42_) );
  DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf41), .D(core_v0_reg_43__FF_INPUT), .Q(core_v0_reg_43_) );
  DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf40), .D(core_v0_reg_44__FF_INPUT), .Q(core_v0_reg_44_) );
  DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf39), .D(core_v0_reg_45__FF_INPUT), .Q(core_v0_reg_45_) );
  DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf38), .D(core_v0_reg_46__FF_INPUT), .Q(core_v0_reg_46_) );
  DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf37), .D(core_v0_reg_47__FF_INPUT), .Q(core_v0_reg_47_) );
  DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf36), .D(core_v0_reg_48__FF_INPUT), .Q(core_v0_reg_48_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf46), .D(key0_reg_26__FF_INPUT), .Q(core_key_26_) );
  DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf35), .D(core_v0_reg_49__FF_INPUT), .Q(core_v0_reg_49_) );
  DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf34), .D(core_v0_reg_50__FF_INPUT), .Q(core_v0_reg_50_) );
  DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf33), .D(core_v0_reg_51__FF_INPUT), .Q(core_v0_reg_51_) );
  DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf32), .D(core_v0_reg_52__FF_INPUT), .Q(core_v0_reg_52_) );
  DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf31), .D(core_v0_reg_53__FF_INPUT), .Q(core_v0_reg_53_) );
  DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf30), .D(core_v0_reg_54__FF_INPUT), .Q(core_v0_reg_54_) );
  DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf29), .D(core_v0_reg_55__FF_INPUT), .Q(core_v0_reg_55_) );
  DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf28), .D(core_v0_reg_56__FF_INPUT), .Q(core_v0_reg_56_) );
  DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf27), .D(core_v0_reg_57__FF_INPUT), .Q(core_v0_reg_57_) );
  DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf26), .D(core_v0_reg_58__FF_INPUT), .Q(core_v0_reg_58_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf81), .D(long_reg_FF_INPUT), .Q(core_long) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf45), .D(key0_reg_27__FF_INPUT), .Q(core_key_27_) );
  DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf25), .D(core_v0_reg_59__FF_INPUT), .Q(core_v0_reg_59_) );
  DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf24), .D(core_v0_reg_60__FF_INPUT), .Q(core_v0_reg_60_) );
  DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf23), .D(core_v0_reg_61__FF_INPUT), .Q(core_v0_reg_61_) );
  DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf22), .D(core_v0_reg_62__FF_INPUT), .Q(core_v0_reg_62_) );
  DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf21), .D(core_v0_reg_63__FF_INPUT), .Q(core_v0_reg_63_) );
  DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf20), .D(core_v1_reg_0__FF_INPUT), .Q(core_v1_reg_0_) );
  DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf19), .D(core_v1_reg_1__FF_INPUT), .Q(core_v1_reg_1_) );
  DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf18), .D(core_v1_reg_2__FF_INPUT), .Q(core_v1_reg_2_) );
  DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf17), .D(core_v1_reg_3__FF_INPUT), .Q(core_v1_reg_3_) );
  DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf16), .D(core_v1_reg_4__FF_INPUT), .Q(core_v1_reg_4_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf44), .D(key0_reg_28__FF_INPUT), .Q(core_key_28_) );
  DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf15), .D(core_v1_reg_5__FF_INPUT), .Q(core_v1_reg_5_) );
  DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf14), .D(core_v1_reg_6__FF_INPUT), .Q(core_v1_reg_6_) );
  DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf13), .D(core_v1_reg_7__FF_INPUT), .Q(core_v1_reg_7_) );
  DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf12), .D(core_v1_reg_8__FF_INPUT), .Q(core_v1_reg_8_) );
  DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf11), .D(core_v1_reg_9__FF_INPUT), .Q(core_v1_reg_9_) );
  DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf10), .D(core_v1_reg_10__FF_INPUT), .Q(core_v1_reg_10_) );
  DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf9), .D(core_v1_reg_11__FF_INPUT), .Q(core_v1_reg_11_) );
  DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf8), .D(core_v1_reg_12__FF_INPUT), .Q(core_v1_reg_12_) );
  DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf7), .D(core_v1_reg_13__FF_INPUT), .Q(core_v1_reg_13_) );
  DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf6), .D(core_v1_reg_14__FF_INPUT), .Q(core_v1_reg_14_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf43), .D(key0_reg_29__FF_INPUT), .Q(core_key_29_) );
  DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf5), .D(core_v1_reg_15__FF_INPUT), .Q(core_v1_reg_15_) );
  DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf4), .D(core_v1_reg_16__FF_INPUT), .Q(core_v1_reg_16_) );
  DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf3), .D(core_v1_reg_17__FF_INPUT), .Q(core_v1_reg_17_) );
  DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf2), .D(core_v1_reg_18__FF_INPUT), .Q(core_v1_reg_18_) );
  DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf1), .D(core_v1_reg_19__FF_INPUT), .Q(core_v1_reg_19_) );
  DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf0), .D(core_v1_reg_20__FF_INPUT), .Q(core_v1_reg_20_) );
  DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf84), .D(core_v1_reg_21__FF_INPUT), .Q(core_v1_reg_21_) );
  DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf83), .D(core_v1_reg_22__FF_INPUT), .Q(core_v1_reg_22_) );
  DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf82), .D(core_v1_reg_23__FF_INPUT), .Q(core_v1_reg_23_) );
  DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf81), .D(core_v1_reg_24__FF_INPUT), .Q(core_v1_reg_24_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf42), .D(key0_reg_30__FF_INPUT), .Q(core_key_30_) );
  DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf80), .D(core_v1_reg_25__FF_INPUT), .Q(core_v1_reg_25_) );
  DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf79), .D(core_v1_reg_26__FF_INPUT), .Q(core_v1_reg_26_) );
  DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf78), .D(core_v1_reg_27__FF_INPUT), .Q(core_v1_reg_27_) );
  DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf77), .D(core_v1_reg_28__FF_INPUT), .Q(core_v1_reg_28_) );
  DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf76), .D(core_v1_reg_29__FF_INPUT), .Q(core_v1_reg_29_) );
  DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf75), .D(core_v1_reg_30__FF_INPUT), .Q(core_v1_reg_30_) );
  DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf74), .D(core_v1_reg_31__FF_INPUT), .Q(core_v1_reg_31_) );
  DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf73), .D(core_v1_reg_32__FF_INPUT), .Q(core_v1_reg_32_) );
  DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf72), .D(core_v1_reg_33__FF_INPUT), .Q(core_v1_reg_33_) );
  DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf71), .D(core_v1_reg_34__FF_INPUT), .Q(core_v1_reg_34_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf41), .D(key0_reg_31__FF_INPUT), .Q(core_key_31_) );
  DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf70), .D(core_v1_reg_35__FF_INPUT), .Q(core_v1_reg_35_) );
  DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf69), .D(core_v1_reg_36__FF_INPUT), .Q(core_v1_reg_36_) );
  DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf68), .D(core_v1_reg_37__FF_INPUT), .Q(core_v1_reg_37_) );
  DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf67), .D(core_v1_reg_38__FF_INPUT), .Q(core_v1_reg_38_) );
  DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf66), .D(core_v1_reg_39__FF_INPUT), .Q(core_v1_reg_39_) );
  DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf65), .D(core_v1_reg_40__FF_INPUT), .Q(core_v1_reg_40_) );
  DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf64), .D(core_v1_reg_41__FF_INPUT), .Q(core_v1_reg_41_) );
  DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf63), .D(core_v1_reg_42__FF_INPUT), .Q(core_v1_reg_42_) );
  DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf62), .D(core_v1_reg_43__FF_INPUT), .Q(core_v1_reg_43_) );
  DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf61), .D(core_v1_reg_44__FF_INPUT), .Q(core_v1_reg_44_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf40), .D(key1_reg_0__FF_INPUT), .Q(core_key_32_) );
  DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf60), .D(core_v1_reg_45__FF_INPUT), .Q(core_v1_reg_45_) );
  DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf59), .D(core_v1_reg_46__FF_INPUT), .Q(core_v1_reg_46_) );
  DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf58), .D(core_v1_reg_47__FF_INPUT), .Q(core_v1_reg_47_) );
  DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf57), .D(core_v1_reg_48__FF_INPUT), .Q(core_v1_reg_48_) );
  DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf56), .D(core_v1_reg_49__FF_INPUT), .Q(core_v1_reg_49_) );
  DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf55), .D(core_v1_reg_50__FF_INPUT), .Q(core_v1_reg_50_) );
  DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf54), .D(core_v1_reg_51__FF_INPUT), .Q(core_v1_reg_51_) );
  DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf53), .D(core_v1_reg_52__FF_INPUT), .Q(core_v1_reg_52_) );
  DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf52), .D(core_v1_reg_53__FF_INPUT), .Q(core_v1_reg_53_) );
  DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf51), .D(core_v1_reg_54__FF_INPUT), .Q(core_v1_reg_54_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf39), .D(key1_reg_1__FF_INPUT), .Q(core_key_33_) );
  DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf50), .D(core_v1_reg_55__FF_INPUT), .Q(core_v1_reg_55_) );
  DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf49), .D(core_v1_reg_56__FF_INPUT), .Q(core_v1_reg_56_) );
  DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf48), .D(core_v1_reg_57__FF_INPUT), .Q(core_v1_reg_57_) );
  DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf47), .D(core_v1_reg_58__FF_INPUT), .Q(core_v1_reg_58_) );
  DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf46), .D(core_v1_reg_59__FF_INPUT), .Q(core_v1_reg_59_) );
  DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf45), .D(core_v1_reg_60__FF_INPUT), .Q(core_v1_reg_60_) );
  DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf44), .D(core_v1_reg_61__FF_INPUT), .Q(core_v1_reg_61_) );
  DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf43), .D(core_v1_reg_62__FF_INPUT), .Q(core_v1_reg_62_) );
  DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf42), .D(core_v1_reg_63__FF_INPUT), .Q(core_v1_reg_63_) );
  DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf41), .D(core_v2_reg_0__FF_INPUT), .Q(core_v2_reg_0_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf38), .D(key1_reg_2__FF_INPUT), .Q(core_key_34_) );
  DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf40), .D(core_v2_reg_1__FF_INPUT), .Q(core_v2_reg_1_) );
  DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf39), .D(core_v2_reg_2__FF_INPUT), .Q(core_v2_reg_2_) );
  DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf38), .D(core_v2_reg_3__FF_INPUT), .Q(core_v2_reg_3_) );
  DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf37), .D(core_v2_reg_4__FF_INPUT), .Q(core_v2_reg_4_) );
  DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf36), .D(core_v2_reg_5__FF_INPUT), .Q(core_v2_reg_5_) );
  DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf35), .D(core_v2_reg_6__FF_INPUT), .Q(core_v2_reg_6_) );
  DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf34), .D(core_v2_reg_7__FF_INPUT), .Q(core_v2_reg_7_) );
  DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf33), .D(core_v2_reg_8__FF_INPUT), .Q(core_v2_reg_8_) );
  DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf32), .D(core_v2_reg_9__FF_INPUT), .Q(core_v2_reg_9_) );
  DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf31), .D(core_v2_reg_10__FF_INPUT), .Q(core_v2_reg_10_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf37), .D(key1_reg_3__FF_INPUT), .Q(core_key_35_) );
  DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf30), .D(core_v2_reg_11__FF_INPUT), .Q(core_v2_reg_11_) );
  DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf29), .D(core_v2_reg_12__FF_INPUT), .Q(core_v2_reg_12_) );
  DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf28), .D(core_v2_reg_13__FF_INPUT), .Q(core_v2_reg_13_) );
  DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf27), .D(core_v2_reg_14__FF_INPUT), .Q(core_v2_reg_14_) );
  DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf26), .D(core_v2_reg_15__FF_INPUT), .Q(core_v2_reg_15_) );
  DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf25), .D(core_v2_reg_16__FF_INPUT), .Q(core_v2_reg_16_) );
  DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf24), .D(core_v2_reg_17__FF_INPUT), .Q(core_v2_reg_17_) );
  DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf23), .D(core_v2_reg_18__FF_INPUT), .Q(core_v2_reg_18_) );
  DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf22), .D(core_v2_reg_19__FF_INPUT), .Q(core_v2_reg_19_) );
  DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf21), .D(core_v2_reg_20__FF_INPUT), .Q(core_v2_reg_20_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf36), .D(key1_reg_4__FF_INPUT), .Q(core_key_36_) );
  DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf20), .D(core_v2_reg_21__FF_INPUT), .Q(core_v2_reg_21_) );
  DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf19), .D(core_v2_reg_22__FF_INPUT), .Q(core_v2_reg_22_) );
  DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf18), .D(core_v2_reg_23__FF_INPUT), .Q(core_v2_reg_23_) );
  DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf17), .D(core_v2_reg_24__FF_INPUT), .Q(core_v2_reg_24_) );
  DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf16), .D(core_v2_reg_25__FF_INPUT), .Q(core_v2_reg_25_) );
  DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf15), .D(core_v2_reg_26__FF_INPUT), .Q(core_v2_reg_26_) );
  DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf14), .D(core_v2_reg_27__FF_INPUT), .Q(core_v2_reg_27_) );
  DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf13), .D(core_v2_reg_28__FF_INPUT), .Q(core_v2_reg_28_) );
  DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf12), .D(core_v2_reg_29__FF_INPUT), .Q(core_v2_reg_29_) );
  DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf11), .D(core_v2_reg_30__FF_INPUT), .Q(core_v2_reg_30_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf80), .D(param_reg_0__FF_INPUT), .Q(core_compression_rounds_0_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf35), .D(key1_reg_5__FF_INPUT), .Q(core_key_37_) );
  DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf10), .D(core_v2_reg_31__FF_INPUT), .Q(core_v2_reg_31_) );
  DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf9), .D(core_v2_reg_32__FF_INPUT), .Q(core_v2_reg_32_) );
  DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf8), .D(core_v2_reg_33__FF_INPUT), .Q(core_v2_reg_33_) );
  DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf7), .D(core_v2_reg_34__FF_INPUT), .Q(core_v2_reg_34_) );
  DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf6), .D(core_v2_reg_35__FF_INPUT), .Q(core_v2_reg_35_) );
  DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf5), .D(core_v2_reg_36__FF_INPUT), .Q(core_v2_reg_36_) );
  DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf4), .D(core_v2_reg_37__FF_INPUT), .Q(core_v2_reg_37_) );
  DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf3), .D(core_v2_reg_38__FF_INPUT), .Q(core_v2_reg_38_) );
  DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf2), .D(core_v2_reg_39__FF_INPUT), .Q(core_v2_reg_39_) );
  DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf1), .D(core_v2_reg_40__FF_INPUT), .Q(core_v2_reg_40_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf34), .D(key1_reg_6__FF_INPUT), .Q(core_key_38_) );
  DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf0), .D(core_v2_reg_41__FF_INPUT), .Q(core_v2_reg_41_) );
  DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf84), .D(core_v2_reg_42__FF_INPUT), .Q(core_v2_reg_42_) );
  DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf83), .D(core_v2_reg_43__FF_INPUT), .Q(core_v2_reg_43_) );
  DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf82), .D(core_v2_reg_44__FF_INPUT), .Q(core_v2_reg_44_) );
  DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf81), .D(core_v2_reg_45__FF_INPUT), .Q(core_v2_reg_45_) );
  DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf80), .D(core_v2_reg_46__FF_INPUT), .Q(core_v2_reg_46_) );
  DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf79), .D(core_v2_reg_47__FF_INPUT), .Q(core_v2_reg_47_) );
  DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf78), .D(core_v2_reg_48__FF_INPUT), .Q(core_v2_reg_48_) );
  DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf77), .D(core_v2_reg_49__FF_INPUT), .Q(core_v2_reg_49_) );
  DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf76), .D(core_v2_reg_50__FF_INPUT), .Q(core_v2_reg_50_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf33), .D(key1_reg_7__FF_INPUT), .Q(core_key_39_) );
  DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf75), .D(core_v2_reg_51__FF_INPUT), .Q(core_v2_reg_51_) );
  DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf74), .D(core_v2_reg_52__FF_INPUT), .Q(core_v2_reg_52_) );
  DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf73), .D(core_v2_reg_53__FF_INPUT), .Q(core_v2_reg_53_) );
  DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf72), .D(core_v2_reg_54__FF_INPUT), .Q(core_v2_reg_54_) );
  DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf71), .D(core_v2_reg_55__FF_INPUT), .Q(core_v2_reg_55_) );
  DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf70), .D(core_v2_reg_56__FF_INPUT), .Q(core_v2_reg_56_) );
  DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf69), .D(core_v2_reg_57__FF_INPUT), .Q(core_v2_reg_57_) );
  DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf68), .D(core_v2_reg_58__FF_INPUT), .Q(core_v2_reg_58_) );
  DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf67), .D(core_v2_reg_59__FF_INPUT), .Q(core_v2_reg_59_) );
  DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf66), .D(core_v2_reg_60__FF_INPUT), .Q(core_v2_reg_60_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf32), .D(key1_reg_8__FF_INPUT), .Q(core_key_40_) );
  DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf65), .D(core_v2_reg_61__FF_INPUT), .Q(core_v2_reg_61_) );
  DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf64), .D(core_v2_reg_62__FF_INPUT), .Q(core_v2_reg_62_) );
  DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf63), .D(core_v2_reg_63__FF_INPUT), .Q(core_v2_reg_63_) );
  DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf62), .D(core_v3_reg_0__FF_INPUT), .Q(core_v3_reg_0_) );
  DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf61), .D(core_v3_reg_1__FF_INPUT), .Q(core_v3_reg_1_) );
  DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf60), .D(core_v3_reg_2__FF_INPUT), .Q(core_v3_reg_2_) );
  DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf59), .D(core_v3_reg_3__FF_INPUT), .Q(core_v3_reg_3_) );
  DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf58), .D(core_v3_reg_4__FF_INPUT), .Q(core_v3_reg_4_) );
  DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf57), .D(core_v3_reg_5__FF_INPUT), .Q(core_v3_reg_5_) );
  DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf56), .D(core_v3_reg_6__FF_INPUT), .Q(core_v3_reg_6_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf31), .D(key1_reg_9__FF_INPUT), .Q(core_key_41_) );
  DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf55), .D(core_v3_reg_7__FF_INPUT), .Q(core_v3_reg_7_) );
  DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf54), .D(core_v3_reg_8__FF_INPUT), .Q(core_v3_reg_8_) );
  DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf53), .D(core_v3_reg_9__FF_INPUT), .Q(core_v3_reg_9_) );
  DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf52), .D(core_v3_reg_10__FF_INPUT), .Q(core_v3_reg_10_) );
  DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf51), .D(core_v3_reg_11__FF_INPUT), .Q(core_v3_reg_11_) );
  DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf50), .D(core_v3_reg_12__FF_INPUT), .Q(core_v3_reg_12_) );
  DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf49), .D(core_v3_reg_13__FF_INPUT), .Q(core_v3_reg_13_) );
  DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf48), .D(core_v3_reg_14__FF_INPUT), .Q(core_v3_reg_14_) );
  DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf47), .D(core_v3_reg_15__FF_INPUT), .Q(core_v3_reg_15_) );
  DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf46), .D(core_v3_reg_16__FF_INPUT), .Q(core_v3_reg_16_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf30), .D(key1_reg_10__FF_INPUT), .Q(core_key_42_) );
  DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf45), .D(core_v3_reg_17__FF_INPUT), .Q(core_v3_reg_17_) );
  DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf44), .D(core_v3_reg_18__FF_INPUT), .Q(core_v3_reg_18_) );
  DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf43), .D(core_v3_reg_19__FF_INPUT), .Q(core_v3_reg_19_) );
  DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf42), .D(core_v3_reg_20__FF_INPUT), .Q(core_v3_reg_20_) );
  DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf41), .D(core_v3_reg_21__FF_INPUT), .Q(core_v3_reg_21_) );
  DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf40), .D(core_v3_reg_22__FF_INPUT), .Q(core_v3_reg_22_) );
  DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf39), .D(core_v3_reg_23__FF_INPUT), .Q(core_v3_reg_23_) );
  DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf38), .D(core_v3_reg_24__FF_INPUT), .Q(core_v3_reg_24_) );
  DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf37), .D(core_v3_reg_25__FF_INPUT), .Q(core_v3_reg_25_) );
  DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf36), .D(core_v3_reg_26__FF_INPUT), .Q(core_v3_reg_26_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf29), .D(key1_reg_11__FF_INPUT), .Q(core_key_43_) );
  DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf35), .D(core_v3_reg_27__FF_INPUT), .Q(core_v3_reg_27_) );
  DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf34), .D(core_v3_reg_28__FF_INPUT), .Q(core_v3_reg_28_) );
  DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf33), .D(core_v3_reg_29__FF_INPUT), .Q(core_v3_reg_29_) );
  DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf32), .D(core_v3_reg_30__FF_INPUT), .Q(core_v3_reg_30_) );
  DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf31), .D(core_v3_reg_31__FF_INPUT), .Q(core_v3_reg_31_) );
  DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf30), .D(core_v3_reg_32__FF_INPUT), .Q(core_v3_reg_32_) );
  DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf29), .D(core_v3_reg_33__FF_INPUT), .Q(core_v3_reg_33_) );
  DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf28), .D(core_v3_reg_34__FF_INPUT), .Q(core_v3_reg_34_) );
  DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf27), .D(core_v3_reg_35__FF_INPUT), .Q(core_v3_reg_35_) );
  DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf26), .D(core_v3_reg_36__FF_INPUT), .Q(core_v3_reg_36_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf28), .D(key1_reg_12__FF_INPUT), .Q(core_key_44_) );
  DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf25), .D(core_v3_reg_37__FF_INPUT), .Q(core_v3_reg_37_) );
  DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf24), .D(core_v3_reg_38__FF_INPUT), .Q(core_v3_reg_38_) );
  DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf23), .D(core_v3_reg_39__FF_INPUT), .Q(core_v3_reg_39_) );
  DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf22), .D(core_v3_reg_40__FF_INPUT), .Q(core_v3_reg_40_) );
  DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf21), .D(core_v3_reg_41__FF_INPUT), .Q(core_v3_reg_41_) );
  DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf20), .D(core_v3_reg_42__FF_INPUT), .Q(core_v3_reg_42_) );
  DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf19), .D(core_v3_reg_43__FF_INPUT), .Q(core_v3_reg_43_) );
  DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf18), .D(core_v3_reg_44__FF_INPUT), .Q(core_v3_reg_44_) );
  DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf17), .D(core_v3_reg_45__FF_INPUT), .Q(core_v3_reg_45_) );
  DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf16), .D(core_v3_reg_46__FF_INPUT), .Q(core_v3_reg_46_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf27), .D(key1_reg_13__FF_INPUT), .Q(core_key_45_) );
  DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf15), .D(core_v3_reg_47__FF_INPUT), .Q(core_v3_reg_47_) );
  DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf14), .D(core_v3_reg_48__FF_INPUT), .Q(core_v3_reg_48_) );
  DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf13), .D(core_v3_reg_49__FF_INPUT), .Q(core_v3_reg_49_) );
  DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf12), .D(core_v3_reg_50__FF_INPUT), .Q(core_v3_reg_50_) );
  DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf11), .D(core_v3_reg_51__FF_INPUT), .Q(core_v3_reg_51_) );
  DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf10), .D(core_v3_reg_52__FF_INPUT), .Q(core_v3_reg_52_) );
  DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf9), .D(core_v3_reg_53__FF_INPUT), .Q(core_v3_reg_53_) );
  DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf8), .D(core_v3_reg_54__FF_INPUT), .Q(core_v3_reg_54_) );
  DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf7), .D(core_v3_reg_55__FF_INPUT), .Q(core_v3_reg_55_) );
  DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf6), .D(core_v3_reg_56__FF_INPUT), .Q(core_v3_reg_56_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf26), .D(key1_reg_14__FF_INPUT), .Q(core_key_46_) );
  DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf5), .D(core_v3_reg_57__FF_INPUT), .Q(core_v3_reg_57_) );
  DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf4), .D(core_v3_reg_58__FF_INPUT), .Q(core_v3_reg_58_) );
  DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf3), .D(core_v3_reg_59__FF_INPUT), .Q(core_v3_reg_59_) );
  DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf2), .D(core_v3_reg_60__FF_INPUT), .Q(core_v3_reg_60_) );
  DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf1), .D(core_v3_reg_61__FF_INPUT), .Q(core_v3_reg_61_) );
  DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf0), .D(core_v3_reg_62__FF_INPUT), .Q(core_v3_reg_62_) );
  DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf84), .D(core_v3_reg_63__FF_INPUT), .Q(core_v3_reg_63_) );
  DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf83), .D(core_mi_reg_0__FF_INPUT), .Q(core_mi_reg_0_) );
  DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf82), .D(core_mi_reg_1__FF_INPUT), .Q(core_mi_reg_1_) );
  DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf81), .D(core_mi_reg_2__FF_INPUT), .Q(core_mi_reg_2_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf79), .D(param_reg_1__FF_INPUT), .Q(core_compression_rounds_1_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf25), .D(key1_reg_15__FF_INPUT), .Q(core_key_47_) );
  DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf80), .D(core_mi_reg_3__FF_INPUT), .Q(core_mi_reg_3_) );
  DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf79), .D(core_mi_reg_4__FF_INPUT), .Q(core_mi_reg_4_) );
  DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf78), .D(core_mi_reg_5__FF_INPUT), .Q(core_mi_reg_5_) );
  DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf77), .D(core_mi_reg_6__FF_INPUT), .Q(core_mi_reg_6_) );
  DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf76), .D(core_mi_reg_7__FF_INPUT), .Q(core_mi_reg_7_) );
  DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf75), .D(core_mi_reg_8__FF_INPUT), .Q(core_mi_reg_8_) );
  DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf74), .D(core_mi_reg_9__FF_INPUT), .Q(core_mi_reg_9_) );
  DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf73), .D(core_mi_reg_10__FF_INPUT), .Q(core_mi_reg_10_) );
  DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf72), .D(core_mi_reg_11__FF_INPUT), .Q(core_mi_reg_11_) );
  DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf71), .D(core_mi_reg_12__FF_INPUT), .Q(core_mi_reg_12_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf24), .D(key1_reg_16__FF_INPUT), .Q(core_key_48_) );
  DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf70), .D(core_mi_reg_13__FF_INPUT), .Q(core_mi_reg_13_) );
  DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf69), .D(core_mi_reg_14__FF_INPUT), .Q(core_mi_reg_14_) );
  DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf68), .D(core_mi_reg_15__FF_INPUT), .Q(core_mi_reg_15_) );
  DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf67), .D(core_mi_reg_16__FF_INPUT), .Q(core_mi_reg_16_) );
  DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf66), .D(core_mi_reg_17__FF_INPUT), .Q(core_mi_reg_17_) );
  DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf65), .D(core_mi_reg_18__FF_INPUT), .Q(core_mi_reg_18_) );
  DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf64), .D(core_mi_reg_19__FF_INPUT), .Q(core_mi_reg_19_) );
  DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf63), .D(core_mi_reg_20__FF_INPUT), .Q(core_mi_reg_20_) );
  DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf62), .D(core_mi_reg_21__FF_INPUT), .Q(core_mi_reg_21_) );
  DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf61), .D(core_mi_reg_22__FF_INPUT), .Q(core_mi_reg_22_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf23), .D(key1_reg_17__FF_INPUT), .Q(core_key_49_) );
  DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf60), .D(core_mi_reg_23__FF_INPUT), .Q(core_mi_reg_23_) );
  DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf59), .D(core_mi_reg_24__FF_INPUT), .Q(core_mi_reg_24_) );
  DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf58), .D(core_mi_reg_25__FF_INPUT), .Q(core_mi_reg_25_) );
  DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf57), .D(core_mi_reg_26__FF_INPUT), .Q(core_mi_reg_26_) );
  DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf56), .D(core_mi_reg_27__FF_INPUT), .Q(core_mi_reg_27_) );
  DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf55), .D(core_mi_reg_28__FF_INPUT), .Q(core_mi_reg_28_) );
  DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf54), .D(core_mi_reg_29__FF_INPUT), .Q(core_mi_reg_29_) );
  DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf53), .D(core_mi_reg_30__FF_INPUT), .Q(core_mi_reg_30_) );
  DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf52), .D(core_mi_reg_31__FF_INPUT), .Q(core_mi_reg_31_) );
  DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf51), .D(core_mi_reg_32__FF_INPUT), .Q(core_mi_reg_32_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf22), .D(key1_reg_18__FF_INPUT), .Q(core_key_50_) );
  DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf50), .D(core_mi_reg_33__FF_INPUT), .Q(core_mi_reg_33_) );
  DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf49), .D(core_mi_reg_34__FF_INPUT), .Q(core_mi_reg_34_) );
  DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf48), .D(core_mi_reg_35__FF_INPUT), .Q(core_mi_reg_35_) );
  DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf47), .D(core_mi_reg_36__FF_INPUT), .Q(core_mi_reg_36_) );
  DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf46), .D(core_mi_reg_37__FF_INPUT), .Q(core_mi_reg_37_) );
  DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf45), .D(core_mi_reg_38__FF_INPUT), .Q(core_mi_reg_38_) );
  DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf44), .D(core_mi_reg_39__FF_INPUT), .Q(core_mi_reg_39_) );
  DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf43), .D(core_mi_reg_40__FF_INPUT), .Q(core_mi_reg_40_) );
  DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf42), .D(core_mi_reg_41__FF_INPUT), .Q(core_mi_reg_41_) );
  DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf41), .D(core_mi_reg_42__FF_INPUT), .Q(core_mi_reg_42_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf21), .D(key1_reg_19__FF_INPUT), .Q(core_key_51_) );
  DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf40), .D(core_mi_reg_43__FF_INPUT), .Q(core_mi_reg_43_) );
  DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf39), .D(core_mi_reg_44__FF_INPUT), .Q(core_mi_reg_44_) );
  DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf38), .D(core_mi_reg_45__FF_INPUT), .Q(core_mi_reg_45_) );
  DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf37), .D(core_mi_reg_46__FF_INPUT), .Q(core_mi_reg_46_) );
  DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf36), .D(core_mi_reg_47__FF_INPUT), .Q(core_mi_reg_47_) );
  DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf35), .D(core_mi_reg_48__FF_INPUT), .Q(core_mi_reg_48_) );
  DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf34), .D(core_mi_reg_49__FF_INPUT), .Q(core_mi_reg_49_) );
  DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf33), .D(core_mi_reg_50__FF_INPUT), .Q(core_mi_reg_50_) );
  DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf32), .D(core_mi_reg_51__FF_INPUT), .Q(core_mi_reg_51_) );
  DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf31), .D(core_mi_reg_52__FF_INPUT), .Q(core_mi_reg_52_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf20), .D(key1_reg_20__FF_INPUT), .Q(core_key_52_) );
  DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf30), .D(core_mi_reg_53__FF_INPUT), .Q(core_mi_reg_53_) );
  DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf29), .D(core_mi_reg_54__FF_INPUT), .Q(core_mi_reg_54_) );
  DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf28), .D(core_mi_reg_55__FF_INPUT), .Q(core_mi_reg_55_) );
  DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf27), .D(core_mi_reg_56__FF_INPUT), .Q(core_mi_reg_56_) );
  DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf26), .D(core_mi_reg_57__FF_INPUT), .Q(core_mi_reg_57_) );
  DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf25), .D(core_mi_reg_58__FF_INPUT), .Q(core_mi_reg_58_) );
  DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf24), .D(core_mi_reg_59__FF_INPUT), .Q(core_mi_reg_59_) );
  DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf23), .D(core_mi_reg_60__FF_INPUT), .Q(core_mi_reg_60_) );
  DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf22), .D(core_mi_reg_61__FF_INPUT), .Q(core_mi_reg_61_) );
  DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf21), .D(core_mi_reg_62__FF_INPUT), .Q(core_mi_reg_62_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf19), .D(key1_reg_21__FF_INPUT), .Q(core_key_53_) );
  DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf20), .D(core_mi_reg_63__FF_INPUT), .Q(core_mi_reg_63_) );
  DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf19), .D(core_loop_ctr_reg_0__FF_INPUT), .Q(core_loop_ctr_reg_0_) );
  DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf18), .D(core_loop_ctr_reg_1__FF_INPUT), .Q(core_loop_ctr_reg_1_) );
  DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf17), .D(core_loop_ctr_reg_2__FF_INPUT), .Q(core_loop_ctr_reg_2_) );
  DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf16), .D(core_loop_ctr_reg_3__FF_INPUT), .Q(core_loop_ctr_reg_3_) );
  DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf15), .D(core_ready_reg_FF_INPUT), .Q(core_ready) );
  DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf14), .D(core_siphash_word0_reg_0__FF_INPUT), .Q(core_siphash_word_0_) );
  DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf13), .D(core_siphash_word0_reg_1__FF_INPUT), .Q(core_siphash_word_1_) );
  DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf12), .D(core_siphash_word0_reg_2__FF_INPUT), .Q(core_siphash_word_2_) );
  DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf11), .D(core_siphash_word0_reg_3__FF_INPUT), .Q(core_siphash_word_3_) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf18), .D(key1_reg_22__FF_INPUT), .Q(core_key_54_) );
  DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf10), .D(core_siphash_word0_reg_4__FF_INPUT), .Q(core_siphash_word_4_) );
  DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf9), .D(core_siphash_word0_reg_5__FF_INPUT), .Q(core_siphash_word_5_) );
  DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf8), .D(core_siphash_word0_reg_6__FF_INPUT), .Q(core_siphash_word_6_) );
  DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf7), .D(core_siphash_word0_reg_7__FF_INPUT), .Q(core_siphash_word_7_) );
  DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf6), .D(core_siphash_word0_reg_8__FF_INPUT), .Q(core_siphash_word_8_) );
  DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf5), .D(core_siphash_word0_reg_9__FF_INPUT), .Q(core_siphash_word_9_) );
  DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf4), .D(core_siphash_word0_reg_10__FF_INPUT), .Q(core_siphash_word_10_) );
  DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf3), .D(core_siphash_word0_reg_11__FF_INPUT), .Q(core_siphash_word_11_) );
  DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf2), .D(core_siphash_word0_reg_12__FF_INPUT), .Q(core_siphash_word_12_) );
  DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf1), .D(core_siphash_word0_reg_13__FF_INPUT), .Q(core_siphash_word_13_) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf17), .D(key1_reg_23__FF_INPUT), .Q(core_key_55_) );
  DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf0), .D(core_siphash_word0_reg_14__FF_INPUT), .Q(core_siphash_word_14_) );
  DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_bF_buf84), .D(core_siphash_word0_reg_15__FF_INPUT), .Q(core_siphash_word_15_) );
  DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_bF_buf83), .D(core_siphash_word0_reg_16__FF_INPUT), .Q(core_siphash_word_16_) );
  DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_bF_buf82), .D(core_siphash_word0_reg_17__FF_INPUT), .Q(core_siphash_word_17_) );
  DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_bF_buf81), .D(core_siphash_word0_reg_18__FF_INPUT), .Q(core_siphash_word_18_) );
  DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_bF_buf80), .D(core_siphash_word0_reg_19__FF_INPUT), .Q(core_siphash_word_19_) );
  DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_bF_buf79), .D(core_siphash_word0_reg_20__FF_INPUT), .Q(core_siphash_word_20_) );
  DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_bF_buf78), .D(core_siphash_word0_reg_21__FF_INPUT), .Q(core_siphash_word_21_) );
  DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_bF_buf77), .D(core_siphash_word0_reg_22__FF_INPUT), .Q(core_siphash_word_22_) );
  DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_bF_buf76), .D(core_siphash_word0_reg_23__FF_INPUT), .Q(core_siphash_word_23_) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf16), .D(key1_reg_24__FF_INPUT), .Q(core_key_56_) );
  DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_bF_buf75), .D(core_siphash_word0_reg_24__FF_INPUT), .Q(core_siphash_word_24_) );
  DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_bF_buf74), .D(core_siphash_word0_reg_25__FF_INPUT), .Q(core_siphash_word_25_) );
  DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_bF_buf73), .D(core_siphash_word0_reg_26__FF_INPUT), .Q(core_siphash_word_26_) );
  DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_bF_buf72), .D(core_siphash_word0_reg_27__FF_INPUT), .Q(core_siphash_word_27_) );
  DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_bF_buf71), .D(core_siphash_word0_reg_28__FF_INPUT), .Q(core_siphash_word_28_) );
  DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_bF_buf70), .D(core_siphash_word0_reg_29__FF_INPUT), .Q(core_siphash_word_29_) );
  DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_bF_buf69), .D(core_siphash_word0_reg_30__FF_INPUT), .Q(core_siphash_word_30_) );
  DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_bF_buf68), .D(core_siphash_word0_reg_31__FF_INPUT), .Q(core_siphash_word_31_) );
  DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_bF_buf67), .D(core_siphash_word0_reg_32__FF_INPUT), .Q(core_siphash_word_32_) );
  DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_bF_buf66), .D(core_siphash_word0_reg_33__FF_INPUT), .Q(core_siphash_word_33_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf78), .D(param_reg_2__FF_INPUT), .Q(core_compression_rounds_2_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf15), .D(key1_reg_25__FF_INPUT), .Q(core_key_57_) );
  DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_bF_buf65), .D(core_siphash_word0_reg_34__FF_INPUT), .Q(core_siphash_word_34_) );
  DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_bF_buf64), .D(core_siphash_word0_reg_35__FF_INPUT), .Q(core_siphash_word_35_) );
  DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_bF_buf63), .D(core_siphash_word0_reg_36__FF_INPUT), .Q(core_siphash_word_36_) );
  DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_bF_buf62), .D(core_siphash_word0_reg_37__FF_INPUT), .Q(core_siphash_word_37_) );
  DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_bF_buf61), .D(core_siphash_word0_reg_38__FF_INPUT), .Q(core_siphash_word_38_) );
  DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_bF_buf60), .D(core_siphash_word0_reg_39__FF_INPUT), .Q(core_siphash_word_39_) );
  DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_bF_buf59), .D(core_siphash_word0_reg_40__FF_INPUT), .Q(core_siphash_word_40_) );
  DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_bF_buf58), .D(core_siphash_word0_reg_41__FF_INPUT), .Q(core_siphash_word_41_) );
  DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_bF_buf57), .D(core_siphash_word0_reg_42__FF_INPUT), .Q(core_siphash_word_42_) );
  DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_bF_buf56), .D(core_siphash_word0_reg_43__FF_INPUT), .Q(core_siphash_word_43_) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf14), .D(key1_reg_26__FF_INPUT), .Q(core_key_58_) );
  DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_bF_buf55), .D(core_siphash_word0_reg_44__FF_INPUT), .Q(core_siphash_word_44_) );
  DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_bF_buf54), .D(core_siphash_word0_reg_45__FF_INPUT), .Q(core_siphash_word_45_) );
  DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_bF_buf53), .D(core_siphash_word0_reg_46__FF_INPUT), .Q(core_siphash_word_46_) );
  DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_bF_buf52), .D(core_siphash_word0_reg_47__FF_INPUT), .Q(core_siphash_word_47_) );
  DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_bF_buf51), .D(core_siphash_word0_reg_48__FF_INPUT), .Q(core_siphash_word_48_) );
  DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_bF_buf50), .D(core_siphash_word0_reg_49__FF_INPUT), .Q(core_siphash_word_49_) );
  DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_bF_buf49), .D(core_siphash_word0_reg_50__FF_INPUT), .Q(core_siphash_word_50_) );
  DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_bF_buf48), .D(core_siphash_word0_reg_51__FF_INPUT), .Q(core_siphash_word_51_) );
  DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_bF_buf47), .D(core_siphash_word0_reg_52__FF_INPUT), .Q(core_siphash_word_52_) );
  DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_bF_buf46), .D(core_siphash_word0_reg_53__FF_INPUT), .Q(core_siphash_word_53_) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf13), .D(key1_reg_27__FF_INPUT), .Q(core_key_59_) );
  DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_bF_buf45), .D(core_siphash_word0_reg_54__FF_INPUT), .Q(core_siphash_word_54_) );
  DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_bF_buf44), .D(core_siphash_word0_reg_55__FF_INPUT), .Q(core_siphash_word_55_) );
  DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_bF_buf43), .D(core_siphash_word0_reg_56__FF_INPUT), .Q(core_siphash_word_56_) );
  DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_bF_buf42), .D(core_siphash_word0_reg_57__FF_INPUT), .Q(core_siphash_word_57_) );
  DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_bF_buf41), .D(core_siphash_word0_reg_58__FF_INPUT), .Q(core_siphash_word_58_) );
  DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_bF_buf40), .D(core_siphash_word0_reg_59__FF_INPUT), .Q(core_siphash_word_59_) );
  DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_bF_buf39), .D(core_siphash_word0_reg_60__FF_INPUT), .Q(core_siphash_word_60_) );
  DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_bF_buf38), .D(core_siphash_word0_reg_61__FF_INPUT), .Q(core_siphash_word_61_) );
  DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_bF_buf37), .D(core_siphash_word0_reg_62__FF_INPUT), .Q(core_siphash_word_62_) );
  DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_bF_buf36), .D(core_siphash_word0_reg_63__FF_INPUT), .Q(core_siphash_word_63_) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf12), .D(key1_reg_28__FF_INPUT), .Q(core_key_60_) );
  DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_bF_buf35), .D(core_siphash_word1_reg_0__FF_INPUT), .Q(core_siphash_word_64_) );
  DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_bF_buf34), .D(core_siphash_word1_reg_1__FF_INPUT), .Q(core_siphash_word_65_) );
  DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_bF_buf33), .D(core_siphash_word1_reg_2__FF_INPUT), .Q(core_siphash_word_66_) );
  DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_bF_buf32), .D(core_siphash_word1_reg_3__FF_INPUT), .Q(core_siphash_word_67_) );
  DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_bF_buf31), .D(core_siphash_word1_reg_4__FF_INPUT), .Q(core_siphash_word_68_) );
  DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_bF_buf30), .D(core_siphash_word1_reg_5__FF_INPUT), .Q(core_siphash_word_69_) );
  DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_bF_buf29), .D(core_siphash_word1_reg_6__FF_INPUT), .Q(core_siphash_word_70_) );
  DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_bF_buf28), .D(core_siphash_word1_reg_7__FF_INPUT), .Q(core_siphash_word_71_) );
  DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_bF_buf27), .D(core_siphash_word1_reg_8__FF_INPUT), .Q(core_siphash_word_72_) );
  DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_bF_buf26), .D(core_siphash_word1_reg_9__FF_INPUT), .Q(core_siphash_word_73_) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf11), .D(key1_reg_29__FF_INPUT), .Q(core_key_61_) );
  DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_bF_buf25), .D(core_siphash_word1_reg_10__FF_INPUT), .Q(core_siphash_word_74_) );
  DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_bF_buf24), .D(core_siphash_word1_reg_11__FF_INPUT), .Q(core_siphash_word_75_) );
  DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_bF_buf23), .D(core_siphash_word1_reg_12__FF_INPUT), .Q(core_siphash_word_76_) );
  DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_bF_buf22), .D(core_siphash_word1_reg_13__FF_INPUT), .Q(core_siphash_word_77_) );
  DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_bF_buf21), .D(core_siphash_word1_reg_14__FF_INPUT), .Q(core_siphash_word_78_) );
  DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_bF_buf20), .D(core_siphash_word1_reg_15__FF_INPUT), .Q(core_siphash_word_79_) );
  DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_bF_buf19), .D(core_siphash_word1_reg_16__FF_INPUT), .Q(core_siphash_word_80_) );
  DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_bF_buf18), .D(core_siphash_word1_reg_17__FF_INPUT), .Q(core_siphash_word_81_) );
  DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_bF_buf17), .D(core_siphash_word1_reg_18__FF_INPUT), .Q(core_siphash_word_82_) );
  DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_bF_buf16), .D(core_siphash_word1_reg_19__FF_INPUT), .Q(core_siphash_word_83_) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf10), .D(key1_reg_30__FF_INPUT), .Q(core_key_62_) );
  DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_bF_buf15), .D(core_siphash_word1_reg_20__FF_INPUT), .Q(core_siphash_word_84_) );
  DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_bF_buf14), .D(core_siphash_word1_reg_21__FF_INPUT), .Q(core_siphash_word_85_) );
  DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_bF_buf13), .D(core_siphash_word1_reg_22__FF_INPUT), .Q(core_siphash_word_86_) );
  DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_bF_buf12), .D(core_siphash_word1_reg_23__FF_INPUT), .Q(core_siphash_word_87_) );
  DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_bF_buf11), .D(core_siphash_word1_reg_24__FF_INPUT), .Q(core_siphash_word_88_) );
  DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_bF_buf10), .D(core_siphash_word1_reg_25__FF_INPUT), .Q(core_siphash_word_89_) );
  DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_bF_buf9), .D(core_siphash_word1_reg_26__FF_INPUT), .Q(core_siphash_word_90_) );
  DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_bF_buf8), .D(core_siphash_word1_reg_27__FF_INPUT), .Q(core_siphash_word_91_) );
  DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_bF_buf7), .D(core_siphash_word1_reg_28__FF_INPUT), .Q(core_siphash_word_92_) );
  DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_bF_buf6), .D(core_siphash_word1_reg_29__FF_INPUT), .Q(core_siphash_word_93_) );
  DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf9), .D(key1_reg_31__FF_INPUT), .Q(core_key_63_) );
  DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_bF_buf5), .D(core_siphash_word1_reg_30__FF_INPUT), .Q(core_siphash_word_94_) );
  DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_bF_buf4), .D(core_siphash_word1_reg_31__FF_INPUT), .Q(core_siphash_word_95_) );
  DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_bF_buf3), .D(core_siphash_word1_reg_32__FF_INPUT), .Q(core_siphash_word_96_) );
  DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_bF_buf2), .D(core_siphash_word1_reg_33__FF_INPUT), .Q(core_siphash_word_97_) );
  DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_bF_buf1), .D(core_siphash_word1_reg_34__FF_INPUT), .Q(core_siphash_word_98_) );
  DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_bF_buf0), .D(core_siphash_word1_reg_35__FF_INPUT), .Q(core_siphash_word_99_) );
  DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_bF_buf84), .D(core_siphash_word1_reg_36__FF_INPUT), .Q(core_siphash_word_100_) );
  DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_bF_buf83), .D(core_siphash_word1_reg_37__FF_INPUT), .Q(core_siphash_word_101_) );
  DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_bF_buf82), .D(core_siphash_word1_reg_38__FF_INPUT), .Q(core_siphash_word_102_) );
  DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_bF_buf81), .D(core_siphash_word1_reg_39__FF_INPUT), .Q(core_siphash_word_103_) );
  DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf8), .D(key2_reg_0__FF_INPUT), .Q(core_key_64_) );
  DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_bF_buf80), .D(core_siphash_word1_reg_40__FF_INPUT), .Q(core_siphash_word_104_) );
  DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_bF_buf79), .D(core_siphash_word1_reg_41__FF_INPUT), .Q(core_siphash_word_105_) );
  DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_bF_buf78), .D(core_siphash_word1_reg_42__FF_INPUT), .Q(core_siphash_word_106_) );
  DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_bF_buf77), .D(core_siphash_word1_reg_43__FF_INPUT), .Q(core_siphash_word_107_) );
  DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_bF_buf76), .D(core_siphash_word1_reg_44__FF_INPUT), .Q(core_siphash_word_108_) );
  DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_bF_buf75), .D(core_siphash_word1_reg_45__FF_INPUT), .Q(core_siphash_word_109_) );
  DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_bF_buf74), .D(core_siphash_word1_reg_46__FF_INPUT), .Q(core_siphash_word_110_) );
  DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_bF_buf73), .D(core_siphash_word1_reg_47__FF_INPUT), .Q(core_siphash_word_111_) );
  DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_bF_buf72), .D(core_siphash_word1_reg_48__FF_INPUT), .Q(core_siphash_word_112_) );
  DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_bF_buf71), .D(core_siphash_word1_reg_49__FF_INPUT), .Q(core_siphash_word_113_) );
  DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf7), .D(key2_reg_1__FF_INPUT), .Q(core_key_65_) );
  DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_bF_buf70), .D(core_siphash_word1_reg_50__FF_INPUT), .Q(core_siphash_word_114_) );
  DFFPOSX1 DFFPOSX1_781 ( .CLK(clk_bF_buf69), .D(core_siphash_word1_reg_51__FF_INPUT), .Q(core_siphash_word_115_) );
  DFFPOSX1 DFFPOSX1_782 ( .CLK(clk_bF_buf68), .D(core_siphash_word1_reg_52__FF_INPUT), .Q(core_siphash_word_116_) );
  DFFPOSX1 DFFPOSX1_783 ( .CLK(clk_bF_buf67), .D(core_siphash_word1_reg_53__FF_INPUT), .Q(core_siphash_word_117_) );
  DFFPOSX1 DFFPOSX1_784 ( .CLK(clk_bF_buf66), .D(core_siphash_word1_reg_54__FF_INPUT), .Q(core_siphash_word_118_) );
  DFFPOSX1 DFFPOSX1_785 ( .CLK(clk_bF_buf65), .D(core_siphash_word1_reg_55__FF_INPUT), .Q(core_siphash_word_119_) );
  DFFPOSX1 DFFPOSX1_786 ( .CLK(clk_bF_buf64), .D(core_siphash_word1_reg_56__FF_INPUT), .Q(core_siphash_word_120_) );
  DFFPOSX1 DFFPOSX1_787 ( .CLK(clk_bF_buf63), .D(core_siphash_word1_reg_57__FF_INPUT), .Q(core_siphash_word_121_) );
  DFFPOSX1 DFFPOSX1_788 ( .CLK(clk_bF_buf62), .D(core_siphash_word1_reg_58__FF_INPUT), .Q(core_siphash_word_122_) );
  DFFPOSX1 DFFPOSX1_789 ( .CLK(clk_bF_buf61), .D(core_siphash_word1_reg_59__FF_INPUT), .Q(core_siphash_word_123_) );
  DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf6), .D(key2_reg_2__FF_INPUT), .Q(core_key_66_) );
  DFFPOSX1 DFFPOSX1_790 ( .CLK(clk_bF_buf60), .D(core_siphash_word1_reg_60__FF_INPUT), .Q(core_siphash_word_124_) );
  DFFPOSX1 DFFPOSX1_791 ( .CLK(clk_bF_buf59), .D(core_siphash_word1_reg_61__FF_INPUT), .Q(core_siphash_word_125_) );
  DFFPOSX1 DFFPOSX1_792 ( .CLK(clk_bF_buf58), .D(core_siphash_word1_reg_62__FF_INPUT), .Q(core_siphash_word_126_) );
  DFFPOSX1 DFFPOSX1_793 ( .CLK(clk_bF_buf57), .D(core_siphash_word1_reg_63__FF_INPUT), .Q(core_siphash_word_127_) );
  DFFPOSX1 DFFPOSX1_794 ( .CLK(clk_bF_buf56), .D(core_siphash_valid_reg_FF_INPUT), .Q(core_siphash_valid_reg) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf77), .D(param_reg_3__FF_INPUT), .Q(core_compression_rounds_3_) );
  DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf5), .D(key2_reg_3__FF_INPUT), .Q(core_key_67_) );
  DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf4), .D(key2_reg_4__FF_INPUT), .Q(core_key_68_) );
  DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf3), .D(key2_reg_5__FF_INPUT), .Q(core_key_69_) );
  DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf2), .D(key2_reg_6__FF_INPUT), .Q(core_key_70_) );
  DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf1), .D(key2_reg_7__FF_INPUT), .Q(core_key_71_) );
  DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf0), .D(key2_reg_8__FF_INPUT), .Q(core_key_72_) );
  DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf84), .D(key2_reg_9__FF_INPUT), .Q(core_key_73_) );
  DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf83), .D(key2_reg_10__FF_INPUT), .Q(core_key_74_) );
  DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf82), .D(key2_reg_11__FF_INPUT), .Q(core_key_75_) );
  DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf81), .D(key2_reg_12__FF_INPUT), .Q(core_key_76_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf76), .D(param_reg_4__FF_INPUT), .Q(core_final_rounds_0_) );
  DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf80), .D(key2_reg_13__FF_INPUT), .Q(core_key_77_) );
  DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf79), .D(key2_reg_14__FF_INPUT), .Q(core_key_78_) );
  DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf78), .D(key2_reg_15__FF_INPUT), .Q(core_key_79_) );
  DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf77), .D(key2_reg_16__FF_INPUT), .Q(core_key_80_) );
  DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf76), .D(key2_reg_17__FF_INPUT), .Q(core_key_81_) );
  DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf75), .D(key2_reg_18__FF_INPUT), .Q(core_key_82_) );
  DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf74), .D(key2_reg_19__FF_INPUT), .Q(core_key_83_) );
  DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf73), .D(key2_reg_20__FF_INPUT), .Q(core_key_84_) );
  DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf72), .D(key2_reg_21__FF_INPUT), .Q(core_key_85_) );
  DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf71), .D(key2_reg_22__FF_INPUT), .Q(core_key_86_) );
  INVX1 INVX1_1 ( .A(\addr[2] ), .Y(_abc_19068_n870_1) );
  INVX1 INVX1_10 ( .A(_abc_19068_n2136), .Y(_abc_19068_n2137) );
  INVX1 INVX1_100 ( .A(_abc_19068_n2619), .Y(_abc_19068_n2620) );
  INVX1 INVX1_1000 ( .A(core_key_85_), .Y(core__abc_21380_n4736) );
  INVX1 INVX1_1001 ( .A(core__abc_21380_n4739), .Y(core__abc_21380_n4740) );
  INVX1 INVX1_1002 ( .A(core__abc_21380_n4722_1), .Y(core__abc_21380_n4751) );
  INVX1 INVX1_1003 ( .A(core__abc_21380_n4756), .Y(core__abc_21380_n4757_1) );
  INVX1 INVX1_1004 ( .A(core__abc_21380_n4760), .Y(core__abc_21380_n4761) );
  INVX1 INVX1_1005 ( .A(core__abc_21380_n4764), .Y(core__abc_21380_n4765) );
  INVX1 INVX1_1006 ( .A(core__abc_21380_n4767_1), .Y(core__abc_21380_n4768) );
  INVX1 INVX1_1007 ( .A(core__abc_21380_n4771), .Y(core__abc_21380_n4772_1) );
  INVX1 INVX1_1008 ( .A(core__abc_21380_n4775), .Y(core__abc_21380_n4776) );
  INVX1 INVX1_1009 ( .A(core__abc_21380_n4781), .Y(core__abc_21380_n4782) );
  INVX1 INVX1_101 ( .A(_abc_19068_n2624), .Y(_abc_19068_n2625) );
  INVX1 INVX1_1010 ( .A(core__abc_21380_n4783_1), .Y(core__abc_21380_n4784) );
  INVX1 INVX1_1011 ( .A(core_key_86_), .Y(core__abc_21380_n4789) );
  INVX1 INVX1_1012 ( .A(core__abc_21380_n4792), .Y(core__abc_21380_n4793_1) );
  INVX1 INVX1_1013 ( .A(core__abc_21380_n4777_1), .Y(core__abc_21380_n4802) );
  INVX1 INVX1_1014 ( .A(core__abc_21380_n4803_1), .Y(core__abc_21380_n4804) );
  INVX1 INVX1_1015 ( .A(core__abc_21380_n4805), .Y(core__abc_21380_n4806) );
  INVX1 INVX1_1016 ( .A(core__abc_21380_n4810), .Y(core__abc_21380_n4811) );
  INVX1 INVX1_1017 ( .A(core__abc_21380_n4816), .Y(core__abc_21380_n4817) );
  INVX1 INVX1_1018 ( .A(core__abc_21380_n4807), .Y(core__abc_21380_n4820_1) );
  INVX1 INVX1_1019 ( .A(core__abc_21380_n4808_1), .Y(core__abc_21380_n4821) );
  INVX1 INVX1_102 ( .A(_abc_19068_n2629), .Y(_abc_19068_n2630) );
  INVX1 INVX1_1020 ( .A(core__abc_21380_n4815), .Y(core__abc_21380_n4823) );
  INVX1 INVX1_1021 ( .A(core__abc_21380_n4832), .Y(core__abc_21380_n4834) );
  INVX1 INVX1_1022 ( .A(core__abc_21380_n4840_1), .Y(core__abc_21380_n4841) );
  INVX1 INVX1_1023 ( .A(core__abc_21380_n4749), .Y(core__abc_21380_n4850) );
  INVX1 INVX1_1024 ( .A(core__abc_21380_n4779), .Y(core__abc_21380_n4851_1) );
  INVX1 INVX1_1025 ( .A(core__abc_21380_n4854), .Y(core__abc_21380_n4855) );
  INVX1 INVX1_1026 ( .A(core__abc_21380_n4862_1), .Y(core__abc_21380_n4863) );
  INVX1 INVX1_1027 ( .A(core__abc_21380_n4866), .Y(core__abc_21380_n4867_1) );
  INVX1 INVX1_1028 ( .A(core__abc_21380_n4870), .Y(core__abc_21380_n4871) );
  INVX1 INVX1_1029 ( .A(core__abc_21380_n4878_1), .Y(core__abc_21380_n4879) );
  INVX1 INVX1_103 ( .A(_abc_19068_n2634), .Y(_abc_19068_n2635) );
  INVX1 INVX1_1030 ( .A(core__abc_21380_n4885), .Y(core__abc_21380_n4886) );
  INVX1 INVX1_1031 ( .A(core_v3_reg_8_), .Y(core__abc_21380_n4887) );
  INVX1 INVX1_1032 ( .A(core__abc_21380_n3094), .Y(core__abc_21380_n4888_1) );
  INVX1 INVX1_1033 ( .A(core__abc_21380_n3074), .Y(core__abc_21380_n4889) );
  INVX1 INVX1_1034 ( .A(core__abc_21380_n4891), .Y(core__abc_21380_n4893_1) );
  INVX1 INVX1_1035 ( .A(core__abc_21380_n4895), .Y(core__abc_21380_n4896_1) );
  INVX1 INVX1_1036 ( .A(core__abc_21380_n4899), .Y(core__abc_21380_n4900_1) );
  INVX1 INVX1_1037 ( .A(core__abc_21380_n4903), .Y(core__abc_21380_n4904) );
  INVX1 INVX1_1038 ( .A(core__abc_21380_n4907), .Y(core__abc_21380_n4908) );
  INVX1 INVX1_1039 ( .A(core_key_88_), .Y(core__abc_21380_n4913) );
  INVX1 INVX1_104 ( .A(_abc_19068_n2639), .Y(_abc_19068_n2640) );
  INVX1 INVX1_1040 ( .A(core__abc_21380_n4916), .Y(core__abc_21380_n4917) );
  INVX1 INVX1_1041 ( .A(core__abc_21380_n4901), .Y(core__abc_21380_n4926) );
  INVX1 INVX1_1042 ( .A(core__abc_21380_n4905), .Y(core__abc_21380_n4927) );
  INVX1 INVX1_1043 ( .A(core__abc_21380_n4930), .Y(core__abc_21380_n4931) );
  INVX1 INVX1_1044 ( .A(core_v3_reg_9_), .Y(core__abc_21380_n4937) );
  INVX1 INVX1_1045 ( .A(core__abc_21380_n4938), .Y(core__abc_21380_n4939) );
  INVX1 INVX1_1046 ( .A(core__abc_21380_n4942), .Y(core__abc_21380_n4944) );
  INVX1 INVX1_1047 ( .A(core__abc_21380_n4948), .Y(core__abc_21380_n4949) );
  INVX1 INVX1_1048 ( .A(core__abc_21380_n4928), .Y(core__abc_21380_n4952) );
  INVX1 INVX1_1049 ( .A(core__abc_21380_n4950), .Y(core__abc_21380_n4953) );
  INVX1 INVX1_105 ( .A(_abc_19068_n2644), .Y(_abc_19068_n2645) );
  INVX1 INVX1_1050 ( .A(core__abc_21380_n4955), .Y(core__abc_21380_n4956) );
  INVX1 INVX1_1051 ( .A(core__abc_21380_n4963), .Y(core__abc_21380_n4964) );
  INVX1 INVX1_1052 ( .A(core__abc_21380_n4974), .Y(core__abc_21380_n4976) );
  INVX1 INVX1_1053 ( .A(core__abc_21380_n4978), .Y(core__abc_21380_n4979) );
  INVX1 INVX1_1054 ( .A(core_v3_reg_10_), .Y(core__abc_21380_n4980) );
  INVX1 INVX1_1055 ( .A(core__abc_21380_n4982), .Y(core__abc_21380_n4983) );
  INVX1 INVX1_1056 ( .A(core__abc_21380_n4986), .Y(core__abc_21380_n4987) );
  INVX1 INVX1_1057 ( .A(core__abc_21380_n4990), .Y(core__abc_21380_n4991) );
  INVX1 INVX1_1058 ( .A(core__abc_21380_n4997), .Y(core__abc_21380_n4998) );
  INVX1 INVX1_1059 ( .A(core__abc_21380_n5002), .Y(core__abc_21380_n5003) );
  INVX1 INVX1_106 ( .A(_abc_19068_n2650), .Y(_abc_19068_n2651) );
  INVX1 INVX1_1060 ( .A(core__abc_21380_n5004), .Y(core__abc_21380_n5006) );
  INVX1 INVX1_1061 ( .A(core__abc_21380_n5012), .Y(core__abc_21380_n5013) );
  INVX1 INVX1_1062 ( .A(core__abc_21380_n3697), .Y(core__abc_21380_n5022) );
  INVX1 INVX1_1063 ( .A(core__abc_21380_n4992), .Y(core__abc_21380_n5023) );
  INVX1 INVX1_1064 ( .A(core__abc_21380_n5025), .Y(core__abc_21380_n5026) );
  INVX1 INVX1_1065 ( .A(core__abc_21380_n5027), .Y(core__abc_21380_n5028) );
  INVX1 INVX1_1066 ( .A(core__abc_21380_n5029), .Y(core__abc_21380_n5030) );
  INVX1 INVX1_1067 ( .A(core_v3_reg_11_), .Y(core__abc_21380_n5032) );
  INVX1 INVX1_1068 ( .A(core__abc_21380_n5033), .Y(core__abc_21380_n5034) );
  INVX1 INVX1_1069 ( .A(core__abc_21380_n5038), .Y(core__abc_21380_n5039) );
  INVX1 INVX1_107 ( .A(_abc_19068_n2655), .Y(_abc_19068_n2656) );
  INVX1 INVX1_1070 ( .A(core__abc_21380_n5040), .Y(core__abc_21380_n5044) );
  INVX1 INVX1_1071 ( .A(core__abc_21380_n5024), .Y(core__abc_21380_n5049) );
  INVX1 INVX1_1072 ( .A(core__abc_21380_n5054), .Y(core__abc_21380_n5056) );
  INVX1 INVX1_1073 ( .A(core_key_91_), .Y(core__abc_21380_n5060) );
  INVX1 INVX1_1074 ( .A(core__abc_21380_n5063), .Y(core__abc_21380_n5064) );
  INVX1 INVX1_1075 ( .A(core__abc_21380_n4996), .Y(core__abc_21380_n5073) );
  INVX1 INVX1_1076 ( .A(core__abc_21380_n4994), .Y(core__abc_21380_n5074) );
  INVX1 INVX1_1077 ( .A(core__abc_21380_n5082), .Y(core__abc_21380_n5083) );
  INVX1 INVX1_1078 ( .A(core__abc_21380_n5085), .Y(core__abc_21380_n5093) );
  INVX1 INVX1_1079 ( .A(core__abc_21380_n5090), .Y(core__abc_21380_n5095) );
  INVX1 INVX1_108 ( .A(_abc_19068_n2660), .Y(_abc_19068_n2661) );
  INVX1 INVX1_1080 ( .A(core__abc_21380_n5098), .Y(core__abc_21380_n5099) );
  INVX1 INVX1_1081 ( .A(core_v3_reg_12_), .Y(core__abc_21380_n5100) );
  INVX1 INVX1_1082 ( .A(core__abc_21380_n3102), .Y(core__abc_21380_n5101) );
  INVX1 INVX1_1083 ( .A(core__abc_21380_n3066), .Y(core__abc_21380_n5102) );
  INVX1 INVX1_1084 ( .A(core__abc_21380_n5104), .Y(core__abc_21380_n5105) );
  INVX1 INVX1_1085 ( .A(core__abc_21380_n5108), .Y(core__abc_21380_n5109) );
  INVX1 INVX1_1086 ( .A(core__abc_21380_n5112), .Y(core__abc_21380_n5113) );
  INVX1 INVX1_1087 ( .A(core__abc_21380_n5116), .Y(core__abc_21380_n5118) );
  INVX1 INVX1_1088 ( .A(core__abc_21380_n5120), .Y(core__abc_21380_n5122) );
  INVX1 INVX1_1089 ( .A(core_key_92_), .Y(core__abc_21380_n5126) );
  INVX1 INVX1_109 ( .A(_abc_19068_n2665), .Y(_abc_19068_n2666) );
  INVX1 INVX1_1090 ( .A(core__abc_21380_n5129), .Y(core__abc_21380_n5130) );
  INVX1 INVX1_1091 ( .A(core__abc_21380_n5119), .Y(core__abc_21380_n5139) );
  INVX1 INVX1_1092 ( .A(core__abc_21380_n5114), .Y(core__abc_21380_n5140) );
  INVX1 INVX1_1093 ( .A(core__abc_21380_n5146), .Y(core__abc_21380_n5147) );
  INVX1 INVX1_1094 ( .A(core__abc_21380_n5148), .Y(core__abc_21380_n5149) );
  INVX1 INVX1_1095 ( .A(core_v3_reg_13_), .Y(core__abc_21380_n5150) );
  INVX1 INVX1_1096 ( .A(core__abc_21380_n5151), .Y(core__abc_21380_n5152) );
  INVX1 INVX1_1097 ( .A(core__abc_21380_n5156), .Y(core__abc_21380_n5157) );
  INVX1 INVX1_1098 ( .A(core__abc_21380_n5158), .Y(core__abc_21380_n5161) );
  INVX1 INVX1_1099 ( .A(core__abc_21380_n5166), .Y(core__abc_21380_n5167) );
  INVX1 INVX1_11 ( .A(_abc_19068_n2142), .Y(_abc_19068_n2143) );
  INVX1 INVX1_110 ( .A(_abc_19068_n2670), .Y(_abc_19068_n2671) );
  INVX1 INVX1_1100 ( .A(core__abc_21380_n5173), .Y(core__abc_21380_n5174) );
  INVX1 INVX1_1101 ( .A(core__abc_21380_n5176), .Y(core__abc_21380_n5178) );
  INVX1 INVX1_1102 ( .A(core_key_93_), .Y(core__abc_21380_n5182) );
  INVX1 INVX1_1103 ( .A(core__abc_21380_n5185), .Y(core__abc_21380_n5186) );
  INVX1 INVX1_1104 ( .A(core__abc_21380_n3900), .Y(core__abc_21380_n5195) );
  INVX1 INVX1_1105 ( .A(core__abc_21380_n5142), .Y(core__abc_21380_n5198) );
  INVX1 INVX1_1106 ( .A(core__abc_21380_n5200), .Y(core__abc_21380_n5201) );
  INVX1 INVX1_1107 ( .A(core__abc_21380_n5206), .Y(core__abc_21380_n5207) );
  INVX1 INVX1_1108 ( .A(core__abc_21380_n3062), .Y(core__abc_21380_n5208) );
  INVX1 INVX1_1109 ( .A(core__abc_21380_n5212), .Y(core__abc_21380_n5213) );
  INVX1 INVX1_111 ( .A(_abc_19068_n2675), .Y(_abc_19068_n2676) );
  INVX1 INVX1_1110 ( .A(core__abc_21380_n5214), .Y(core__abc_21380_n5215) );
  INVX1 INVX1_1111 ( .A(core_v3_reg_14_), .Y(core__abc_21380_n5217) );
  INVX1 INVX1_1112 ( .A(core__abc_21380_n5219), .Y(core__abc_21380_n5221) );
  INVX1 INVX1_1113 ( .A(core__abc_21380_n5225), .Y(core__abc_21380_n5226) );
  INVX1 INVX1_1114 ( .A(core__abc_21380_n5227), .Y(core__abc_21380_n5228) );
  INVX1 INVX1_1115 ( .A(core_key_94_), .Y(core__abc_21380_n5233) );
  INVX1 INVX1_1116 ( .A(core__abc_21380_n5236), .Y(core__abc_21380_n5237) );
  INVX1 INVX1_1117 ( .A(core__abc_21380_n5220), .Y(core__abc_21380_n5246) );
  INVX1 INVX1_1118 ( .A(core__abc_21380_n5247), .Y(core__abc_21380_n5248) );
  INVX1 INVX1_1119 ( .A(core__abc_21380_n2415), .Y(core__abc_21380_n5249) );
  INVX1 INVX1_112 ( .A(_abc_19068_n2680), .Y(_abc_19068_n2681) );
  INVX1 INVX1_1120 ( .A(core_v3_reg_15_), .Y(core__abc_21380_n5256) );
  INVX1 INVX1_1121 ( .A(core__abc_21380_n5259), .Y(core__abc_21380_n5260) );
  INVX1 INVX1_1122 ( .A(core__abc_21380_n5258), .Y(core__abc_21380_n5263) );
  INVX1 INVX1_1123 ( .A(core__abc_21380_n5265), .Y(core__abc_21380_n5272) );
  INVX1 INVX1_1124 ( .A(core__abc_21380_n5281), .Y(core__abc_21380_n5283) );
  INVX1 INVX1_1125 ( .A(core__abc_21380_n5289), .Y(core__abc_21380_n5290) );
  INVX1 INVX1_1126 ( .A(core__abc_21380_n5080), .Y(core__abc_21380_n5299) );
  INVX1 INVX1_1127 ( .A(core__abc_21380_n5172), .Y(core__abc_21380_n5300) );
  INVX1 INVX1_1128 ( .A(core__abc_21380_n5078), .Y(core__abc_21380_n5308) );
  INVX1 INVX1_1129 ( .A(core__abc_21380_n5267), .Y(core__abc_21380_n5312) );
  INVX1 INVX1_113 ( .A(_abc_19068_n2685), .Y(_abc_19068_n2686) );
  INVX1 INVX1_1130 ( .A(core__abc_21380_n5314), .Y(core__abc_21380_n5315) );
  INVX1 INVX1_1131 ( .A(core_v3_reg_16_), .Y(core__abc_21380_n5320) );
  INVX1 INVX1_1132 ( .A(core__abc_21380_n3115), .Y(core__abc_21380_n5321) );
  INVX1 INVX1_1133 ( .A(core__abc_21380_n5324), .Y(core__abc_21380_n5325) );
  INVX1 INVX1_1134 ( .A(core__abc_21380_n5328), .Y(core__abc_21380_n5329) );
  INVX1 INVX1_1135 ( .A(core__abc_21380_n5223), .Y(core__abc_21380_n5335) );
  INVX1 INVX1_1136 ( .A(core__abc_21380_n4753), .Y(core__abc_21380_n5341) );
  INVX1 INVX1_1137 ( .A(core__abc_21380_n5332), .Y(core__abc_21380_n5354) );
  INVX1 INVX1_1138 ( .A(core__abc_21380_n5356), .Y(core__abc_21380_n5358) );
  INVX1 INVX1_1139 ( .A(core__abc_21380_n5364), .Y(core__abc_21380_n5365) );
  INVX1 INVX1_114 ( .A(_abc_19068_n2690), .Y(_abc_19068_n2691) );
  INVX1 INVX1_1140 ( .A(core__abc_21380_n5375), .Y(core__abc_21380_n5376) );
  INVX1 INVX1_1141 ( .A(core_v3_reg_17_), .Y(core__abc_21380_n5377) );
  INVX1 INVX1_1142 ( .A(core__abc_21380_n5378), .Y(core__abc_21380_n5379) );
  INVX1 INVX1_1143 ( .A(core__abc_21380_n5382), .Y(core__abc_21380_n5384) );
  INVX1 INVX1_1144 ( .A(core__abc_21380_n5386), .Y(core__abc_21380_n5387) );
  INVX1 INVX1_1145 ( .A(core__abc_21380_n5330), .Y(core__abc_21380_n5391) );
  INVX1 INVX1_1146 ( .A(core__abc_21380_n5355), .Y(core__abc_21380_n5392) );
  INVX1 INVX1_1147 ( .A(core__abc_21380_n5395), .Y(core__abc_21380_n5396) );
  INVX1 INVX1_1148 ( .A(core__abc_21380_n5397), .Y(core__abc_21380_n5398) );
  INVX1 INVX1_1149 ( .A(core_key_97_), .Y(core__abc_21380_n5403) );
  INVX1 INVX1_115 ( .A(_abc_19068_n2695), .Y(_abc_19068_n2696) );
  INVX1 INVX1_1150 ( .A(core__abc_21380_n5406), .Y(core__abc_21380_n5407) );
  INVX1 INVX1_1151 ( .A(core__abc_21380_n5390), .Y(core__abc_21380_n5416) );
  INVX1 INVX1_1152 ( .A(core__abc_21380_n5418), .Y(core__abc_21380_n5419) );
  INVX1 INVX1_1153 ( .A(core__abc_21380_n5421), .Y(core__abc_21380_n5422) );
  INVX1 INVX1_1154 ( .A(core__abc_21380_n5426), .Y(core__abc_21380_n5427) );
  INVX1 INVX1_1155 ( .A(core_v3_reg_18_), .Y(core__abc_21380_n5428) );
  INVX1 INVX1_1156 ( .A(core__abc_21380_n3119), .Y(core__abc_21380_n5429) );
  INVX1 INVX1_1157 ( .A(core__abc_21380_n5433), .Y(core__abc_21380_n5434) );
  INVX1 INVX1_1158 ( .A(core__abc_21380_n5435), .Y(core__abc_21380_n5436) );
  INVX1 INVX1_1159 ( .A(core__abc_21380_n5439), .Y(core__abc_21380_n5440) );
  INVX1 INVX1_116 ( .A(_abc_19068_n2700), .Y(_abc_19068_n2701) );
  INVX1 INVX1_1160 ( .A(core__abc_21380_n5445), .Y(core__abc_21380_n5446) );
  INVX1 INVX1_1161 ( .A(core__abc_21380_n5447), .Y(core__abc_21380_n5449) );
  INVX1 INVX1_1162 ( .A(core__abc_21380_n5455), .Y(core__abc_21380_n5456) );
  INVX1 INVX1_1163 ( .A(core__abc_21380_n5441), .Y(core__abc_21380_n5465) );
  INVX1 INVX1_1164 ( .A(core__abc_21380_n5466), .Y(core__abc_21380_n5467) );
  INVX1 INVX1_1165 ( .A(core__abc_21380_n5468), .Y(core__abc_21380_n5469) );
  INVX1 INVX1_1166 ( .A(core__abc_21380_n5472), .Y(core__abc_21380_n5473) );
  INVX1 INVX1_1167 ( .A(core_v3_reg_19_), .Y(core__abc_21380_n5474) );
  INVX1 INVX1_1168 ( .A(core__abc_21380_n5476), .Y(core__abc_21380_n5477) );
  INVX1 INVX1_1169 ( .A(core__abc_21380_n5479), .Y(core__abc_21380_n5480) );
  INVX1 INVX1_117 ( .A(_abc_19068_n2705), .Y(_abc_19068_n2706) );
  INVX1 INVX1_1170 ( .A(core__abc_21380_n5483), .Y(core__abc_21380_n5484) );
  INVX1 INVX1_1171 ( .A(core__abc_21380_n5487), .Y(core__abc_21380_n5488) );
  INVX1 INVX1_1172 ( .A(core__abc_21380_n5491), .Y(core__abc_21380_n5493) );
  INVX1 INVX1_1173 ( .A(core__abc_21380_n5499), .Y(core__abc_21380_n5500) );
  INVX1 INVX1_1174 ( .A(core__abc_21380_n5509), .Y(core__abc_21380_n5510) );
  INVX1 INVX1_1175 ( .A(core__abc_21380_n5485), .Y(core__abc_21380_n5512) );
  INVX1 INVX1_1176 ( .A(core__abc_21380_n5514), .Y(core__abc_21380_n5515) );
  INVX1 INVX1_1177 ( .A(core__abc_21380_n5522), .Y(core__abc_21380_n5523) );
  INVX1 INVX1_1178 ( .A(core_v3_reg_20_), .Y(core__abc_21380_n5524) );
  INVX1 INVX1_1179 ( .A(core__abc_21380_n5526), .Y(core__abc_21380_n5528) );
  INVX1 INVX1_118 ( .A(_abc_19068_n2710), .Y(_abc_19068_n2711) );
  INVX1 INVX1_1180 ( .A(core__abc_21380_n5530), .Y(core__abc_21380_n5531) );
  INVX1 INVX1_1181 ( .A(core__abc_21380_n5534), .Y(core__abc_21380_n5535) );
  INVX1 INVX1_1182 ( .A(core__abc_21380_n5538), .Y(core__abc_21380_n5539) );
  INVX1 INVX1_1183 ( .A(core__abc_21380_n5519), .Y(core__abc_21380_n5541) );
  INVX1 INVX1_1184 ( .A(core__abc_21380_n5543), .Y(core__abc_21380_n5545) );
  INVX1 INVX1_1185 ( .A(core__abc_21380_n5551), .Y(core__abc_21380_n5552) );
  INVX1 INVX1_1186 ( .A(core__abc_21380_n5562), .Y(core__abc_21380_n5563) );
  INVX1 INVX1_1187 ( .A(core__abc_21380_n5566), .Y(core__abc_21380_n5567) );
  INVX1 INVX1_1188 ( .A(core__abc_21380_n5568), .Y(core__abc_21380_n5569) );
  INVX1 INVX1_1189 ( .A(core__abc_21380_n5573), .Y(core__abc_21380_n5574) );
  INVX1 INVX1_119 ( .A(_abc_19068_n2715), .Y(_abc_19068_n2716) );
  INVX1 INVX1_1190 ( .A(core__abc_21380_n5576), .Y(core__abc_21380_n5577) );
  INVX1 INVX1_1191 ( .A(core__abc_21380_n5578), .Y(core__abc_21380_n5579) );
  INVX1 INVX1_1192 ( .A(core__abc_21380_n5580), .Y(core__abc_21380_n5581) );
  INVX1 INVX1_1193 ( .A(core__abc_21380_n5561), .Y(core__abc_21380_n5584) );
  INVX1 INVX1_1194 ( .A(core__abc_21380_n5582), .Y(core__abc_21380_n5585) );
  INVX1 INVX1_1195 ( .A(core__abc_21380_n5587), .Y(core__abc_21380_n5588) );
  INVX1 INVX1_1196 ( .A(core_key_101_), .Y(core__abc_21380_n5593) );
  INVX1 INVX1_1197 ( .A(core__abc_21380_n5596), .Y(core__abc_21380_n5597) );
  INVX1 INVX1_1198 ( .A(core__abc_21380_n5610), .Y(core__abc_21380_n5611) );
  INVX1 INVX1_1199 ( .A(core__abc_21380_n5614), .Y(core__abc_21380_n5615) );
  INVX1 INVX1_12 ( .A(_abc_19068_n2148), .Y(_abc_19068_n2149) );
  INVX1 INVX1_120 ( .A(_abc_19068_n2720), .Y(_abc_19068_n2721) );
  INVX1 INVX1_1200 ( .A(core__abc_21380_n5619), .Y(core__abc_21380_n5620) );
  INVX1 INVX1_1201 ( .A(core__abc_21380_n5623), .Y(core__abc_21380_n5624) );
  INVX1 INVX1_1202 ( .A(core_v3_reg_22_), .Y(core__abc_21380_n5626) );
  INVX1 INVX1_1203 ( .A(core__abc_21380_n5617), .Y(core__abc_21380_n5630) );
  INVX1 INVX1_1204 ( .A(core__abc_21380_n5628), .Y(core__abc_21380_n5631) );
  INVX1 INVX1_1205 ( .A(core__abc_21380_n5633), .Y(core__abc_21380_n5635) );
  INVX1 INVX1_1206 ( .A(core__abc_21380_n5637), .Y(core__abc_21380_n5639) );
  INVX1 INVX1_1207 ( .A(core_key_102_), .Y(core__abc_21380_n5643) );
  INVX1 INVX1_1208 ( .A(core__abc_21380_n5646), .Y(core__abc_21380_n5647) );
  INVX1 INVX1_1209 ( .A(core__abc_21380_n1376), .Y(core__abc_21380_n5657) );
  INVX1 INVX1_121 ( .A(_abc_19068_n2725), .Y(_abc_19068_n2726) );
  INVX1 INVX1_1210 ( .A(core__abc_21380_n5659), .Y(core__abc_21380_n5660) );
  INVX1 INVX1_1211 ( .A(core_v3_reg_23_), .Y(core__abc_21380_n5663) );
  INVX1 INVX1_1212 ( .A(core__abc_21380_n5664), .Y(core__abc_21380_n5665) );
  INVX1 INVX1_1213 ( .A(core__abc_21380_n5669), .Y(core__abc_21380_n5670) );
  INVX1 INVX1_1214 ( .A(core__abc_21380_n5673), .Y(core__abc_21380_n5674) );
  INVX1 INVX1_1215 ( .A(core__abc_21380_n5656), .Y(core__abc_21380_n5678) );
  INVX1 INVX1_1216 ( .A(core__abc_21380_n5662), .Y(core__abc_21380_n5679) );
  INVX1 INVX1_1217 ( .A(core__abc_21380_n5671), .Y(core__abc_21380_n5680) );
  INVX1 INVX1_1218 ( .A(core__abc_21380_n5685), .Y(core__abc_21380_n5687) );
  INVX1 INVX1_1219 ( .A(core__abc_21380_n5693), .Y(core__abc_21380_n5694) );
  INVX1 INVX1_122 ( .A(_abc_19068_n2730), .Y(_abc_19068_n2731) );
  INVX1 INVX1_1220 ( .A(core__abc_21380_n5716), .Y(core__abc_21380_n5717) );
  INVX1 INVX1_1221 ( .A(core_v3_reg_24_), .Y(core__abc_21380_n5718) );
  INVX1 INVX1_1222 ( .A(core__abc_21380_n5721), .Y(core__abc_21380_n5722) );
  INVX1 INVX1_1223 ( .A(core__abc_21380_n5725), .Y(core__abc_21380_n5726) );
  INVX1 INVX1_1224 ( .A(core__abc_21380_n5729), .Y(core__abc_21380_n5730) );
  INVX1 INVX1_1225 ( .A(core__abc_21380_n5713), .Y(core__abc_21380_n5732) );
  INVX1 INVX1_1226 ( .A(core__abc_21380_n5734), .Y(core__abc_21380_n5735) );
  INVX1 INVX1_1227 ( .A(core__abc_21380_n5742), .Y(core__abc_21380_n5743) );
  INVX1 INVX1_1228 ( .A(core__abc_21380_n5727), .Y(core__abc_21380_n5752) );
  INVX1 INVX1_1229 ( .A(core__abc_21380_n5731), .Y(core__abc_21380_n5753) );
  INVX1 INVX1_123 ( .A(_abc_19068_n2735), .Y(_abc_19068_n2736) );
  INVX1 INVX1_1230 ( .A(core__abc_21380_n5755), .Y(core__abc_21380_n5756) );
  INVX1 INVX1_1231 ( .A(core__abc_21380_n5759), .Y(core__abc_21380_n5760) );
  INVX1 INVX1_1232 ( .A(core_v3_reg_25_), .Y(core__abc_21380_n5761) );
  INVX1 INVX1_1233 ( .A(core__abc_21380_n5762), .Y(core__abc_21380_n5763) );
  INVX1 INVX1_1234 ( .A(core__abc_21380_n5766), .Y(core__abc_21380_n5768) );
  INVX1 INVX1_1235 ( .A(core__abc_21380_n5770), .Y(core__abc_21380_n5771) );
  INVX1 INVX1_1236 ( .A(core__abc_21380_n5772), .Y(core__abc_21380_n5773) );
  INVX1 INVX1_1237 ( .A(core__abc_21380_n5774), .Y(core__abc_21380_n5775) );
  INVX1 INVX1_1238 ( .A(core__abc_21380_n5754), .Y(core__abc_21380_n5778) );
  INVX1 INVX1_1239 ( .A(core__abc_21380_n5776), .Y(core__abc_21380_n5779) );
  INVX1 INVX1_124 ( .A(_abc_19068_n2740), .Y(_abc_19068_n2741) );
  INVX1 INVX1_1240 ( .A(core__abc_21380_n5781), .Y(core__abc_21380_n5782) );
  INVX1 INVX1_1241 ( .A(core__abc_21380_n5789), .Y(core__abc_21380_n5790) );
  INVX1 INVX1_1242 ( .A(core__abc_21380_n5801), .Y(core__abc_21380_n5802) );
  INVX1 INVX1_1243 ( .A(core_v3_reg_26_), .Y(core__abc_21380_n5805) );
  INVX1 INVX1_1244 ( .A(core__abc_21380_n5807), .Y(core__abc_21380_n5809) );
  INVX1 INVX1_1245 ( .A(core__abc_21380_n5811), .Y(core__abc_21380_n5812) );
  INVX1 INVX1_1246 ( .A(core__abc_21380_n5804), .Y(core__abc_21380_n5814) );
  INVX1 INVX1_1247 ( .A(core__abc_21380_n5821), .Y(core__abc_21380_n5822) );
  INVX1 INVX1_1248 ( .A(core__abc_21380_n5823), .Y(core__abc_21380_n5825) );
  INVX1 INVX1_1249 ( .A(core_key_106_), .Y(core__abc_21380_n5829) );
  INVX1 INVX1_125 ( .A(_abc_19068_n2745), .Y(_abc_19068_n2746) );
  INVX1 INVX1_1250 ( .A(core__abc_21380_n5832), .Y(core__abc_21380_n5833) );
  INVX1 INVX1_1251 ( .A(core__abc_21380_n5813), .Y(core__abc_21380_n5842) );
  INVX1 INVX1_1252 ( .A(core__abc_21380_n5845), .Y(core__abc_21380_n5846) );
  INVX1 INVX1_1253 ( .A(core__abc_21380_n5848), .Y(core__abc_21380_n5849) );
  INVX1 INVX1_1254 ( .A(core__abc_21380_n5852), .Y(core__abc_21380_n5853) );
  INVX1 INVX1_1255 ( .A(core__abc_21380_n5843), .Y(core__abc_21380_n5855) );
  INVX1 INVX1_1256 ( .A(core__abc_21380_n5857), .Y(core__abc_21380_n5858) );
  INVX1 INVX1_1257 ( .A(core__abc_21380_n5865), .Y(core__abc_21380_n5866) );
  INVX1 INVX1_1258 ( .A(core__abc_21380_n5875), .Y(core__abc_21380_n5876) );
  INVX1 INVX1_1259 ( .A(core__abc_21380_n5816), .Y(core__abc_21380_n5877) );
  INVX1 INVX1_126 ( .A(_abc_19068_n2750), .Y(_abc_19068_n2751) );
  INVX1 INVX1_1260 ( .A(core__abc_21380_n5882), .Y(core__abc_21380_n5883) );
  INVX1 INVX1_1261 ( .A(core__abc_21380_n5888), .Y(core__abc_21380_n5889) );
  INVX1 INVX1_1262 ( .A(core__abc_21380_n5891), .Y(core__abc_21380_n5892) );
  INVX1 INVX1_1263 ( .A(core__abc_21380_n5895), .Y(core__abc_21380_n5896) );
  INVX1 INVX1_1264 ( .A(core__abc_21380_n5899), .Y(core__abc_21380_n5901) );
  INVX1 INVX1_1265 ( .A(core__abc_21380_n5903), .Y(core__abc_21380_n5905) );
  INVX1 INVX1_1266 ( .A(core__abc_21380_n5911), .Y(core__abc_21380_n5912) );
  INVX1 INVX1_1267 ( .A(core__abc_21380_n5921), .Y(core__abc_21380_n5922) );
  INVX1 INVX1_1268 ( .A(core__abc_21380_n5925), .Y(core__abc_21380_n5927) );
  INVX1 INVX1_1269 ( .A(core__abc_21380_n5929), .Y(core__abc_21380_n5930) );
  INVX1 INVX1_127 ( .A(_abc_19068_n2755), .Y(_abc_19068_n2756) );
  INVX1 INVX1_1270 ( .A(core__abc_21380_n5897), .Y(core__abc_21380_n5931) );
  INVX1 INVX1_1271 ( .A(core__abc_21380_n5902), .Y(core__abc_21380_n5932) );
  INVX1 INVX1_1272 ( .A(core__abc_21380_n5935), .Y(core__abc_21380_n5936) );
  INVX1 INVX1_1273 ( .A(core__abc_21380_n5937), .Y(core__abc_21380_n5938) );
  INVX1 INVX1_1274 ( .A(core_key_109_), .Y(core__abc_21380_n5943) );
  INVX1 INVX1_1275 ( .A(core__abc_21380_n5946), .Y(core__abc_21380_n5947) );
  INVX1 INVX1_1276 ( .A(core__abc_21380_n5926), .Y(core__abc_21380_n5958) );
  INVX1 INVX1_1277 ( .A(core__abc_21380_n5961), .Y(core__abc_21380_n5962) );
  INVX1 INVX1_1278 ( .A(core__abc_21380_n5965), .Y(core__abc_21380_n5966) );
  INVX1 INVX1_1279 ( .A(core__abc_21380_n5968), .Y(core__abc_21380_n5970) );
  INVX1 INVX1_128 ( .A(_abc_19068_n2760), .Y(_abc_19068_n2761) );
  INVX1 INVX1_1280 ( .A(core__abc_21380_n5972), .Y(core__abc_21380_n5974) );
  INVX1 INVX1_1281 ( .A(core__abc_21380_n4946), .Y(core__abc_21380_n5978) );
  INVX1 INVX1_1282 ( .A(core__abc_21380_n5976), .Y(core__abc_21380_n5979) );
  INVX1 INVX1_1283 ( .A(core_key_110_), .Y(core__abc_21380_n5983) );
  INVX1 INVX1_1284 ( .A(core__abc_21380_n5986), .Y(core__abc_21380_n5987) );
  INVX1 INVX1_1285 ( .A(core__abc_21380_n5997), .Y(core__abc_21380_n5998) );
  INVX1 INVX1_1286 ( .A(core__abc_21380_n6001), .Y(core__abc_21380_n6002) );
  INVX1 INVX1_1287 ( .A(core__abc_21380_n5996), .Y(core__abc_21380_n6007) );
  INVX1 INVX1_1288 ( .A(core__abc_21380_n6012), .Y(core__abc_21380_n6013) );
  INVX1 INVX1_1289 ( .A(core__abc_21380_n6020), .Y(core__abc_21380_n6021) );
  INVX1 INVX1_129 ( .A(_abc_19068_n2765), .Y(_abc_19068_n2766) );
  INVX1 INVX1_1290 ( .A(core__abc_21380_n5969), .Y(core__abc_21380_n6038) );
  INVX1 INVX1_1291 ( .A(core__abc_21380_n6040), .Y(core__abc_21380_n6041) );
  INVX1 INVX1_1292 ( .A(core__abc_21380_n6048), .Y(core__abc_21380_n6049) );
  INVX1 INVX1_1293 ( .A(core__abc_21380_n6052), .Y(core__abc_21380_n6053) );
  INVX1 INVX1_1294 ( .A(core__abc_21380_n6033), .Y(core__abc_21380_n6055) );
  INVX1 INVX1_1295 ( .A(core__abc_21380_n5516), .Y(core__abc_21380_n6057) );
  INVX1 INVX1_1296 ( .A(core__abc_21380_n5608), .Y(core__abc_21380_n6058) );
  INVX1 INVX1_1297 ( .A(core__abc_21380_n5607), .Y(core__abc_21380_n6062) );
  INVX1 INVX1_1298 ( .A(core__abc_21380_n5708), .Y(core__abc_21380_n6064) );
  INVX1 INVX1_1299 ( .A(core__abc_21380_n6032), .Y(core__abc_21380_n6067) );
  INVX1 INVX1_13 ( .A(_abc_19068_n2154), .Y(_abc_19068_n2155) );
  INVX1 INVX1_130 ( .A(_abc_19068_n2770), .Y(_abc_19068_n2771) );
  INVX1 INVX1_1300 ( .A(core__abc_21380_n6036), .Y(core__abc_21380_n6069) );
  INVX1 INVX1_1301 ( .A(core__abc_21380_n6042), .Y(core__abc_21380_n6070) );
  INVX1 INVX1_1302 ( .A(core__abc_21380_n6075), .Y(core__abc_21380_n6076) );
  INVX1 INVX1_1303 ( .A(core_key_112_), .Y(core__abc_21380_n6081) );
  INVX1 INVX1_1304 ( .A(core__abc_21380_n6084), .Y(core__abc_21380_n6085) );
  INVX1 INVX1_1305 ( .A(core__abc_21380_n6050), .Y(core__abc_21380_n6094) );
  INVX1 INVX1_1306 ( .A(core__abc_21380_n6054), .Y(core__abc_21380_n6095) );
  INVX1 INVX1_1307 ( .A(core__abc_21380_n6096), .Y(core__abc_21380_n6097) );
  INVX1 INVX1_1308 ( .A(core__abc_21380_n6098), .Y(core__abc_21380_n6099) );
  INVX1 INVX1_1309 ( .A(core__abc_21380_n6102), .Y(core__abc_21380_n6103) );
  INVX1 INVX1_131 ( .A(_abc_19068_n2775), .Y(_abc_19068_n2776) );
  INVX1 INVX1_1310 ( .A(core__abc_21380_n6104), .Y(core__abc_21380_n6105) );
  INVX1 INVX1_1311 ( .A(core__abc_21380_n6106), .Y(core__abc_21380_n6107) );
  INVX1 INVX1_1312 ( .A(core__abc_21380_n6108), .Y(core__abc_21380_n6110) );
  INVX1 INVX1_1313 ( .A(core__abc_21380_n6112), .Y(core__abc_21380_n6114) );
  INVX1 INVX1_1314 ( .A(core__abc_21380_n6120), .Y(core__abc_21380_n6121) );
  INVX1 INVX1_1315 ( .A(core__abc_21380_n6131), .Y(core__abc_21380_n6132) );
  INVX1 INVX1_1316 ( .A(core__abc_21380_n6135), .Y(core__abc_21380_n6136) );
  INVX1 INVX1_1317 ( .A(core__abc_21380_n6139), .Y(core__abc_21380_n6140) );
  INVX1 INVX1_1318 ( .A(core__abc_21380_n6142), .Y(core__abc_21380_n6144) );
  INVX1 INVX1_1319 ( .A(core__abc_21380_n6146), .Y(core__abc_21380_n6148) );
  INVX1 INVX1_132 ( .A(_abc_19068_n2780), .Y(_abc_19068_n2781) );
  INVX1 INVX1_1320 ( .A(core__abc_21380_n6150), .Y(core__abc_21380_n6152) );
  INVX1 INVX1_1321 ( .A(core_key_114_), .Y(core__abc_21380_n6156) );
  INVX1 INVX1_1322 ( .A(core__abc_21380_n6159), .Y(core__abc_21380_n6160) );
  INVX1 INVX1_1323 ( .A(core__abc_21380_n6171), .Y(core__abc_21380_n6172) );
  INVX1 INVX1_1324 ( .A(core__abc_21380_n6174), .Y(core__abc_21380_n6175) );
  INVX1 INVX1_1325 ( .A(core__abc_21380_n6169), .Y(core__abc_21380_n6180) );
  INVX1 INVX1_1326 ( .A(core__abc_21380_n6185), .Y(core__abc_21380_n6186) );
  INVX1 INVX1_1327 ( .A(core__abc_21380_n6193), .Y(core__abc_21380_n6194) );
  INVX1 INVX1_1328 ( .A(core__abc_21380_n6210), .Y(core__abc_21380_n6211) );
  INVX1 INVX1_1329 ( .A(core__abc_21380_n6213), .Y(core__abc_21380_n6214) );
  INVX1 INVX1_133 ( .A(_abc_19068_n2785), .Y(_abc_19068_n2786) );
  INVX1 INVX1_1330 ( .A(core__abc_21380_n6217), .Y(core__abc_21380_n6218) );
  INVX1 INVX1_1331 ( .A(core__abc_21380_n6221), .Y(core__abc_21380_n6223) );
  INVX1 INVX1_1332 ( .A(core__abc_21380_n6225), .Y(core__abc_21380_n6227) );
  INVX1 INVX1_1333 ( .A(core__abc_21380_n6233), .Y(core__abc_21380_n6234) );
  INVX1 INVX1_1334 ( .A(core__abc_21380_n6244), .Y(core__abc_21380_n6245) );
  INVX1 INVX1_1335 ( .A(core__abc_21380_n6248), .Y(core__abc_21380_n6249) );
  INVX1 INVX1_1336 ( .A(core__abc_21380_n6252), .Y(core__abc_21380_n6253) );
  INVX1 INVX1_1337 ( .A(core__abc_21380_n6243), .Y(core__abc_21380_n6255) );
  INVX1 INVX1_1338 ( .A(core__abc_21380_n6257), .Y(core__abc_21380_n6259) );
  INVX1 INVX1_1339 ( .A(core_key_117_), .Y(core__abc_21380_n6263) );
  INVX1 INVX1_134 ( .A(_abc_19068_n2790), .Y(_abc_19068_n2791) );
  INVX1 INVX1_1340 ( .A(core__abc_21380_n6266), .Y(core__abc_21380_n6267) );
  INVX1 INVX1_1341 ( .A(core__abc_21380_n6250), .Y(core__abc_21380_n6276) );
  INVX1 INVX1_1342 ( .A(core__abc_21380_n6219), .Y(core__abc_21380_n6277) );
  INVX1 INVX1_1343 ( .A(core__abc_21380_n6279), .Y(core__abc_21380_n6280) );
  INVX1 INVX1_1344 ( .A(core__abc_21380_n6281), .Y(core__abc_21380_n6282) );
  INVX1 INVX1_1345 ( .A(core__abc_21380_n6284), .Y(core__abc_21380_n6285) );
  INVX1 INVX1_1346 ( .A(core__abc_21380_n6288), .Y(core__abc_21380_n6289) );
  INVX1 INVX1_1347 ( .A(core__abc_21380_n6291), .Y(core__abc_21380_n6293) );
  INVX1 INVX1_1348 ( .A(core__abc_21380_n6295), .Y(core__abc_21380_n6297) );
  INVX1 INVX1_1349 ( .A(core__abc_21380_n6299), .Y(core__abc_21380_n6301) );
  INVX1 INVX1_135 ( .A(_abc_19068_n2795), .Y(_abc_19068_n2796) );
  INVX1 INVX1_1350 ( .A(core_key_118_), .Y(core__abc_21380_n6305) );
  INVX1 INVX1_1351 ( .A(core__abc_21380_n6308), .Y(core__abc_21380_n6309) );
  INVX1 INVX1_1352 ( .A(core__abc_21380_n6321), .Y(core__abc_21380_n6322) );
  INVX1 INVX1_1353 ( .A(core__abc_21380_n6323), .Y(core__abc_21380_n6325) );
  INVX1 INVX1_1354 ( .A(core__abc_21380_n6318), .Y(core__abc_21380_n6329) );
  INVX1 INVX1_1355 ( .A(core__abc_21380_n6334), .Y(core__abc_21380_n6335) );
  INVX1 INVX1_1356 ( .A(core__abc_21380_n6342), .Y(core__abc_21380_n6343) );
  INVX1 INVX1_1357 ( .A(core__abc_21380_n6208), .Y(core__abc_21380_n6352) );
  INVX1 INVX1_1358 ( .A(core__abc_21380_n6206), .Y(core__abc_21380_n6359) );
  INVX1 INVX1_1359 ( .A(core__abc_21380_n6292), .Y(core__abc_21380_n6364) );
  INVX1 INVX1_136 ( .A(_abc_19068_n2800), .Y(_abc_19068_n2801) );
  INVX1 INVX1_1360 ( .A(core__abc_21380_n6366), .Y(core__abc_21380_n6367) );
  INVX1 INVX1_1361 ( .A(core__abc_21380_n6368), .Y(core__abc_21380_n6369) );
  INVX1 INVX1_1362 ( .A(core__abc_21380_n3248), .Y(core__abc_21380_n6375) );
  INVX1 INVX1_1363 ( .A(core__abc_21380_n3230_1), .Y(core__abc_21380_n6376) );
  INVX1 INVX1_1364 ( .A(core__abc_21380_n6380), .Y(core__abc_21380_n6381) );
  INVX1 INVX1_1365 ( .A(core__abc_21380_n6384), .Y(core__abc_21380_n6392) );
  INVX1 INVX1_1366 ( .A(core__abc_21380_n6394), .Y(core__abc_21380_n6395) );
  INVX1 INVX1_1367 ( .A(core__abc_21380_n6402), .Y(core__abc_21380_n6403) );
  INVX1 INVX1_1368 ( .A(core__abc_21380_n6382), .Y(core__abc_21380_n6412) );
  INVX1 INVX1_1369 ( .A(core__abc_21380_n6393), .Y(core__abc_21380_n6413) );
  INVX1 INVX1_137 ( .A(_abc_19068_n2805), .Y(_abc_19068_n2806) );
  INVX1 INVX1_1370 ( .A(core__abc_21380_n6414), .Y(core__abc_21380_n6415) );
  INVX1 INVX1_1371 ( .A(core__abc_21380_n6416), .Y(core__abc_21380_n6417) );
  INVX1 INVX1_1372 ( .A(core__abc_21380_n6420), .Y(core__abc_21380_n6421) );
  INVX1 INVX1_1373 ( .A(core__abc_21380_n6422), .Y(core__abc_21380_n6423) );
  INVX1 INVX1_1374 ( .A(core__abc_21380_n6424), .Y(core__abc_21380_n6425) );
  INVX1 INVX1_1375 ( .A(core__abc_21380_n6426), .Y(core__abc_21380_n6428) );
  INVX1 INVX1_1376 ( .A(core__abc_21380_n6430), .Y(core__abc_21380_n6432) );
  INVX1 INVX1_1377 ( .A(core__abc_21380_n6438), .Y(core__abc_21380_n6439) );
  INVX1 INVX1_1378 ( .A(core__abc_21380_n6449), .Y(core__abc_21380_n6450) );
  INVX1 INVX1_1379 ( .A(core__abc_21380_n6453), .Y(core__abc_21380_n6454) );
  INVX1 INVX1_138 ( .A(_abc_19068_n2811), .Y(_abc_19068_n2812) );
  INVX1 INVX1_1380 ( .A(core__abc_21380_n3219), .Y(core__abc_21380_n6455) );
  INVX1 INVX1_1381 ( .A(core__abc_21380_n6457), .Y(core__abc_21380_n6458) );
  INVX1 INVX1_1382 ( .A(core__abc_21380_n6461), .Y(core__abc_21380_n6462) );
  INVX1 INVX1_1383 ( .A(core__abc_21380_n6465), .Y(core__abc_21380_n6467) );
  INVX1 INVX1_1384 ( .A(core__abc_21380_n6469), .Y(core__abc_21380_n6470) );
  INVX1 INVX1_1385 ( .A(core_key_122_), .Y(core__abc_21380_n6475) );
  INVX1 INVX1_1386 ( .A(core__abc_21380_n6478), .Y(core__abc_21380_n6479) );
  INVX1 INVX1_1387 ( .A(core__abc_21380_n6489), .Y(core__abc_21380_n6490) );
  INVX1 INVX1_1388 ( .A(core__abc_21380_n6493), .Y(core__abc_21380_n6494) );
  INVX1 INVX1_1389 ( .A(core__abc_21380_n6495), .Y(core__abc_21380_n6496) );
  INVX1 INVX1_139 ( .A(_abc_19068_n2816), .Y(_abc_19068_n2817) );
  INVX1 INVX1_1390 ( .A(core__abc_21380_n6488), .Y(core__abc_21380_n6500) );
  INVX1 INVX1_1391 ( .A(core__abc_21380_n6504), .Y(core__abc_21380_n6505) );
  INVX1 INVX1_1392 ( .A(core__abc_21380_n6512), .Y(core__abc_21380_n6513) );
  INVX1 INVX1_1393 ( .A(core__abc_21380_n6463), .Y(core__abc_21380_n6526) );
  INVX1 INVX1_1394 ( .A(core__abc_21380_n6528), .Y(core__abc_21380_n6529) );
  INVX1 INVX1_1395 ( .A(core__abc_21380_n6533), .Y(core__abc_21380_n6534) );
  INVX1 INVX1_1396 ( .A(core__abc_21380_n6537), .Y(core__abc_21380_n6539) );
  INVX1 INVX1_1397 ( .A(core__abc_21380_n6541), .Y(core__abc_21380_n6542) );
  INVX1 INVX1_1398 ( .A(core__abc_21380_n6451), .Y(core__abc_21380_n6544) );
  INVX1 INVX1_1399 ( .A(core__abc_21380_n6552), .Y(core__abc_21380_n6553) );
  INVX1 INVX1_14 ( .A(_abc_19068_n2160), .Y(_abc_19068_n2161) );
  INVX1 INVX1_140 ( .A(_abc_19068_n2821), .Y(_abc_19068_n2822) );
  INVX1 INVX1_1400 ( .A(core_key_124_), .Y(core__abc_21380_n6558) );
  INVX1 INVX1_1401 ( .A(core__abc_21380_n6561), .Y(core__abc_21380_n6562) );
  INVX1 INVX1_1402 ( .A(core__abc_21380_n6572), .Y(core__abc_21380_n6573) );
  INVX1 INVX1_1403 ( .A(core__abc_21380_n6576), .Y(core__abc_21380_n6577) );
  INVX1 INVX1_1404 ( .A(core__abc_21380_n6579), .Y(core__abc_21380_n6580) );
  INVX1 INVX1_1405 ( .A(core__abc_21380_n6571), .Y(core__abc_21380_n6583) );
  INVX1 INVX1_1406 ( .A(core__abc_21380_n6578), .Y(core__abc_21380_n6584) );
  INVX1 INVX1_1407 ( .A(core__abc_21380_n6587), .Y(core__abc_21380_n6588) );
  INVX1 INVX1_1408 ( .A(core_key_125_), .Y(core__abc_21380_n6593) );
  INVX1 INVX1_1409 ( .A(core__abc_21380_n6596), .Y(core__abc_21380_n6597) );
  INVX1 INVX1_141 ( .A(_abc_19068_n2826), .Y(_abc_19068_n2827) );
  INVX1 INVX1_1410 ( .A(core__abc_21380_n6613), .Y(core__abc_21380_n6614) );
  INVX1 INVX1_1411 ( .A(core__abc_21380_n6616), .Y(core__abc_21380_n6618) );
  INVX1 INVX1_1412 ( .A(core__abc_21380_n6620), .Y(core__abc_21380_n6621) );
  INVX1 INVX1_1413 ( .A(core__abc_21380_n6608), .Y(core__abc_21380_n6625) );
  INVX1 INVX1_1414 ( .A(core__abc_21380_n6629), .Y(core__abc_21380_n6630) );
  INVX1 INVX1_1415 ( .A(core_key_126_), .Y(core__abc_21380_n6635) );
  INVX1 INVX1_1416 ( .A(core__abc_21380_n6638), .Y(core__abc_21380_n6639) );
  INVX1 INVX1_1417 ( .A(core__abc_21380_n6652), .Y(core__abc_21380_n6653) );
  INVX1 INVX1_1418 ( .A(core__abc_21380_n6655), .Y(core__abc_21380_n6656) );
  INVX1 INVX1_1419 ( .A(core__abc_21380_n6654), .Y(core__abc_21380_n6657) );
  INVX1 INVX1_142 ( .A(_abc_19068_n2831), .Y(_abc_19068_n2832) );
  INVX1 INVX1_1420 ( .A(core__abc_21380_n6658), .Y(core__abc_21380_n6659) );
  INVX1 INVX1_1421 ( .A(core__abc_21380_n6617), .Y(core__abc_21380_n6662) );
  INVX1 INVX1_1422 ( .A(core__abc_21380_n6666), .Y(core__abc_21380_n6667) );
  INVX1 INVX1_1423 ( .A(core__abc_21380_n6674), .Y(core__abc_21380_n6675) );
  INVX1 INVX1_1424 ( .A(core_v1_reg_18_), .Y(core__abc_21380_n6684) );
  INVX1 INVX1_1425 ( .A(core__abc_21380_n6686), .Y(core__abc_21380_n6687) );
  INVX1 INVX1_1426 ( .A(core__abc_21380_n6685), .Y(core__abc_21380_n6690) );
  INVX1 INVX1_1427 ( .A(core__abc_21380_n6696), .Y(core__abc_21380_n6697) );
  INVX1 INVX1_1428 ( .A(core__abc_21380_n6700), .Y(core__abc_21380_n6701) );
  INVX1 INVX1_1429 ( .A(core__abc_21380_n5155), .Y(core__abc_21380_n6703) );
  INVX1 INVX1_143 ( .A(_abc_19068_n2836), .Y(_abc_19068_n2837) );
  INVX1 INVX1_1430 ( .A(core__abc_21380_n6706), .Y(core__abc_21380_n6707) );
  INVX1 INVX1_1431 ( .A(core__abc_21380_n6708), .Y(core__abc_21380_n6709) );
  INVX1 INVX1_1432 ( .A(core__abc_21380_n6710), .Y(core__abc_21380_n6711) );
  INVX1 INVX1_1433 ( .A(core__abc_21380_n6715), .Y(core__abc_21380_n6716) );
  INVX1 INVX1_1434 ( .A(core__abc_21380_n6719), .Y(core__abc_21380_n6720) );
  INVX1 INVX1_1435 ( .A(core__abc_21380_n6723), .Y(core__abc_21380_n6724) );
  INVX1 INVX1_1436 ( .A(core__abc_21380_n6728), .Y(core__abc_21380_n6729) );
  INVX1 INVX1_1437 ( .A(core__abc_21380_n6733), .Y(core__abc_21380_n6734) );
  INVX1 INVX1_1438 ( .A(core__abc_21380_n6737), .Y(core__abc_21380_n6738) );
  INVX1 INVX1_1439 ( .A(core__abc_21380_n6743), .Y(core__abc_21380_n6744) );
  INVX1 INVX1_144 ( .A(_abc_19068_n2841), .Y(_abc_19068_n2842) );
  INVX1 INVX1_1440 ( .A(core__abc_21380_n6742), .Y(core__abc_21380_n6745) );
  INVX1 INVX1_1441 ( .A(core__abc_21380_n6746), .Y(core__abc_21380_n6747) );
  INVX1 INVX1_1442 ( .A(core_v1_reg_11_), .Y(core__abc_21380_n6748) );
  INVX1 INVX1_1443 ( .A(core__abc_21380_n6751), .Y(core__abc_21380_n6752) );
  INVX1 INVX1_1444 ( .A(core__abc_21380_n6753), .Y(core__abc_21380_n6754) );
  INVX1 INVX1_1445 ( .A(core__abc_21380_n6755), .Y(core__abc_21380_n6756) );
  INVX1 INVX1_1446 ( .A(core__abc_21380_n6735), .Y(core__abc_21380_n6759) );
  INVX1 INVX1_1447 ( .A(core__abc_21380_n6761), .Y(core__abc_21380_n6762) );
  INVX1 INVX1_1448 ( .A(core__abc_21380_n6717), .Y(core__abc_21380_n6765) );
  INVX1 INVX1_1449 ( .A(core__abc_21380_n6766), .Y(core__abc_21380_n6767) );
  INVX1 INVX1_145 ( .A(_abc_19068_n2846), .Y(_abc_19068_n2847) );
  INVX1 INVX1_1450 ( .A(core__abc_21380_n6698), .Y(core__abc_21380_n6771) );
  INVX1 INVX1_1451 ( .A(core__abc_21380_n6773), .Y(core__abc_21380_n6774) );
  INVX1 INVX1_1452 ( .A(core__abc_21380_n6779), .Y(core__abc_21380_n6780) );
  INVX1 INVX1_1453 ( .A(core_v1_reg_10_), .Y(core__abc_21380_n6784) );
  INVX1 INVX1_1454 ( .A(core__abc_21380_n6786), .Y(core__abc_21380_n6787) );
  INVX1 INVX1_1455 ( .A(core__abc_21380_n4814_1), .Y(core__abc_21380_n6790) );
  INVX1 INVX1_1456 ( .A(core__abc_21380_n6797), .Y(core__abc_21380_n6798) );
  INVX1 INVX1_1457 ( .A(core__abc_21380_n6801), .Y(core__abc_21380_n6802) );
  INVX1 INVX1_1458 ( .A(core_v1_reg_8_), .Y(core__abc_21380_n6804) );
  INVX1 INVX1_1459 ( .A(core__abc_21380_n6807), .Y(core__abc_21380_n6808) );
  INVX1 INVX1_146 ( .A(_abc_19068_n2851), .Y(_abc_19068_n2852) );
  INVX1 INVX1_1460 ( .A(core__abc_21380_n6809), .Y(core__abc_21380_n6810) );
  INVX1 INVX1_1461 ( .A(core__abc_21380_n6811), .Y(core__abc_21380_n6812) );
  INVX1 INVX1_1462 ( .A(core__abc_21380_n6816), .Y(core__abc_21380_n6817) );
  INVX1 INVX1_1463 ( .A(core__abc_21380_n6820), .Y(core__abc_21380_n6821) );
  INVX1 INVX1_1464 ( .A(core__abc_21380_n6827), .Y(core__abc_21380_n6828) );
  INVX1 INVX1_1465 ( .A(core__abc_21380_n6833), .Y(core__abc_21380_n6834) );
  INVX1 INVX1_1466 ( .A(core__abc_21380_n6837), .Y(core__abc_21380_n6838) );
  INVX1 INVX1_1467 ( .A(core_v1_reg_4_), .Y(core__abc_21380_n6840) );
  INVX1 INVX1_1468 ( .A(core__abc_21380_n6843), .Y(core__abc_21380_n6844) );
  INVX1 INVX1_1469 ( .A(core__abc_21380_n6848), .Y(core__abc_21380_n6849) );
  INVX1 INVX1_147 ( .A(_abc_19068_n2856), .Y(_abc_19068_n2857) );
  INVX1 INVX1_1470 ( .A(core__abc_21380_n6851), .Y(core__abc_21380_n6852) );
  INVX1 INVX1_1471 ( .A(core__abc_21380_n6829), .Y(core__abc_21380_n6856) );
  INVX1 INVX1_1472 ( .A(core__abc_21380_n6835), .Y(core__abc_21380_n6857) );
  INVX1 INVX1_1473 ( .A(core__abc_21380_n6859), .Y(core__abc_21380_n6860) );
  INVX1 INVX1_1474 ( .A(core__abc_21380_n6818), .Y(core__abc_21380_n6863) );
  INVX1 INVX1_1475 ( .A(core__abc_21380_n6864), .Y(core__abc_21380_n6865) );
  INVX1 INVX1_1476 ( .A(core__abc_21380_n6799), .Y(core__abc_21380_n6869) );
  INVX1 INVX1_1477 ( .A(core__abc_21380_n6871), .Y(core__abc_21380_n6872) );
  INVX1 INVX1_1478 ( .A(core__abc_21380_n6878), .Y(core__abc_21380_n6879) );
  INVX1 INVX1_1479 ( .A(core__abc_21380_n6884), .Y(core__abc_21380_n6885) );
  INVX1 INVX1_148 ( .A(_abc_19068_n2861), .Y(_abc_19068_n2862) );
  INVX1 INVX1_1480 ( .A(core__abc_21380_n6888), .Y(core__abc_21380_n6889) );
  INVX1 INVX1_1481 ( .A(core_v1_reg_0_), .Y(core__abc_21380_n6891) );
  INVX1 INVX1_1482 ( .A(core__abc_21380_n6894), .Y(core__abc_21380_n6896) );
  INVX1 INVX1_1483 ( .A(core__abc_21380_n6897), .Y(core__abc_21380_n6898) );
  INVX1 INVX1_1484 ( .A(core__abc_21380_n6901), .Y(core__abc_21380_n6902) );
  INVX1 INVX1_1485 ( .A(core__abc_21380_n6903), .Y(core__abc_21380_n6904) );
  INVX1 INVX1_1486 ( .A(core__abc_21380_n6906), .Y(core__abc_21380_n6907) );
  INVX1 INVX1_1487 ( .A(core__abc_21380_n6895), .Y(core__abc_21380_n6912) );
  INVX1 INVX1_1488 ( .A(core__abc_21380_n6915), .Y(core__abc_21380_n6916) );
  INVX1 INVX1_1489 ( .A(core__abc_21380_n6920), .Y(core__abc_21380_n6921) );
  INVX1 INVX1_149 ( .A(_abc_19068_n2866), .Y(_abc_19068_n2867) );
  INVX1 INVX1_1490 ( .A(core__abc_21380_n6926), .Y(core__abc_21380_n6927) );
  INVX1 INVX1_1491 ( .A(core__abc_21380_n6928), .Y(core__abc_21380_n6929) );
  INVX1 INVX1_1492 ( .A(core__abc_21380_n6932), .Y(core__abc_21380_n6933) );
  INVX1 INVX1_1493 ( .A(core__abc_21380_n6936), .Y(core__abc_21380_n6937) );
  INVX1 INVX1_1494 ( .A(core__abc_21380_n6938), .Y(core__abc_21380_n6939) );
  INVX1 INVX1_1495 ( .A(core__abc_21380_n6943), .Y(core__abc_21380_n6944) );
  INVX1 INVX1_1496 ( .A(core__abc_21380_n6945), .Y(core__abc_21380_n6946) );
  INVX1 INVX1_1497 ( .A(core__abc_21380_n6948), .Y(core__abc_21380_n6949) );
  INVX1 INVX1_1498 ( .A(core__abc_21380_n6923), .Y(core__abc_21380_n6950) );
  INVX1 INVX1_1499 ( .A(core__abc_21380_n6953), .Y(core__abc_21380_n6954) );
  INVX1 INVX1_15 ( .A(_abc_19068_n2166), .Y(_abc_19068_n2167) );
  INVX1 INVX1_150 ( .A(_abc_19068_n2871), .Y(_abc_19068_n2872) );
  INVX1 INVX1_1500 ( .A(core__abc_21380_n6960), .Y(core__abc_21380_n6962) );
  INVX1 INVX1_1501 ( .A(core__abc_21380_n6963), .Y(core__abc_21380_n6964) );
  INVX1 INVX1_1502 ( .A(core__abc_21380_n6967), .Y(core__abc_21380_n6968) );
  INVX1 INVX1_1503 ( .A(core__abc_21380_n6961), .Y(core__abc_21380_n6972) );
  INVX1 INVX1_1504 ( .A(core__abc_21380_n6975), .Y(core__abc_21380_n6976) );
  INVX1 INVX1_1505 ( .A(core__abc_21380_n6980), .Y(core__abc_21380_n6981) );
  INVX1 INVX1_1506 ( .A(core__abc_21380_n6984), .Y(core__abc_21380_n6985) );
  INVX1 INVX1_1507 ( .A(core__abc_21380_n6988), .Y(core__abc_21380_n6989) );
  INVX1 INVX1_1508 ( .A(core__abc_21380_n6994), .Y(core__abc_21380_n6995) );
  INVX1 INVX1_1509 ( .A(core__abc_21380_n6996), .Y(core__abc_21380_n6997) );
  INVX1 INVX1_151 ( .A(_abc_19068_n2876), .Y(_abc_19068_n2877) );
  INVX1 INVX1_1510 ( .A(core__abc_21380_n7001), .Y(core__abc_21380_n7002) );
  INVX1 INVX1_1511 ( .A(core_v1_reg_52_), .Y(core__abc_21380_n7004) );
  INVX1 INVX1_1512 ( .A(core__abc_21380_n7007), .Y(core__abc_21380_n7008) );
  INVX1 INVX1_1513 ( .A(core__abc_21380_n7009), .Y(core__abc_21380_n7014) );
  INVX1 INVX1_1514 ( .A(core__abc_21380_n7015), .Y(core__abc_21380_n7016) );
  INVX1 INVX1_1515 ( .A(core__abc_21380_n7003), .Y(core__abc_21380_n7020) );
  INVX1 INVX1_1516 ( .A(core__abc_21380_n7021), .Y(core__abc_21380_n7022) );
  INVX1 INVX1_1517 ( .A(core__abc_21380_n7029), .Y(core__abc_21380_n7030) );
  INVX1 INVX1_1518 ( .A(core__abc_21380_n6940), .Y(core__abc_21380_n7037) );
  INVX1 INVX1_1519 ( .A(core__abc_21380_n7040), .Y(core__abc_21380_n7041) );
  INVX1 INVX1_152 ( .A(_abc_19068_n2881), .Y(_abc_19068_n2882) );
  INVX1 INVX1_1520 ( .A(core__abc_21380_n6845), .Y(core__abc_21380_n7048) );
  INVX1 INVX1_1521 ( .A(core__abc_21380_n7051), .Y(core__abc_21380_n7052) );
  INVX1 INVX1_1522 ( .A(core__abc_21380_n7059), .Y(core__abc_21380_n7060) );
  INVX1 INVX1_1523 ( .A(core_v1_reg_19_), .Y(core__abc_21380_n7061) );
  INVX1 INVX1_1524 ( .A(core__abc_21380_n7064), .Y(core__abc_21380_n7065) );
  INVX1 INVX1_1525 ( .A(core__abc_21380_n7068), .Y(core__abc_21380_n7070) );
  INVX1 INVX1_1526 ( .A(core__abc_21380_n7072), .Y(core__abc_21380_n7073) );
  INVX1 INVX1_1527 ( .A(core_key_0_), .Y(core__abc_21380_n7077) );
  INVX1 INVX1_1528 ( .A(core__abc_21380_n7093), .Y(core__abc_21380_n7095) );
  INVX1 INVX1_1529 ( .A(core__abc_21380_n7066), .Y(core__abc_21380_n7098) );
  INVX1 INVX1_153 ( .A(_abc_19068_n2886), .Y(_abc_19068_n2887) );
  INVX1 INVX1_1530 ( .A(core__abc_21380_n7071), .Y(core__abc_21380_n7099) );
  INVX1 INVX1_1531 ( .A(core__abc_21380_n7102), .Y(core__abc_21380_n7103) );
  INVX1 INVX1_1532 ( .A(core__abc_21380_n7104), .Y(core__abc_21380_n7105) );
  INVX1 INVX1_1533 ( .A(core__abc_21380_n7097), .Y(core__abc_21380_n7115) );
  INVX1 INVX1_1534 ( .A(core__abc_21380_n7120), .Y(core__abc_21380_n7121) );
  INVX1 INVX1_1535 ( .A(core__abc_21380_n7124), .Y(core__abc_21380_n7125) );
  INVX1 INVX1_1536 ( .A(core__abc_21380_n7128), .Y(core__abc_21380_n7130) );
  INVX1 INVX1_1537 ( .A(core__abc_21380_n7132), .Y(core__abc_21380_n7133) );
  INVX1 INVX1_1538 ( .A(core__abc_21380_n7143), .Y(core__abc_21380_n7144) );
  INVX1 INVX1_1539 ( .A(core__abc_21380_n7147), .Y(core__abc_21380_n7148) );
  INVX1 INVX1_154 ( .A(_abc_19068_n2891), .Y(_abc_19068_n2892) );
  INVX1 INVX1_1540 ( .A(core__abc_21380_n7149), .Y(core__abc_21380_n7150) );
  INVX1 INVX1_1541 ( .A(core__abc_21380_n7151), .Y(core__abc_21380_n7152) );
  INVX1 INVX1_1542 ( .A(core__abc_21380_n7153), .Y(core__abc_21380_n7154) );
  INVX1 INVX1_1543 ( .A(core__abc_21380_n7157), .Y(core__abc_21380_n7158) );
  INVX1 INVX1_1544 ( .A(core__abc_21380_n7178), .Y(core__abc_21380_n7179) );
  INVX1 INVX1_1545 ( .A(core__abc_21380_n7182), .Y(core__abc_21380_n7183) );
  INVX1 INVX1_1546 ( .A(core__abc_21380_n7184), .Y(core__abc_21380_n7185) );
  INVX1 INVX1_1547 ( .A(core__abc_21380_n7180), .Y(core__abc_21380_n7200) );
  INVX1 INVX1_1548 ( .A(core__abc_21380_n7201), .Y(core__abc_21380_n7202) );
  INVX1 INVX1_1549 ( .A(core__abc_21380_n5572), .Y(core__abc_21380_n7203) );
  INVX1 INVX1_155 ( .A(_abc_19068_n2896), .Y(_abc_19068_n2897) );
  INVX1 INVX1_1550 ( .A(core__abc_21380_n7206), .Y(core__abc_21380_n7207) );
  INVX1 INVX1_1551 ( .A(core__abc_21380_n7208), .Y(core__abc_21380_n7209) );
  INVX1 INVX1_1552 ( .A(core__abc_21380_n7210), .Y(core__abc_21380_n7211) );
  INVX1 INVX1_1553 ( .A(core__abc_21380_n7212), .Y(core__abc_21380_n7213) );
  INVX1 INVX1_1554 ( .A(core_key_5_), .Y(core__abc_21380_n7218) );
  INVX1 INVX1_1555 ( .A(core__abc_21380_n3686), .Y(core__abc_21380_n7227) );
  INVX1 INVX1_1556 ( .A(core__abc_21380_n7230), .Y(core__abc_21380_n7231) );
  INVX1 INVX1_1557 ( .A(core__abc_21380_n7239), .Y(core__abc_21380_n7240) );
  INVX1 INVX1_1558 ( .A(core__abc_21380_n7241), .Y(core__abc_21380_n7242) );
  INVX1 INVX1_1559 ( .A(core_key_6_), .Y(core__abc_21380_n7244) );
  INVX1 INVX1_156 ( .A(_abc_19068_n2901), .Y(_abc_19068_n2902) );
  INVX1 INVX1_1560 ( .A(core__abc_21380_n7232), .Y(core__abc_21380_n7253) );
  INVX1 INVX1_1561 ( .A(core__abc_21380_n5668), .Y(core__abc_21380_n7255) );
  INVX1 INVX1_1562 ( .A(core_v1_reg_26_), .Y(core__abc_21380_n7256) );
  INVX1 INVX1_1563 ( .A(core__abc_21380_n7259), .Y(core__abc_21380_n7260) );
  INVX1 INVX1_1564 ( .A(core__abc_21380_n7264), .Y(core__abc_21380_n7265) );
  INVX1 INVX1_1565 ( .A(core__abc_21380_n7278), .Y(core__abc_21380_n7279) );
  INVX1 INVX1_1566 ( .A(core__abc_21380_n7283), .Y(core__abc_21380_n7284) );
  INVX1 INVX1_1567 ( .A(core__abc_21380_n7262), .Y(core__abc_21380_n7287) );
  INVX1 INVX1_1568 ( .A(core__abc_21380_n7289), .Y(core__abc_21380_n7290) );
  INVX1 INVX1_1569 ( .A(core__abc_21380_n7292), .Y(core__abc_21380_n7293) );
  INVX1 INVX1_157 ( .A(_abc_19068_n2906), .Y(_abc_19068_n2907) );
  INVX1 INVX1_1570 ( .A(core__abc_21380_n7297), .Y(core__abc_21380_n7298) );
  INVX1 INVX1_1571 ( .A(core__abc_21380_n7301), .Y(core__abc_21380_n7302) );
  INVX1 INVX1_1572 ( .A(core__abc_21380_n7294), .Y(core__abc_21380_n7304) );
  INVX1 INVX1_1573 ( .A(core__abc_21380_n7306), .Y(core__abc_21380_n7307) );
  INVX1 INVX1_1574 ( .A(core__abc_21380_n7299), .Y(core__abc_21380_n7317) );
  INVX1 INVX1_1575 ( .A(core__abc_21380_n7303), .Y(core__abc_21380_n7318) );
  INVX1 INVX1_1576 ( .A(core__abc_21380_n7320), .Y(core__abc_21380_n7321) );
  INVX1 INVX1_1577 ( .A(core__abc_21380_n7324), .Y(core__abc_21380_n7325) );
  INVX1 INVX1_1578 ( .A(core__abc_21380_n7323), .Y(core__abc_21380_n7326) );
  INVX1 INVX1_1579 ( .A(core__abc_21380_n7327), .Y(core__abc_21380_n7328) );
  INVX1 INVX1_158 ( .A(_abc_19068_n2911), .Y(_abc_19068_n2912) );
  INVX1 INVX1_1580 ( .A(core__abc_21380_n7329), .Y(core__abc_21380_n7330) );
  INVX1 INVX1_1581 ( .A(core__abc_21380_n7331), .Y(core__abc_21380_n7332) );
  INVX1 INVX1_1582 ( .A(core_key_9_), .Y(core__abc_21380_n7336) );
  INVX1 INVX1_1583 ( .A(core__abc_21380_n7346), .Y(core__abc_21380_n7347) );
  INVX1 INVX1_1584 ( .A(core__abc_21380_n7350), .Y(core__abc_21380_n7351) );
  INVX1 INVX1_1585 ( .A(core__abc_21380_n7354), .Y(core__abc_21380_n7355) );
  INVX1 INVX1_1586 ( .A(core__abc_21380_n7358), .Y(core__abc_21380_n7360) );
  INVX1 INVX1_1587 ( .A(core__abc_21380_n7362), .Y(core__abc_21380_n7363) );
  INVX1 INVX1_1588 ( .A(core__abc_21380_n7373), .Y(core__abc_21380_n7374) );
  INVX1 INVX1_1589 ( .A(core__abc_21380_n7377), .Y(core__abc_21380_n7379) );
  INVX1 INVX1_159 ( .A(_abc_19068_n2916), .Y(_abc_19068_n2917) );
  INVX1 INVX1_1590 ( .A(core__abc_21380_n7381), .Y(core__abc_21380_n7383) );
  INVX1 INVX1_1591 ( .A(core__abc_21380_n7385), .Y(core__abc_21380_n7386) );
  INVX1 INVX1_1592 ( .A(core__abc_21380_n7403), .Y(core__abc_21380_n7404) );
  INVX1 INVX1_1593 ( .A(core__abc_21380_n7407), .Y(core__abc_21380_n7408) );
  INVX1 INVX1_1594 ( .A(core__abc_21380_n7411), .Y(core__abc_21380_n7413) );
  INVX1 INVX1_1595 ( .A(core__abc_21380_n7415), .Y(core__abc_21380_n7416) );
  INVX1 INVX1_1596 ( .A(core_key_12_), .Y(core__abc_21380_n7418) );
  INVX1 INVX1_1597 ( .A(core__abc_21380_n7431), .Y(core__abc_21380_n7432) );
  INVX1 INVX1_1598 ( .A(core__abc_21380_n7433), .Y(core__abc_21380_n7434) );
  INVX1 INVX1_1599 ( .A(core__abc_21380_n7409), .Y(core__abc_21380_n7435) );
  INVX1 INVX1_16 ( .A(_abc_19068_n2172), .Y(_abc_19068_n2173) );
  INVX1 INVX1_160 ( .A(_abc_19068_n2921), .Y(_abc_19068_n2922) );
  INVX1 INVX1_1600 ( .A(core__abc_21380_n7414), .Y(core__abc_21380_n7436) );
  INVX1 INVX1_1601 ( .A(core__abc_21380_n7439), .Y(core__abc_21380_n7440) );
  INVX1 INVX1_1602 ( .A(core__abc_21380_n7441), .Y(core__abc_21380_n7442) );
  INVX1 INVX1_1603 ( .A(core_key_13_), .Y(core__abc_21380_n7444) );
  INVX1 INVX1_1604 ( .A(core__abc_21380_n7430), .Y(core__abc_21380_n7455) );
  INVX1 INVX1_1605 ( .A(core__abc_21380_n7458), .Y(core__abc_21380_n7459) );
  INVX1 INVX1_1606 ( .A(core__abc_21380_n7462), .Y(core__abc_21380_n7463) );
  INVX1 INVX1_1607 ( .A(core__abc_21380_n7466), .Y(core__abc_21380_n7468) );
  INVX1 INVX1_1608 ( .A(core__abc_21380_n7470), .Y(core__abc_21380_n7471) );
  INVX1 INVX1_1609 ( .A(core_key_14_), .Y(core__abc_21380_n7473) );
  INVX1 INVX1_161 ( .A(_abc_19068_n2926), .Y(_abc_19068_n2927) );
  INVX1 INVX1_1610 ( .A(core__abc_21380_n7482), .Y(core__abc_21380_n7483) );
  INVX1 INVX1_1611 ( .A(core__abc_21380_n7486), .Y(core__abc_21380_n7487) );
  INVX1 INVX1_1612 ( .A(core__abc_21380_n7490), .Y(core__abc_21380_n7492) );
  INVX1 INVX1_1613 ( .A(core__abc_21380_n7494), .Y(core__abc_21380_n7495) );
  INVX1 INVX1_1614 ( .A(core__abc_21380_n7489), .Y(core__abc_21380_n7509) );
  INVX1 INVX1_1615 ( .A(core__abc_21380_n7519), .Y(core__abc_21380_n7521) );
  INVX1 INVX1_1616 ( .A(core__abc_21380_n7523), .Y(core__abc_21380_n7524) );
  INVX1 INVX1_1617 ( .A(core__abc_21380_n7513), .Y(core__abc_21380_n7526) );
  INVX1 INVX1_1618 ( .A(core__abc_21380_n7514), .Y(core__abc_21380_n7527) );
  INVX1 INVX1_1619 ( .A(core__abc_21380_n7531), .Y(core__abc_21380_n7532) );
  INVX1 INVX1_162 ( .A(_abc_19068_n2931), .Y(_abc_19068_n2932) );
  INVX1 INVX1_1620 ( .A(core__abc_21380_n7535), .Y(core__abc_21380_n7536) );
  INVX1 INVX1_1621 ( .A(core_key_16_), .Y(core__abc_21380_n7538) );
  INVX1 INVX1_1622 ( .A(core__abc_21380_n7522), .Y(core__abc_21380_n7547) );
  INVX1 INVX1_1623 ( .A(core__abc_21380_n7525), .Y(core__abc_21380_n7548) );
  INVX1 INVX1_1624 ( .A(core__abc_21380_n7549), .Y(core__abc_21380_n7550) );
  INVX1 INVX1_1625 ( .A(core__abc_21380_n7553), .Y(core__abc_21380_n7554) );
  INVX1 INVX1_1626 ( .A(core__abc_21380_n7555), .Y(core__abc_21380_n7556) );
  INVX1 INVX1_1627 ( .A(core__abc_21380_n7557), .Y(core__abc_21380_n7558) );
  INVX1 INVX1_1628 ( .A(core__abc_21380_n7559), .Y(core__abc_21380_n7561) );
  INVX1 INVX1_1629 ( .A(core__abc_21380_n7577), .Y(core__abc_21380_n7578) );
  INVX1 INVX1_163 ( .A(_abc_19068_n2936), .Y(_abc_19068_n2937) );
  INVX1 INVX1_1630 ( .A(core__abc_21380_n7581), .Y(core__abc_21380_n7583) );
  INVX1 INVX1_1631 ( .A(core__abc_21380_n7585), .Y(core__abc_21380_n7587) );
  INVX1 INVX1_1632 ( .A(core__abc_21380_n7589), .Y(core__abc_21380_n7590) );
  INVX1 INVX1_1633 ( .A(core_key_18_), .Y(core__abc_21380_n7592) );
  INVX1 INVX1_1634 ( .A(core__abc_21380_n7604), .Y(core__abc_21380_n7605) );
  INVX1 INVX1_1635 ( .A(core__abc_21380_n7606), .Y(core__abc_21380_n7607) );
  INVX1 INVX1_1636 ( .A(core__abc_21380_n7601), .Y(core__abc_21380_n7611) );
  INVX1 INVX1_1637 ( .A(core__abc_21380_n7609), .Y(core__abc_21380_n7612) );
  INVX1 INVX1_1638 ( .A(core__abc_21380_n7628), .Y(core__abc_21380_n7629) );
  INVX1 INVX1_1639 ( .A(core__abc_21380_n7630), .Y(core__abc_21380_n7631) );
  INVX1 INVX1_164 ( .A(_abc_19068_n2941), .Y(_abc_19068_n2942) );
  INVX1 INVX1_1640 ( .A(core__abc_21380_n7636), .Y(core__abc_21380_n7637) );
  INVX1 INVX1_1641 ( .A(core__abc_21380_n7642), .Y(core__abc_21380_n7643) );
  INVX1 INVX1_1642 ( .A(core__abc_21380_n7644), .Y(core__abc_21380_n7645) );
  INVX1 INVX1_1643 ( .A(core__abc_21380_n7657), .Y(core__abc_21380_n7658) );
  INVX1 INVX1_1644 ( .A(core__abc_21380_n7638), .Y(core__abc_21380_n7662) );
  INVX1 INVX1_1645 ( .A(core__abc_21380_n7664), .Y(core__abc_21380_n7665) );
  INVX1 INVX1_1646 ( .A(core_key_21_), .Y(core__abc_21380_n7669) );
  INVX1 INVX1_1647 ( .A(core__abc_21380_n7661), .Y(core__abc_21380_n7678) );
  INVX1 INVX1_1648 ( .A(core__abc_21380_n7682), .Y(core__abc_21380_n7683) );
  INVX1 INVX1_1649 ( .A(core__abc_21380_n7686), .Y(core__abc_21380_n7687) );
  INVX1 INVX1_165 ( .A(_abc_19068_n2946), .Y(_abc_19068_n2947) );
  INVX1 INVX1_1650 ( .A(core__abc_21380_n7690), .Y(core__abc_21380_n7692) );
  INVX1 INVX1_1651 ( .A(core__abc_21380_n7694), .Y(core__abc_21380_n7695) );
  INVX1 INVX1_1652 ( .A(core_key_22_), .Y(core__abc_21380_n7697) );
  INVX1 INVX1_1653 ( .A(core__abc_21380_n7709), .Y(core__abc_21380_n7710) );
  INVX1 INVX1_1654 ( .A(core__abc_21380_n7711), .Y(core__abc_21380_n7712) );
  INVX1 INVX1_1655 ( .A(core__abc_21380_n7713), .Y(core__abc_21380_n7714) );
  INVX1 INVX1_1656 ( .A(core__abc_21380_n7715), .Y(core__abc_21380_n7716) );
  INVX1 INVX1_1657 ( .A(core__abc_21380_n7706), .Y(core__abc_21380_n7718) );
  INVX1 INVX1_1658 ( .A(core__abc_21380_n7720), .Y(core__abc_21380_n7721) );
  INVX1 INVX1_1659 ( .A(core__abc_21380_n7732), .Y(core__abc_21380_n7733) );
  INVX1 INVX1_166 ( .A(_abc_19068_n2951), .Y(_abc_19068_n2952) );
  INVX1 INVX1_1660 ( .A(core__abc_21380_n7734), .Y(core__abc_21380_n7735) );
  INVX1 INVX1_1661 ( .A(core__abc_21380_n7736), .Y(core__abc_21380_n7737) );
  INVX1 INVX1_1662 ( .A(core__abc_21380_n7744), .Y(core__abc_21380_n7745) );
  INVX1 INVX1_1663 ( .A(core__abc_21380_n7749), .Y(core__abc_21380_n7751) );
  INVX1 INVX1_1664 ( .A(core__abc_21380_n7755), .Y(core__abc_21380_n7756) );
  INVX1 INVX1_1665 ( .A(core__abc_21380_n7757), .Y(core__abc_21380_n7758) );
  INVX1 INVX1_1666 ( .A(core__abc_21380_n7752), .Y(core__abc_21380_n7768) );
  INVX1 INVX1_1667 ( .A(core__abc_21380_n7770), .Y(core__abc_21380_n7771) );
  INVX1 INVX1_1668 ( .A(core__abc_21380_n7774), .Y(core__abc_21380_n7775) );
  INVX1 INVX1_1669 ( .A(core__abc_21380_n7773), .Y(core__abc_21380_n7776) );
  INVX1 INVX1_167 ( .A(_abc_19068_n2956), .Y(_abc_19068_n2957) );
  INVX1 INVX1_1670 ( .A(core__abc_21380_n7777), .Y(core__abc_21380_n7778) );
  INVX1 INVX1_1671 ( .A(core__abc_21380_n7769), .Y(core__abc_21380_n7781) );
  INVX1 INVX1_1672 ( .A(core__abc_21380_n7779), .Y(core__abc_21380_n7782) );
  INVX1 INVX1_1673 ( .A(core__abc_21380_n7784), .Y(core__abc_21380_n7785) );
  INVX1 INVX1_1674 ( .A(core_key_25_), .Y(core__abc_21380_n7787) );
  INVX1 INVX1_1675 ( .A(core__abc_21380_n7798), .Y(core__abc_21380_n7800) );
  INVX1 INVX1_1676 ( .A(core__abc_21380_n7809), .Y(core__abc_21380_n7810) );
  INVX1 INVX1_1677 ( .A(core__abc_21380_n7811), .Y(core__abc_21380_n7812) );
  INVX1 INVX1_1678 ( .A(core_key_26_), .Y(core__abc_21380_n7814) );
  INVX1 INVX1_1679 ( .A(core__abc_21380_n7801), .Y(core__abc_21380_n7823) );
  INVX1 INVX1_168 ( .A(_abc_19068_n2961), .Y(_abc_19068_n2962) );
  INVX1 INVX1_1680 ( .A(core__abc_21380_n7827), .Y(core__abc_21380_n7828) );
  INVX1 INVX1_1681 ( .A(core__abc_21380_n7829), .Y(core__abc_21380_n7830) );
  INVX1 INVX1_1682 ( .A(core__abc_21380_n4422_1), .Y(core__abc_21380_n7831) );
  INVX1 INVX1_1683 ( .A(core__abc_21380_n7832), .Y(core__abc_21380_n7833) );
  INVX1 INVX1_1684 ( .A(core__abc_21380_n7834), .Y(core__abc_21380_n7835) );
  INVX1 INVX1_1685 ( .A(core__abc_21380_n7824), .Y(core__abc_21380_n7837) );
  INVX1 INVX1_1686 ( .A(core__abc_21380_n7839), .Y(core__abc_21380_n7840) );
  INVX1 INVX1_1687 ( .A(core_key_27_), .Y(core__abc_21380_n7842) );
  INVX1 INVX1_1688 ( .A(core__abc_21380_n7854), .Y(core__abc_21380_n7855) );
  INVX1 INVX1_1689 ( .A(core__abc_21380_n7859), .Y(core__abc_21380_n7860) );
  INVX1 INVX1_169 ( .A(_abc_19068_n2966), .Y(_abc_19068_n2967) );
  INVX1 INVX1_1690 ( .A(core__abc_21380_n7861), .Y(core__abc_21380_n7862) );
  INVX1 INVX1_1691 ( .A(core__abc_21380_n7866), .Y(core__abc_21380_n7868) );
  INVX1 INVX1_1692 ( .A(core__abc_21380_n7870), .Y(core__abc_21380_n7871) );
  INVX1 INVX1_1693 ( .A(core__abc_21380_n7876), .Y(core__abc_21380_n7877) );
  INVX1 INVX1_1694 ( .A(core__abc_21380_n4550), .Y(core__abc_21380_n7888) );
  INVX1 INVX1_1695 ( .A(core__abc_21380_n7891), .Y(core__abc_21380_n7893) );
  INVX1 INVX1_1696 ( .A(core__abc_21380_n7887), .Y(core__abc_21380_n7897) );
  INVX1 INVX1_1697 ( .A(core__abc_21380_n7895), .Y(core__abc_21380_n7898) );
  INVX1 INVX1_1698 ( .A(core__abc_21380_n7900), .Y(core__abc_21380_n7901) );
  INVX1 INVX1_1699 ( .A(core_key_29_), .Y(core__abc_21380_n7903) );
  INVX1 INVX1_17 ( .A(_abc_19068_n2178), .Y(_abc_19068_n2179) );
  INVX1 INVX1_170 ( .A(_abc_19068_n2972), .Y(_abc_19068_n2973) );
  INVX1 INVX1_1700 ( .A(core__abc_21380_n7912), .Y(core__abc_21380_n7913) );
  INVX1 INVX1_1701 ( .A(core__abc_21380_n7916), .Y(core__abc_21380_n7917) );
  INVX1 INVX1_1702 ( .A(core__abc_21380_n7921), .Y(core__abc_21380_n7922) );
  INVX1 INVX1_1703 ( .A(core__abc_21380_n7925), .Y(core__abc_21380_n7929) );
  INVX1 INVX1_1704 ( .A(core__abc_21380_n7931), .Y(core__abc_21380_n7932) );
  INVX1 INVX1_1705 ( .A(core_key_30_), .Y(core__abc_21380_n7934) );
  INVX1 INVX1_1706 ( .A(core__abc_21380_n7923), .Y(core__abc_21380_n7943) );
  INVX1 INVX1_1707 ( .A(core__abc_21380_n7948), .Y(core__abc_21380_n7949) );
  INVX1 INVX1_1708 ( .A(core__abc_21380_n7952), .Y(core__abc_21380_n7953) );
  INVX1 INVX1_1709 ( .A(core__abc_21380_n7954), .Y(core__abc_21380_n7955) );
  INVX1 INVX1_171 ( .A(_abc_19068_n2977), .Y(_abc_19068_n2978) );
  INVX1 INVX1_1710 ( .A(core_key_32_), .Y(core__abc_21380_n7967) );
  INVX1 INVX1_1711 ( .A(core__abc_21380_n7012), .Y(core__abc_21380_n7969) );
  INVX1 INVX1_1712 ( .A(core__abc_21380_n7971), .Y(core__abc_21380_n7972) );
  INVX1 INVX1_1713 ( .A(core__abc_21380_n7018), .Y(core__abc_21380_n7980) );
  INVX1 INVX1_1714 ( .A(core__abc_21380_n7024), .Y(core__abc_21380_n7991) );
  INVX1 INVX1_1715 ( .A(core_key_34_), .Y(core__abc_21380_n7995) );
  INVX1 INVX1_1716 ( .A(core__abc_21380_n7026), .Y(core__abc_21380_n8001) );
  INVX1 INVX1_1717 ( .A(core__abc_21380_n7031), .Y(core__abc_21380_n8013) );
  INVX1 INVX1_1718 ( .A(core__abc_21380_n7033), .Y(core__abc_21380_n8025) );
  INVX1 INVX1_1719 ( .A(core_key_37_), .Y(core__abc_21380_n8029) );
  INVX1 INVX1_172 ( .A(_abc_19068_n2982), .Y(_abc_19068_n2983) );
  INVX1 INVX1_1720 ( .A(core__abc_21380_n8038), .Y(core__abc_21380_n8039) );
  INVX1 INVX1_1721 ( .A(core_key_38_), .Y(core__abc_21380_n8043) );
  INVX1 INVX1_1722 ( .A(core__abc_21380_n6973), .Y(core__abc_21380_n8054) );
  INVX1 INVX1_1723 ( .A(core__abc_21380_n8052), .Y(core__abc_21380_n8055) );
  INVX1 INVX1_1724 ( .A(core__abc_21380_n7036), .Y(core__abc_21380_n8067) );
  INVX1 INVX1_1725 ( .A(core__abc_21380_n8070), .Y(core__abc_21380_n8071) );
  INVX1 INVX1_1726 ( .A(core_key_40_), .Y(core__abc_21380_n8073) );
  INVX1 INVX1_1727 ( .A(core__abc_21380_n7038), .Y(core__abc_21380_n8082) );
  INVX1 INVX1_1728 ( .A(core__abc_21380_n8083), .Y(core__abc_21380_n8084) );
  INVX1 INVX1_1729 ( .A(core__abc_21380_n8087), .Y(core__abc_21380_n8088) );
  INVX1 INVX1_173 ( .A(_abc_19068_n2987), .Y(_abc_19068_n2988) );
  INVX1 INVX1_1730 ( .A(core_key_41_), .Y(core__abc_21380_n8090) );
  INVX1 INVX1_1731 ( .A(core__abc_21380_n8101), .Y(core__abc_21380_n8102) );
  INVX1 INVX1_1732 ( .A(core_key_42_), .Y(core__abc_21380_n8106) );
  INVX1 INVX1_1733 ( .A(core__abc_21380_n6951), .Y(core__abc_21380_n8115) );
  INVX1 INVX1_1734 ( .A(core__abc_21380_n8117), .Y(core__abc_21380_n8118) );
  INVX1 INVX1_1735 ( .A(core__abc_21380_n7045), .Y(core__abc_21380_n8131) );
  INVX1 INVX1_1736 ( .A(core__abc_21380_n8133), .Y(core__abc_21380_n8134) );
  INVX1 INVX1_1737 ( .A(core__abc_21380_n6913), .Y(core__abc_21380_n8144) );
  INVX1 INVX1_1738 ( .A(core__abc_21380_n8146), .Y(core__abc_21380_n8147) );
  INVX1 INVX1_1739 ( .A(core__abc_21380_n8149), .Y(core__abc_21380_n8150) );
  INVX1 INVX1_174 ( .A(_abc_19068_n2992), .Y(_abc_19068_n2993) );
  INVX1 INVX1_1740 ( .A(core_key_45_), .Y(core__abc_21380_n8152) );
  INVX1 INVX1_1741 ( .A(core__abc_21380_n8163), .Y(core__abc_21380_n8164) );
  INVX1 INVX1_1742 ( .A(core_key_46_), .Y(core__abc_21380_n8168) );
  INVX1 INVX1_1743 ( .A(core__abc_21380_n6881), .Y(core__abc_21380_n8177) );
  INVX1 INVX1_1744 ( .A(core__abc_21380_n8178), .Y(core__abc_21380_n8179) );
  INVX1 INVX1_1745 ( .A(core__abc_21380_n8182), .Y(core__abc_21380_n8183) );
  INVX1 INVX1_1746 ( .A(core__abc_21380_n7047), .Y(core__abc_21380_n8193) );
  INVX1 INVX1_1747 ( .A(core__abc_21380_n8196), .Y(core__abc_21380_n8197) );
  INVX1 INVX1_1748 ( .A(core_key_48_), .Y(core__abc_21380_n8199) );
  INVX1 INVX1_1749 ( .A(core__abc_21380_n7049), .Y(core__abc_21380_n8208) );
  INVX1 INVX1_175 ( .A(_abc_19068_n2997), .Y(_abc_19068_n2998) );
  INVX1 INVX1_1750 ( .A(core__abc_21380_n8209), .Y(core__abc_21380_n8211) );
  INVX1 INVX1_1751 ( .A(core__abc_21380_n8224), .Y(core__abc_21380_n8225) );
  INVX1 INVX1_1752 ( .A(core__abc_21380_n8228), .Y(core__abc_21380_n8229) );
  INVX1 INVX1_1753 ( .A(core__abc_21380_n6830), .Y(core__abc_21380_n8239) );
  INVX1 INVX1_1754 ( .A(core__abc_21380_n8240), .Y(core__abc_21380_n8241) );
  INVX1 INVX1_1755 ( .A(core__abc_21380_n8244), .Y(core__abc_21380_n8245) );
  INVX1 INVX1_1756 ( .A(core_key_51_), .Y(core__abc_21380_n8247) );
  INVX1 INVX1_1757 ( .A(core__abc_21380_n8258), .Y(core__abc_21380_n8259) );
  INVX1 INVX1_1758 ( .A(core_key_52_), .Y(core__abc_21380_n8263) );
  INVX1 INVX1_1759 ( .A(core__abc_21380_n6813), .Y(core__abc_21380_n8272) );
  INVX1 INVX1_176 ( .A(_abc_19068_n3002), .Y(_abc_19068_n3003) );
  INVX1 INVX1_1760 ( .A(core__abc_21380_n8273), .Y(core__abc_21380_n8274) );
  INVX1 INVX1_1761 ( .A(core_key_53_), .Y(core__abc_21380_n8279) );
  INVX1 INVX1_1762 ( .A(core__abc_21380_n8291), .Y(core__abc_21380_n8292) );
  INVX1 INVX1_1763 ( .A(core__abc_21380_n8293), .Y(core__abc_21380_n8294) );
  INVX1 INVX1_1764 ( .A(core_key_54_), .Y(core__abc_21380_n8296) );
  INVX1 INVX1_1765 ( .A(core__abc_21380_n6794), .Y(core__abc_21380_n8305) );
  INVX1 INVX1_1766 ( .A(core__abc_21380_n8307), .Y(core__abc_21380_n8308) );
  INVX1 INVX1_1767 ( .A(core__abc_21380_n7057), .Y(core__abc_21380_n8321) );
  INVX1 INVX1_1768 ( .A(core__abc_21380_n8323), .Y(core__abc_21380_n8324) );
  INVX1 INVX1_1769 ( .A(core__abc_21380_n6777), .Y(core__abc_21380_n8334) );
  INVX1 INVX1_177 ( .A(_abc_19068_n3007), .Y(_abc_19068_n3008) );
  INVX1 INVX1_1770 ( .A(core__abc_21380_n8320), .Y(core__abc_21380_n8335) );
  INVX1 INVX1_1771 ( .A(core__abc_21380_n8336), .Y(core__abc_21380_n8337) );
  INVX1 INVX1_1772 ( .A(core__abc_21380_n8353), .Y(core__abc_21380_n8354) );
  INVX1 INVX1_1773 ( .A(core__abc_21380_n8355), .Y(core__abc_21380_n8356) );
  INVX1 INVX1_1774 ( .A(core_key_58_), .Y(core__abc_21380_n8358) );
  INVX1 INVX1_1775 ( .A(core__abc_21380_n6730), .Y(core__abc_21380_n8367) );
  INVX1 INVX1_1776 ( .A(core__abc_21380_n8369), .Y(core__abc_21380_n8370) );
  INVX1 INVX1_1777 ( .A(core_key_59_), .Y(core__abc_21380_n8374) );
  INVX1 INVX1_1778 ( .A(core__abc_21380_n8384), .Y(core__abc_21380_n8385) );
  INVX1 INVX1_1779 ( .A(core__abc_21380_n8388), .Y(core__abc_21380_n8389) );
  INVX1 INVX1_178 ( .A(_abc_19068_n3012), .Y(_abc_19068_n3013) );
  INVX1 INVX1_1780 ( .A(core__abc_21380_n6712), .Y(core__abc_21380_n8399) );
  INVX1 INVX1_1781 ( .A(core__abc_21380_n8387), .Y(core__abc_21380_n8400) );
  INVX1 INVX1_1782 ( .A(core__abc_21380_n8401), .Y(core__abc_21380_n8402) );
  INVX1 INVX1_1783 ( .A(core_key_61_), .Y(core__abc_21380_n8407) );
  INVX1 INVX1_1784 ( .A(core__abc_21380_n8419), .Y(core__abc_21380_n8420) );
  INVX1 INVX1_1785 ( .A(core__abc_21380_n8421), .Y(core__abc_21380_n8422) );
  INVX1 INVX1_1786 ( .A(core_key_62_), .Y(core__abc_21380_n8424) );
  INVX1 INVX1_1787 ( .A(core__abc_21380_n6693), .Y(core__abc_21380_n8433) );
  INVX1 INVX1_1788 ( .A(core__abc_21380_n8435), .Y(core__abc_21380_n8436) );
  INVX1 INVX1_1789 ( .A(core__abc_21380_n3311), .Y(core__abc_21380_n8452) );
  INVX1 INVX1_179 ( .A(_abc_19068_n3017), .Y(_abc_19068_n3018) );
  INVX1 INVX1_1790 ( .A(core__abc_21380_n7982), .Y(core__abc_21380_n8465) );
  INVX1 INVX1_1791 ( .A(core__abc_21380_n7993), .Y(core__abc_21380_n8480) );
  INVX1 INVX1_1792 ( .A(core_key_66_), .Y(core__abc_21380_n8487) );
  INVX1 INVX1_1793 ( .A(core__abc_21380_n8003), .Y(core__abc_21380_n8498) );
  INVX1 INVX1_1794 ( .A(core_key_67_), .Y(core__abc_21380_n8504) );
  INVX1 INVX1_1795 ( .A(core__abc_21380_n8015), .Y(core__abc_21380_n8514) );
  INVX1 INVX1_1796 ( .A(core__abc_21380_n8027), .Y(core__abc_21380_n8528) );
  INVX1 INVX1_1797 ( .A(core__abc_21380_n8041), .Y(core__abc_21380_n8543) );
  INVX1 INVX1_1798 ( .A(core__abc_21380_n8057), .Y(core__abc_21380_n8560) );
  INVX1 INVX1_1799 ( .A(core__abc_21380_n8565), .Y(core__abc_21380_n8566) );
  INVX1 INVX1_18 ( .A(_abc_19068_n2184), .Y(_abc_19068_n2185) );
  INVX1 INVX1_180 ( .A(_abc_19068_n3022), .Y(_abc_19068_n3023) );
  INVX1 INVX1_1800 ( .A(core_key_73_), .Y(core__abc_21380_n8592) );
  INVX1 INVX1_1801 ( .A(core__abc_21380_n8104), .Y(core__abc_21380_n8600) );
  INVX1 INVX1_1802 ( .A(core__abc_21380_n8120), .Y(core__abc_21380_n8613) );
  INVX1 INVX1_1803 ( .A(core_key_75_), .Y(core__abc_21380_n8618) );
  INVX1 INVX1_1804 ( .A(core__abc_21380_n8166), .Y(core__abc_21380_n8648) );
  INVX1 INVX1_1805 ( .A(core__abc_21380_n8213), .Y(core__abc_21380_n8683) );
  INVX1 INVX1_1806 ( .A(core__abc_21380_n8261), .Y(core__abc_21380_n8716) );
  INVX1 INVX1_1807 ( .A(core__abc_21380_n6993), .Y(core__abc_21380_n8718) );
  INVX1 INVX1_1808 ( .A(core__abc_21380_n8277), .Y(core__abc_21380_n8731) );
  INVX1 INVX1_1809 ( .A(core__abc_21380_n8310), .Y(core__abc_21380_n8754) );
  INVX1 INVX1_181 ( .A(_abc_19068_n3027), .Y(_abc_19068_n3028) );
  INVX1 INVX1_1810 ( .A(core__abc_21380_n8340), .Y(core__abc_21380_n8778) );
  INVX1 INVX1_1811 ( .A(core_key_89_), .Y(core__abc_21380_n8783) );
  INVX1 INVX1_1812 ( .A(core_key_90_), .Y(core__abc_21380_n8796) );
  INVX1 INVX1_1813 ( .A(core__abc_21380_n8372), .Y(core__abc_21380_n8805) );
  INVX1 INVX1_1814 ( .A(core__abc_21380_n6922), .Y(core__abc_21380_n8816) );
  INVX1 INVX1_1815 ( .A(core__abc_21380_n8405), .Y(core__abc_21380_n8830) );
  INVX1 INVX1_1816 ( .A(core__abc_21380_n8438), .Y(core__abc_21380_n8853) );
  INVX1 INVX1_1817 ( .A(core__abc_21380_n6877), .Y(core__abc_21380_n8865) );
  INVX1 INVX1_1818 ( .A(core_key_96_), .Y(core__abc_21380_n8870) );
  INVX1 INVX1_1819 ( .A(core__abc_21380_n6826), .Y(core__abc_21380_n8913) );
  INVX1 INVX1_182 ( .A(_abc_19068_n3032), .Y(_abc_19068_n3033) );
  INVX1 INVX1_1820 ( .A(core__abc_21380_n7187), .Y(core__abc_21380_n8914) );
  INVX1 INVX1_1821 ( .A(core__abc_21380_n7216), .Y(core__abc_21380_n8926) );
  INVX1 INVX1_1822 ( .A(core__abc_21380_n7267), .Y(core__abc_21380_n8949) );
  INVX1 INVX1_1823 ( .A(core__abc_21380_n7334), .Y(core__abc_21380_n8972) );
  INVX1 INVX1_1824 ( .A(core_key_105_), .Y(core__abc_21380_n8977) );
  INVX1 INVX1_1825 ( .A(core__abc_21380_n6725), .Y(core__abc_21380_n9008) );
  INVX1 INVX1_1826 ( .A(core_key_108_), .Y(core__abc_21380_n9015) );
  INVX1 INVX1_1827 ( .A(core__abc_21380_n7563), .Y(core__abc_21380_n9068) );
  INVX1 INVX1_1828 ( .A(core_key_113_), .Y(core__abc_21380_n9073) );
  INVX1 INVX1_1829 ( .A(core__abc_21380_n7614), .Y(core__abc_21380_n9093) );
  INVX1 INVX1_183 ( .A(_abc_19068_n3037), .Y(_abc_19068_n3038) );
  INVX1 INVX1_1830 ( .A(core_key_115_), .Y(core__abc_21380_n9098) );
  INVX1 INVX1_1831 ( .A(core__abc_21380_n7667), .Y(core__abc_21380_n9118) );
  INVX1 INVX1_1832 ( .A(core__abc_21380_n7429), .Y(core__abc_21380_n9219) );
  INVX1 INVX1_1833 ( .A(core__abc_21380_n3165), .Y(core__abc_21380_n9247) );
  INVX1 INVX1_1834 ( .A(core__abc_21380_n9249), .Y(core__abc_21380_n9250) );
  INVX1 INVX1_1835 ( .A(core_mi_reg_1_), .Y(core__abc_21380_n9261) );
  INVX1 INVX1_1836 ( .A(core_key_2_), .Y(core__abc_21380_n9273) );
  INVX1 INVX1_1837 ( .A(core_mi_reg_2_), .Y(core__abc_21380_n9275) );
  INVX1 INVX1_1838 ( .A(core_mi_reg_3_), .Y(core__abc_21380_n9287) );
  INVX1 INVX1_1839 ( .A(core_key_4_), .Y(core__abc_21380_n9299) );
  INVX1 INVX1_184 ( .A(_abc_19068_n3042), .Y(_abc_19068_n3043) );
  INVX1 INVX1_1840 ( .A(core__abc_21380_n9301), .Y(core__abc_21380_n9302) );
  INVX1 INVX1_1841 ( .A(core_mi_reg_5_), .Y(core__abc_21380_n9313) );
  INVX1 INVX1_1842 ( .A(core_mi_reg_6_), .Y(core__abc_21380_n9325) );
  INVX1 INVX1_1843 ( .A(core_mi_reg_7_), .Y(core__abc_21380_n9337) );
  INVX1 INVX1_1844 ( .A(core_key_8_), .Y(core__abc_21380_n9349) );
  INVX1 INVX1_1845 ( .A(core__abc_21380_n9351), .Y(core__abc_21380_n9352) );
  INVX1 INVX1_1846 ( .A(core_mi_reg_9_), .Y(core__abc_21380_n9364) );
  INVX1 INVX1_1847 ( .A(core_key_10_), .Y(core__abc_21380_n9376) );
  INVX1 INVX1_1848 ( .A(core__abc_21380_n9378), .Y(core__abc_21380_n9379) );
  INVX1 INVX1_1849 ( .A(core_mi_reg_11_), .Y(core__abc_21380_n9390) );
  INVX1 INVX1_185 ( .A(_abc_19068_n3047), .Y(_abc_19068_n3048) );
  INVX1 INVX1_1850 ( .A(core_v0_reg_11_), .Y(core__abc_21380_n9392) );
  INVX1 INVX1_1851 ( .A(core_mi_reg_12_), .Y(core__abc_21380_n9404) );
  INVX1 INVX1_1852 ( .A(core_mi_reg_13_), .Y(core__abc_21380_n9416) );
  INVX1 INVX1_1853 ( .A(core_mi_reg_14_), .Y(core__abc_21380_n9428) );
  INVX1 INVX1_1854 ( .A(core_mi_reg_15_), .Y(core__abc_21380_n9440) );
  INVX1 INVX1_1855 ( .A(core_mi_reg_16_), .Y(core__abc_21380_n9452) );
  INVX1 INVX1_1856 ( .A(core_key_17_), .Y(core__abc_21380_n9464) );
  INVX1 INVX1_1857 ( .A(core_mi_reg_17_), .Y(core__abc_21380_n9466) );
  INVX1 INVX1_1858 ( .A(core_mi_reg_18_), .Y(core__abc_21380_n9479) );
  INVX1 INVX1_1859 ( .A(core_v0_reg_18_), .Y(core__abc_21380_n9481) );
  INVX1 INVX1_186 ( .A(_abc_19068_n3052), .Y(_abc_19068_n3053) );
  INVX1 INVX1_1860 ( .A(core_mi_reg_19_), .Y(core__abc_21380_n9491) );
  INVX1 INVX1_1861 ( .A(core_v0_reg_19_), .Y(core__abc_21380_n9493) );
  INVX1 INVX1_1862 ( .A(core_key_20_), .Y(core__abc_21380_n9504) );
  INVX1 INVX1_1863 ( .A(core_mi_reg_20_), .Y(core__abc_21380_n9506) );
  INVX1 INVX1_1864 ( .A(core_mi_reg_21_), .Y(core__abc_21380_n9518) );
  INVX1 INVX1_1865 ( .A(core_mi_reg_22_), .Y(core__abc_21380_n9530) );
  INVX1 INVX1_1866 ( .A(core_mi_reg_23_), .Y(core__abc_21380_n9542) );
  INVX1 INVX1_1867 ( .A(core_mi_reg_24_), .Y(core__abc_21380_n9554) );
  INVX1 INVX1_1868 ( .A(core_mi_reg_25_), .Y(core__abc_21380_n9567) );
  INVX1 INVX1_1869 ( .A(core__abc_21380_n9580), .Y(core__abc_21380_n9581) );
  INVX1 INVX1_187 ( .A(_abc_19068_n3057), .Y(_abc_19068_n3058) );
  INVX1 INVX1_1870 ( .A(core_mi_reg_27_), .Y(core__abc_21380_n9593) );
  INVX1 INVX1_1871 ( .A(core_key_28_), .Y(core__abc_21380_n9605) );
  INVX1 INVX1_1872 ( .A(core_mi_reg_28_), .Y(core__abc_21380_n9607) );
  INVX1 INVX1_1873 ( .A(core_mi_reg_29_), .Y(core__abc_21380_n9619) );
  INVX1 INVX1_1874 ( .A(core_mi_reg_30_), .Y(core__abc_21380_n9631) );
  INVX1 INVX1_1875 ( .A(core_mi_reg_31_), .Y(core__abc_21380_n9643) );
  INVX1 INVX1_1876 ( .A(core_mi_reg_32_), .Y(core__abc_21380_n9655) );
  INVX1 INVX1_1877 ( .A(core_mi_reg_33_), .Y(core__abc_21380_n9667) );
  INVX1 INVX1_1878 ( .A(core_mi_reg_34_), .Y(core__abc_21380_n9679) );
  INVX1 INVX1_1879 ( .A(core_mi_reg_35_), .Y(core__abc_21380_n9691) );
  INVX1 INVX1_188 ( .A(_abc_19068_n3062), .Y(_abc_19068_n3063) );
  INVX1 INVX1_1880 ( .A(core_mi_reg_36_), .Y(core__abc_21380_n9703) );
  INVX1 INVX1_1881 ( .A(core_mi_reg_37_), .Y(core__abc_21380_n9715) );
  INVX1 INVX1_1882 ( .A(core_mi_reg_38_), .Y(core__abc_21380_n9727) );
  INVX1 INVX1_1883 ( .A(core_mi_reg_39_), .Y(core__abc_21380_n9739) );
  INVX1 INVX1_1884 ( .A(core_mi_reg_40_), .Y(core__abc_21380_n9751) );
  INVX1 INVX1_1885 ( .A(core_mi_reg_41_), .Y(core__abc_21380_n9764) );
  INVX1 INVX1_1886 ( .A(core_mi_reg_42_), .Y(core__abc_21380_n9776) );
  INVX1 INVX1_1887 ( .A(core_key_43_), .Y(core__abc_21380_n9788) );
  INVX1 INVX1_1888 ( .A(core_mi_reg_43_), .Y(core__abc_21380_n9790) );
  INVX1 INVX1_1889 ( .A(core_mi_reg_44_), .Y(core__abc_21380_n9802) );
  INVX1 INVX1_189 ( .A(_abc_19068_n3067), .Y(_abc_19068_n3068) );
  INVX1 INVX1_1890 ( .A(core_mi_reg_45_), .Y(core__abc_21380_n9814) );
  INVX1 INVX1_1891 ( .A(core_mi_reg_46_), .Y(core__abc_21380_n9826) );
  INVX1 INVX1_1892 ( .A(core_mi_reg_47_), .Y(core__abc_21380_n9838) );
  INVX1 INVX1_1893 ( .A(core_mi_reg_48_), .Y(core__abc_21380_n9850) );
  INVX1 INVX1_1894 ( .A(core_key_49_), .Y(core__abc_21380_n9862) );
  INVX1 INVX1_1895 ( .A(core_mi_reg_49_), .Y(core__abc_21380_n9864) );
  INVX1 INVX1_1896 ( .A(core_key_50_), .Y(core__abc_21380_n9876) );
  INVX1 INVX1_1897 ( .A(core_mi_reg_50_), .Y(core__abc_21380_n9878) );
  INVX1 INVX1_1898 ( .A(core_mi_reg_51_), .Y(core__abc_21380_n9890) );
  INVX1 INVX1_1899 ( .A(core__abc_21380_n9903), .Y(core__abc_21380_n9904) );
  INVX1 INVX1_19 ( .A(_abc_19068_n2190), .Y(_abc_19068_n2191) );
  INVX1 INVX1_190 ( .A(_abc_19068_n3072), .Y(_abc_19068_n3073) );
  INVX1 INVX1_1900 ( .A(core_mi_reg_53_), .Y(core__abc_21380_n9915) );
  INVX1 INVX1_1901 ( .A(core_mi_reg_54_), .Y(core__abc_21380_n9927) );
  INVX1 INVX1_1902 ( .A(core_mi_reg_55_), .Y(core__abc_21380_n9939) );
  INVX1 INVX1_1903 ( .A(core_mi_reg_56_), .Y(core__abc_21380_n9951) );
  INVX1 INVX1_1904 ( .A(core_key_56_), .Y(core__abc_21380_n9956) );
  INVX1 INVX1_1905 ( .A(core_key_57_), .Y(core__abc_21380_n9965) );
  INVX1 INVX1_1906 ( .A(core_mi_reg_57_), .Y(core__abc_21380_n9967) );
  INVX1 INVX1_1907 ( .A(core_mi_reg_58_), .Y(core__abc_21380_n9980) );
  INVX1 INVX1_1908 ( .A(core_mi_reg_59_), .Y(core__abc_21380_n9993) );
  INVX1 INVX1_1909 ( .A(core_key_60_), .Y(core__abc_21380_n10005) );
  INVX1 INVX1_191 ( .A(_abc_19068_n3077), .Y(_abc_19068_n3078) );
  INVX1 INVX1_1910 ( .A(core_mi_reg_60_), .Y(core__abc_21380_n10007) );
  INVX1 INVX1_1911 ( .A(core_mi_reg_61_), .Y(core__abc_21380_n10019) );
  INVX1 INVX1_1912 ( .A(core_mi_reg_62_), .Y(core__abc_21380_n10031) );
  INVX1 INVX1_1913 ( .A(core_mi_reg_63_), .Y(core__abc_21380_n10043) );
  INVX1 INVX1_1914 ( .A(core__abc_21380_n1143), .Y(core__abc_21380_n10061) );
  INVX1 INVX1_192 ( .A(_abc_19068_n3082), .Y(_abc_19068_n3083) );
  INVX1 INVX1_193 ( .A(_abc_19068_n3087), .Y(_abc_19068_n3088) );
  INVX1 INVX1_194 ( .A(_abc_19068_n3092), .Y(_abc_19068_n3093) );
  INVX1 INVX1_195 ( .A(_abc_19068_n3097), .Y(_abc_19068_n3098) );
  INVX1 INVX1_196 ( .A(_abc_19068_n3102), .Y(_abc_19068_n3103) );
  INVX1 INVX1_197 ( .A(_abc_19068_n3107), .Y(_abc_19068_n3108) );
  INVX1 INVX1_198 ( .A(_abc_19068_n3112), .Y(_abc_19068_n3113) );
  INVX1 INVX1_199 ( .A(_abc_19068_n3117), .Y(_abc_19068_n3118) );
  INVX1 INVX1_2 ( .A(\addr[1] ), .Y(_abc_19068_n872) );
  INVX1 INVX1_20 ( .A(_abc_19068_n2196), .Y(_abc_19068_n2197) );
  INVX1 INVX1_200 ( .A(_abc_19068_n3122), .Y(_abc_19068_n3123) );
  INVX1 INVX1_201 ( .A(_abc_19068_n3127), .Y(_abc_19068_n3128) );
  INVX1 INVX1_202 ( .A(reset_n_bF_buf18), .Y(_abc_19068_n3138) );
  INVX1 INVX1_203 ( .A(_abc_19068_n3176), .Y(_abc_19068_n3177) );
  INVX1 INVX1_204 ( .A(core_finalize), .Y(core__abc_21380_n1130_1) );
  INVX1 INVX1_205 ( .A(core_compress), .Y(core__abc_21380_n1131) );
  INVX1 INVX1_206 ( .A(core_siphash_ctrl_reg_1_), .Y(core__abc_21380_n1133_1) );
  INVX1 INVX1_207 ( .A(core_siphash_ctrl_reg_2_), .Y(core__abc_21380_n1136_1) );
  INVX1 INVX1_208 ( .A(core_siphash_ctrl_reg_5_), .Y(core__abc_21380_n1137_1) );
  INVX1 INVX1_209 ( .A(core__abc_21380_n1132_1), .Y(core__abc_21380_n1145_1) );
  INVX1 INVX1_21 ( .A(_abc_19068_n2202), .Y(_abc_19068_n2203) );
  INVX1 INVX1_210 ( .A(core_compression_rounds_3_), .Y(core__abc_21380_n1148_1) );
  INVX1 INVX1_211 ( .A(core_compression_rounds_2_), .Y(core__abc_21380_n1149_1) );
  INVX1 INVX1_212 ( .A(core_compression_rounds_1_), .Y(core__abc_21380_n1150_1) );
  INVX1 INVX1_213 ( .A(core_compression_rounds_0_), .Y(core__abc_21380_n1151) );
  INVX1 INVX1_214 ( .A(core_loop_ctr_reg_0_), .Y(core__abc_21380_n1155) );
  INVX1 INVX1_215 ( .A(core_loop_ctr_reg_1_), .Y(core__abc_21380_n1157_1) );
  INVX1 INVX1_216 ( .A(core__abc_21380_n1159), .Y(core__abc_21380_n1160_1) );
  INVX1 INVX1_217 ( .A(core__abc_21380_n1166_1), .Y(core__abc_21380_n1167) );
  INVX1 INVX1_218 ( .A(core__abc_21380_n1153_1), .Y(core__abc_21380_n1168_1) );
  INVX1 INVX1_219 ( .A(core__abc_21380_n1171), .Y(core__abc_21380_n1172_1) );
  INVX1 INVX1_22 ( .A(_abc_19068_n2208), .Y(_abc_19068_n2209) );
  INVX1 INVX1_220 ( .A(core__abc_21380_n1177_1), .Y(core__abc_21380_n1178_1) );
  INVX1 INVX1_221 ( .A(core_loop_ctr_reg_3_), .Y(core__abc_21380_n1180_1) );
  INVX1 INVX1_222 ( .A(core__abc_21380_n1182_1), .Y(core__abc_21380_n1183) );
  INVX1 INVX1_223 ( .A(core_final_rounds_3_), .Y(core__abc_21380_n1186_1) );
  INVX1 INVX1_224 ( .A(core_final_rounds_2_), .Y(core__abc_21380_n1187) );
  INVX1 INVX1_225 ( .A(core_final_rounds_1_), .Y(core__abc_21380_n1188_1) );
  INVX1 INVX1_226 ( .A(core_final_rounds_0_), .Y(core__abc_21380_n1189_1) );
  INVX1 INVX1_227 ( .A(core__abc_21380_n1197_1), .Y(core__abc_21380_n1198_1) );
  INVX1 INVX1_228 ( .A(core__abc_21380_n1202_1), .Y(core__abc_21380_n1203) );
  INVX1 INVX1_229 ( .A(core_loop_ctr_reg_2_), .Y(core__abc_21380_n1204_1) );
  INVX1 INVX1_23 ( .A(_abc_19068_n2214), .Y(_abc_19068_n2215) );
  INVX1 INVX1_230 ( .A(core__abc_21380_n1191), .Y(core__abc_21380_n1205_1) );
  INVX1 INVX1_231 ( .A(core__abc_21380_n1207), .Y(core__abc_21380_n1208_1) );
  INVX1 INVX1_232 ( .A(core__abc_21380_n1214_1), .Y(core__abc_21380_n1215) );
  INVX1 INVX1_233 ( .A(core__abc_21380_n1218_1), .Y(core__abc_21380_n1219) );
  INVX1 INVX1_234 ( .A(core__abc_21380_n1139), .Y(core__abc_21380_n1222_1) );
  INVX1 INVX1_235 ( .A(core__abc_21380_n1220_1), .Y(core__abc_21380_n1230_1) );
  INVX1 INVX1_236 ( .A(core__abc_21380_n1184_1), .Y(core__abc_21380_n1232_1) );
  INVX1 INVX1_237 ( .A(core__abc_21380_n1225_1), .Y(core__abc_21380_n1238_1) );
  INVX1 INVX1_238 ( .A(core__abc_21380_n1135), .Y(core__abc_21380_n1241_1) );
  INVX1 INVX1_239 ( .A(reset_n_bF_buf8), .Y(core__abc_21380_n1242_1) );
  INVX1 INVX1_24 ( .A(_abc_19068_n2220), .Y(_abc_19068_n2221) );
  INVX1 INVX1_240 ( .A(core__abc_21380_n1260_1), .Y(core__abc_21380_n1261_1) );
  INVX1 INVX1_241 ( .A(core_v3_reg_0_), .Y(core__abc_21380_n1263) );
  INVX1 INVX1_242 ( .A(core_v2_reg_0_), .Y(core__abc_21380_n1264_1) );
  INVX1 INVX1_243 ( .A(core__abc_21380_n1267), .Y(core__abc_21380_n1268_1) );
  INVX1 INVX1_244 ( .A(core__abc_21380_n1262_1), .Y(core__abc_21380_n1270_1) );
  INVX1 INVX1_245 ( .A(core__abc_21380_n1278_1), .Y(core__abc_21380_n1279) );
  INVX1 INVX1_246 ( .A(core_v3_reg_1_), .Y(core__abc_21380_n1282_1) );
  INVX1 INVX1_247 ( .A(core_v2_reg_1_), .Y(core__abc_21380_n1283) );
  INVX1 INVX1_248 ( .A(core__abc_21380_n1285_1), .Y(core__abc_21380_n1286_1) );
  INVX1 INVX1_249 ( .A(core_v0_reg_1_), .Y(core__abc_21380_n1288_1) );
  INVX1 INVX1_25 ( .A(_abc_19068_n2226), .Y(_abc_19068_n2227) );
  INVX1 INVX1_250 ( .A(core_v1_reg_1_), .Y(core__abc_21380_n1289) );
  INVX1 INVX1_251 ( .A(core_v0_reg_2_), .Y(core__abc_21380_n1298) );
  INVX1 INVX1_252 ( .A(core_v1_reg_2_), .Y(core__abc_21380_n1299) );
  INVX1 INVX1_253 ( .A(core__abc_21380_n1302), .Y(core__abc_21380_n1303) );
  INVX1 INVX1_254 ( .A(core_v3_reg_2_), .Y(core__abc_21380_n1305) );
  INVX1 INVX1_255 ( .A(core_v2_reg_2_), .Y(core__abc_21380_n1306) );
  INVX1 INVX1_256 ( .A(core__abc_21380_n1308), .Y(core__abc_21380_n1309) );
  INVX1 INVX1_257 ( .A(core_v0_reg_3_), .Y(core__abc_21380_n1318) );
  INVX1 INVX1_258 ( .A(core_v1_reg_3_), .Y(core__abc_21380_n1319) );
  INVX1 INVX1_259 ( .A(core__abc_21380_n1321), .Y(core__abc_21380_n1322) );
  INVX1 INVX1_26 ( .A(_abc_19068_n2232), .Y(_abc_19068_n2233) );
  INVX1 INVX1_260 ( .A(core_v2_reg_3_), .Y(core__abc_21380_n1324) );
  INVX1 INVX1_261 ( .A(core_v3_reg_3_), .Y(core__abc_21380_n1325) );
  INVX1 INVX1_262 ( .A(core__abc_21380_n1327), .Y(core__abc_21380_n1329) );
  INVX1 INVX1_263 ( .A(core__abc_21380_n1337), .Y(core__abc_21380_n1338) );
  INVX1 INVX1_264 ( .A(core_v3_reg_4_), .Y(core__abc_21380_n1341) );
  INVX1 INVX1_265 ( .A(core_v2_reg_4_), .Y(core__abc_21380_n1342) );
  INVX1 INVX1_266 ( .A(core__abc_21380_n1344), .Y(core__abc_21380_n1345) );
  INVX1 INVX1_267 ( .A(core__abc_21380_n1339), .Y(core__abc_21380_n1347) );
  INVX1 INVX1_268 ( .A(core_v0_reg_5_), .Y(core__abc_21380_n1355) );
  INVX1 INVX1_269 ( .A(core_v1_reg_5_), .Y(core__abc_21380_n1356) );
  INVX1 INVX1_27 ( .A(_abc_19068_n2238), .Y(_abc_19068_n2239) );
  INVX1 INVX1_270 ( .A(core__abc_21380_n1358), .Y(core__abc_21380_n1359) );
  INVX1 INVX1_271 ( .A(core_v2_reg_5_), .Y(core__abc_21380_n1361) );
  INVX1 INVX1_272 ( .A(core_v3_reg_5_), .Y(core__abc_21380_n1362) );
  INVX1 INVX1_273 ( .A(core__abc_21380_n1364), .Y(core__abc_21380_n1366) );
  INVX1 INVX1_274 ( .A(core_v0_reg_6_), .Y(core__abc_21380_n1373) );
  INVX1 INVX1_275 ( .A(core_v1_reg_6_), .Y(core__abc_21380_n1374) );
  INVX1 INVX1_276 ( .A(core__abc_21380_n1377), .Y(core__abc_21380_n1378) );
  INVX1 INVX1_277 ( .A(core_v3_reg_6_), .Y(core__abc_21380_n1380) );
  INVX1 INVX1_278 ( .A(core_v2_reg_6_), .Y(core__abc_21380_n1381) );
  INVX1 INVX1_279 ( .A(core__abc_21380_n1383), .Y(core__abc_21380_n1384) );
  INVX1 INVX1_28 ( .A(_abc_19068_n2244), .Y(_abc_19068_n2245) );
  INVX1 INVX1_280 ( .A(core_v0_reg_7_), .Y(core__abc_21380_n1392) );
  INVX1 INVX1_281 ( .A(core_v1_reg_7_), .Y(core__abc_21380_n1393) );
  INVX1 INVX1_282 ( .A(core__abc_21380_n1396), .Y(core__abc_21380_n1397) );
  INVX1 INVX1_283 ( .A(core_v3_reg_7_), .Y(core__abc_21380_n1399) );
  INVX1 INVX1_284 ( .A(core_v2_reg_7_), .Y(core__abc_21380_n1400) );
  INVX1 INVX1_285 ( .A(core__abc_21380_n1402), .Y(core__abc_21380_n1403) );
  INVX1 INVX1_286 ( .A(core__abc_21380_n1411), .Y(core__abc_21380_n1412) );
  INVX1 INVX1_287 ( .A(core__abc_21380_n1415), .Y(core__abc_21380_n1416) );
  INVX1 INVX1_288 ( .A(core__abc_21380_n1418), .Y(core__abc_21380_n1419) );
  INVX1 INVX1_289 ( .A(core__abc_21380_n1414), .Y(core__abc_21380_n1421) );
  INVX1 INVX1_29 ( .A(_abc_19068_n2250), .Y(_abc_19068_n2251) );
  INVX1 INVX1_290 ( .A(core__abc_21380_n1428), .Y(core__abc_21380_n1429) );
  INVX1 INVX1_291 ( .A(core_v0_reg_9_), .Y(core__abc_21380_n1430) );
  INVX1 INVX1_292 ( .A(core_v1_reg_9_), .Y(core__abc_21380_n1431) );
  INVX1 INVX1_293 ( .A(core__abc_21380_n1432), .Y(core__abc_21380_n1433) );
  INVX1 INVX1_294 ( .A(core__abc_21380_n1435), .Y(core__abc_21380_n1436) );
  INVX1 INVX1_295 ( .A(core__abc_21380_n1438), .Y(core__abc_21380_n1439) );
  INVX1 INVX1_296 ( .A(core__abc_21380_n1434), .Y(core__abc_21380_n1441) );
  INVX1 INVX1_297 ( .A(core__abc_21380_n1449), .Y(core__abc_21380_n1450) );
  INVX1 INVX1_298 ( .A(core__abc_21380_n1452), .Y(core__abc_21380_n1453) );
  INVX1 INVX1_299 ( .A(core__abc_21380_n1451), .Y(core__abc_21380_n1457) );
  INVX1 INVX1_3 ( .A(\addr[7] ), .Y(_abc_19068_n875) );
  INVX1 INVX1_30 ( .A(_abc_19068_n2256), .Y(_abc_19068_n2257) );
  INVX1 INVX1_300 ( .A(core__abc_21380_n1455), .Y(core__abc_21380_n1458) );
  INVX1 INVX1_301 ( .A(core__abc_21380_n1466), .Y(core__abc_21380_n1467) );
  INVX1 INVX1_302 ( .A(core__abc_21380_n1469), .Y(core__abc_21380_n1470) );
  INVX1 INVX1_303 ( .A(core__abc_21380_n1468), .Y(core__abc_21380_n1474) );
  INVX1 INVX1_304 ( .A(core__abc_21380_n1472), .Y(core__abc_21380_n1475) );
  INVX1 INVX1_305 ( .A(core_v0_reg_12_), .Y(core__abc_21380_n1483) );
  INVX1 INVX1_306 ( .A(core_v1_reg_12_), .Y(core__abc_21380_n1484) );
  INVX1 INVX1_307 ( .A(core__abc_21380_n1486), .Y(core__abc_21380_n1487) );
  INVX1 INVX1_308 ( .A(core__abc_21380_n1488), .Y(core__abc_21380_n1489) );
  INVX1 INVX1_309 ( .A(core__abc_21380_n1491), .Y(core__abc_21380_n1492) );
  INVX1 INVX1_31 ( .A(_abc_19068_n2262), .Y(_abc_19068_n2263) );
  INVX1 INVX1_310 ( .A(core_v0_reg_13_), .Y(core__abc_21380_n1500) );
  INVX1 INVX1_311 ( .A(core_v1_reg_13_), .Y(core__abc_21380_n1501) );
  INVX1 INVX1_312 ( .A(core__abc_21380_n1504), .Y(core__abc_21380_n1505) );
  INVX1 INVX1_313 ( .A(core__abc_21380_n1506), .Y(core__abc_21380_n1507) );
  INVX1 INVX1_314 ( .A(core__abc_21380_n1509), .Y(core__abc_21380_n1511) );
  INVX1 INVX1_315 ( .A(core_v0_reg_14_), .Y(core__abc_21380_n1518) );
  INVX1 INVX1_316 ( .A(core_v1_reg_14_), .Y(core__abc_21380_n1519) );
  INVX1 INVX1_317 ( .A(core__abc_21380_n1522), .Y(core__abc_21380_n1523) );
  INVX1 INVX1_318 ( .A(core__abc_21380_n1524), .Y(core__abc_21380_n1525) );
  INVX1 INVX1_319 ( .A(core__abc_21380_n1527), .Y(core__abc_21380_n1529) );
  INVX1 INVX1_32 ( .A(_abc_19068_n2268), .Y(_abc_19068_n2269) );
  INVX1 INVX1_320 ( .A(core_v0_reg_15_), .Y(core__abc_21380_n1536) );
  INVX1 INVX1_321 ( .A(core_v1_reg_15_), .Y(core__abc_21380_n1537) );
  INVX1 INVX1_322 ( .A(core__abc_21380_n1538), .Y(core__abc_21380_n1539) );
  INVX1 INVX1_323 ( .A(core__abc_21380_n1540), .Y(core__abc_21380_n1541) );
  INVX1 INVX1_324 ( .A(core__abc_21380_n1543), .Y(core__abc_21380_n1544) );
  INVX1 INVX1_325 ( .A(core__abc_21380_n1542), .Y(core__abc_21380_n1548) );
  INVX1 INVX1_326 ( .A(core__abc_21380_n1546), .Y(core__abc_21380_n1549) );
  INVX1 INVX1_327 ( .A(core_v0_reg_16_), .Y(core__abc_21380_n1557) );
  INVX1 INVX1_328 ( .A(core_v1_reg_16_), .Y(core__abc_21380_n1558) );
  INVX1 INVX1_329 ( .A(core__abc_21380_n1560), .Y(core__abc_21380_n1561) );
  INVX1 INVX1_33 ( .A(_abc_19068_n2274), .Y(_abc_19068_n2275) );
  INVX1 INVX1_330 ( .A(core__abc_21380_n1562), .Y(core__abc_21380_n1563) );
  INVX1 INVX1_331 ( .A(core__abc_21380_n1565), .Y(core__abc_21380_n1566) );
  INVX1 INVX1_332 ( .A(core__abc_21380_n1574), .Y(core__abc_21380_n1575) );
  INVX1 INVX1_333 ( .A(core_v0_reg_17_), .Y(core__abc_21380_n1576) );
  INVX1 INVX1_334 ( .A(core_v1_reg_17_), .Y(core__abc_21380_n1577) );
  INVX1 INVX1_335 ( .A(core__abc_21380_n1578), .Y(core__abc_21380_n1579) );
  INVX1 INVX1_336 ( .A(core__abc_21380_n1581), .Y(core__abc_21380_n1582) );
  INVX1 INVX1_337 ( .A(core__abc_21380_n1584), .Y(core__abc_21380_n1585) );
  INVX1 INVX1_338 ( .A(core__abc_21380_n1580), .Y(core__abc_21380_n1587) );
  INVX1 INVX1_339 ( .A(core__abc_21380_n1595), .Y(core__abc_21380_n1596) );
  INVX1 INVX1_34 ( .A(_abc_19068_n2280), .Y(_abc_19068_n2281) );
  INVX1 INVX1_340 ( .A(core__abc_21380_n1598), .Y(core__abc_21380_n1599) );
  INVX1 INVX1_341 ( .A(core__abc_21380_n1597), .Y(core__abc_21380_n1603) );
  INVX1 INVX1_342 ( .A(core__abc_21380_n1601), .Y(core__abc_21380_n1604) );
  INVX1 INVX1_343 ( .A(core__abc_21380_n1611), .Y(core__abc_21380_n1612) );
  INVX1 INVX1_344 ( .A(core__abc_21380_n1615), .Y(core__abc_21380_n1616) );
  INVX1 INVX1_345 ( .A(core__abc_21380_n1618), .Y(core__abc_21380_n1619) );
  INVX1 INVX1_346 ( .A(core__abc_21380_n1614), .Y(core__abc_21380_n1621) );
  INVX1 INVX1_347 ( .A(core_v0_reg_20_), .Y(core__abc_21380_n1628) );
  INVX1 INVX1_348 ( .A(core_v1_reg_20_), .Y(core__abc_21380_n1629) );
  INVX1 INVX1_349 ( .A(core__abc_21380_n1632), .Y(core__abc_21380_n1633) );
  INVX1 INVX1_35 ( .A(_abc_19068_n2286), .Y(_abc_19068_n2287) );
  INVX1 INVX1_350 ( .A(core__abc_21380_n1634), .Y(core__abc_21380_n1635) );
  INVX1 INVX1_351 ( .A(core__abc_21380_n1637), .Y(core__abc_21380_n1639) );
  INVX1 INVX1_352 ( .A(core_v0_reg_21_), .Y(core__abc_21380_n1646) );
  INVX1 INVX1_353 ( .A(core_v1_reg_21_), .Y(core__abc_21380_n1647) );
  INVX1 INVX1_354 ( .A(core__abc_21380_n1650), .Y(core__abc_21380_n1651) );
  INVX1 INVX1_355 ( .A(core__abc_21380_n1652), .Y(core__abc_21380_n1653) );
  INVX1 INVX1_356 ( .A(core__abc_21380_n1655_1), .Y(core__abc_21380_n1657) );
  INVX1 INVX1_357 ( .A(core_v0_reg_22_), .Y(core__abc_21380_n1664) );
  INVX1 INVX1_358 ( .A(core_v1_reg_22_), .Y(core__abc_21380_n1665) );
  INVX1 INVX1_359 ( .A(core__abc_21380_n1668), .Y(core__abc_21380_n1669) );
  INVX1 INVX1_36 ( .A(_abc_19068_n2292), .Y(_abc_19068_n2293) );
  INVX1 INVX1_360 ( .A(core__abc_21380_n1670), .Y(core__abc_21380_n1671) );
  INVX1 INVX1_361 ( .A(core__abc_21380_n1673), .Y(core__abc_21380_n1675) );
  INVX1 INVX1_362 ( .A(core_v0_reg_23_), .Y(core__abc_21380_n1682) );
  INVX1 INVX1_363 ( .A(core_v1_reg_23_), .Y(core__abc_21380_n1683) );
  INVX1 INVX1_364 ( .A(core__abc_21380_n1684), .Y(core__abc_21380_n1685) );
  INVX1 INVX1_365 ( .A(core__abc_21380_n1686), .Y(core__abc_21380_n1687) );
  INVX1 INVX1_366 ( .A(core__abc_21380_n1689), .Y(core__abc_21380_n1690) );
  INVX1 INVX1_367 ( .A(core__abc_21380_n1688), .Y(core__abc_21380_n1694) );
  INVX1 INVX1_368 ( .A(core__abc_21380_n1692), .Y(core__abc_21380_n1695) );
  INVX1 INVX1_369 ( .A(core_v0_reg_24_), .Y(core__abc_21380_n1702) );
  INVX1 INVX1_37 ( .A(_abc_19068_n2298), .Y(_abc_19068_n2299) );
  INVX1 INVX1_370 ( .A(core_v1_reg_24_), .Y(core__abc_21380_n1703) );
  INVX1 INVX1_371 ( .A(core__abc_21380_n1706), .Y(core__abc_21380_n1707) );
  INVX1 INVX1_372 ( .A(core__abc_21380_n1708), .Y(core__abc_21380_n1709) );
  INVX1 INVX1_373 ( .A(core__abc_21380_n1711), .Y(core__abc_21380_n1713) );
  INVX1 INVX1_374 ( .A(core_v0_reg_25_), .Y(core__abc_21380_n1720) );
  INVX1 INVX1_375 ( .A(core_v1_reg_25_), .Y(core__abc_21380_n1721) );
  INVX1 INVX1_376 ( .A(core__abc_21380_n1722), .Y(core__abc_21380_n1723) );
  INVX1 INVX1_377 ( .A(core__abc_21380_n1724), .Y(core__abc_21380_n1725) );
  INVX1 INVX1_378 ( .A(core__abc_21380_n1727), .Y(core__abc_21380_n1728) );
  INVX1 INVX1_379 ( .A(core__abc_21380_n1726), .Y(core__abc_21380_n1732) );
  INVX1 INVX1_38 ( .A(_abc_19068_n2304), .Y(_abc_19068_n2305) );
  INVX1 INVX1_380 ( .A(core__abc_21380_n1730), .Y(core__abc_21380_n1733) );
  INVX1 INVX1_381 ( .A(core__abc_21380_n1741), .Y(core__abc_21380_n1742) );
  INVX1 INVX1_382 ( .A(core__abc_21380_n1744), .Y(core__abc_21380_n1745) );
  INVX1 INVX1_383 ( .A(core__abc_21380_n1743), .Y(core__abc_21380_n1749) );
  INVX1 INVX1_384 ( .A(core__abc_21380_n1747), .Y(core__abc_21380_n1750) );
  INVX1 INVX1_385 ( .A(core_v0_reg_27_), .Y(core__abc_21380_n1757) );
  INVX1 INVX1_386 ( .A(core_v1_reg_27_), .Y(core__abc_21380_n1758) );
  INVX1 INVX1_387 ( .A(core__abc_21380_n1759), .Y(core__abc_21380_n1760_1) );
  INVX1 INVX1_388 ( .A(core__abc_21380_n1761), .Y(core__abc_21380_n1762) );
  INVX1 INVX1_389 ( .A(core__abc_21380_n1764), .Y(core__abc_21380_n1765) );
  INVX1 INVX1_39 ( .A(_abc_19068_n2310), .Y(_abc_19068_n2311) );
  INVX1 INVX1_390 ( .A(core__abc_21380_n1763), .Y(core__abc_21380_n1769) );
  INVX1 INVX1_391 ( .A(core__abc_21380_n1767), .Y(core__abc_21380_n1770) );
  INVX1 INVX1_392 ( .A(core_v0_reg_28_), .Y(core__abc_21380_n1777) );
  INVX1 INVX1_393 ( .A(core_v1_reg_28_), .Y(core__abc_21380_n1778) );
  INVX1 INVX1_394 ( .A(core__abc_21380_n1781), .Y(core__abc_21380_n1782_1) );
  INVX1 INVX1_395 ( .A(core__abc_21380_n1783), .Y(core__abc_21380_n1784) );
  INVX1 INVX1_396 ( .A(core__abc_21380_n1786_1), .Y(core__abc_21380_n1788) );
  INVX1 INVX1_397 ( .A(core_v0_reg_29_), .Y(core__abc_21380_n1795) );
  INVX1 INVX1_398 ( .A(core_v1_reg_29_), .Y(core__abc_21380_n1796) );
  INVX1 INVX1_399 ( .A(core__abc_21380_n1797), .Y(core__abc_21380_n1798) );
  INVX1 INVX1_4 ( .A(\addr[6] ), .Y(_abc_19068_n876_1) );
  INVX1 INVX1_40 ( .A(_abc_19068_n2316), .Y(_abc_19068_n2317) );
  INVX1 INVX1_400 ( .A(core__abc_21380_n1799), .Y(core__abc_21380_n1800) );
  INVX1 INVX1_401 ( .A(core__abc_21380_n1802), .Y(core__abc_21380_n1803) );
  INVX1 INVX1_402 ( .A(core__abc_21380_n1801), .Y(core__abc_21380_n1807) );
  INVX1 INVX1_403 ( .A(core__abc_21380_n1805), .Y(core__abc_21380_n1808) );
  INVX1 INVX1_404 ( .A(core_v0_reg_30_), .Y(core__abc_21380_n1815) );
  INVX1 INVX1_405 ( .A(core_v1_reg_30_), .Y(core__abc_21380_n1816_1) );
  INVX1 INVX1_406 ( .A(core__abc_21380_n1819), .Y(core__abc_21380_n1820) );
  INVX1 INVX1_407 ( .A(core__abc_21380_n1821), .Y(core__abc_21380_n1822) );
  INVX1 INVX1_408 ( .A(core__abc_21380_n1824), .Y(core__abc_21380_n1826) );
  INVX1 INVX1_409 ( .A(core_v0_reg_31_), .Y(core__abc_21380_n1833) );
  INVX1 INVX1_41 ( .A(_abc_19068_n2322), .Y(_abc_19068_n2323) );
  INVX1 INVX1_410 ( .A(core_v1_reg_31_), .Y(core__abc_21380_n1834) );
  INVX1 INVX1_411 ( .A(core__abc_21380_n1835), .Y(core__abc_21380_n1836) );
  INVX1 INVX1_412 ( .A(core__abc_21380_n1837), .Y(core__abc_21380_n1838) );
  INVX1 INVX1_413 ( .A(core__abc_21380_n1840), .Y(core__abc_21380_n1841) );
  INVX1 INVX1_414 ( .A(core__abc_21380_n1839), .Y(core__abc_21380_n1845) );
  INVX1 INVX1_415 ( .A(core__abc_21380_n1843), .Y(core__abc_21380_n1846_1) );
  INVX1 INVX1_416 ( .A(core_v0_reg_32_), .Y(core__abc_21380_n1853) );
  INVX1 INVX1_417 ( .A(core_v1_reg_32_), .Y(core__abc_21380_n1854) );
  INVX1 INVX1_418 ( .A(core__abc_21380_n1857), .Y(core__abc_21380_n1858) );
  INVX1 INVX1_419 ( .A(core__abc_21380_n1859), .Y(core__abc_21380_n1860) );
  INVX1 INVX1_42 ( .A(_abc_19068_n2328), .Y(_abc_19068_n2329) );
  INVX1 INVX1_420 ( .A(core__abc_21380_n1862), .Y(core__abc_21380_n1864) );
  INVX1 INVX1_421 ( .A(core_v0_reg_33_), .Y(core__abc_21380_n1871) );
  INVX1 INVX1_422 ( .A(core_v1_reg_33_), .Y(core__abc_21380_n1872) );
  INVX1 INVX1_423 ( .A(core__abc_21380_n1877), .Y(core__abc_21380_n1878) );
  INVX1 INVX1_424 ( .A(core__abc_21380_n1880), .Y(core__abc_21380_n1882) );
  INVX1 INVX1_425 ( .A(core_v0_reg_34_), .Y(core__abc_21380_n1889) );
  INVX1 INVX1_426 ( .A(core_v1_reg_34_), .Y(core__abc_21380_n1890) );
  INVX1 INVX1_427 ( .A(core__abc_21380_n1893), .Y(core__abc_21380_n1894_1) );
  INVX1 INVX1_428 ( .A(core__abc_21380_n1895), .Y(core__abc_21380_n1896) );
  INVX1 INVX1_429 ( .A(core__abc_21380_n1898), .Y(core__abc_21380_n1900) );
  INVX1 INVX1_43 ( .A(_abc_19068_n2333), .Y(_abc_19068_n2334) );
  INVX1 INVX1_430 ( .A(core_v0_reg_35_), .Y(core__abc_21380_n1907) );
  INVX1 INVX1_431 ( .A(core_v1_reg_35_), .Y(core__abc_21380_n1908) );
  INVX1 INVX1_432 ( .A(core__abc_21380_n1909), .Y(core__abc_21380_n1910) );
  INVX1 INVX1_433 ( .A(core__abc_21380_n1911), .Y(core__abc_21380_n1912) );
  INVX1 INVX1_434 ( .A(core__abc_21380_n1914), .Y(core__abc_21380_n1915) );
  INVX1 INVX1_435 ( .A(core__abc_21380_n1913), .Y(core__abc_21380_n1919) );
  INVX1 INVX1_436 ( .A(core__abc_21380_n1917), .Y(core__abc_21380_n1920) );
  INVX1 INVX1_437 ( .A(core_v0_reg_36_), .Y(core__abc_21380_n1928_1) );
  INVX1 INVX1_438 ( .A(core_v1_reg_36_), .Y(core__abc_21380_n1929) );
  INVX1 INVX1_439 ( .A(core__abc_21380_n1932), .Y(core__abc_21380_n1933) );
  INVX1 INVX1_44 ( .A(_abc_19068_n2338), .Y(_abc_19068_n2339) );
  INVX1 INVX1_440 ( .A(core__abc_21380_n1931), .Y(core__abc_21380_n1937) );
  INVX1 INVX1_441 ( .A(core__abc_21380_n1935), .Y(core__abc_21380_n1938) );
  INVX1 INVX1_442 ( .A(core__abc_21380_n1945), .Y(core__abc_21380_n1946) );
  INVX1 INVX1_443 ( .A(core_v0_reg_37_), .Y(core__abc_21380_n1947) );
  INVX1 INVX1_444 ( .A(core_v1_reg_37_), .Y(core__abc_21380_n1948) );
  INVX1 INVX1_445 ( .A(core__abc_21380_n1949), .Y(core__abc_21380_n1950) );
  INVX1 INVX1_446 ( .A(core__abc_21380_n1952), .Y(core__abc_21380_n1953) );
  INVX1 INVX1_447 ( .A(core__abc_21380_n1955), .Y(core__abc_21380_n1956) );
  INVX1 INVX1_448 ( .A(core__abc_21380_n1951), .Y(core__abc_21380_n1958) );
  INVX1 INVX1_449 ( .A(core_v0_reg_38_), .Y(core__abc_21380_n1965_1) );
  INVX1 INVX1_45 ( .A(_abc_19068_n2343), .Y(_abc_19068_n2344) );
  INVX1 INVX1_450 ( .A(core_v1_reg_38_), .Y(core__abc_21380_n1966) );
  INVX1 INVX1_451 ( .A(core__abc_21380_n1969), .Y(core__abc_21380_n1970) );
  INVX1 INVX1_452 ( .A(core__abc_21380_n1971), .Y(core__abc_21380_n1972) );
  INVX1 INVX1_453 ( .A(core__abc_21380_n1974), .Y(core__abc_21380_n1976) );
  INVX1 INVX1_454 ( .A(core_v0_reg_39_), .Y(core__abc_21380_n1983) );
  INVX1 INVX1_455 ( .A(core_v1_reg_39_), .Y(core__abc_21380_n1984) );
  INVX1 INVX1_456 ( .A(core__abc_21380_n1985), .Y(core__abc_21380_n1986) );
  INVX1 INVX1_457 ( .A(core__abc_21380_n1987), .Y(core__abc_21380_n1988) );
  INVX1 INVX1_458 ( .A(core__abc_21380_n1990), .Y(core__abc_21380_n1991) );
  INVX1 INVX1_459 ( .A(core__abc_21380_n1989), .Y(core__abc_21380_n1995_1) );
  INVX1 INVX1_46 ( .A(_abc_19068_n2348), .Y(_abc_19068_n2349) );
  INVX1 INVX1_460 ( .A(core__abc_21380_n1993), .Y(core__abc_21380_n1996) );
  INVX1 INVX1_461 ( .A(core_v0_reg_40_), .Y(core__abc_21380_n2004) );
  INVX1 INVX1_462 ( .A(core_v1_reg_40_), .Y(core__abc_21380_n2005) );
  INVX1 INVX1_463 ( .A(core__abc_21380_n2007), .Y(core__abc_21380_n2008) );
  INVX1 INVX1_464 ( .A(core__abc_21380_n2009), .Y(core__abc_21380_n2010) );
  INVX1 INVX1_465 ( .A(core__abc_21380_n2012), .Y(core__abc_21380_n2013) );
  INVX1 INVX1_466 ( .A(core_v0_reg_41_), .Y(core__abc_21380_n2022) );
  INVX1 INVX1_467 ( .A(core_v1_reg_41_), .Y(core__abc_21380_n2023) );
  INVX1 INVX1_468 ( .A(core__abc_21380_n2026), .Y(core__abc_21380_n2027) );
  INVX1 INVX1_469 ( .A(core__abc_21380_n2025), .Y(core__abc_21380_n2031) );
  INVX1 INVX1_47 ( .A(_abc_19068_n2353), .Y(_abc_19068_n2354) );
  INVX1 INVX1_470 ( .A(core__abc_21380_n2029), .Y(core__abc_21380_n2032) );
  INVX1 INVX1_471 ( .A(core_v0_reg_42_), .Y(core__abc_21380_n2039_1) );
  INVX1 INVX1_472 ( .A(core_v1_reg_42_), .Y(core__abc_21380_n2040) );
  INVX1 INVX1_473 ( .A(core__abc_21380_n2043), .Y(core__abc_21380_n2044) );
  INVX1 INVX1_474 ( .A(core__abc_21380_n2045), .Y(core__abc_21380_n2046) );
  INVX1 INVX1_475 ( .A(core__abc_21380_n2048), .Y(core__abc_21380_n2050) );
  INVX1 INVX1_476 ( .A(core_v0_reg_43_), .Y(core__abc_21380_n2057) );
  INVX1 INVX1_477 ( .A(core_v1_reg_43_), .Y(core__abc_21380_n2058) );
  INVX1 INVX1_478 ( .A(core__abc_21380_n2059), .Y(core__abc_21380_n2060) );
  INVX1 INVX1_479 ( .A(core__abc_21380_n2061), .Y(core__abc_21380_n2062) );
  INVX1 INVX1_48 ( .A(_abc_19068_n2358), .Y(_abc_19068_n2359) );
  INVX1 INVX1_480 ( .A(core__abc_21380_n2065), .Y(core__abc_21380_n2066) );
  INVX1 INVX1_481 ( .A(core__abc_21380_n2063), .Y(core__abc_21380_n2069) );
  INVX1 INVX1_482 ( .A(core__abc_21380_n2067_1), .Y(core__abc_21380_n2070) );
  INVX1 INVX1_483 ( .A(core_v0_reg_44_), .Y(core__abc_21380_n2078) );
  INVX1 INVX1_484 ( .A(core_v1_reg_44_), .Y(core__abc_21380_n2079) );
  INVX1 INVX1_485 ( .A(core__abc_21380_n2083), .Y(core__abc_21380_n2084) );
  INVX1 INVX1_486 ( .A(core__abc_21380_n2081), .Y(core__abc_21380_n2087) );
  INVX1 INVX1_487 ( .A(core__abc_21380_n2085), .Y(core__abc_21380_n2088) );
  INVX1 INVX1_488 ( .A(core_v0_reg_45_), .Y(core__abc_21380_n2095) );
  INVX1 INVX1_489 ( .A(core_v1_reg_45_), .Y(core__abc_21380_n2096) );
  INVX1 INVX1_49 ( .A(_abc_19068_n2363), .Y(_abc_19068_n2364) );
  INVX1 INVX1_490 ( .A(core__abc_21380_n2097), .Y(core__abc_21380_n2098) );
  INVX1 INVX1_491 ( .A(core__abc_21380_n2099_1), .Y(core__abc_21380_n2100) );
  INVX1 INVX1_492 ( .A(core__abc_21380_n2103_1), .Y(core__abc_21380_n2104) );
  INVX1 INVX1_493 ( .A(core__abc_21380_n2101), .Y(core__abc_21380_n2107) );
  INVX1 INVX1_494 ( .A(core__abc_21380_n2105), .Y(core__abc_21380_n2108) );
  INVX1 INVX1_495 ( .A(core_v0_reg_46_), .Y(core__abc_21380_n2116) );
  INVX1 INVX1_496 ( .A(core_v1_reg_46_), .Y(core__abc_21380_n2117) );
  INVX1 INVX1_497 ( .A(core__abc_21380_n2121), .Y(core__abc_21380_n2122) );
  INVX1 INVX1_498 ( .A(core__abc_21380_n2119), .Y(core__abc_21380_n2125) );
  INVX1 INVX1_499 ( .A(core__abc_21380_n2123), .Y(core__abc_21380_n2126) );
  INVX1 INVX1_5 ( .A(\addr[4] ), .Y(_abc_19068_n878) );
  INVX1 INVX1_50 ( .A(_abc_19068_n2368), .Y(_abc_19068_n2369) );
  INVX1 INVX1_500 ( .A(core__abc_21380_n2133), .Y(core__abc_21380_n2134) );
  INVX1 INVX1_501 ( .A(core_v0_reg_47_), .Y(core__abc_21380_n2135) );
  INVX1 INVX1_502 ( .A(core_v1_reg_47_), .Y(core__abc_21380_n2136) );
  INVX1 INVX1_503 ( .A(core__abc_21380_n2137), .Y(core__abc_21380_n2138) );
  INVX1 INVX1_504 ( .A(core__abc_21380_n2139_1), .Y(core__abc_21380_n2140) );
  INVX1 INVX1_505 ( .A(core__abc_21380_n2142), .Y(core__abc_21380_n2143_1) );
  INVX1 INVX1_506 ( .A(core__abc_21380_n2144), .Y(core__abc_21380_n2146) );
  INVX1 INVX1_507 ( .A(core_v0_reg_48_), .Y(core__abc_21380_n2153) );
  INVX1 INVX1_508 ( .A(core_v1_reg_48_), .Y(core__abc_21380_n2154) );
  INVX1 INVX1_509 ( .A(core__abc_21380_n2157), .Y(core__abc_21380_n2158) );
  INVX1 INVX1_51 ( .A(_abc_19068_n2373), .Y(_abc_19068_n2374) );
  INVX1 INVX1_510 ( .A(core__abc_21380_n2160), .Y(core__abc_21380_n2161) );
  INVX1 INVX1_511 ( .A(core__abc_21380_n2162), .Y(core__abc_21380_n2164) );
  INVX1 INVX1_512 ( .A(core_v0_reg_49_), .Y(core__abc_21380_n2172) );
  INVX1 INVX1_513 ( .A(core_v1_reg_49_), .Y(core__abc_21380_n2173) );
  INVX1 INVX1_514 ( .A(core__abc_21380_n2177), .Y(core__abc_21380_n2178) );
  INVX1 INVX1_515 ( .A(core__abc_21380_n2175), .Y(core__abc_21380_n2181) );
  INVX1 INVX1_516 ( .A(core__abc_21380_n2179_1), .Y(core__abc_21380_n2182) );
  INVX1 INVX1_517 ( .A(core_v0_reg_50_), .Y(core__abc_21380_n2190) );
  INVX1 INVX1_518 ( .A(core_v1_reg_50_), .Y(core__abc_21380_n2191) );
  INVX1 INVX1_519 ( .A(core__abc_21380_n2195), .Y(core__abc_21380_n2196) );
  INVX1 INVX1_52 ( .A(_abc_19068_n2378), .Y(_abc_19068_n2379) );
  INVX1 INVX1_520 ( .A(core__abc_21380_n2193), .Y(core__abc_21380_n2199) );
  INVX1 INVX1_521 ( .A(core__abc_21380_n2197), .Y(core__abc_21380_n2200) );
  INVX1 INVX1_522 ( .A(core__abc_21380_n2207), .Y(core__abc_21380_n2208) );
  INVX1 INVX1_523 ( .A(core_v0_reg_51_), .Y(core__abc_21380_n2209) );
  INVX1 INVX1_524 ( .A(core_v1_reg_51_), .Y(core__abc_21380_n2210) );
  INVX1 INVX1_525 ( .A(core__abc_21380_n2211), .Y(core__abc_21380_n2212) );
  INVX1 INVX1_526 ( .A(core__abc_21380_n2213_1), .Y(core__abc_21380_n2214) );
  INVX1 INVX1_527 ( .A(core__abc_21380_n2216), .Y(core__abc_21380_n2217) );
  INVX1 INVX1_528 ( .A(core__abc_21380_n2218), .Y(core__abc_21380_n2220) );
  INVX1 INVX1_529 ( .A(core__abc_21380_n2228), .Y(core__abc_21380_n2229) );
  INVX1 INVX1_53 ( .A(_abc_19068_n2383), .Y(_abc_19068_n2384) );
  INVX1 INVX1_530 ( .A(core__abc_21380_n2232), .Y(core__abc_21380_n2233) );
  INVX1 INVX1_531 ( .A(core__abc_21380_n2230), .Y(core__abc_21380_n2236) );
  INVX1 INVX1_532 ( .A(core__abc_21380_n2234), .Y(core__abc_21380_n2237) );
  INVX1 INVX1_533 ( .A(core__abc_21380_n2244), .Y(core__abc_21380_n2245) );
  INVX1 INVX1_534 ( .A(core_v0_reg_53_), .Y(core__abc_21380_n2246) );
  INVX1 INVX1_535 ( .A(core_v1_reg_53_), .Y(core__abc_21380_n2247_1) );
  INVX1 INVX1_536 ( .A(core__abc_21380_n2248), .Y(core__abc_21380_n2249) );
  INVX1 INVX1_537 ( .A(core__abc_21380_n2250), .Y(core__abc_21380_n2251) );
  INVX1 INVX1_538 ( .A(core__abc_21380_n2253), .Y(core__abc_21380_n2254) );
  INVX1 INVX1_539 ( .A(core__abc_21380_n2255), .Y(core__abc_21380_n2257) );
  INVX1 INVX1_54 ( .A(_abc_19068_n2388), .Y(_abc_19068_n2389) );
  INVX1 INVX1_540 ( .A(core_v0_reg_54_), .Y(core__abc_21380_n2264) );
  INVX1 INVX1_541 ( .A(core_v1_reg_54_), .Y(core__abc_21380_n2265) );
  INVX1 INVX1_542 ( .A(core__abc_21380_n2268), .Y(core__abc_21380_n2269) );
  INVX1 INVX1_543 ( .A(core__abc_21380_n2271), .Y(core__abc_21380_n2272) );
  INVX1 INVX1_544 ( .A(core__abc_21380_n2273), .Y(core__abc_21380_n2275) );
  INVX1 INVX1_545 ( .A(core_v0_reg_55_), .Y(core__abc_21380_n2282) );
  INVX1 INVX1_546 ( .A(core_v1_reg_55_), .Y(core__abc_21380_n2283) );
  INVX1 INVX1_547 ( .A(core__abc_21380_n2284), .Y(core__abc_21380_n2285) );
  INVX1 INVX1_548 ( .A(core__abc_21380_n2286), .Y(core__abc_21380_n2287) );
  INVX1 INVX1_549 ( .A(core__abc_21380_n2290), .Y(core__abc_21380_n2291) );
  INVX1 INVX1_55 ( .A(_abc_19068_n2393), .Y(_abc_19068_n2394) );
  INVX1 INVX1_550 ( .A(core__abc_21380_n2288), .Y(core__abc_21380_n2294_1) );
  INVX1 INVX1_551 ( .A(core__abc_21380_n2292), .Y(core__abc_21380_n2295) );
  INVX1 INVX1_552 ( .A(core_v0_reg_56_), .Y(core__abc_21380_n2302) );
  INVX1 INVX1_553 ( .A(core_v1_reg_56_), .Y(core__abc_21380_n2303) );
  INVX1 INVX1_554 ( .A(core__abc_21380_n2306), .Y(core__abc_21380_n2307) );
  INVX1 INVX1_555 ( .A(core__abc_21380_n2309), .Y(core__abc_21380_n2310) );
  INVX1 INVX1_556 ( .A(core__abc_21380_n2311), .Y(core__abc_21380_n2313) );
  INVX1 INVX1_557 ( .A(core_v0_reg_57_), .Y(core__abc_21380_n2320) );
  INVX1 INVX1_558 ( .A(core_v1_reg_57_), .Y(core__abc_21380_n2321) );
  INVX1 INVX1_559 ( .A(core__abc_21380_n2324), .Y(core__abc_21380_n2325) );
  INVX1 INVX1_56 ( .A(_abc_19068_n2398), .Y(_abc_19068_n2399) );
  INVX1 INVX1_560 ( .A(core__abc_21380_n2327), .Y(core__abc_21380_n2328_1) );
  INVX1 INVX1_561 ( .A(core__abc_21380_n2329), .Y(core__abc_21380_n2331) );
  INVX1 INVX1_562 ( .A(core_v0_reg_58_), .Y(core__abc_21380_n2338) );
  INVX1 INVX1_563 ( .A(core_v1_reg_58_), .Y(core__abc_21380_n2339) );
  INVX1 INVX1_564 ( .A(core__abc_21380_n2342), .Y(core__abc_21380_n2343) );
  INVX1 INVX1_565 ( .A(core__abc_21380_n2345), .Y(core__abc_21380_n2346) );
  INVX1 INVX1_566 ( .A(core__abc_21380_n2347), .Y(core__abc_21380_n2349) );
  INVX1 INVX1_567 ( .A(core_v0_reg_59_), .Y(core__abc_21380_n2356) );
  INVX1 INVX1_568 ( .A(core_v1_reg_59_), .Y(core__abc_21380_n2357) );
  INVX1 INVX1_569 ( .A(core__abc_21380_n2358), .Y(core__abc_21380_n2359) );
  INVX1 INVX1_57 ( .A(_abc_19068_n2403), .Y(_abc_19068_n2404) );
  INVX1 INVX1_570 ( .A(core__abc_21380_n2360), .Y(core__abc_21380_n2361) );
  INVX1 INVX1_571 ( .A(core__abc_21380_n2364), .Y(core__abc_21380_n2365) );
  INVX1 INVX1_572 ( .A(core__abc_21380_n2362), .Y(core__abc_21380_n2368) );
  INVX1 INVX1_573 ( .A(core__abc_21380_n2366), .Y(core__abc_21380_n2369_1) );
  INVX1 INVX1_574 ( .A(core_v0_reg_60_), .Y(core__abc_21380_n2376) );
  INVX1 INVX1_575 ( .A(core_v1_reg_60_), .Y(core__abc_21380_n2377) );
  INVX1 INVX1_576 ( .A(core__abc_21380_n2380), .Y(core__abc_21380_n2381) );
  INVX1 INVX1_577 ( .A(core__abc_21380_n2383), .Y(core__abc_21380_n2384) );
  INVX1 INVX1_578 ( .A(core__abc_21380_n2385), .Y(core__abc_21380_n2387) );
  INVX1 INVX1_579 ( .A(core_v0_reg_61_), .Y(core__abc_21380_n2394) );
  INVX1 INVX1_58 ( .A(_abc_19068_n2408), .Y(_abc_19068_n2409) );
  INVX1 INVX1_580 ( .A(core_v1_reg_61_), .Y(core__abc_21380_n2395_1) );
  INVX1 INVX1_581 ( .A(core__abc_21380_n2398), .Y(core__abc_21380_n2399) );
  INVX1 INVX1_582 ( .A(core__abc_21380_n2401), .Y(core__abc_21380_n2402) );
  INVX1 INVX1_583 ( .A(core__abc_21380_n2403), .Y(core__abc_21380_n2405) );
  INVX1 INVX1_584 ( .A(core_v0_reg_62_), .Y(core__abc_21380_n2412) );
  INVX1 INVX1_585 ( .A(core_v1_reg_62_), .Y(core__abc_21380_n2413) );
  INVX1 INVX1_586 ( .A(core__abc_21380_n2416), .Y(core__abc_21380_n2417) );
  INVX1 INVX1_587 ( .A(core__abc_21380_n2419), .Y(core__abc_21380_n2420) );
  INVX1 INVX1_588 ( .A(core__abc_21380_n2421), .Y(core__abc_21380_n2423) );
  INVX1 INVX1_589 ( .A(core_v0_reg_63_), .Y(core__abc_21380_n2430_1) );
  INVX1 INVX1_59 ( .A(_abc_19068_n2413), .Y(_abc_19068_n2414) );
  INVX1 INVX1_590 ( .A(core_v1_reg_63_), .Y(core__abc_21380_n2432) );
  INVX1 INVX1_591 ( .A(core__abc_21380_n2434), .Y(core__abc_21380_n2435) );
  INVX1 INVX1_592 ( .A(core__abc_21380_n2437), .Y(core__abc_21380_n2438) );
  INVX1 INVX1_593 ( .A(core__abc_21380_n2439), .Y(core__abc_21380_n2440) );
  INVX1 INVX1_594 ( .A(core_siphash_ctrl_reg_0_), .Y(core__abc_21380_n2449) );
  INVX1 INVX1_595 ( .A(core__abc_21380_n1146_1), .Y(core__abc_21380_n2709) );
  INVX1 INVX1_596 ( .A(core__abc_21380_n2710), .Y(core__abc_21380_n2711) );
  INVX1 INVX1_597 ( .A(core__abc_21380_n1147), .Y(core__abc_21380_n2715) );
  INVX1 INVX1_598 ( .A(core__abc_21380_n2716), .Y(core__abc_21380_n2717) );
  INVX1 INVX1_599 ( .A(core__abc_21380_n2725), .Y(core__abc_21380_n2726) );
  INVX1 INVX1_6 ( .A(\addr[5] ), .Y(_abc_19068_n879_1) );
  INVX1 INVX1_60 ( .A(_abc_19068_n2418), .Y(_abc_19068_n2419) );
  INVX1 INVX1_600 ( .A(core__abc_21380_n2733), .Y(core__abc_21380_n2734) );
  INVX1 INVX1_601 ( .A(core_v3_reg_27_), .Y(core__abc_21380_n3007) );
  INVX1 INVX1_602 ( .A(core__abc_21380_n3009), .Y(core__abc_21380_n3010) );
  INVX1 INVX1_603 ( .A(core__abc_21380_n3020), .Y(core__abc_21380_n3021) );
  INVX1 INVX1_604 ( .A(core__abc_21380_n3022), .Y(core__abc_21380_n3023) );
  INVX1 INVX1_605 ( .A(core__abc_21380_n3024_1), .Y(core__abc_21380_n3025) );
  INVX1 INVX1_606 ( .A(core__abc_21380_n3029), .Y(core__abc_21380_n3030_1) );
  INVX1 INVX1_607 ( .A(core__abc_21380_n3039), .Y(core__abc_21380_n3040_1) );
  INVX1 INVX1_608 ( .A(core__abc_21380_n1437), .Y(core__abc_21380_n3042) );
  INVX1 INVX1_609 ( .A(core__abc_21380_n3044_1), .Y(core__abc_21380_n3045) );
  INVX1 INVX1_61 ( .A(_abc_19068_n2423), .Y(_abc_19068_n2424) );
  INVX1 INVX1_610 ( .A(core__abc_21380_n3052), .Y(core__abc_21380_n3053) );
  INVX1 INVX1_611 ( .A(core__abc_21380_n3058), .Y(core__abc_21380_n3059) );
  INVX1 INVX1_612 ( .A(core__abc_21380_n3075), .Y(core__abc_21380_n3076) );
  INVX1 INVX1_613 ( .A(core__abc_21380_n1583), .Y(core__abc_21380_n3078) );
  INVX1 INVX1_614 ( .A(core__abc_21380_n3080), .Y(core__abc_21380_n3081) );
  INVX1 INVX1_615 ( .A(core__abc_21380_n3088), .Y(core__abc_21380_n3089) );
  INVX1 INVX1_616 ( .A(core__abc_21380_n3097), .Y(core__abc_21380_n3098) );
  INVX1 INVX1_617 ( .A(core__abc_21380_n1804), .Y(core__abc_21380_n3106) );
  INVX1 INVX1_618 ( .A(core__abc_21380_n3108), .Y(core__abc_21380_n3109) );
  INVX1 INVX1_619 ( .A(core__abc_21380_n3113), .Y(core__abc_21380_n3114) );
  INVX1 INVX1_62 ( .A(_abc_19068_n2428), .Y(_abc_19068_n2429) );
  INVX1 INVX1_620 ( .A(core__abc_21380_n3122_1), .Y(core__abc_21380_n3123) );
  INVX1 INVX1_621 ( .A(core__abc_21380_n1879), .Y(core__abc_21380_n3125) );
  INVX1 INVX1_622 ( .A(core__abc_21380_n3127), .Y(core__abc_21380_n3128_1) );
  INVX1 INVX1_623 ( .A(core__abc_21380_n3135), .Y(core__abc_21380_n3136) );
  INVX1 INVX1_624 ( .A(core__abc_21380_n3141_1), .Y(core__abc_21380_n3142) );
  INVX1 INVX1_625 ( .A(core__abc_21380_n3143), .Y(core__abc_21380_n3144) );
  INVX1 INVX1_626 ( .A(core__abc_21380_n3148), .Y(core__abc_21380_n3149) );
  INVX1 INVX1_627 ( .A(core__abc_21380_n3151), .Y(core__abc_21380_n3152) );
  INVX1 INVX1_628 ( .A(core__abc_21380_n3153), .Y(core__abc_21380_n3156) );
  INVX1 INVX1_629 ( .A(core__abc_21380_n3160), .Y(core__abc_21380_n3161) );
  INVX1 INVX1_63 ( .A(_abc_19068_n2433), .Y(_abc_19068_n2434) );
  INVX1 INVX1_630 ( .A(core__abc_21380_n3163_1_bF_buf6), .Y(core__abc_21380_n3164) );
  INVX1 INVX1_631 ( .A(core__abc_21380_n3170), .Y(core__abc_21380_n3171) );
  INVX1 INVX1_632 ( .A(core__abc_21380_n1320), .Y(core__abc_21380_n3173) );
  INVX1 INVX1_633 ( .A(core__abc_21380_n1357), .Y(core__abc_21380_n3181_1) );
  INVX1 INVX1_634 ( .A(core__abc_21380_n1394), .Y(core__abc_21380_n3185) );
  INVX1 INVX1_635 ( .A(core__abc_21380_n3191), .Y(core__abc_21380_n3192) );
  INVX1 INVX1_636 ( .A(core__abc_21380_n3206), .Y(core__abc_21380_n3207) );
  INVX1 INVX1_637 ( .A(core__abc_21380_n3208), .Y(core__abc_21380_n3209) );
  INVX1 INVX1_638 ( .A(core__abc_21380_n3224), .Y(core__abc_21380_n3225) );
  INVX1 INVX1_639 ( .A(core__abc_21380_n3240), .Y(core__abc_21380_n3241) );
  INVX1 INVX1_64 ( .A(_abc_19068_n2438), .Y(_abc_19068_n2439) );
  INVX1 INVX1_640 ( .A(core__abc_21380_n3242), .Y(core__abc_21380_n3243) );
  INVX1 INVX1_641 ( .A(core__abc_21380_n1705), .Y(core__abc_21380_n3250) );
  INVX1 INVX1_642 ( .A(core__abc_21380_n3252), .Y(core__abc_21380_n3253) );
  INVX1 INVX1_643 ( .A(core__abc_21380_n1780), .Y(core__abc_21380_n3261) );
  INVX1 INVX1_644 ( .A(core__abc_21380_n3263), .Y(core__abc_21380_n3264) );
  INVX1 INVX1_645 ( .A(core__abc_21380_n3175), .Y(core__abc_21380_n3274) );
  INVX1 INVX1_646 ( .A(core__abc_21380_n3179), .Y(core__abc_21380_n3276) );
  INVX1 INVX1_647 ( .A(core__abc_21380_n3188), .Y(core__abc_21380_n3278) );
  INVX1 INVX1_648 ( .A(core__abc_21380_n3197), .Y(core__abc_21380_n3280) );
  INVX1 INVX1_649 ( .A(core__abc_21380_n3214), .Y(core__abc_21380_n3282) );
  INVX1 INVX1_65 ( .A(_abc_19068_n2443), .Y(_abc_19068_n2444) );
  INVX1 INVX1_650 ( .A(core__abc_21380_n3231), .Y(core__abc_21380_n3284) );
  INVX1 INVX1_651 ( .A(core__abc_21380_n3268_1), .Y(core__abc_21380_n3286) );
  INVX1 INVX1_652 ( .A(core__abc_21380_n3289), .Y(core__abc_21380_n3290) );
  INVX1 INVX1_653 ( .A(core__abc_21380_n3291), .Y(core__abc_21380_n3292) );
  INVX1 INVX1_654 ( .A(core__abc_21380_n3294), .Y(core__abc_21380_n3295) );
  INVX1 INVX1_655 ( .A(core__abc_21380_n3298), .Y(core__abc_21380_n3304) );
  INVX1 INVX1_656 ( .A(core__abc_21380_n3314), .Y(core__abc_21380_n3315) );
  INVX1 INVX1_657 ( .A(core_key_64_), .Y(core__abc_21380_n3318) );
  INVX1 INVX1_658 ( .A(core__abc_21380_n3321), .Y(core__abc_21380_n3322) );
  INVX1 INVX1_659 ( .A(core__abc_21380_n3332), .Y(core__abc_21380_n3333) );
  INVX1 INVX1_66 ( .A(_abc_19068_n2448), .Y(_abc_19068_n2449) );
  INVX1 INVX1_660 ( .A(core__abc_21380_n3337), .Y(core__abc_21380_n3338) );
  INVX1 INVX1_661 ( .A(core_v3_reg_49_), .Y(core__abc_21380_n3341) );
  INVX1 INVX1_662 ( .A(core__abc_21380_n1266_1), .Y(core__abc_21380_n3342) );
  INVX1 INVX1_663 ( .A(core__abc_21380_n3344), .Y(core__abc_21380_n3345) );
  INVX1 INVX1_664 ( .A(core__abc_21380_n3348), .Y(core__abc_21380_n3349) );
  INVX1 INVX1_665 ( .A(core__abc_21380_n3350), .Y(core__abc_21380_n3351) );
  INVX1 INVX1_666 ( .A(core__abc_21380_n3296), .Y(core__abc_21380_n3355) );
  INVX1 INVX1_667 ( .A(core__abc_21380_n3335), .Y(core__abc_21380_n3356) );
  INVX1 INVX1_668 ( .A(core__abc_21380_n3363), .Y(core__abc_21380_n3364) );
  INVX1 INVX1_669 ( .A(core_v3_reg_28_), .Y(core__abc_21380_n3365) );
  INVX1 INVX1_67 ( .A(_abc_19068_n2453), .Y(_abc_19068_n2454) );
  INVX1 INVX1_670 ( .A(core__abc_21380_n3370), .Y(core__abc_21380_n3371) );
  INVX1 INVX1_671 ( .A(core__abc_21380_n3372), .Y(core__abc_21380_n3373) );
  INVX1 INVX1_672 ( .A(core__abc_21380_n3375), .Y(core__abc_21380_n3376) );
  INVX1 INVX1_673 ( .A(core__abc_21380_n3379), .Y(core__abc_21380_n3380) );
  INVX1 INVX1_674 ( .A(core__abc_21380_n3383), .Y(core__abc_21380_n3384) );
  INVX1 INVX1_675 ( .A(core_key_65_), .Y(core__abc_21380_n3389) );
  INVX1 INVX1_676 ( .A(core__abc_21380_n3392), .Y(core__abc_21380_n3393) );
  INVX1 INVX1_677 ( .A(core__abc_21380_n3405), .Y(core__abc_21380_n3406) );
  INVX1 INVX1_678 ( .A(core__abc_21380_n3409), .Y(core__abc_21380_n3410) );
  INVX1 INVX1_679 ( .A(core_v3_reg_50_), .Y(core__abc_21380_n3411) );
  INVX1 INVX1_68 ( .A(_abc_19068_n2458), .Y(_abc_19068_n2459) );
  INVX1 INVX1_680 ( .A(core__abc_21380_n3014), .Y(core__abc_21380_n3413) );
  INVX1 INVX1_681 ( .A(core__abc_21380_n3415), .Y(core__abc_21380_n3416) );
  INVX1 INVX1_682 ( .A(core__abc_21380_n3419), .Y(core__abc_21380_n3420) );
  INVX1 INVX1_683 ( .A(core__abc_21380_n3423), .Y(core__abc_21380_n3426) );
  INVX1 INVX1_684 ( .A(core_v3_reg_29_), .Y(core__abc_21380_n3429) );
  INVX1 INVX1_685 ( .A(core__abc_21380_n3430), .Y(core__abc_21380_n3431) );
  INVX1 INVX1_686 ( .A(core__abc_21380_n3434), .Y(core__abc_21380_n3436) );
  INVX1 INVX1_687 ( .A(core__abc_21380_n3428), .Y(core__abc_21380_n3440) );
  INVX1 INVX1_688 ( .A(core__abc_21380_n3435), .Y(core__abc_21380_n3441) );
  INVX1 INVX1_689 ( .A(core__abc_21380_n3449), .Y(core__abc_21380_n3450) );
  INVX1 INVX1_69 ( .A(_abc_19068_n2463), .Y(_abc_19068_n2464) );
  INVX1 INVX1_690 ( .A(core__abc_21380_n3459), .Y(core__abc_21380_n3460) );
  INVX1 INVX1_691 ( .A(core__abc_21380_n1304), .Y(core__abc_21380_n3464) );
  INVX1 INVX1_692 ( .A(core__abc_21380_n3412), .Y(core__abc_21380_n3465) );
  INVX1 INVX1_693 ( .A(core__abc_21380_n3466), .Y(core__abc_21380_n3467) );
  INVX1 INVX1_694 ( .A(core__abc_21380_n3470), .Y(core__abc_21380_n3471) );
  INVX1 INVX1_695 ( .A(core_v3_reg_51_), .Y(core__abc_21380_n3473) );
  INVX1 INVX1_696 ( .A(core__abc_21380_n3463), .Y(core__abc_21380_n3477) );
  INVX1 INVX1_697 ( .A(core__abc_21380_n3475), .Y(core__abc_21380_n3478) );
  INVX1 INVX1_698 ( .A(core__abc_21380_n3480), .Y(core__abc_21380_n3481) );
  INVX1 INVX1_699 ( .A(core__abc_21380_n3421), .Y(core__abc_21380_n3482) );
  INVX1 INVX1_7 ( .A(\addr[0] ), .Y(_abc_19068_n886_1) );
  INVX1 INVX1_70 ( .A(_abc_19068_n2468), .Y(_abc_19068_n2469) );
  INVX1 INVX1_700 ( .A(core__abc_21380_n3486), .Y(core__abc_21380_n3487) );
  INVX1 INVX1_701 ( .A(core__abc_21380_n3488), .Y(core__abc_21380_n3489) );
  INVX1 INVX1_702 ( .A(core__abc_21380_n3490_1), .Y(core__abc_21380_n3491) );
  INVX1 INVX1_703 ( .A(core__abc_21380_n2102), .Y(core__abc_21380_n3493) );
  INVX1 INVX1_704 ( .A(core__abc_21380_n3496), .Y(core__abc_21380_n3498) );
  INVX1 INVX1_705 ( .A(core__abc_21380_n3500), .Y(core__abc_21380_n3501_1) );
  INVX1 INVX1_706 ( .A(core_v3_reg_30_), .Y(core__abc_21380_n3503) );
  INVX1 INVX1_707 ( .A(core__abc_21380_n3505_1), .Y(core__abc_21380_n3507) );
  INVX1 INVX1_708 ( .A(core__abc_21380_n3513), .Y(core__abc_21380_n3514) );
  INVX1 INVX1_709 ( .A(core__abc_21380_n3527), .Y(core__abc_21380_n3532) );
  INVX1 INVX1_71 ( .A(_abc_19068_n2473), .Y(_abc_19068_n2474) );
  INVX1 INVX1_710 ( .A(core__abc_21380_n3528), .Y(core__abc_21380_n3533) );
  INVX1 INVX1_711 ( .A(core__abc_21380_n3537), .Y(core__abc_21380_n3538) );
  INVX1 INVX1_712 ( .A(core_v3_reg_52_), .Y(core__abc_21380_n3539) );
  INVX1 INVX1_713 ( .A(core__abc_21380_n3017), .Y(core__abc_21380_n3541) );
  INVX1 INVX1_714 ( .A(core__abc_21380_n3543), .Y(core__abc_21380_n3545) );
  INVX1 INVX1_715 ( .A(core__abc_21380_n3547), .Y(core__abc_21380_n3548_1) );
  INVX1 INVX1_716 ( .A(core__abc_21380_n3551), .Y(core__abc_21380_n3552_1) );
  INVX1 INVX1_717 ( .A(core__abc_21380_n3553), .Y(core__abc_21380_n3554) );
  INVX1 INVX1_718 ( .A(core__abc_21380_n3479), .Y(core__abc_21380_n3558) );
  INVX1 INVX1_719 ( .A(core__abc_21380_n3562), .Y(core__abc_21380_n3563) );
  INVX1 INVX1_72 ( .A(_abc_19068_n2478), .Y(_abc_19068_n2479) );
  INVX1 INVX1_720 ( .A(core__abc_21380_n3565), .Y(core__abc_21380_n3567) );
  INVX1 INVX1_721 ( .A(core_v3_reg_31_), .Y(core__abc_21380_n3571) );
  INVX1 INVX1_722 ( .A(core__abc_21380_n3566), .Y(core__abc_21380_n3572) );
  INVX1 INVX1_723 ( .A(core_key_68_), .Y(core__abc_21380_n3584) );
  INVX1 INVX1_724 ( .A(core__abc_21380_n3587), .Y(core__abc_21380_n3588) );
  INVX1 INVX1_725 ( .A(core__abc_21380_n3597), .Y(core__abc_21380_n3598) );
  INVX1 INVX1_726 ( .A(core__abc_21380_n3599), .Y(core__abc_21380_n3600_1) );
  INVX1 INVX1_727 ( .A(core__abc_21380_n3603), .Y(core__abc_21380_n3604_1) );
  INVX1 INVX1_728 ( .A(core_v3_reg_53_), .Y(core__abc_21380_n3605) );
  INVX1 INVX1_729 ( .A(core__abc_21380_n3606), .Y(core__abc_21380_n3607) );
  INVX1 INVX1_73 ( .A(_abc_19068_n2483), .Y(_abc_19068_n2484) );
  INVX1 INVX1_730 ( .A(core__abc_21380_n3610), .Y(core__abc_21380_n3612) );
  INVX1 INVX1_731 ( .A(core__abc_21380_n3614), .Y(core__abc_21380_n3615) );
  INVX1 INVX1_732 ( .A(core__abc_21380_n3618), .Y(core__abc_21380_n3620) );
  INVX1 INVX1_733 ( .A(core__abc_21380_n3622), .Y(core__abc_21380_n3623_1) );
  INVX1 INVX1_734 ( .A(core_v3_reg_32_), .Y(core__abc_21380_n3624) );
  INVX1 INVX1_735 ( .A(core__abc_21380_n3495), .Y(core__abc_21380_n3628) );
  INVX1 INVX1_736 ( .A(core__abc_21380_n3633), .Y(core__abc_21380_n3638) );
  INVX1 INVX1_737 ( .A(core__abc_21380_n3626), .Y(core__abc_21380_n3639) );
  INVX1 INVX1_738 ( .A(core__abc_21380_n3643), .Y(core__abc_21380_n3644) );
  INVX1 INVX1_739 ( .A(core__abc_21380_n3647_1), .Y(core__abc_21380_n3648) );
  INVX1 INVX1_74 ( .A(_abc_19068_n2489), .Y(_abc_19068_n2490) );
  INVX1 INVX1_740 ( .A(core_key_69_), .Y(core__abc_21380_n3653) );
  INVX1 INVX1_741 ( .A(core__abc_21380_n3656), .Y(core__abc_21380_n3657) );
  INVX1 INVX1_742 ( .A(core__abc_21380_n3617), .Y(core__abc_21380_n3668) );
  INVX1 INVX1_743 ( .A(core__abc_21380_n3670), .Y(core__abc_21380_n3671) );
  INVX1 INVX1_744 ( .A(core__abc_21380_n3672), .Y(core__abc_21380_n3673) );
  INVX1 INVX1_745 ( .A(core__abc_21380_n3674), .Y(core__abc_21380_n3675) );
  INVX1 INVX1_746 ( .A(core__abc_21380_n1927), .Y(core__abc_21380_n3677) );
  INVX1 INVX1_747 ( .A(core__abc_21380_n3679), .Y(core__abc_21380_n3683) );
  INVX1 INVX1_748 ( .A(core_v3_reg_54_), .Y(core__abc_21380_n3687) );
  INVX1 INVX1_749 ( .A(core__abc_21380_n3691), .Y(core__abc_21380_n3692) );
  INVX1 INVX1_75 ( .A(_abc_19068_n2494), .Y(_abc_19068_n2495) );
  INVX1 INVX1_750 ( .A(core__abc_21380_n3693_1), .Y(core__abc_21380_n3694) );
  INVX1 INVX1_751 ( .A(core__abc_21380_n3698), .Y(core__abc_21380_n3699) );
  INVX1 INVX1_752 ( .A(core__abc_21380_n3701), .Y(core__abc_21380_n3702) );
  INVX1 INVX1_753 ( .A(core__abc_21380_n3705), .Y(core__abc_21380_n3706) );
  INVX1 INVX1_754 ( .A(core_v3_reg_33_), .Y(core__abc_21380_n3707) );
  INVX1 INVX1_755 ( .A(core__abc_21380_n3637), .Y(core__abc_21380_n3708_1) );
  INVX1 INVX1_756 ( .A(core__abc_21380_n3715), .Y(core__abc_21380_n3717) );
  INVX1 INVX1_757 ( .A(core__abc_21380_n3719), .Y(core__abc_21380_n3720_1) );
  INVX1 INVX1_758 ( .A(core_key_70_), .Y(core__abc_21380_n3725) );
  INVX1 INVX1_759 ( .A(core__abc_21380_n3728), .Y(core__abc_21380_n3729) );
  INVX1 INVX1_76 ( .A(_abc_19068_n2499), .Y(_abc_19068_n2500) );
  INVX1 INVX1_760 ( .A(core__abc_21380_n3738), .Y(core__abc_21380_n3739) );
  INVX1 INVX1_761 ( .A(core__abc_21380_n1968), .Y(core__abc_21380_n3740_1) );
  INVX1 INVX1_762 ( .A(core_v3_reg_55_), .Y(core__abc_21380_n3747) );
  INVX1 INVX1_763 ( .A(core__abc_21380_n3748), .Y(core__abc_21380_n3749) );
  INVX1 INVX1_764 ( .A(core__abc_21380_n3752_1), .Y(core__abc_21380_n3754) );
  INVX1 INVX1_765 ( .A(core__abc_21380_n3756_1), .Y(core__abc_21380_n3761) );
  INVX1 INVX1_766 ( .A(core__abc_21380_n3763), .Y(core__abc_21380_n3764) );
  INVX1 INVX1_767 ( .A(core__abc_21380_n3767_1), .Y(core__abc_21380_n3768) );
  INVX1 INVX1_768 ( .A(core_v3_reg_34_), .Y(core__abc_21380_n3769) );
  INVX1 INVX1_769 ( .A(core__abc_21380_n3772_1), .Y(core__abc_21380_n3773) );
  INVX1 INVX1_77 ( .A(_abc_19068_n2504), .Y(_abc_19068_n2505) );
  INVX1 INVX1_770 ( .A(core__abc_21380_n3775), .Y(core__abc_21380_n3777) );
  INVX1 INVX1_771 ( .A(core__abc_21380_n3779_1), .Y(core__abc_21380_n3780) );
  INVX1 INVX1_772 ( .A(core__abc_21380_n3787), .Y(core__abc_21380_n3788) );
  INVX1 INVX1_773 ( .A(core__abc_21380_n3804), .Y(core__abc_21380_n3809_1) );
  INVX1 INVX1_774 ( .A(core__abc_21380_n3805), .Y(core__abc_21380_n3810) );
  INVX1 INVX1_775 ( .A(core__abc_21380_n3814_1), .Y(core__abc_21380_n3815) );
  INVX1 INVX1_776 ( .A(core_v3_reg_56_), .Y(core__abc_21380_n3816) );
  INVX1 INVX1_777 ( .A(core__abc_21380_n3032), .Y(core__abc_21380_n3818) );
  INVX1 INVX1_778 ( .A(core__abc_21380_n3820), .Y(core__abc_21380_n3821) );
  INVX1 INVX1_779 ( .A(core__abc_21380_n3824), .Y(core__abc_21380_n3825) );
  INVX1 INVX1_78 ( .A(_abc_19068_n2509), .Y(_abc_19068_n2510) );
  INVX1 INVX1_780 ( .A(core__abc_21380_n3828_1), .Y(core__abc_21380_n3838_1) );
  INVX1 INVX1_781 ( .A(core__abc_21380_n3831), .Y(core__abc_21380_n3839) );
  INVX1 INVX1_782 ( .A(core__abc_21380_n3666), .Y(core__abc_21380_n3843) );
  INVX1 INVX1_783 ( .A(core__abc_21380_n3848), .Y(core__abc_21380_n3849) );
  INVX1 INVX1_784 ( .A(core_v3_reg_35_), .Y(core__abc_21380_n3850) );
  INVX1 INVX1_785 ( .A(core__abc_21380_n3852), .Y(core__abc_21380_n3853_1) );
  INVX1 INVX1_786 ( .A(core__abc_21380_n3856), .Y(core__abc_21380_n3857_1) );
  INVX1 INVX1_787 ( .A(core__abc_21380_n3858), .Y(core__abc_21380_n3861) );
  INVX1 INVX1_788 ( .A(core_key_72_), .Y(core__abc_21380_n3866) );
  INVX1 INVX1_789 ( .A(core__abc_21380_n3869_1), .Y(core__abc_21380_n3870) );
  INVX1 INVX1_79 ( .A(_abc_19068_n2514), .Y(_abc_19068_n2515) );
  INVX1 INVX1_790 ( .A(core__abc_21380_n3826), .Y(core__abc_21380_n3879) );
  INVX1 INVX1_791 ( .A(core__abc_21380_n3847), .Y(core__abc_21380_n3880) );
  INVX1 INVX1_792 ( .A(core__abc_21380_n3881_1), .Y(core__abc_21380_n3882) );
  INVX1 INVX1_793 ( .A(core__abc_21380_n3884), .Y(core__abc_21380_n3885) );
  INVX1 INVX1_794 ( .A(core_v3_reg_57_), .Y(core__abc_21380_n3891) );
  INVX1 INVX1_795 ( .A(core__abc_21380_n3892), .Y(core__abc_21380_n3893_1) );
  INVX1 INVX1_796 ( .A(core__abc_21380_n3896), .Y(core__abc_21380_n3898_1) );
  INVX1 INVX1_797 ( .A(core__abc_21380_n3902), .Y(core__abc_21380_n3903) );
  INVX1 INVX1_798 ( .A(core__abc_21380_n3904), .Y(core__abc_21380_n3905) );
  INVX1 INVX1_799 ( .A(core_v3_reg_36_), .Y(core__abc_21380_n3909) );
  INVX1 INVX1_8 ( .A(\addr[3] ), .Y(_abc_19068_n892_1) );
  INVX1 INVX1_80 ( .A(_abc_19068_n2519), .Y(_abc_19068_n2520) );
  INVX1 INVX1_800 ( .A(core__abc_21380_n3911), .Y(core__abc_21380_n3912) );
  INVX1 INVX1_801 ( .A(core__abc_21380_n3917), .Y(core__abc_21380_n3918) );
  INVX1 INVX1_802 ( .A(core__abc_21380_n3919), .Y(core__abc_21380_n3920) );
  INVX1 INVX1_803 ( .A(core__abc_21380_n3923), .Y(core__abc_21380_n3924) );
  INVX1 INVX1_804 ( .A(core__abc_21380_n3927_1), .Y(core__abc_21380_n3928) );
  INVX1 INVX1_805 ( .A(core__abc_21380_n3908), .Y(core__abc_21380_n3930) );
  INVX1 INVX1_806 ( .A(core__abc_21380_n3936), .Y(core__abc_21380_n3937_1) );
  INVX1 INVX1_807 ( .A(core__abc_21380_n3947), .Y(core__abc_21380_n3949) );
  INVX1 INVX1_808 ( .A(core__abc_21380_n3951), .Y(core__abc_21380_n3952_1) );
  INVX1 INVX1_809 ( .A(core_v3_reg_58_), .Y(core__abc_21380_n3953) );
  INVX1 INVX1_81 ( .A(_abc_19068_n2524), .Y(_abc_19068_n2525) );
  INVX1 INVX1_810 ( .A(core__abc_21380_n3954), .Y(core__abc_21380_n3955_1) );
  INVX1 INVX1_811 ( .A(core__abc_21380_n3958), .Y(core__abc_21380_n3959) );
  INVX1 INVX1_812 ( .A(core__abc_21380_n3960), .Y(core__abc_21380_n3961_1) );
  INVX1 INVX1_813 ( .A(core__abc_21380_n3964), .Y(core__abc_21380_n3965_1) );
  INVX1 INVX1_814 ( .A(core__abc_21380_n3968), .Y(core__abc_21380_n3969_1) );
  INVX1 INVX1_815 ( .A(core__abc_21380_n3972), .Y(core__abc_21380_n3973) );
  INVX1 INVX1_816 ( .A(core__abc_21380_n3976), .Y(core__abc_21380_n3977) );
  INVX1 INVX1_817 ( .A(core_v3_reg_37_), .Y(core__abc_21380_n3978) );
  INVX1 INVX1_818 ( .A(core__abc_21380_n3979_1), .Y(core__abc_21380_n3980) );
  INVX1 INVX1_819 ( .A(core__abc_21380_n3983), .Y(core__abc_21380_n3985) );
  INVX1 INVX1_82 ( .A(_abc_19068_n2529), .Y(_abc_19068_n2530) );
  INVX1 INVX1_820 ( .A(core__abc_21380_n3987), .Y(core__abc_21380_n3988_1) );
  INVX1 INVX1_821 ( .A(core_key_74_), .Y(core__abc_21380_n3993) );
  INVX1 INVX1_822 ( .A(core__abc_21380_n3996), .Y(core__abc_21380_n3997) );
  INVX1 INVX1_823 ( .A(core__abc_21380_n4007), .Y(core__abc_21380_n4008_1) );
  INVX1 INVX1_824 ( .A(core_v3_reg_59_), .Y(core__abc_21380_n4012_1) );
  INVX1 INVX1_825 ( .A(core__abc_21380_n4014), .Y(core__abc_21380_n4015) );
  INVX1 INVX1_826 ( .A(core__abc_21380_n4017), .Y(core__abc_21380_n4018_1) );
  INVX1 INVX1_827 ( .A(core__abc_21380_n4023_1), .Y(core__abc_21380_n4024) );
  INVX1 INVX1_828 ( .A(core__abc_21380_n4026_1), .Y(core__abc_21380_n4027) );
  INVX1 INVX1_829 ( .A(core__abc_21380_n4029), .Y(core__abc_21380_n4030) );
  INVX1 INVX1_83 ( .A(_abc_19068_n2534), .Y(_abc_19068_n2535) );
  INVX1 INVX1_830 ( .A(core__abc_21380_n4031_1), .Y(core__abc_21380_n4032) );
  INVX1 INVX1_831 ( .A(core__abc_21380_n2252), .Y(core__abc_21380_n4034_1) );
  INVX1 INVX1_832 ( .A(core__abc_21380_n4037), .Y(core__abc_21380_n4038) );
  INVX1 INVX1_833 ( .A(core__abc_21380_n4041), .Y(core__abc_21380_n4042) );
  INVX1 INVX1_834 ( .A(core_v3_reg_38_), .Y(core__abc_21380_n4044) );
  INVX1 INVX1_835 ( .A(core__abc_21380_n4046), .Y(core__abc_21380_n4047_1) );
  INVX1 INVX1_836 ( .A(core__abc_21380_n4054_1), .Y(core__abc_21380_n4055) );
  INVX1 INVX1_837 ( .A(core__abc_21380_n4066), .Y(core__abc_21380_n4067_1) );
  INVX1 INVX1_838 ( .A(core__abc_21380_n4009), .Y(core__abc_21380_n4070) );
  INVX1 INVX1_839 ( .A(core__abc_21380_n4010), .Y(core__abc_21380_n4071) );
  INVX1 INVX1_84 ( .A(_abc_19068_n2539), .Y(_abc_19068_n2540) );
  INVX1 INVX1_840 ( .A(core__abc_21380_n4021), .Y(core__abc_21380_n4073) );
  INVX1 INVX1_841 ( .A(core__abc_21380_n4079), .Y(core__abc_21380_n4080_1) );
  INVX1 INVX1_842 ( .A(core__abc_21380_n4082_1), .Y(core__abc_21380_n4083) );
  INVX1 INVX1_843 ( .A(core__abc_21380_n4088), .Y(core__abc_21380_n4093) );
  INVX1 INVX1_844 ( .A(core__abc_21380_n4089), .Y(core__abc_21380_n4094) );
  INVX1 INVX1_845 ( .A(core__abc_21380_n4098_1), .Y(core__abc_21380_n4099) );
  INVX1 INVX1_846 ( .A(core_v3_reg_60_), .Y(core__abc_21380_n4100) );
  INVX1 INVX1_847 ( .A(core__abc_21380_n4102_1), .Y(core__abc_21380_n4104) );
  INVX1 INVX1_848 ( .A(core__abc_21380_n4106_1), .Y(core__abc_21380_n4107) );
  INVX1 INVX1_849 ( .A(core__abc_21380_n4110), .Y(core__abc_21380_n4111_1) );
  INVX1 INVX1_85 ( .A(_abc_19068_n2544), .Y(_abc_19068_n2545) );
  INVX1 INVX1_850 ( .A(core__abc_21380_n4114), .Y(core__abc_21380_n4115_1) );
  INVX1 INVX1_851 ( .A(core__abc_21380_n4118), .Y(core__abc_21380_n4119) );
  INVX1 INVX1_852 ( .A(core__abc_21380_n4121), .Y(core__abc_21380_n4123) );
  INVX1 INVX1_853 ( .A(core_v3_reg_39_), .Y(core__abc_21380_n4127) );
  INVX1 INVX1_854 ( .A(core__abc_21380_n4122), .Y(core__abc_21380_n4128) );
  INVX1 INVX1_855 ( .A(core__abc_21380_n4142), .Y(core__abc_21380_n4143) );
  INVX1 INVX1_856 ( .A(core__abc_21380_n4112), .Y(core__abc_21380_n4152) );
  INVX1 INVX1_857 ( .A(core__abc_21380_n4116), .Y(core__abc_21380_n4153_1) );
  INVX1 INVX1_858 ( .A(core__abc_21380_n4154), .Y(core__abc_21380_n4155) );
  INVX1 INVX1_859 ( .A(core__abc_21380_n4158), .Y(core__abc_21380_n4159) );
  INVX1 INVX1_86 ( .A(_abc_19068_n2549), .Y(_abc_19068_n2550) );
  INVX1 INVX1_860 ( .A(core_v3_reg_61_), .Y(core__abc_21380_n4161_1) );
  INVX1 INVX1_861 ( .A(core__abc_21380_n4162), .Y(core__abc_21380_n4163) );
  INVX1 INVX1_862 ( .A(core__abc_21380_n4166), .Y(core__abc_21380_n4168) );
  INVX1 INVX1_863 ( .A(core__abc_21380_n4170_1), .Y(core__abc_21380_n4171) );
  INVX1 INVX1_864 ( .A(core__abc_21380_n4172), .Y(core__abc_21380_n4173_1) );
  INVX1 INVX1_865 ( .A(core__abc_21380_n4160), .Y(core__abc_21380_n4174) );
  INVX1 INVX1_866 ( .A(core__abc_21380_n4175), .Y(core__abc_21380_n4176) );
  INVX1 INVX1_867 ( .A(core__abc_21380_n4177), .Y(core__abc_21380_n4178_1) );
  INVX1 INVX1_868 ( .A(core_v3_reg_40_), .Y(core__abc_21380_n4182_1) );
  INVX1 INVX1_869 ( .A(core__abc_21380_n4036), .Y(core__abc_21380_n4186_1) );
  INVX1 INVX1_87 ( .A(_abc_19068_n2554), .Y(_abc_19068_n2555) );
  INVX1 INVX1_870 ( .A(core__abc_21380_n4194_1), .Y(core__abc_21380_n4195) );
  INVX1 INVX1_871 ( .A(core__abc_21380_n4198_1), .Y(core__abc_21380_n4199) );
  INVX1 INVX1_872 ( .A(core__abc_21380_n4202), .Y(core__abc_21380_n4203_1) );
  INVX1 INVX1_873 ( .A(core__abc_21380_n4181), .Y(core__abc_21380_n4205) );
  INVX1 INVX1_874 ( .A(core_key_77_), .Y(core__abc_21380_n4209) );
  INVX1 INVX1_875 ( .A(core__abc_21380_n4212), .Y(core__abc_21380_n4213) );
  INVX1 INVX1_876 ( .A(core__abc_21380_n4222), .Y(core__abc_21380_n4223) );
  INVX1 INVX1_877 ( .A(core__abc_21380_n2077), .Y(core__abc_21380_n4225) );
  INVX1 INVX1_878 ( .A(core__abc_21380_n4227), .Y(core__abc_21380_n4231) );
  INVX1 INVX1_879 ( .A(core__abc_21380_n4234), .Y(core__abc_21380_n4235) );
  INVX1 INVX1_88 ( .A(_abc_19068_n2559), .Y(_abc_19068_n2560) );
  INVX1 INVX1_880 ( .A(core_v3_reg_62_), .Y(core__abc_21380_n4236) );
  INVX1 INVX1_881 ( .A(core__abc_21380_n4238), .Y(core__abc_21380_n4239) );
  INVX1 INVX1_882 ( .A(core__abc_21380_n4242), .Y(core__abc_21380_n4243_1) );
  INVX1 INVX1_883 ( .A(core__abc_21380_n4246), .Y(core__abc_21380_n4247) );
  INVX1 INVX1_884 ( .A(core__abc_21380_n4253), .Y(core__abc_21380_n4254) );
  INVX1 INVX1_885 ( .A(core__abc_21380_n4258), .Y(core__abc_21380_n4259) );
  INVX1 INVX1_886 ( .A(core_v3_reg_41_), .Y(core__abc_21380_n4261) );
  INVX1 INVX1_887 ( .A(core__abc_21380_n4197), .Y(core__abc_21380_n4263) );
  INVX1 INVX1_888 ( .A(core__abc_21380_n4268), .Y(core__abc_21380_n4270) );
  INVX1 INVX1_889 ( .A(core__abc_21380_n4260), .Y(core__abc_21380_n4274) );
  INVX1 INVX1_89 ( .A(_abc_19068_n2564), .Y(_abc_19068_n2565) );
  INVX1 INVX1_890 ( .A(core__abc_21380_n4272), .Y(core__abc_21380_n4275) );
  INVX1 INVX1_891 ( .A(core_key_78_), .Y(core__abc_21380_n4279) );
  INVX1 INVX1_892 ( .A(core__abc_21380_n4282), .Y(core__abc_21380_n4283) );
  INVX1 INVX1_893 ( .A(core__abc_21380_n4248), .Y(core__abc_21380_n4292) );
  INVX1 INVX1_894 ( .A(core__abc_21380_n2115), .Y(core__abc_21380_n4294_1) );
  INVX1 INVX1_895 ( .A(core_v3_reg_63_), .Y(core__abc_21380_n4301) );
  INVX1 INVX1_896 ( .A(core__abc_21380_n4302), .Y(core__abc_21380_n4303) );
  INVX1 INVX1_897 ( .A(core__abc_21380_n4306), .Y(core__abc_21380_n4308) );
  INVX1 INVX1_898 ( .A(core__abc_21380_n4310), .Y(core__abc_21380_n4311) );
  INVX1 INVX1_899 ( .A(core__abc_21380_n4318), .Y(core__abc_21380_n4319_1) );
  INVX1 INVX1_9 ( .A(we), .Y(_abc_19068_n921_1) );
  INVX1 INVX1_90 ( .A(_abc_19068_n2569), .Y(_abc_19068_n2570) );
  INVX1 INVX1_900 ( .A(core__abc_21380_n4321), .Y(core__abc_21380_n4322) );
  INVX1 INVX1_901 ( .A(core__abc_21380_n4325), .Y(core__abc_21380_n4326) );
  INVX1 INVX1_902 ( .A(core_v3_reg_42_), .Y(core__abc_21380_n4330) );
  INVX1 INVX1_903 ( .A(core__abc_21380_n4328), .Y(core__abc_21380_n4331) );
  INVX1 INVX1_904 ( .A(core__abc_21380_n4333), .Y(core__abc_21380_n4334_1) );
  INVX1 INVX1_905 ( .A(core__abc_21380_n4341), .Y(core__abc_21380_n4342) );
  INVX1 INVX1_906 ( .A(core__abc_21380_n4250), .Y(core__abc_21380_n4352) );
  INVX1 INVX1_907 ( .A(core__abc_21380_n4069), .Y(core__abc_21380_n4359) );
  INVX1 INVX1_908 ( .A(core__abc_21380_n4252), .Y(core__abc_21380_n4363) );
  INVX1 INVX1_909 ( .A(core__abc_21380_n4353), .Y(core__abc_21380_n4365) );
  INVX1 INVX1_91 ( .A(_abc_19068_n2574), .Y(_abc_19068_n2575) );
  INVX1 INVX1_910 ( .A(core__abc_21380_n4374), .Y(core__abc_21380_n4386_1) );
  INVX1 INVX1_911 ( .A(core__abc_21380_n4383), .Y(core__abc_21380_n4388) );
  INVX1 INVX1_912 ( .A(core__abc_21380_n4391), .Y(core__abc_21380_n4392_1) );
  INVX1 INVX1_913 ( .A(core__abc_21380_n3060), .Y(core__abc_21380_n4394) );
  INVX1 INVX1_914 ( .A(core__abc_21380_n4396), .Y(core__abc_21380_n4397_1) );
  INVX1 INVX1_915 ( .A(core__abc_21380_n4400), .Y(core__abc_21380_n4402_1) );
  INVX1 INVX1_916 ( .A(core__abc_21380_n4404), .Y(core__abc_21380_n4405) );
  INVX1 INVX1_917 ( .A(core__abc_21380_n4367), .Y(core__abc_21380_n4412_1) );
  INVX1 INVX1_918 ( .A(core__abc_21380_n4419), .Y(core__abc_21380_n4420) );
  INVX1 INVX1_919 ( .A(core__abc_21380_n4423), .Y(core__abc_21380_n4424) );
  INVX1 INVX1_92 ( .A(_abc_19068_n2579), .Y(_abc_19068_n2580) );
  INVX1 INVX1_920 ( .A(core__abc_21380_n4417_1), .Y(core__abc_21380_n4428) );
  INVX1 INVX1_921 ( .A(core__abc_21380_n4425), .Y(core__abc_21380_n4429) );
  INVX1 INVX1_922 ( .A(core__abc_21380_n4436), .Y(core__abc_21380_n4437) );
  INVX1 INVX1_923 ( .A(core__abc_21380_n4401), .Y(core__abc_21380_n4446) );
  INVX1 INVX1_924 ( .A(core__abc_21380_n4406), .Y(core__abc_21380_n4447) );
  INVX1 INVX1_925 ( .A(core__abc_21380_n4448_1), .Y(core__abc_21380_n4449) );
  INVX1 INVX1_926 ( .A(core__abc_21380_n4385), .Y(core__abc_21380_n4450) );
  INVX1 INVX1_927 ( .A(core__abc_21380_n2156), .Y(core__abc_21380_n4451) );
  INVX1 INVX1_928 ( .A(core__abc_21380_n4453), .Y(core__abc_21380_n4454_1) );
  INVX1 INVX1_929 ( .A(core__abc_21380_n4455), .Y(core__abc_21380_n4456) );
  INVX1 INVX1_93 ( .A(_abc_19068_n2584), .Y(_abc_19068_n2585) );
  INVX1 INVX1_930 ( .A(core__abc_21380_n4458), .Y(core__abc_21380_n4459_1) );
  INVX1 INVX1_931 ( .A(core__abc_21380_n4462), .Y(core__abc_21380_n4463) );
  INVX1 INVX1_932 ( .A(core__abc_21380_n4466), .Y(core__abc_21380_n4468) );
  INVX1 INVX1_933 ( .A(core__abc_21380_n4470), .Y(core__abc_21380_n4471) );
  INVX1 INVX1_934 ( .A(core__abc_21380_n4472), .Y(core__abc_21380_n4473) );
  INVX1 INVX1_935 ( .A(core__abc_21380_n4461), .Y(core__abc_21380_n4474_1) );
  INVX1 INVX1_936 ( .A(core__abc_21380_n4475), .Y(core__abc_21380_n4476) );
  INVX1 INVX1_937 ( .A(core__abc_21380_n4477), .Y(core__abc_21380_n4479) );
  INVX1 INVX1_938 ( .A(core__abc_21380_n4481), .Y(core__abc_21380_n4482) );
  INVX1 INVX1_939 ( .A(core__abc_21380_n4486), .Y(core__abc_21380_n4487) );
  INVX1 INVX1_94 ( .A(_abc_19068_n2589), .Y(_abc_19068_n2590) );
  INVX1 INVX1_940 ( .A(core__abc_21380_n4490), .Y(core__abc_21380_n4491_1) );
  INVX1 INVX1_941 ( .A(core_v3_reg_44_), .Y(core__abc_21380_n4493) );
  INVX1 INVX1_942 ( .A(core__abc_21380_n4495), .Y(core__abc_21380_n4496_1) );
  INVX1 INVX1_943 ( .A(core__abc_21380_n4503), .Y(core__abc_21380_n4504) );
  INVX1 INVX1_944 ( .A(core__abc_21380_n4514), .Y(core__abc_21380_n4515) );
  INVX1 INVX1_945 ( .A(core__abc_21380_n4518), .Y(core__abc_21380_n4519) );
  INVX1 INVX1_946 ( .A(core__abc_21380_n4521), .Y(core__abc_21380_n4522_1) );
  INVX1 INVX1_947 ( .A(core__abc_21380_n4525), .Y(core__abc_21380_n4526) );
  INVX1 INVX1_948 ( .A(core__abc_21380_n3071), .Y(core__abc_21380_n4527_1) );
  INVX1 INVX1_949 ( .A(core__abc_21380_n4531), .Y(core__abc_21380_n4532_1) );
  INVX1 INVX1_95 ( .A(_abc_19068_n2594), .Y(_abc_19068_n2595) );
  INVX1 INVX1_950 ( .A(core__abc_21380_n4533), .Y(core__abc_21380_n4534) );
  INVX1 INVX1_951 ( .A(core__abc_21380_n4537_1), .Y(core__abc_21380_n4538) );
  INVX1 INVX1_952 ( .A(core__abc_21380_n4541), .Y(core__abc_21380_n4543) );
  INVX1 INVX1_953 ( .A(core__abc_21380_n4546), .Y(core__abc_21380_n4548) );
  INVX1 INVX1_954 ( .A(core__abc_21380_n4551), .Y(core__abc_21380_n4552_1) );
  INVX1 INVX1_955 ( .A(core__abc_21380_n4554), .Y(core__abc_21380_n4555) );
  INVX1 INVX1_956 ( .A(core__abc_21380_n4545), .Y(core__abc_21380_n4557) );
  INVX1 INVX1_957 ( .A(core_key_82_), .Y(core__abc_21380_n4561) );
  INVX1 INVX1_958 ( .A(core__abc_21380_n4564), .Y(core__abc_21380_n4565_1) );
  INVX1 INVX1_959 ( .A(core_v3_reg_46_), .Y(core__abc_21380_n4574) );
  INVX1 INVX1_96 ( .A(_abc_19068_n2599), .Y(_abc_19068_n2600) );
  INVX1 INVX1_960 ( .A(core__abc_21380_n2400), .Y(core__abc_21380_n4575) );
  INVX1 INVX1_961 ( .A(core__abc_21380_n4577), .Y(core__abc_21380_n4578) );
  INVX1 INVX1_962 ( .A(core__abc_21380_n4581), .Y(core__abc_21380_n4583) );
  INVX1 INVX1_963 ( .A(core__abc_21380_n4539), .Y(core__abc_21380_n4586) );
  INVX1 INVX1_964 ( .A(core__abc_21380_n4544), .Y(core__abc_21380_n4587_1) );
  INVX1 INVX1_965 ( .A(core__abc_21380_n4588), .Y(core__abc_21380_n4589) );
  INVX1 INVX1_966 ( .A(core__abc_21380_n4592_1), .Y(core__abc_21380_n4593) );
  INVX1 INVX1_967 ( .A(core__abc_21380_n4596), .Y(core__abc_21380_n4597_1) );
  INVX1 INVX1_968 ( .A(core__abc_21380_n4599), .Y(core__abc_21380_n4600) );
  INVX1 INVX1_969 ( .A(core__abc_21380_n4603_1), .Y(core__abc_21380_n4604) );
  INVX1 INVX1_97 ( .A(_abc_19068_n2604), .Y(_abc_19068_n2605) );
  INVX1 INVX1_970 ( .A(core__abc_21380_n4594), .Y(core__abc_21380_n4606) );
  INVX1 INVX1_971 ( .A(core__abc_21380_n4608_1), .Y(core__abc_21380_n4609) );
  INVX1 INVX1_972 ( .A(core__abc_21380_n4612), .Y(core__abc_21380_n4613) );
  INVX1 INVX1_973 ( .A(core__abc_21380_n4585), .Y(core__abc_21380_n4616) );
  INVX1 INVX1_974 ( .A(core__abc_21380_n4621), .Y(core__abc_21380_n4622) );
  INVX1 INVX1_975 ( .A(core__abc_21380_n4639_1), .Y(core__abc_21380_n4640) );
  INVX1 INVX1_976 ( .A(core__abc_21380_n4643), .Y(core__abc_21380_n4644_1) );
  INVX1 INVX1_977 ( .A(core__abc_21380_n4646), .Y(core__abc_21380_n4648) );
  INVX1 INVX1_978 ( .A(core__abc_21380_n4650_1), .Y(core__abc_21380_n4651) );
  INVX1 INVX1_979 ( .A(core__abc_21380_n4654), .Y(core__abc_21380_n4655_1) );
  INVX1 INVX1_98 ( .A(_abc_19068_n2609), .Y(_abc_19068_n2610) );
  INVX1 INVX1_980 ( .A(core__abc_21380_n4605), .Y(core__abc_21380_n4659) );
  INVX1 INVX1_981 ( .A(core__abc_21380_n4661), .Y(core__abc_21380_n4662) );
  INVX1 INVX1_982 ( .A(core__abc_21380_n4665), .Y(core__abc_21380_n4666_1) );
  INVX1 INVX1_983 ( .A(core__abc_21380_n4667), .Y(core__abc_21380_n4668) );
  INVX1 INVX1_984 ( .A(core__abc_21380_n4672), .Y(core__abc_21380_n4673) );
  INVX1 INVX1_985 ( .A(core_v3_reg_47_), .Y(core__abc_21380_n4675) );
  INVX1 INVX1_986 ( .A(core__abc_21380_n4676_1), .Y(core__abc_21380_n4677) );
  INVX1 INVX1_987 ( .A(core__abc_21380_n4680), .Y(core__abc_21380_n4682) );
  INVX1 INVX1_988 ( .A(core__abc_21380_n4674), .Y(core__abc_21380_n4686_1) );
  INVX1 INVX1_989 ( .A(core__abc_21380_n4681_1), .Y(core__abc_21380_n4687) );
  INVX1 INVX1_99 ( .A(_abc_19068_n2614), .Y(_abc_19068_n2615) );
  INVX1 INVX1_990 ( .A(core_key_84_), .Y(core__abc_21380_n4693) );
  INVX1 INVX1_991 ( .A(core__abc_21380_n4696_1), .Y(core__abc_21380_n4697) );
  INVX1 INVX1_992 ( .A(core__abc_21380_n4706), .Y(core__abc_21380_n4707_1) );
  INVX1 INVX1_993 ( .A(core__abc_21380_n4710), .Y(core__abc_21380_n4711) );
  INVX1 INVX1_994 ( .A(core__abc_21380_n4712_1), .Y(core__abc_21380_n4713) );
  INVX1 INVX1_995 ( .A(core__abc_21380_n4716), .Y(core__abc_21380_n4718) );
  INVX1 INVX1_996 ( .A(core__abc_21380_n4720), .Y(core__abc_21380_n4721) );
  INVX1 INVX1_997 ( .A(core__abc_21380_n4656), .Y(core__abc_21380_n4725) );
  INVX1 INVX1_998 ( .A(core__abc_21380_n4728), .Y(core__abc_21380_n4729) );
  INVX1 INVX1_999 ( .A(core__abc_21380_n4730), .Y(core__abc_21380_n4731) );
  INVX2 INVX2_1 ( .A(\write_data[0] ), .Y(_abc_19068_n2135) );
  INVX2 INVX2_10 ( .A(\write_data[9] ), .Y(_abc_19068_n2189) );
  INVX2 INVX2_11 ( .A(\write_data[10] ), .Y(_abc_19068_n2195) );
  INVX2 INVX2_12 ( .A(\write_data[11] ), .Y(_abc_19068_n2201) );
  INVX2 INVX2_13 ( .A(\write_data[12] ), .Y(_abc_19068_n2207) );
  INVX2 INVX2_14 ( .A(\write_data[13] ), .Y(_abc_19068_n2213) );
  INVX2 INVX2_15 ( .A(\write_data[14] ), .Y(_abc_19068_n2219) );
  INVX2 INVX2_16 ( .A(\write_data[15] ), .Y(_abc_19068_n2225) );
  INVX2 INVX2_17 ( .A(\write_data[16] ), .Y(_abc_19068_n2231) );
  INVX2 INVX2_18 ( .A(\write_data[17] ), .Y(_abc_19068_n2237) );
  INVX2 INVX2_19 ( .A(\write_data[18] ), .Y(_abc_19068_n2243) );
  INVX2 INVX2_2 ( .A(\write_data[1] ), .Y(_abc_19068_n2141) );
  INVX2 INVX2_20 ( .A(\write_data[19] ), .Y(_abc_19068_n2249) );
  INVX2 INVX2_21 ( .A(\write_data[20] ), .Y(_abc_19068_n2255) );
  INVX2 INVX2_22 ( .A(\write_data[21] ), .Y(_abc_19068_n2261) );
  INVX2 INVX2_23 ( .A(\write_data[22] ), .Y(_abc_19068_n2267) );
  INVX2 INVX2_24 ( .A(\write_data[23] ), .Y(_abc_19068_n2273) );
  INVX2 INVX2_25 ( .A(\write_data[24] ), .Y(_abc_19068_n2279) );
  INVX2 INVX2_26 ( .A(\write_data[25] ), .Y(_abc_19068_n2285) );
  INVX2 INVX2_27 ( .A(\write_data[26] ), .Y(_abc_19068_n2291) );
  INVX2 INVX2_28 ( .A(\write_data[27] ), .Y(_abc_19068_n2297) );
  INVX2 INVX2_29 ( .A(\write_data[28] ), .Y(_abc_19068_n2303) );
  INVX2 INVX2_3 ( .A(\write_data[2] ), .Y(_abc_19068_n2147) );
  INVX2 INVX2_30 ( .A(\write_data[29] ), .Y(_abc_19068_n2309) );
  INVX2 INVX2_31 ( .A(\write_data[30] ), .Y(_abc_19068_n2315) );
  INVX2 INVX2_32 ( .A(\write_data[31] ), .Y(_abc_19068_n2321) );
  INVX2 INVX2_33 ( .A(_abc_19068_n3131), .Y(_abc_19068_n3133) );
  INVX2 INVX2_34 ( .A(core__abc_21380_n1141_1), .Y(core__abc_21380_n1142_1) );
  INVX2 INVX2_35 ( .A(core_initalize), .Y(core__abc_21380_n1144_1) );
  INVX2 INVX2_36 ( .A(core__abc_21380_n1875), .Y(core__abc_21380_n1876) );
  INVX2 INVX2_37 ( .A(core_long), .Y(core__abc_21380_n7079) );
  INVX2 INVX2_4 ( .A(\write_data[3] ), .Y(_abc_19068_n2153) );
  INVX2 INVX2_5 ( .A(\write_data[4] ), .Y(_abc_19068_n2159) );
  INVX2 INVX2_6 ( .A(\write_data[5] ), .Y(_abc_19068_n2165) );
  INVX2 INVX2_7 ( .A(\write_data[6] ), .Y(_abc_19068_n2171) );
  INVX2 INVX2_8 ( .A(\write_data[7] ), .Y(_abc_19068_n2177) );
  INVX2 INVX2_9 ( .A(\write_data[8] ), .Y(_abc_19068_n2183) );
  INVX8 INVX8_1 ( .A(core_siphash_valid_reg_bF_buf8), .Y(_abc_19068_n1620) );
  INVX8 INVX8_2 ( .A(core_siphash_word1_we_bF_buf7), .Y(core__abc_21380_n1134_1) );
  INVX8 INVX8_3 ( .A(core__abc_21380_n2451_1_bF_buf7), .Y(core__abc_21380_n2452) );
  INVX8 INVX8_4 ( .A(core__abc_21380_n2749_bF_buf10), .Y(core__abc_21380_n2750) );
  INVX8 INVX8_5 ( .A(core__abc_21380_n3317_bF_buf6), .Y(core__abc_21380_n3328) );
  INVX8 INVX8_6 ( .A(core__abc_21380_n7076_bF_buf5), .Y(core__abc_21380_n7087) );
  INVX8 INVX8_7 ( .A(core__abc_21380_n8454_bF_buf7), .Y(core__abc_21380_n8455) );
  INVX8 INVX8_8 ( .A(core__abc_21380_n9245_bF_buf7), .Y(core__abc_21380_n9246) );
  OR2X2 OR2X2_1 ( .A(_abc_19068_n885_1), .B(_abc_19068_n889_1), .Y(_abc_19068_n890) );
  OR2X2 OR2X2_10 ( .A(_abc_19068_n917), .B(_abc_19068_n914), .Y(_abc_19068_n918_1) );
  OR2X2 OR2X2_100 ( .A(_abc_19068_n1116_1), .B(_abc_19068_n1109), .Y(_abc_19068_n1117_1) );
  OR2X2 OR2X2_1000 ( .A(core__abc_21380_n2297), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n2298_1) );
  OR2X2 OR2X2_1001 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_119_), .Y(core__abc_21380_n2299) );
  OR2X2 OR2X2_1002 ( .A(core__abc_21380_n2304), .B(core__abc_21380_n2305), .Y(core__abc_21380_n2306) );
  OR2X2 OR2X2_1003 ( .A(core_v2_reg_56_), .B(core_v3_reg_56_), .Y(core__abc_21380_n2308) );
  OR2X2 OR2X2_1004 ( .A(core__abc_21380_n2307), .B(core__abc_21380_n2311), .Y(core__abc_21380_n2312) );
  OR2X2 OR2X2_1005 ( .A(core__abc_21380_n2313), .B(core__abc_21380_n2306), .Y(core__abc_21380_n2314) );
  OR2X2 OR2X2_1006 ( .A(core__abc_21380_n2315), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n2316) );
  OR2X2 OR2X2_1007 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_120_), .Y(core__abc_21380_n2317) );
  OR2X2 OR2X2_1008 ( .A(core__abc_21380_n2322), .B(core__abc_21380_n2323), .Y(core__abc_21380_n2324) );
  OR2X2 OR2X2_1009 ( .A(core_v2_reg_57_), .B(core_v3_reg_57_), .Y(core__abc_21380_n2326) );
  OR2X2 OR2X2_101 ( .A(_abc_19068_n1117_1), .B(_abc_19068_n1104_1), .Y(_abc_19068_n1118) );
  OR2X2 OR2X2_1010 ( .A(core__abc_21380_n2325), .B(core__abc_21380_n2329), .Y(core__abc_21380_n2330) );
  OR2X2 OR2X2_1011 ( .A(core__abc_21380_n2331), .B(core__abc_21380_n2324), .Y(core__abc_21380_n2332_1) );
  OR2X2 OR2X2_1012 ( .A(core__abc_21380_n2333), .B(core__abc_21380_n1134_1_bF_buf5), .Y(core__abc_21380_n2334) );
  OR2X2 OR2X2_1013 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_121_), .Y(core__abc_21380_n2335) );
  OR2X2 OR2X2_1014 ( .A(core__abc_21380_n2340), .B(core__abc_21380_n2341), .Y(core__abc_21380_n2342) );
  OR2X2 OR2X2_1015 ( .A(core_v3_reg_58_), .B(core_v2_reg_58_), .Y(core__abc_21380_n2344) );
  OR2X2 OR2X2_1016 ( .A(core__abc_21380_n2343), .B(core__abc_21380_n2347), .Y(core__abc_21380_n2348) );
  OR2X2 OR2X2_1017 ( .A(core__abc_21380_n2349), .B(core__abc_21380_n2342), .Y(core__abc_21380_n2350) );
  OR2X2 OR2X2_1018 ( .A(core__abc_21380_n2351), .B(core__abc_21380_n1134_1_bF_buf4), .Y(core__abc_21380_n2352) );
  OR2X2 OR2X2_1019 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_122_), .Y(core__abc_21380_n2353) );
  OR2X2 OR2X2_102 ( .A(_abc_19068_n1120_1), .B(_abc_19068_n1121), .Y(_abc_19068_n1122_1) );
  OR2X2 OR2X2_1020 ( .A(core_v3_reg_59_), .B(core_v2_reg_59_), .Y(core__abc_21380_n2363_1) );
  OR2X2 OR2X2_1021 ( .A(core__abc_21380_n2362), .B(core__abc_21380_n2366), .Y(core__abc_21380_n2367) );
  OR2X2 OR2X2_1022 ( .A(core__abc_21380_n2368), .B(core__abc_21380_n2369_1), .Y(core__abc_21380_n2370) );
  OR2X2 OR2X2_1023 ( .A(core__abc_21380_n2371), .B(core__abc_21380_n1134_1_bF_buf3), .Y(core__abc_21380_n2372) );
  OR2X2 OR2X2_1024 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_123_), .Y(core__abc_21380_n2373) );
  OR2X2 OR2X2_1025 ( .A(core__abc_21380_n2378), .B(core__abc_21380_n2379), .Y(core__abc_21380_n2380) );
  OR2X2 OR2X2_1026 ( .A(core_v3_reg_60_), .B(core_v2_reg_60_), .Y(core__abc_21380_n2382) );
  OR2X2 OR2X2_1027 ( .A(core__abc_21380_n2381), .B(core__abc_21380_n2385), .Y(core__abc_21380_n2386) );
  OR2X2 OR2X2_1028 ( .A(core__abc_21380_n2387), .B(core__abc_21380_n2380), .Y(core__abc_21380_n2388) );
  OR2X2 OR2X2_1029 ( .A(core__abc_21380_n2389), .B(core__abc_21380_n1134_1_bF_buf2), .Y(core__abc_21380_n2390) );
  OR2X2 OR2X2_103 ( .A(_abc_19068_n1124), .B(_abc_19068_n1125_1), .Y(_abc_19068_n1126_1) );
  OR2X2 OR2X2_1030 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_124_), .Y(core__abc_21380_n2391_1) );
  OR2X2 OR2X2_1031 ( .A(core__abc_21380_n2396), .B(core__abc_21380_n2397), .Y(core__abc_21380_n2398) );
  OR2X2 OR2X2_1032 ( .A(core_v3_reg_61_), .B(core_v2_reg_61_), .Y(core__abc_21380_n2400) );
  OR2X2 OR2X2_1033 ( .A(core__abc_21380_n2399), .B(core__abc_21380_n2403), .Y(core__abc_21380_n2404) );
  OR2X2 OR2X2_1034 ( .A(core__abc_21380_n2405), .B(core__abc_21380_n2398), .Y(core__abc_21380_n2406) );
  OR2X2 OR2X2_1035 ( .A(core__abc_21380_n2407), .B(core__abc_21380_n1134_1_bF_buf1), .Y(core__abc_21380_n2408) );
  OR2X2 OR2X2_1036 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_125_), .Y(core__abc_21380_n2409) );
  OR2X2 OR2X2_1037 ( .A(core__abc_21380_n2414), .B(core__abc_21380_n2415), .Y(core__abc_21380_n2416) );
  OR2X2 OR2X2_1038 ( .A(core_v3_reg_62_), .B(core_v2_reg_62_), .Y(core__abc_21380_n2418) );
  OR2X2 OR2X2_1039 ( .A(core__abc_21380_n2417), .B(core__abc_21380_n2421), .Y(core__abc_21380_n2422) );
  OR2X2 OR2X2_104 ( .A(_abc_19068_n1126_1), .B(_abc_19068_n1123_1), .Y(_abc_19068_n1127) );
  OR2X2 OR2X2_1040 ( .A(core__abc_21380_n2423), .B(core__abc_21380_n2416), .Y(core__abc_21380_n2424_1) );
  OR2X2 OR2X2_1041 ( .A(core__abc_21380_n2425), .B(core__abc_21380_n1134_1_bF_buf0), .Y(core__abc_21380_n2426) );
  OR2X2 OR2X2_1042 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_126_), .Y(core__abc_21380_n2427) );
  OR2X2 OR2X2_1043 ( .A(core__abc_21380_n2430_1), .B(core_v1_reg_63_), .Y(core__abc_21380_n2431) );
  OR2X2 OR2X2_1044 ( .A(core__abc_21380_n2432), .B(core_v0_reg_63_), .Y(core__abc_21380_n2433) );
  OR2X2 OR2X2_1045 ( .A(core_v3_reg_63_), .B(core_v2_reg_63_), .Y(core__abc_21380_n2436) );
  OR2X2 OR2X2_1046 ( .A(core__abc_21380_n2441), .B(core__abc_21380_n2442), .Y(core__abc_21380_n2443) );
  OR2X2 OR2X2_1047 ( .A(core__abc_21380_n2443), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n2444) );
  OR2X2 OR2X2_1048 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_127_), .Y(core__abc_21380_n2445_1) );
  OR2X2 OR2X2_1049 ( .A(core__abc_21380_n2452_bF_buf7), .B(core__abc_21380_n1272_1), .Y(core__abc_21380_n2453) );
  OR2X2 OR2X2_105 ( .A(_abc_19068_n1127), .B(_abc_19068_n1122_1), .Y(_abc_19068_n1128_1) );
  OR2X2 OR2X2_1050 ( .A(core__abc_21380_n2451_1_bF_buf6), .B(core_siphash_word_0_), .Y(core__abc_21380_n2454) );
  OR2X2 OR2X2_1051 ( .A(core__abc_21380_n2452_bF_buf6), .B(core__abc_21380_n1293), .Y(core__abc_21380_n2457) );
  OR2X2 OR2X2_1052 ( .A(core__abc_21380_n2451_1_bF_buf5), .B(core_siphash_word_1_), .Y(core__abc_21380_n2458) );
  OR2X2 OR2X2_1053 ( .A(core__abc_21380_n1312), .B(core__abc_21380_n2452_bF_buf5), .Y(core__abc_21380_n2461) );
  OR2X2 OR2X2_1054 ( .A(core__abc_21380_n2451_1_bF_buf4), .B(core_siphash_word_2_), .Y(core__abc_21380_n2462) );
  OR2X2 OR2X2_1055 ( .A(core__abc_21380_n2465), .B(core__abc_21380_n2466), .Y(core__abc_21380_n2467) );
  OR2X2 OR2X2_1056 ( .A(core__abc_21380_n2452_bF_buf3), .B(core__abc_21380_n1349), .Y(core__abc_21380_n2469) );
  OR2X2 OR2X2_1057 ( .A(core__abc_21380_n2451_1_bF_buf2), .B(core_siphash_word_4_), .Y(core__abc_21380_n2470) );
  OR2X2 OR2X2_1058 ( .A(core__abc_21380_n2473), .B(core__abc_21380_n2474), .Y(core__abc_21380_n2475) );
  OR2X2 OR2X2_1059 ( .A(core__abc_21380_n1387), .B(core__abc_21380_n2452_bF_buf1), .Y(core__abc_21380_n2477_1) );
  OR2X2 OR2X2_106 ( .A(_abc_19068_n1130), .B(_abc_19068_n1131_1), .Y(_abc_19068_n1132) );
  OR2X2 OR2X2_1060 ( .A(core__abc_21380_n2451_1_bF_buf0), .B(core_siphash_word_6_), .Y(core__abc_21380_n2478) );
  OR2X2 OR2X2_1061 ( .A(core__abc_21380_n1406), .B(core__abc_21380_n2452_bF_buf0), .Y(core__abc_21380_n2481) );
  OR2X2 OR2X2_1062 ( .A(core__abc_21380_n2451_1_bF_buf7), .B(core_siphash_word_7_), .Y(core__abc_21380_n2482) );
  OR2X2 OR2X2_1063 ( .A(core__abc_21380_n2486), .B(core__abc_21380_n2485), .Y(core__abc_21380_n2487) );
  OR2X2 OR2X2_1064 ( .A(core__abc_21380_n1443), .B(core__abc_21380_n2452_bF_buf6), .Y(core__abc_21380_n2489) );
  OR2X2 OR2X2_1065 ( .A(core__abc_21380_n2451_1_bF_buf5), .B(core_siphash_word_9_), .Y(core__abc_21380_n2490) );
  OR2X2 OR2X2_1066 ( .A(core__abc_21380_n2452_bF_buf5), .B(core__abc_21380_n1460), .Y(core__abc_21380_n2493_1) );
  OR2X2 OR2X2_1067 ( .A(core__abc_21380_n2451_1_bF_buf4), .B(core_siphash_word_10_), .Y(core__abc_21380_n2494) );
  OR2X2 OR2X2_1068 ( .A(core__abc_21380_n2452_bF_buf4), .B(core__abc_21380_n1477), .Y(core__abc_21380_n2497_1) );
  OR2X2 OR2X2_1069 ( .A(core__abc_21380_n2451_1_bF_buf3), .B(core_siphash_word_11_), .Y(core__abc_21380_n2498) );
  OR2X2 OR2X2_107 ( .A(_abc_19068_n1133), .B(_abc_19068_n1134_1), .Y(_abc_19068_n1135) );
  OR2X2 OR2X2_1070 ( .A(core__abc_21380_n2502), .B(core__abc_21380_n2501), .Y(core__abc_21380_n2503) );
  OR2X2 OR2X2_1071 ( .A(core__abc_21380_n2452_bF_buf2), .B(core__abc_21380_n1513), .Y(core__abc_21380_n2505) );
  OR2X2 OR2X2_1072 ( .A(core__abc_21380_n2451_1_bF_buf1), .B(core_siphash_word_13_), .Y(core__abc_21380_n2506) );
  OR2X2 OR2X2_1073 ( .A(core__abc_21380_n2452_bF_buf1), .B(core__abc_21380_n1531), .Y(core__abc_21380_n2509) );
  OR2X2 OR2X2_1074 ( .A(core__abc_21380_n2451_1_bF_buf0), .B(core_siphash_word_14_), .Y(core__abc_21380_n2510) );
  OR2X2 OR2X2_1075 ( .A(core__abc_21380_n1551), .B(core__abc_21380_n2452_bF_buf0), .Y(core__abc_21380_n2513) );
  OR2X2 OR2X2_1076 ( .A(core__abc_21380_n2451_1_bF_buf7), .B(core_siphash_word_15_), .Y(core__abc_21380_n2514) );
  OR2X2 OR2X2_1077 ( .A(core__abc_21380_n2518), .B(core__abc_21380_n2517), .Y(core__abc_21380_n2519) );
  OR2X2 OR2X2_1078 ( .A(core__abc_21380_n1589), .B(core__abc_21380_n2452_bF_buf6), .Y(core__abc_21380_n2521) );
  OR2X2 OR2X2_1079 ( .A(core__abc_21380_n2451_1_bF_buf5), .B(core_siphash_word_17_), .Y(core__abc_21380_n2522) );
  OR2X2 OR2X2_108 ( .A(_abc_19068_n1132), .B(_abc_19068_n1135), .Y(_abc_19068_n1136_1) );
  OR2X2 OR2X2_1080 ( .A(core__abc_21380_n2452_bF_buf5), .B(core__abc_21380_n1606), .Y(core__abc_21380_n2525) );
  OR2X2 OR2X2_1081 ( .A(core__abc_21380_n2451_1_bF_buf4), .B(core_siphash_word_18_), .Y(core__abc_21380_n2526) );
  OR2X2 OR2X2_1082 ( .A(core__abc_21380_n2530), .B(core__abc_21380_n2529), .Y(core__abc_21380_n2531) );
  OR2X2 OR2X2_1083 ( .A(core__abc_21380_n2452_bF_buf3), .B(core__abc_21380_n1641), .Y(core__abc_21380_n2533) );
  OR2X2 OR2X2_1084 ( .A(core__abc_21380_n2451_1_bF_buf2), .B(core_siphash_word_20_), .Y(core__abc_21380_n2534_1) );
  OR2X2 OR2X2_1085 ( .A(core__abc_21380_n2452_bF_buf2), .B(core__abc_21380_n1659), .Y(core__abc_21380_n2537) );
  OR2X2 OR2X2_1086 ( .A(core__abc_21380_n2451_1_bF_buf1), .B(core_siphash_word_21_), .Y(core__abc_21380_n2538) );
  OR2X2 OR2X2_1087 ( .A(core__abc_21380_n2452_bF_buf1), .B(core__abc_21380_n1677), .Y(core__abc_21380_n2541) );
  OR2X2 OR2X2_1088 ( .A(core__abc_21380_n2451_1_bF_buf0), .B(core_siphash_word_22_), .Y(core__abc_21380_n2542) );
  OR2X2 OR2X2_1089 ( .A(core__abc_21380_n1697), .B(core__abc_21380_n2452_bF_buf0), .Y(core__abc_21380_n2545) );
  OR2X2 OR2X2_109 ( .A(_abc_19068_n1136_1), .B(_abc_19068_n1129_1), .Y(_abc_19068_n1137_1) );
  OR2X2 OR2X2_1090 ( .A(core__abc_21380_n2451_1_bF_buf7), .B(core_siphash_word_23_), .Y(core__abc_21380_n2546) );
  OR2X2 OR2X2_1091 ( .A(core__abc_21380_n2452_bF_buf7), .B(core__abc_21380_n1715), .Y(core__abc_21380_n2549) );
  OR2X2 OR2X2_1092 ( .A(core__abc_21380_n2451_1_bF_buf6), .B(core_siphash_word_24_), .Y(core__abc_21380_n2550) );
  OR2X2 OR2X2_1093 ( .A(core__abc_21380_n1735), .B(core__abc_21380_n2452_bF_buf6), .Y(core__abc_21380_n2553) );
  OR2X2 OR2X2_1094 ( .A(core__abc_21380_n2451_1_bF_buf5), .B(core_siphash_word_25_), .Y(core__abc_21380_n2554) );
  OR2X2 OR2X2_1095 ( .A(core__abc_21380_n2452_bF_buf5), .B(core__abc_21380_n1752), .Y(core__abc_21380_n2557) );
  OR2X2 OR2X2_1096 ( .A(core__abc_21380_n2451_1_bF_buf4), .B(core_siphash_word_26_), .Y(core__abc_21380_n2558) );
  OR2X2 OR2X2_1097 ( .A(core__abc_21380_n1772), .B(core__abc_21380_n2452_bF_buf4), .Y(core__abc_21380_n2561) );
  OR2X2 OR2X2_1098 ( .A(core__abc_21380_n2451_1_bF_buf3), .B(core_siphash_word_27_), .Y(core__abc_21380_n2562) );
  OR2X2 OR2X2_1099 ( .A(core__abc_21380_n2452_bF_buf3), .B(core__abc_21380_n1790), .Y(core__abc_21380_n2565) );
  OR2X2 OR2X2_11 ( .A(_abc_19068_n918_1), .B(_abc_19068_n910_1), .Y(_abc_19068_n919_1) );
  OR2X2 OR2X2_110 ( .A(_abc_19068_n1137_1), .B(_abc_19068_n1128_1), .Y(_abc_19068_n1138) );
  OR2X2 OR2X2_1100 ( .A(core__abc_21380_n2451_1_bF_buf2), .B(core_siphash_word_28_), .Y(core__abc_21380_n2566) );
  OR2X2 OR2X2_1101 ( .A(core__abc_21380_n1810), .B(core__abc_21380_n2452_bF_buf2), .Y(core__abc_21380_n2569) );
  OR2X2 OR2X2_1102 ( .A(core__abc_21380_n2451_1_bF_buf1), .B(core_siphash_word_29_), .Y(core__abc_21380_n2570) );
  OR2X2 OR2X2_1103 ( .A(core__abc_21380_n2452_bF_buf1), .B(core__abc_21380_n1828), .Y(core__abc_21380_n2573) );
  OR2X2 OR2X2_1104 ( .A(core__abc_21380_n2451_1_bF_buf0), .B(core_siphash_word_30_), .Y(core__abc_21380_n2574) );
  OR2X2 OR2X2_1105 ( .A(core__abc_21380_n1848), .B(core__abc_21380_n2452_bF_buf0), .Y(core__abc_21380_n2577) );
  OR2X2 OR2X2_1106 ( .A(core__abc_21380_n2451_1_bF_buf7), .B(core_siphash_word_31_), .Y(core__abc_21380_n2578_1) );
  OR2X2 OR2X2_1107 ( .A(core__abc_21380_n2452_bF_buf7), .B(core__abc_21380_n1866), .Y(core__abc_21380_n2581) );
  OR2X2 OR2X2_1108 ( .A(core__abc_21380_n2451_1_bF_buf6), .B(core_siphash_word_32_), .Y(core__abc_21380_n2582_1) );
  OR2X2 OR2X2_1109 ( .A(core__abc_21380_n2452_bF_buf6), .B(core__abc_21380_n1884), .Y(core__abc_21380_n2585) );
  OR2X2 OR2X2_111 ( .A(_abc_19068_n1140_1), .B(_abc_19068_n1141), .Y(_abc_19068_n1142_1) );
  OR2X2 OR2X2_1110 ( .A(core__abc_21380_n2451_1_bF_buf5), .B(core_siphash_word_33_), .Y(core__abc_21380_n2586) );
  OR2X2 OR2X2_1111 ( .A(core__abc_21380_n2452_bF_buf5), .B(core__abc_21380_n1902), .Y(core__abc_21380_n2589) );
  OR2X2 OR2X2_1112 ( .A(core__abc_21380_n2451_1_bF_buf4), .B(core_siphash_word_34_), .Y(core__abc_21380_n2590) );
  OR2X2 OR2X2_1113 ( .A(core__abc_21380_n1922), .B(core__abc_21380_n2452_bF_buf4), .Y(core__abc_21380_n2593) );
  OR2X2 OR2X2_1114 ( .A(core__abc_21380_n2451_1_bF_buf3), .B(core_siphash_word_35_), .Y(core__abc_21380_n2594) );
  OR2X2 OR2X2_1115 ( .A(core__abc_21380_n2452_bF_buf3), .B(core__abc_21380_n1940), .Y(core__abc_21380_n2597_1) );
  OR2X2 OR2X2_1116 ( .A(core__abc_21380_n2451_1_bF_buf2), .B(core_siphash_word_36_), .Y(core__abc_21380_n2598) );
  OR2X2 OR2X2_1117 ( .A(core__abc_21380_n2601), .B(core__abc_21380_n2602), .Y(core__abc_21380_n2603_1) );
  OR2X2 OR2X2_1118 ( .A(core__abc_21380_n2452_bF_buf1), .B(core__abc_21380_n1978), .Y(core__abc_21380_n2605) );
  OR2X2 OR2X2_1119 ( .A(core__abc_21380_n2451_1_bF_buf0), .B(core_siphash_word_38_), .Y(core__abc_21380_n2606) );
  OR2X2 OR2X2_112 ( .A(_abc_19068_n1144_1), .B(_abc_19068_n1145), .Y(_abc_19068_n1146_1) );
  OR2X2 OR2X2_1120 ( .A(core__abc_21380_n1998), .B(core__abc_21380_n2452_bF_buf0), .Y(core__abc_21380_n2609) );
  OR2X2 OR2X2_1121 ( .A(core__abc_21380_n2451_1_bF_buf7), .B(core_siphash_word_39_), .Y(core__abc_21380_n2610) );
  OR2X2 OR2X2_1122 ( .A(core__abc_21380_n2614), .B(core__abc_21380_n2613), .Y(core__abc_21380_n2615) );
  OR2X2 OR2X2_1123 ( .A(core__abc_21380_n2452_bF_buf6), .B(core__abc_21380_n2034), .Y(core__abc_21380_n2617) );
  OR2X2 OR2X2_1124 ( .A(core__abc_21380_n2451_1_bF_buf5), .B(core_siphash_word_41_), .Y(core__abc_21380_n2618) );
  OR2X2 OR2X2_1125 ( .A(core__abc_21380_n2452_bF_buf5), .B(core__abc_21380_n2052), .Y(core__abc_21380_n2621) );
  OR2X2 OR2X2_1126 ( .A(core__abc_21380_n2451_1_bF_buf4), .B(core_siphash_word_42_), .Y(core__abc_21380_n2622) );
  OR2X2 OR2X2_1127 ( .A(core__abc_21380_n2072), .B(core__abc_21380_n2452_bF_buf4), .Y(core__abc_21380_n2625) );
  OR2X2 OR2X2_1128 ( .A(core__abc_21380_n2451_1_bF_buf3), .B(core_siphash_word_43_), .Y(core__abc_21380_n2626) );
  OR2X2 OR2X2_1129 ( .A(core__abc_21380_n2630), .B(core__abc_21380_n2629), .Y(core__abc_21380_n2631) );
  OR2X2 OR2X2_113 ( .A(_abc_19068_n1146_1), .B(_abc_19068_n1143), .Y(_abc_19068_n1147_1) );
  OR2X2 OR2X2_1130 ( .A(core__abc_21380_n2110), .B(core__abc_21380_n2452_bF_buf2), .Y(core__abc_21380_n2633_1) );
  OR2X2 OR2X2_1131 ( .A(core__abc_21380_n2451_1_bF_buf1), .B(core_siphash_word_45_), .Y(core__abc_21380_n2634) );
  OR2X2 OR2X2_1132 ( .A(core__abc_21380_n2638), .B(core__abc_21380_n2637), .Y(core__abc_21380_n2639) );
  OR2X2 OR2X2_1133 ( .A(core__abc_21380_n2148), .B(core__abc_21380_n2452_bF_buf0), .Y(core__abc_21380_n2641) );
  OR2X2 OR2X2_1134 ( .A(core__abc_21380_n2451_1_bF_buf7), .B(core_siphash_word_47_), .Y(core__abc_21380_n2642) );
  OR2X2 OR2X2_1135 ( .A(core__abc_21380_n2452_bF_buf7), .B(core__abc_21380_n2166), .Y(core__abc_21380_n2645) );
  OR2X2 OR2X2_1136 ( .A(core__abc_21380_n2451_1_bF_buf6), .B(core_siphash_word_48_), .Y(core__abc_21380_n2646) );
  OR2X2 OR2X2_1137 ( .A(core__abc_21380_n2650), .B(core__abc_21380_n2649), .Y(core__abc_21380_n2651) );
  OR2X2 OR2X2_1138 ( .A(core__abc_21380_n2654_1), .B(core__abc_21380_n2653), .Y(core__abc_21380_n2655) );
  OR2X2 OR2X2_1139 ( .A(core__abc_21380_n2657), .B(core__abc_21380_n2658), .Y(core__abc_21380_n2659) );
  OR2X2 OR2X2_114 ( .A(_abc_19068_n1147_1), .B(_abc_19068_n1142_1), .Y(_abc_19068_n1148) );
  OR2X2 OR2X2_1140 ( .A(core__abc_21380_n2452_bF_buf3), .B(core__abc_21380_n2239), .Y(core__abc_21380_n2661) );
  OR2X2 OR2X2_1141 ( .A(core__abc_21380_n2451_1_bF_buf2), .B(core_siphash_word_52_), .Y(core__abc_21380_n2662) );
  OR2X2 OR2X2_1142 ( .A(core__abc_21380_n2665), .B(core__abc_21380_n2666), .Y(core__abc_21380_n2667) );
  OR2X2 OR2X2_1143 ( .A(core__abc_21380_n2452_bF_buf1), .B(core__abc_21380_n2277), .Y(core__abc_21380_n2669) );
  OR2X2 OR2X2_1144 ( .A(core__abc_21380_n2451_1_bF_buf0), .B(core_siphash_word_54_), .Y(core__abc_21380_n2670) );
  OR2X2 OR2X2_1145 ( .A(core__abc_21380_n2297), .B(core__abc_21380_n2452_bF_buf0), .Y(core__abc_21380_n2673) );
  OR2X2 OR2X2_1146 ( .A(core__abc_21380_n2451_1_bF_buf7), .B(core_siphash_word_55_), .Y(core__abc_21380_n2674) );
  OR2X2 OR2X2_1147 ( .A(core__abc_21380_n2452_bF_buf7), .B(core__abc_21380_n2315), .Y(core__abc_21380_n2677) );
  OR2X2 OR2X2_1148 ( .A(core__abc_21380_n2451_1_bF_buf6), .B(core_siphash_word_56_), .Y(core__abc_21380_n2678) );
  OR2X2 OR2X2_1149 ( .A(core__abc_21380_n2452_bF_buf6), .B(core__abc_21380_n2333), .Y(core__abc_21380_n2681) );
  OR2X2 OR2X2_115 ( .A(_abc_19068_n1150_1), .B(_abc_19068_n1151), .Y(_abc_19068_n1152_1) );
  OR2X2 OR2X2_1150 ( .A(core__abc_21380_n2451_1_bF_buf5), .B(core_siphash_word_57_), .Y(core__abc_21380_n2682_1) );
  OR2X2 OR2X2_1151 ( .A(core__abc_21380_n2452_bF_buf5), .B(core__abc_21380_n2351), .Y(core__abc_21380_n2685) );
  OR2X2 OR2X2_1152 ( .A(core__abc_21380_n2451_1_bF_buf4), .B(core_siphash_word_58_), .Y(core__abc_21380_n2686) );
  OR2X2 OR2X2_1153 ( .A(core__abc_21380_n2371), .B(core__abc_21380_n2452_bF_buf4), .Y(core__abc_21380_n2689) );
  OR2X2 OR2X2_1154 ( .A(core__abc_21380_n2451_1_bF_buf3), .B(core_siphash_word_59_), .Y(core__abc_21380_n2690) );
  OR2X2 OR2X2_1155 ( .A(core__abc_21380_n2452_bF_buf3), .B(core__abc_21380_n2389), .Y(core__abc_21380_n2693) );
  OR2X2 OR2X2_1156 ( .A(core__abc_21380_n2451_1_bF_buf2), .B(core_siphash_word_60_), .Y(core__abc_21380_n2694) );
  OR2X2 OR2X2_1157 ( .A(core__abc_21380_n2452_bF_buf2), .B(core__abc_21380_n2407), .Y(core__abc_21380_n2697) );
  OR2X2 OR2X2_1158 ( .A(core__abc_21380_n2451_1_bF_buf1), .B(core_siphash_word_61_), .Y(core__abc_21380_n2698) );
  OR2X2 OR2X2_1159 ( .A(core__abc_21380_n2452_bF_buf1), .B(core__abc_21380_n2425), .Y(core__abc_21380_n2701) );
  OR2X2 OR2X2_116 ( .A(_abc_19068_n1153_1), .B(_abc_19068_n1154), .Y(_abc_19068_n1155_1) );
  OR2X2 OR2X2_1160 ( .A(core__abc_21380_n2451_1_bF_buf0), .B(core_siphash_word_62_), .Y(core__abc_21380_n2702) );
  OR2X2 OR2X2_1161 ( .A(core__abc_21380_n2706), .B(core__abc_21380_n2705), .Y(core__abc_21380_n2707) );
  OR2X2 OR2X2_1162 ( .A(core__abc_21380_n2711), .B(core__abc_21380_n2709), .Y(core__abc_21380_n2712) );
  OR2X2 OR2X2_1163 ( .A(core__abc_21380_n2713), .B(core__abc_21380_n1244_1), .Y(core_ready_reg_FF_INPUT) );
  OR2X2 OR2X2_1164 ( .A(core__abc_21380_n2719), .B(core__abc_21380_n1155), .Y(core__abc_21380_n2720) );
  OR2X2 OR2X2_1165 ( .A(core__abc_21380_n2716), .B(core_loop_ctr_reg_0_), .Y(core__abc_21380_n2721) );
  OR2X2 OR2X2_1166 ( .A(core__abc_21380_n2724_1), .B(core__abc_21380_n2727), .Y(core__abc_21380_n2728_1) );
  OR2X2 OR2X2_1167 ( .A(core_loop_ctr_reg_1_), .B(core_loop_ctr_reg_0_), .Y(core__abc_21380_n2729) );
  OR2X2 OR2X2_1168 ( .A(core__abc_21380_n2732), .B(core__abc_21380_n2735), .Y(core__abc_21380_n2736) );
  OR2X2 OR2X2_1169 ( .A(core__abc_21380_n2725), .B(core_loop_ctr_reg_2_), .Y(core__abc_21380_n2737) );
  OR2X2 OR2X2_117 ( .A(_abc_19068_n1152_1), .B(_abc_19068_n1155_1), .Y(_abc_19068_n1156_1) );
  OR2X2 OR2X2_1170 ( .A(core__abc_21380_n2735), .B(core__abc_21380_n1180_1), .Y(core__abc_21380_n2740) );
  OR2X2 OR2X2_1171 ( .A(core__abc_21380_n2719), .B(core__abc_21380_n2740), .Y(core__abc_21380_n2741) );
  OR2X2 OR2X2_1172 ( .A(core__abc_21380_n2742), .B(core_loop_ctr_reg_3_), .Y(core__abc_21380_n2743) );
  OR2X2 OR2X2_1173 ( .A(core__abc_21380_n2751), .B(core__abc_21380_n2752), .Y(core__abc_21380_n2753) );
  OR2X2 OR2X2_1174 ( .A(core__abc_21380_n2755), .B(core__abc_21380_n2756), .Y(core__abc_21380_n2757) );
  OR2X2 OR2X2_1175 ( .A(core__abc_21380_n2759), .B(core__abc_21380_n2760), .Y(core__abc_21380_n2761) );
  OR2X2 OR2X2_1176 ( .A(core__abc_21380_n2763), .B(core__abc_21380_n2764), .Y(core__abc_21380_n2765) );
  OR2X2 OR2X2_1177 ( .A(core__abc_21380_n2767), .B(core__abc_21380_n2768), .Y(core__abc_21380_n2769) );
  OR2X2 OR2X2_1178 ( .A(core__abc_21380_n2771), .B(core__abc_21380_n2772), .Y(core__abc_21380_n2773) );
  OR2X2 OR2X2_1179 ( .A(core__abc_21380_n2775), .B(core__abc_21380_n2776), .Y(core__abc_21380_n2777) );
  OR2X2 OR2X2_118 ( .A(_abc_19068_n1156_1), .B(_abc_19068_n1149_1), .Y(_abc_19068_n1157) );
  OR2X2 OR2X2_1180 ( .A(core__abc_21380_n2779), .B(core__abc_21380_n2780), .Y(core__abc_21380_n2781) );
  OR2X2 OR2X2_1181 ( .A(core__abc_21380_n2783), .B(core__abc_21380_n2784), .Y(core__abc_21380_n2785) );
  OR2X2 OR2X2_1182 ( .A(core__abc_21380_n2787), .B(core__abc_21380_n2788), .Y(core__abc_21380_n2789) );
  OR2X2 OR2X2_1183 ( .A(core__abc_21380_n2791), .B(core__abc_21380_n2792), .Y(core__abc_21380_n2793) );
  OR2X2 OR2X2_1184 ( .A(core__abc_21380_n2795), .B(core__abc_21380_n2796), .Y(core__abc_21380_n2797) );
  OR2X2 OR2X2_1185 ( .A(core__abc_21380_n2799), .B(core__abc_21380_n2800_1), .Y(core__abc_21380_n2801) );
  OR2X2 OR2X2_1186 ( .A(core__abc_21380_n2803), .B(core__abc_21380_n2804_1), .Y(core__abc_21380_n2805) );
  OR2X2 OR2X2_1187 ( .A(core__abc_21380_n2807), .B(core__abc_21380_n2808), .Y(core__abc_21380_n2809) );
  OR2X2 OR2X2_1188 ( .A(core__abc_21380_n2811), .B(core__abc_21380_n2812), .Y(core__abc_21380_n2813) );
  OR2X2 OR2X2_1189 ( .A(core__abc_21380_n2815), .B(core__abc_21380_n2816), .Y(core__abc_21380_n2817_1) );
  OR2X2 OR2X2_119 ( .A(_abc_19068_n1157), .B(_abc_19068_n1148), .Y(_abc_19068_n1158_1) );
  OR2X2 OR2X2_1190 ( .A(core__abc_21380_n2819), .B(core__abc_21380_n2820), .Y(core__abc_21380_n2821) );
  OR2X2 OR2X2_1191 ( .A(core__abc_21380_n2823_1), .B(core__abc_21380_n2824), .Y(core__abc_21380_n2825) );
  OR2X2 OR2X2_1192 ( .A(core__abc_21380_n2827), .B(core__abc_21380_n2828), .Y(core__abc_21380_n2829) );
  OR2X2 OR2X2_1193 ( .A(core__abc_21380_n2831), .B(core__abc_21380_n2832), .Y(core__abc_21380_n2833) );
  OR2X2 OR2X2_1194 ( .A(core__abc_21380_n2835), .B(core__abc_21380_n2836), .Y(core__abc_21380_n2837) );
  OR2X2 OR2X2_1195 ( .A(core__abc_21380_n2839_1), .B(core__abc_21380_n2840), .Y(core__abc_21380_n2841) );
  OR2X2 OR2X2_1196 ( .A(core__abc_21380_n2843), .B(core__abc_21380_n2844), .Y(core__abc_21380_n2845_1) );
  OR2X2 OR2X2_1197 ( .A(core__abc_21380_n2847), .B(core__abc_21380_n2848), .Y(core__abc_21380_n2849) );
  OR2X2 OR2X2_1198 ( .A(core__abc_21380_n2851), .B(core__abc_21380_n2852), .Y(core__abc_21380_n2853) );
  OR2X2 OR2X2_1199 ( .A(core__abc_21380_n2855), .B(core__abc_21380_n2856), .Y(core__abc_21380_n2857) );
  OR2X2 OR2X2_12 ( .A(_abc_19068_n905), .B(_abc_19068_n919_1), .Y(_abc_19068_n920) );
  OR2X2 OR2X2_120 ( .A(_abc_19068_n1160), .B(_abc_19068_n1161_1), .Y(_abc_19068_n1162_1) );
  OR2X2 OR2X2_1200 ( .A(core__abc_21380_n2859), .B(core__abc_21380_n2860_1), .Y(core__abc_21380_n2861) );
  OR2X2 OR2X2_1201 ( .A(core__abc_21380_n2863), .B(core__abc_21380_n2864_1), .Y(core__abc_21380_n2865) );
  OR2X2 OR2X2_1202 ( .A(core__abc_21380_n2867), .B(core__abc_21380_n2868), .Y(core__abc_21380_n2869) );
  OR2X2 OR2X2_1203 ( .A(core__abc_21380_n2871), .B(core__abc_21380_n2872), .Y(core__abc_21380_n2873) );
  OR2X2 OR2X2_1204 ( .A(core__abc_21380_n2875), .B(core__abc_21380_n2876), .Y(core__abc_21380_n2877) );
  OR2X2 OR2X2_1205 ( .A(core__abc_21380_n2879), .B(core__abc_21380_n2880), .Y(core__abc_21380_n2881_1) );
  OR2X2 OR2X2_1206 ( .A(core__abc_21380_n2883), .B(core__abc_21380_n2884), .Y(core__abc_21380_n2885_1) );
  OR2X2 OR2X2_1207 ( .A(core__abc_21380_n2887), .B(core__abc_21380_n2888), .Y(core__abc_21380_n2889) );
  OR2X2 OR2X2_1208 ( .A(core__abc_21380_n2891), .B(core__abc_21380_n2892), .Y(core__abc_21380_n2893) );
  OR2X2 OR2X2_1209 ( .A(core__abc_21380_n2895), .B(core__abc_21380_n2896), .Y(core__abc_21380_n2897) );
  OR2X2 OR2X2_121 ( .A(_abc_19068_n1164_1), .B(_abc_19068_n1165_1), .Y(_abc_19068_n1166) );
  OR2X2 OR2X2_1210 ( .A(core__abc_21380_n2899), .B(core__abc_21380_n2900_1), .Y(core__abc_21380_n2901) );
  OR2X2 OR2X2_1211 ( .A(core__abc_21380_n2903), .B(core__abc_21380_n2904_1), .Y(core__abc_21380_n2905) );
  OR2X2 OR2X2_1212 ( .A(core__abc_21380_n2907), .B(core__abc_21380_n2908), .Y(core__abc_21380_n2909) );
  OR2X2 OR2X2_1213 ( .A(core__abc_21380_n2911), .B(core__abc_21380_n2912), .Y(core__abc_21380_n2913) );
  OR2X2 OR2X2_1214 ( .A(core__abc_21380_n2915), .B(core__abc_21380_n2916_1), .Y(core__abc_21380_n2917) );
  OR2X2 OR2X2_1215 ( .A(core__abc_21380_n2919), .B(core__abc_21380_n2920), .Y(core__abc_21380_n2921) );
  OR2X2 OR2X2_1216 ( .A(core__abc_21380_n2923), .B(core__abc_21380_n2924), .Y(core__abc_21380_n2925) );
  OR2X2 OR2X2_1217 ( .A(core__abc_21380_n2927), .B(core__abc_21380_n2928), .Y(core__abc_21380_n2929) );
  OR2X2 OR2X2_1218 ( .A(core__abc_21380_n2931), .B(core__abc_21380_n2932), .Y(core__abc_21380_n2933) );
  OR2X2 OR2X2_1219 ( .A(core__abc_21380_n2935), .B(core__abc_21380_n2936), .Y(core__abc_21380_n2937) );
  OR2X2 OR2X2_122 ( .A(_abc_19068_n1166), .B(_abc_19068_n1163), .Y(_abc_19068_n1167_1) );
  OR2X2 OR2X2_1220 ( .A(core__abc_21380_n2939), .B(core__abc_21380_n2940), .Y(core__abc_21380_n2941) );
  OR2X2 OR2X2_1221 ( .A(core__abc_21380_n2943), .B(core__abc_21380_n2944), .Y(core__abc_21380_n2945) );
  OR2X2 OR2X2_1222 ( .A(core__abc_21380_n2947), .B(core__abc_21380_n2948), .Y(core__abc_21380_n2949) );
  OR2X2 OR2X2_1223 ( .A(core__abc_21380_n2951), .B(core__abc_21380_n2952_1), .Y(core__abc_21380_n2953) );
  OR2X2 OR2X2_1224 ( .A(core__abc_21380_n2955), .B(core__abc_21380_n2956_1), .Y(core__abc_21380_n2957) );
  OR2X2 OR2X2_1225 ( .A(core__abc_21380_n2959), .B(core__abc_21380_n2960), .Y(core__abc_21380_n2961) );
  OR2X2 OR2X2_1226 ( .A(core__abc_21380_n2963), .B(core__abc_21380_n2964), .Y(core__abc_21380_n2965_1) );
  OR2X2 OR2X2_1227 ( .A(core__abc_21380_n2967), .B(core__abc_21380_n2968), .Y(core__abc_21380_n2969) );
  OR2X2 OR2X2_1228 ( .A(core__abc_21380_n2971_1), .B(core__abc_21380_n2972), .Y(core__abc_21380_n2973) );
  OR2X2 OR2X2_1229 ( .A(core__abc_21380_n2975), .B(core__abc_21380_n2976), .Y(core__abc_21380_n2977) );
  OR2X2 OR2X2_123 ( .A(_abc_19068_n1167_1), .B(_abc_19068_n1162_1), .Y(_abc_19068_n1168_1) );
  OR2X2 OR2X2_1230 ( .A(core__abc_21380_n2979), .B(core__abc_21380_n2980), .Y(core__abc_21380_n2981) );
  OR2X2 OR2X2_1231 ( .A(core__abc_21380_n2983), .B(core__abc_21380_n2984), .Y(core__abc_21380_n2985) );
  OR2X2 OR2X2_1232 ( .A(core__abc_21380_n2987), .B(core__abc_21380_n2988_1), .Y(core__abc_21380_n2989) );
  OR2X2 OR2X2_1233 ( .A(core__abc_21380_n2991), .B(core__abc_21380_n2992), .Y(core__abc_21380_n2993) );
  OR2X2 OR2X2_1234 ( .A(core__abc_21380_n2995), .B(core__abc_21380_n2996), .Y(core__abc_21380_n2997) );
  OR2X2 OR2X2_1235 ( .A(core__abc_21380_n2999), .B(core__abc_21380_n3000), .Y(core__abc_21380_n3001_1) );
  OR2X2 OR2X2_1236 ( .A(core__abc_21380_n3003), .B(core__abc_21380_n3004), .Y(core__abc_21380_n3005_1) );
  OR2X2 OR2X2_1237 ( .A(core__abc_21380_n2032), .B(core__abc_21380_n2010), .Y(core__abc_21380_n3008) );
  OR2X2 OR2X2_1238 ( .A(core__abc_21380_n3011), .B(core__abc_21380_n1323), .Y(core__abc_21380_n3012) );
  OR2X2 OR2X2_1239 ( .A(core__abc_21380_n3013), .B(core__abc_21380_n1281_1), .Y(core__abc_21380_n3014) );
  OR2X2 OR2X2_124 ( .A(_abc_19068_n1170_1), .B(_abc_19068_n1171_1), .Y(_abc_19068_n1172) );
  OR2X2 OR2X2_1240 ( .A(core__abc_21380_n3016), .B(core__abc_21380_n3012), .Y(core__abc_21380_n3017) );
  OR2X2 OR2X2_1241 ( .A(core__abc_21380_n1383), .B(core__abc_21380_n1402), .Y(core__abc_21380_n3018) );
  OR2X2 OR2X2_1242 ( .A(core__abc_21380_n1344), .B(core__abc_21380_n1364), .Y(core__abc_21380_n3019) );
  OR2X2 OR2X2_1243 ( .A(core__abc_21380_n3018), .B(core__abc_21380_n3019), .Y(core__abc_21380_n3020) );
  OR2X2 OR2X2_1244 ( .A(core__abc_21380_n1340), .B(core__abc_21380_n1360), .Y(core__abc_21380_n3024_1) );
  OR2X2 OR2X2_1245 ( .A(core__abc_21380_n3025), .B(core__abc_21380_n1363), .Y(core__abc_21380_n3026) );
  OR2X2 OR2X2_1246 ( .A(core__abc_21380_n3018), .B(core__abc_21380_n3026), .Y(core__abc_21380_n3027) );
  OR2X2 OR2X2_1247 ( .A(core__abc_21380_n3028), .B(core__abc_21380_n1398), .Y(core__abc_21380_n3029) );
  OR2X2 OR2X2_1248 ( .A(core__abc_21380_n3032), .B(core__abc_21380_n3040_1), .Y(core__abc_21380_n3041) );
  OR2X2 OR2X2_1249 ( .A(core__abc_21380_n3043), .B(core__abc_21380_n3042), .Y(core__abc_21380_n3044_1) );
  OR2X2 OR2X2_125 ( .A(_abc_19068_n1173_1), .B(_abc_19068_n1174_1), .Y(_abc_19068_n1175) );
  OR2X2 OR2X2_1250 ( .A(core__abc_21380_n3047), .B(core__abc_21380_n1469), .Y(core__abc_21380_n3048) );
  OR2X2 OR2X2_1251 ( .A(core__abc_21380_n3046), .B(core__abc_21380_n3048), .Y(core__abc_21380_n3049) );
  OR2X2 OR2X2_1252 ( .A(core__abc_21380_n1511), .B(core__abc_21380_n1489), .Y(core__abc_21380_n3051) );
  OR2X2 OR2X2_1253 ( .A(core__abc_21380_n3055_1), .B(core__abc_21380_n1543), .Y(core__abc_21380_n3056) );
  OR2X2 OR2X2_1254 ( .A(core__abc_21380_n3054), .B(core__abc_21380_n3056), .Y(core__abc_21380_n3057) );
  OR2X2 OR2X2_1255 ( .A(core__abc_21380_n3057), .B(core__abc_21380_n3050), .Y(core__abc_21380_n3058) );
  OR2X2 OR2X2_1256 ( .A(core__abc_21380_n3060), .B(core__abc_21380_n3076), .Y(core__abc_21380_n3077_1) );
  OR2X2 OR2X2_1257 ( .A(core__abc_21380_n3079), .B(core__abc_21380_n3078), .Y(core__abc_21380_n3080) );
  OR2X2 OR2X2_1258 ( .A(core__abc_21380_n3083), .B(core__abc_21380_n1615), .Y(core__abc_21380_n3084) );
  OR2X2 OR2X2_1259 ( .A(core__abc_21380_n3082), .B(core__abc_21380_n3084), .Y(core__abc_21380_n3085) );
  OR2X2 OR2X2_126 ( .A(_abc_19068_n1172), .B(_abc_19068_n1175), .Y(_abc_19068_n1176_1) );
  OR2X2 OR2X2_1260 ( .A(core__abc_21380_n1657), .B(core__abc_21380_n1635), .Y(core__abc_21380_n3087) );
  OR2X2 OR2X2_1261 ( .A(core__abc_21380_n3091_1), .B(core__abc_21380_n1689), .Y(core__abc_21380_n3092) );
  OR2X2 OR2X2_1262 ( .A(core__abc_21380_n3090), .B(core__abc_21380_n3092), .Y(core__abc_21380_n3093) );
  OR2X2 OR2X2_1263 ( .A(core__abc_21380_n3093), .B(core__abc_21380_n3086), .Y(core__abc_21380_n3094) );
  OR2X2 OR2X2_1264 ( .A(core__abc_21380_n1733), .B(core__abc_21380_n1709), .Y(core__abc_21380_n3096) );
  OR2X2 OR2X2_1265 ( .A(core__abc_21380_n3100), .B(core__abc_21380_n1764), .Y(core__abc_21380_n3101) );
  OR2X2 OR2X2_1266 ( .A(core__abc_21380_n3099), .B(core__abc_21380_n3101), .Y(core__abc_21380_n3102) );
  OR2X2 OR2X2_1267 ( .A(core__abc_21380_n3104_1), .B(core__abc_21380_n1840), .Y(core__abc_21380_n3105) );
  OR2X2 OR2X2_1268 ( .A(core__abc_21380_n3107), .B(core__abc_21380_n3106), .Y(core__abc_21380_n3108) );
  OR2X2 OR2X2_1269 ( .A(core__abc_21380_n3110_1), .B(core__abc_21380_n3105), .Y(core__abc_21380_n3111) );
  OR2X2 OR2X2_127 ( .A(_abc_19068_n1176_1), .B(_abc_19068_n1169), .Y(_abc_19068_n1177_1) );
  OR2X2 OR2X2_1270 ( .A(core__abc_21380_n3103), .B(core__abc_21380_n3111), .Y(core__abc_21380_n3112) );
  OR2X2 OR2X2_1271 ( .A(core__abc_21380_n3095_1), .B(core__abc_21380_n3112), .Y(core__abc_21380_n3113) );
  OR2X2 OR2X2_1272 ( .A(core__abc_21380_n3115), .B(core__abc_21380_n3123), .Y(core__abc_21380_n3124) );
  OR2X2 OR2X2_1273 ( .A(core__abc_21380_n3126), .B(core__abc_21380_n3125), .Y(core__abc_21380_n3127) );
  OR2X2 OR2X2_1274 ( .A(core__abc_21380_n3130), .B(core__abc_21380_n1914), .Y(core__abc_21380_n3131) );
  OR2X2 OR2X2_1275 ( .A(core__abc_21380_n3129), .B(core__abc_21380_n3131), .Y(core__abc_21380_n3132) );
  OR2X2 OR2X2_1276 ( .A(core__abc_21380_n1956), .B(core__abc_21380_n1933), .Y(core__abc_21380_n3134) );
  OR2X2 OR2X2_1277 ( .A(core__abc_21380_n3138), .B(core__abc_21380_n1990), .Y(core__abc_21380_n3139) );
  OR2X2 OR2X2_1278 ( .A(core__abc_21380_n3137), .B(core__abc_21380_n3139), .Y(core__abc_21380_n3140) );
  OR2X2 OR2X2_1279 ( .A(core__abc_21380_n3140), .B(core__abc_21380_n3133), .Y(core__abc_21380_n3141_1) );
  OR2X2 OR2X2_128 ( .A(_abc_19068_n1177_1), .B(_abc_19068_n1168_1), .Y(_abc_19068_n1178) );
  OR2X2 OR2X2_1280 ( .A(core__abc_21380_n3146), .B(core__abc_21380_n3010), .Y(core__abc_21380_n3147) );
  OR2X2 OR2X2_1281 ( .A(core__abc_21380_n3150), .B(core__abc_21380_n2070), .Y(core__abc_21380_n3153) );
  OR2X2 OR2X2_1282 ( .A(core__abc_21380_n3154), .B(core__abc_21380_n3007), .Y(core__abc_21380_n3155) );
  OR2X2 OR2X2_1283 ( .A(core__abc_21380_n3156), .B(core__abc_21380_n3151), .Y(core__abc_21380_n3157) );
  OR2X2 OR2X2_1284 ( .A(core__abc_21380_n3157), .B(core_v3_reg_27_), .Y(core__abc_21380_n3158) );
  OR2X2 OR2X2_1285 ( .A(core__abc_21380_n3168), .B(core__abc_21380_n1278_1), .Y(core__abc_21380_n3169) );
  OR2X2 OR2X2_1286 ( .A(core__abc_21380_n1302), .B(core__abc_21380_n1321), .Y(core__abc_21380_n3170) );
  OR2X2 OR2X2_1287 ( .A(core__abc_21380_n3174), .B(core__abc_21380_n1317), .Y(core__abc_21380_n3175) );
  OR2X2 OR2X2_1288 ( .A(core__abc_21380_n3172), .B(core__abc_21380_n3175), .Y(core__abc_21380_n3176) );
  OR2X2 OR2X2_1289 ( .A(core__abc_21380_n1337), .B(core__abc_21380_n1354), .Y(core__abc_21380_n3182) );
  OR2X2 OR2X2_129 ( .A(_abc_19068_n1181), .B(_abc_19068_n1182_1), .Y(_abc_19068_n1183_1) );
  OR2X2 OR2X2_1290 ( .A(core__abc_21380_n3186), .B(core__abc_21380_n1395), .Y(core__abc_21380_n3187) );
  OR2X2 OR2X2_1291 ( .A(core__abc_21380_n3184), .B(core__abc_21380_n3187), .Y(core__abc_21380_n3188) );
  OR2X2 OR2X2_1292 ( .A(core__abc_21380_n3180), .B(core__abc_21380_n3188), .Y(core__abc_21380_n3189) );
  OR2X2 OR2X2_1293 ( .A(core__abc_21380_n1486), .B(core__abc_21380_n1504), .Y(core__abc_21380_n3191) );
  OR2X2 OR2X2_1294 ( .A(core__abc_21380_n1411), .B(core__abc_21380_n1428), .Y(core__abc_21380_n3199) );
  OR2X2 OR2X2_1295 ( .A(core__abc_21380_n3202), .B(core__abc_21380_n1466), .Y(core__abc_21380_n3203) );
  OR2X2 OR2X2_1296 ( .A(core__abc_21380_n3201), .B(core__abc_21380_n3203), .Y(core__abc_21380_n3204) );
  OR2X2 OR2X2_1297 ( .A(core__abc_21380_n1482), .B(core__abc_21380_n1503), .Y(core__abc_21380_n3206) );
  OR2X2 OR2X2_1298 ( .A(core__abc_21380_n3207), .B(core__abc_21380_n1502), .Y(core__abc_21380_n3208) );
  OR2X2 OR2X2_1299 ( .A(core__abc_21380_n3211_1), .B(core__abc_21380_n1540), .Y(core__abc_21380_n3212) );
  OR2X2 OR2X2_13 ( .A(_abc_19068_n925_1), .B(_abc_19068_n927_1), .Y(_abc_19068_n928_1) );
  OR2X2 OR2X2_130 ( .A(_abc_19068_n1183_1), .B(_abc_19068_n1180_1), .Y(_abc_19068_n1184) );
  OR2X2 OR2X2_1300 ( .A(core__abc_21380_n3210), .B(core__abc_21380_n3212), .Y(core__abc_21380_n3213) );
  OR2X2 OR2X2_1301 ( .A(core__abc_21380_n3205), .B(core__abc_21380_n3213), .Y(core__abc_21380_n3214) );
  OR2X2 OR2X2_1302 ( .A(core__abc_21380_n3198), .B(core__abc_21380_n3214), .Y(core__abc_21380_n3215_1) );
  OR2X2 OR2X2_1303 ( .A(core__abc_21380_n1632), .B(core__abc_21380_n1650), .Y(core__abc_21380_n3224) );
  OR2X2 OR2X2_1304 ( .A(core__abc_21380_n1556), .B(core__abc_21380_n1574), .Y(core__abc_21380_n3233) );
  OR2X2 OR2X2_1305 ( .A(core__abc_21380_n3236_1), .B(core__abc_21380_n1611), .Y(core__abc_21380_n3237) );
  OR2X2 OR2X2_1306 ( .A(core__abc_21380_n3235), .B(core__abc_21380_n3237), .Y(core__abc_21380_n3238) );
  OR2X2 OR2X2_1307 ( .A(core__abc_21380_n1631), .B(core__abc_21380_n1649_1), .Y(core__abc_21380_n3240) );
  OR2X2 OR2X2_1308 ( .A(core__abc_21380_n3241), .B(core__abc_21380_n1648), .Y(core__abc_21380_n3242) );
  OR2X2 OR2X2_1309 ( .A(core__abc_21380_n3245_1), .B(core__abc_21380_n1686), .Y(core__abc_21380_n3246) );
  OR2X2 OR2X2_131 ( .A(_abc_19068_n1186_1), .B(_abc_19068_n1185_1), .Y(_abc_19068_n1187) );
  OR2X2 OR2X2_1310 ( .A(core__abc_21380_n3244), .B(core__abc_21380_n3246), .Y(core__abc_21380_n3247) );
  OR2X2 OR2X2_1311 ( .A(core__abc_21380_n3239), .B(core__abc_21380_n3247), .Y(core__abc_21380_n3248) );
  OR2X2 OR2X2_1312 ( .A(core__abc_21380_n3251_1), .B(core__abc_21380_n1722), .Y(core__abc_21380_n3252) );
  OR2X2 OR2X2_1313 ( .A(core__abc_21380_n3255), .B(core__abc_21380_n1761), .Y(core__abc_21380_n3256) );
  OR2X2 OR2X2_1314 ( .A(core__abc_21380_n3254), .B(core__abc_21380_n3256), .Y(core__abc_21380_n3257) );
  OR2X2 OR2X2_1315 ( .A(core__abc_21380_n3259), .B(core__abc_21380_n1837), .Y(core__abc_21380_n3260) );
  OR2X2 OR2X2_1316 ( .A(core__abc_21380_n3262_1), .B(core__abc_21380_n1797), .Y(core__abc_21380_n3263) );
  OR2X2 OR2X2_1317 ( .A(core__abc_21380_n3265), .B(core__abc_21380_n3260), .Y(core__abc_21380_n3266) );
  OR2X2 OR2X2_1318 ( .A(core__abc_21380_n3258), .B(core__abc_21380_n3266), .Y(core__abc_21380_n3267) );
  OR2X2 OR2X2_1319 ( .A(core__abc_21380_n3249), .B(core__abc_21380_n3267), .Y(core__abc_21380_n3268_1) );
  OR2X2 OR2X2_132 ( .A(_abc_19068_n1188_1), .B(_abc_19068_n1189_1), .Y(_abc_19068_n1190) );
  OR2X2 OR2X2_1320 ( .A(core__abc_21380_n3232), .B(core__abc_21380_n3268_1), .Y(core__abc_21380_n3269) );
  OR2X2 OR2X2_1321 ( .A(core__abc_21380_n1291), .B(core__abc_21380_n1261_1), .Y(core__abc_21380_n3271) );
  OR2X2 OR2X2_1322 ( .A(core__abc_21380_n3272), .B(core__abc_21380_n3170), .Y(core__abc_21380_n3273) );
  OR2X2 OR2X2_1323 ( .A(core__abc_21380_n3275), .B(core__abc_21380_n3276), .Y(core__abc_21380_n3277_1) );
  OR2X2 OR2X2_1324 ( .A(core__abc_21380_n3279), .B(core__abc_21380_n3280), .Y(core__abc_21380_n3281_1) );
  OR2X2 OR2X2_1325 ( .A(core__abc_21380_n3283), .B(core__abc_21380_n3284), .Y(core__abc_21380_n3285) );
  OR2X2 OR2X2_1326 ( .A(core__abc_21380_n3288), .B(core__abc_21380_n3270), .Y(core__abc_21380_n3289) );
  OR2X2 OR2X2_1327 ( .A(core__abc_21380_n1267), .B(core_v3_reg_48_), .Y(core__abc_21380_n3293) );
  OR2X2 OR2X2_1328 ( .A(core__abc_21380_n3296), .B(core__abc_21380_n3297), .Y(core__abc_21380_n3298) );
  OR2X2 OR2X2_1329 ( .A(core__abc_21380_n3159), .B(core__abc_21380_n3299), .Y(core__abc_21380_n3300) );
  OR2X2 OR2X2_133 ( .A(_abc_19068_n1190), .B(_abc_19068_n1187), .Y(_abc_19068_n1191_1) );
  OR2X2 OR2X2_1330 ( .A(core__abc_21380_n3301), .B(core__abc_21380_n3302), .Y(core__abc_21380_n3303) );
  OR2X2 OR2X2_1331 ( .A(core__abc_21380_n3303), .B(core__abc_21380_n3305), .Y(core__abc_21380_n3306) );
  OR2X2 OR2X2_1332 ( .A(core__abc_21380_n3308), .B(core__abc_21380_n3310), .Y(core__abc_21380_n3311) );
  OR2X2 OR2X2_1333 ( .A(core__abc_21380_n3167_1_bF_buf13), .B(core__abc_21380_n3313_bF_buf12), .Y(core__abc_21380_n3314) );
  OR2X2 OR2X2_1334 ( .A(core__abc_21380_n3316), .B(core__abc_21380_n3311), .Y(core__abc_21380_n3317) );
  OR2X2 OR2X2_1335 ( .A(core_v3_reg_0_), .B(core_mi_0_), .Y(core__abc_21380_n3320) );
  OR2X2 OR2X2_1336 ( .A(core__abc_21380_n3319), .B(core__abc_21380_n3324), .Y(core__abc_21380_n3325) );
  OR2X2 OR2X2_1337 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n3325), .Y(core__abc_21380_n3326) );
  OR2X2 OR2X2_1338 ( .A(core__abc_21380_n3307), .B(core__abc_21380_n3326), .Y(core__abc_21380_n3327) );
  OR2X2 OR2X2_1339 ( .A(core__abc_21380_n3328_bF_buf7), .B(core_v3_reg_0_), .Y(core__abc_21380_n3329) );
  OR2X2 OR2X2_134 ( .A(_abc_19068_n1192_1), .B(_abc_19068_n1193), .Y(_abc_19068_n1194_1) );
  OR2X2 OR2X2_1340 ( .A(core__abc_21380_n1876), .B(core__abc_21380_n1856), .Y(core__abc_21380_n3334) );
  OR2X2 OR2X2_1341 ( .A(core__abc_21380_n3270), .B(core__abc_21380_n3334), .Y(core__abc_21380_n3335) );
  OR2X2 OR2X2_1342 ( .A(core__abc_21380_n3013), .B(core__abc_21380_n3343), .Y(core__abc_21380_n3344) );
  OR2X2 OR2X2_1343 ( .A(core__abc_21380_n3345), .B(core__abc_21380_n3341), .Y(core__abc_21380_n3346) );
  OR2X2 OR2X2_1344 ( .A(core__abc_21380_n3344), .B(core_v3_reg_49_), .Y(core__abc_21380_n3347) );
  OR2X2 OR2X2_1345 ( .A(core__abc_21380_n3340), .B(core__abc_21380_n3349), .Y(core__abc_21380_n3352) );
  OR2X2 OR2X2_1346 ( .A(core__abc_21380_n3270), .B(core__abc_21380_n1856), .Y(core__abc_21380_n3357) );
  OR2X2 OR2X2_1347 ( .A(core__abc_21380_n3358), .B(core__abc_21380_n3356), .Y(core__abc_21380_n3359) );
  OR2X2 OR2X2_1348 ( .A(core__abc_21380_n3360), .B(core__abc_21380_n3350), .Y(core__abc_21380_n3361) );
  OR2X2 OR2X2_1349 ( .A(core__abc_21380_n3354), .B(core__abc_21380_n3362), .Y(core__abc_21380_n3363) );
  OR2X2 OR2X2_135 ( .A(_abc_19068_n1195_1), .B(_abc_19068_n1196), .Y(_abc_19068_n1197_1) );
  OR2X2 OR2X2_1350 ( .A(core__abc_21380_n3368), .B(core__abc_21380_n2065), .Y(core__abc_21380_n3369) );
  OR2X2 OR2X2_1351 ( .A(core__abc_21380_n3367), .B(core__abc_21380_n3369), .Y(core__abc_21380_n3370) );
  OR2X2 OR2X2_1352 ( .A(core__abc_21380_n3143), .B(core__abc_21380_n3373), .Y(core__abc_21380_n3374) );
  OR2X2 OR2X2_1353 ( .A(core__abc_21380_n3377), .B(core__abc_21380_n3378), .Y(core__abc_21380_n3379) );
  OR2X2 OR2X2_1354 ( .A(core__abc_21380_n3380), .B(core__abc_21380_n3365), .Y(core__abc_21380_n3381) );
  OR2X2 OR2X2_1355 ( .A(core__abc_21380_n3379), .B(core_v3_reg_28_), .Y(core__abc_21380_n3382) );
  OR2X2 OR2X2_1356 ( .A(core__abc_21380_n3384), .B(core__abc_21380_n3364), .Y(core__abc_21380_n3385) );
  OR2X2 OR2X2_1357 ( .A(core__abc_21380_n3383), .B(core__abc_21380_n3363), .Y(core__abc_21380_n3386) );
  OR2X2 OR2X2_1358 ( .A(core_v3_reg_1_), .B(core_mi_1_), .Y(core__abc_21380_n3391) );
  OR2X2 OR2X2_1359 ( .A(core__abc_21380_n3390), .B(core__abc_21380_n3395), .Y(core__abc_21380_n3396) );
  OR2X2 OR2X2_136 ( .A(_abc_19068_n1194_1), .B(_abc_19068_n1197_1), .Y(_abc_19068_n1198_1) );
  OR2X2 OR2X2_1360 ( .A(core__abc_21380_n3317_bF_buf5), .B(core__abc_21380_n3396), .Y(core__abc_21380_n3397) );
  OR2X2 OR2X2_1361 ( .A(core__abc_21380_n3388), .B(core__abc_21380_n3397), .Y(core__abc_21380_n3398) );
  OR2X2 OR2X2_1362 ( .A(core__abc_21380_n3328_bF_buf6), .B(core_v3_reg_1_), .Y(core__abc_21380_n3399) );
  OR2X2 OR2X2_1363 ( .A(core__abc_21380_n3361), .B(core__abc_21380_n3355), .Y(core__abc_21380_n3402) );
  OR2X2 OR2X2_1364 ( .A(core__abc_21380_n3332), .B(core__abc_21380_n1874), .Y(core__abc_21380_n3404) );
  OR2X2 OR2X2_1365 ( .A(core__abc_21380_n3337), .B(core__abc_21380_n3404), .Y(core__abc_21380_n3405) );
  OR2X2 OR2X2_1366 ( .A(core__abc_21380_n3407), .B(core__abc_21380_n3408), .Y(core__abc_21380_n3409) );
  OR2X2 OR2X2_1367 ( .A(core__abc_21380_n3414), .B(core__abc_21380_n3412), .Y(core__abc_21380_n3415) );
  OR2X2 OR2X2_1368 ( .A(core__abc_21380_n3416), .B(core__abc_21380_n3411), .Y(core__abc_21380_n3417) );
  OR2X2 OR2X2_1369 ( .A(core__abc_21380_n3415), .B(core_v3_reg_50_), .Y(core__abc_21380_n3418) );
  OR2X2 OR2X2_137 ( .A(_abc_19068_n1198_1), .B(_abc_19068_n1191_1), .Y(_abc_19068_n1199) );
  OR2X2 OR2X2_1370 ( .A(core__abc_21380_n3421), .B(core__abc_21380_n3422), .Y(core__abc_21380_n3423) );
  OR2X2 OR2X2_1371 ( .A(core__abc_21380_n3354), .B(core__abc_21380_n3350), .Y(core__abc_21380_n3425) );
  OR2X2 OR2X2_1372 ( .A(core__abc_21380_n3427), .B(core__abc_21380_n3424), .Y(core__abc_21380_n3428) );
  OR2X2 OR2X2_1373 ( .A(core__abc_21380_n3377), .B(core__abc_21380_n2083), .Y(core__abc_21380_n3430) );
  OR2X2 OR2X2_1374 ( .A(core__abc_21380_n3432), .B(core__abc_21380_n3433), .Y(core__abc_21380_n3434) );
  OR2X2 OR2X2_1375 ( .A(core__abc_21380_n3437), .B(core__abc_21380_n3435), .Y(core__abc_21380_n3438) );
  OR2X2 OR2X2_1376 ( .A(core__abc_21380_n3438), .B(core__abc_21380_n3428), .Y(core__abc_21380_n3439) );
  OR2X2 OR2X2_1377 ( .A(core__abc_21380_n3434), .B(core__abc_21380_n3429), .Y(core__abc_21380_n3442) );
  OR2X2 OR2X2_1378 ( .A(core__abc_21380_n3443), .B(core__abc_21380_n3440), .Y(core__abc_21380_n3444) );
  OR2X2 OR2X2_1379 ( .A(core_v3_reg_2_), .B(core_mi_2_), .Y(core__abc_21380_n3448) );
  OR2X2 OR2X2_138 ( .A(_abc_19068_n1199), .B(_abc_19068_n1184), .Y(_abc_19068_n1200_1) );
  OR2X2 OR2X2_1380 ( .A(core__abc_21380_n3447), .B(core__abc_21380_n3452), .Y(core__abc_21380_n3453) );
  OR2X2 OR2X2_1381 ( .A(core__abc_21380_n3317_bF_buf4), .B(core__abc_21380_n3453), .Y(core__abc_21380_n3454) );
  OR2X2 OR2X2_1382 ( .A(core__abc_21380_n3446), .B(core__abc_21380_n3454), .Y(core__abc_21380_n3455) );
  OR2X2 OR2X2_1383 ( .A(core__abc_21380_n3328_bF_buf5), .B(core_v3_reg_2_), .Y(core__abc_21380_n3456) );
  OR2X2 OR2X2_1384 ( .A(core__abc_21380_n3408), .B(core__abc_21380_n1892), .Y(core__abc_21380_n3459) );
  OR2X2 OR2X2_1385 ( .A(core__abc_21380_n3461), .B(core__abc_21380_n3462), .Y(core__abc_21380_n3463) );
  OR2X2 OR2X2_1386 ( .A(core__abc_21380_n3468), .B(core__abc_21380_n3469), .Y(core__abc_21380_n3470) );
  OR2X2 OR2X2_1387 ( .A(core__abc_21380_n3471), .B(core_v3_reg_51_), .Y(core__abc_21380_n3472) );
  OR2X2 OR2X2_1388 ( .A(core__abc_21380_n3470), .B(core__abc_21380_n3473), .Y(core__abc_21380_n3474) );
  OR2X2 OR2X2_1389 ( .A(core__abc_21380_n3463), .B(core__abc_21380_n3475), .Y(core__abc_21380_n3476) );
  OR2X2 OR2X2_139 ( .A(_abc_19068_n1202), .B(_abc_19068_n1203_1), .Y(_abc_19068_n1204_1) );
  OR2X2 OR2X2_1390 ( .A(core__abc_21380_n3477), .B(core__abc_21380_n3478), .Y(core__abc_21380_n3479) );
  OR2X2 OR2X2_1391 ( .A(core__abc_21380_n3403), .B(core__abc_21380_n3423), .Y(core__abc_21380_n3483_1) );
  OR2X2 OR2X2_1392 ( .A(core__abc_21380_n3484), .B(core__abc_21380_n3481), .Y(core__abc_21380_n3486) );
  OR2X2 OR2X2_1393 ( .A(core__abc_21380_n3487), .B(core__abc_21380_n3485_1), .Y(core__abc_21380_n3488) );
  OR2X2 OR2X2_1394 ( .A(core__abc_21380_n3375), .B(core__abc_21380_n3491), .Y(core__abc_21380_n3492) );
  OR2X2 OR2X2_1395 ( .A(core__abc_21380_n3494), .B(core__abc_21380_n3493), .Y(core__abc_21380_n3495) );
  OR2X2 OR2X2_1396 ( .A(core__abc_21380_n3499), .B(core__abc_21380_n3497), .Y(core__abc_21380_n3500) );
  OR2X2 OR2X2_1397 ( .A(core__abc_21380_n3501_1), .B(core_v3_reg_30_), .Y(core__abc_21380_n3502) );
  OR2X2 OR2X2_1398 ( .A(core__abc_21380_n3500), .B(core__abc_21380_n3503), .Y(core__abc_21380_n3504) );
  OR2X2 OR2X2_1399 ( .A(core__abc_21380_n3489), .B(core__abc_21380_n3505_1), .Y(core__abc_21380_n3506) );
  OR2X2 OR2X2_14 ( .A(_abc_19068_n929), .B(_abc_19068_n930_1), .Y(_abc_19068_n931_1) );
  OR2X2 OR2X2_140 ( .A(_abc_19068_n1205), .B(_abc_19068_n1206_1), .Y(_abc_19068_n1207_1) );
  OR2X2 OR2X2_1400 ( .A(core__abc_21380_n3507), .B(core__abc_21380_n3488), .Y(core__abc_21380_n3508) );
  OR2X2 OR2X2_1401 ( .A(core_v3_reg_3_), .B(core_mi_3_), .Y(core__abc_21380_n3512) );
  OR2X2 OR2X2_1402 ( .A(core__abc_21380_n3511), .B(core__abc_21380_n3516), .Y(core__abc_21380_n3517) );
  OR2X2 OR2X2_1403 ( .A(core__abc_21380_n3317_bF_buf3), .B(core__abc_21380_n3517), .Y(core__abc_21380_n3518_1) );
  OR2X2 OR2X2_1404 ( .A(core__abc_21380_n3510), .B(core__abc_21380_n3518_1), .Y(core__abc_21380_n3519) );
  OR2X2 OR2X2_1405 ( .A(core__abc_21380_n3328_bF_buf4), .B(core_v3_reg_3_), .Y(core__abc_21380_n3520) );
  OR2X2 OR2X2_1406 ( .A(core__abc_21380_n3525), .B(core__abc_21380_n1911), .Y(core__abc_21380_n3526) );
  OR2X2 OR2X2_1407 ( .A(core__abc_21380_n3524), .B(core__abc_21380_n3526), .Y(core__abc_21380_n3527) );
  OR2X2 OR2X2_1408 ( .A(core__abc_21380_n3529), .B(core__abc_21380_n3527), .Y(core__abc_21380_n3530) );
  OR2X2 OR2X2_1409 ( .A(core__abc_21380_n3287), .B(core__abc_21380_n3533), .Y(core__abc_21380_n3534) );
  OR2X2 OR2X2_141 ( .A(_abc_19068_n1204_1), .B(_abc_19068_n1207_1), .Y(_abc_19068_n1208) );
  OR2X2 OR2X2_1410 ( .A(core__abc_21380_n3536), .B(core__abc_21380_n3531_1), .Y(core__abc_21380_n3537) );
  OR2X2 OR2X2_1411 ( .A(core__abc_21380_n3542), .B(core__abc_21380_n3540), .Y(core__abc_21380_n3543) );
  OR2X2 OR2X2_1412 ( .A(core__abc_21380_n3546), .B(core__abc_21380_n3544), .Y(core__abc_21380_n3547) );
  OR2X2 OR2X2_1413 ( .A(core__abc_21380_n3549), .B(core__abc_21380_n3550), .Y(core__abc_21380_n3551) );
  OR2X2 OR2X2_1414 ( .A(core__abc_21380_n3427), .B(core__abc_21380_n3554), .Y(core__abc_21380_n3555) );
  OR2X2 OR2X2_1415 ( .A(core__abc_21380_n3559), .B(core__abc_21380_n3558), .Y(core__abc_21380_n3560) );
  OR2X2 OR2X2_1416 ( .A(core__abc_21380_n3557), .B(core__abc_21380_n3561_1), .Y(core__abc_21380_n3562) );
  OR2X2 OR2X2_1417 ( .A(core__abc_21380_n3496), .B(core__abc_21380_n2126), .Y(core__abc_21380_n3564) );
  OR2X2 OR2X2_1418 ( .A(core__abc_21380_n3568), .B(core__abc_21380_n3566), .Y(core__abc_21380_n3569_1) );
  OR2X2 OR2X2_1419 ( .A(core__abc_21380_n3565), .B(core__abc_21380_n2146), .Y(core__abc_21380_n3573) );
  OR2X2 OR2X2_142 ( .A(_abc_19068_n906_1), .B(_abc_19068_n1038_1), .Y(_abc_19068_n1209_1) );
  OR2X2 OR2X2_1420 ( .A(core__abc_21380_n3570), .B(core__abc_21380_n3575), .Y(core__abc_21380_n3576) );
  OR2X2 OR2X2_1421 ( .A(core__abc_21380_n3563), .B(core__abc_21380_n3576), .Y(core__abc_21380_n3577) );
  OR2X2 OR2X2_1422 ( .A(core__abc_21380_n3574), .B(core__abc_21380_n3571), .Y(core__abc_21380_n3578) );
  OR2X2 OR2X2_1423 ( .A(core__abc_21380_n3569_1), .B(core_v3_reg_31_), .Y(core__abc_21380_n3579) );
  OR2X2 OR2X2_1424 ( .A(core__abc_21380_n3580), .B(core__abc_21380_n3562), .Y(core__abc_21380_n3581_1) );
  OR2X2 OR2X2_1425 ( .A(core_v3_reg_4_), .B(core_mi_4_), .Y(core__abc_21380_n3586) );
  OR2X2 OR2X2_1426 ( .A(core__abc_21380_n3585), .B(core__abc_21380_n3590), .Y(core__abc_21380_n3591) );
  OR2X2 OR2X2_1427 ( .A(core__abc_21380_n3317_bF_buf2), .B(core__abc_21380_n3591), .Y(core__abc_21380_n3592) );
  OR2X2 OR2X2_1428 ( .A(core__abc_21380_n3583), .B(core__abc_21380_n3592), .Y(core__abc_21380_n3593) );
  OR2X2 OR2X2_1429 ( .A(core__abc_21380_n3328_bF_buf3), .B(core_v3_reg_4_), .Y(core__abc_21380_n3594) );
  OR2X2 OR2X2_143 ( .A(_abc_19068_n1210_1), .B(_abc_19068_n1211), .Y(_abc_19068_n1212_1) );
  OR2X2 OR2X2_1430 ( .A(core__abc_21380_n3557), .B(core__abc_21380_n3549), .Y(core__abc_21380_n3597) );
  OR2X2 OR2X2_1431 ( .A(core__abc_21380_n3531_1), .B(core__abc_21380_n1927), .Y(core__abc_21380_n3599) );
  OR2X2 OR2X2_1432 ( .A(core__abc_21380_n3601), .B(core__abc_21380_n3602), .Y(core__abc_21380_n3603) );
  OR2X2 OR2X2_1433 ( .A(core__abc_21380_n3540), .B(core__abc_21380_n1340), .Y(core__abc_21380_n3606) );
  OR2X2 OR2X2_1434 ( .A(core__abc_21380_n3608), .B(core__abc_21380_n3609), .Y(core__abc_21380_n3610) );
  OR2X2 OR2X2_1435 ( .A(core__abc_21380_n3613), .B(core__abc_21380_n3611), .Y(core__abc_21380_n3614) );
  OR2X2 OR2X2_1436 ( .A(core__abc_21380_n3616), .B(core__abc_21380_n3617), .Y(core__abc_21380_n3618) );
  OR2X2 OR2X2_1437 ( .A(core__abc_21380_n3619_1), .B(core__abc_21380_n3621), .Y(core__abc_21380_n3622) );
  OR2X2 OR2X2_1438 ( .A(core__abc_21380_n3630), .B(core__abc_21380_n2142), .Y(core__abc_21380_n3631_1) );
  OR2X2 OR2X2_1439 ( .A(core__abc_21380_n3629), .B(core__abc_21380_n3631_1), .Y(core__abc_21380_n3632) );
  OR2X2 OR2X2_144 ( .A(_abc_19068_n1212_1), .B(_abc_19068_n1209_1), .Y(_abc_19068_n1213_1) );
  OR2X2 OR2X2_1440 ( .A(core__abc_21380_n3627), .B(core__abc_21380_n3632), .Y(core__abc_21380_n3633) );
  OR2X2 OR2X2_1441 ( .A(core__abc_21380_n3635), .B(core__abc_21380_n3633), .Y(core__abc_21380_n3636_1) );
  OR2X2 OR2X2_1442 ( .A(core__abc_21380_n3374), .B(core__abc_21380_n3639), .Y(core__abc_21380_n3640) );
  OR2X2 OR2X2_1443 ( .A(core__abc_21380_n3637), .B(core__abc_21380_n3642), .Y(core__abc_21380_n3643) );
  OR2X2 OR2X2_1444 ( .A(core__abc_21380_n3644), .B(core__abc_21380_n3624), .Y(core__abc_21380_n3645) );
  OR2X2 OR2X2_1445 ( .A(core__abc_21380_n3643), .B(core_v3_reg_32_), .Y(core__abc_21380_n3646) );
  OR2X2 OR2X2_1446 ( .A(core__abc_21380_n3623_1), .B(core__abc_21380_n3648), .Y(core__abc_21380_n3649) );
  OR2X2 OR2X2_1447 ( .A(core__abc_21380_n3622), .B(core__abc_21380_n3647_1), .Y(core__abc_21380_n3650) );
  OR2X2 OR2X2_1448 ( .A(core_v3_reg_5_), .B(core_mi_5_), .Y(core__abc_21380_n3655) );
  OR2X2 OR2X2_1449 ( .A(core__abc_21380_n3654), .B(core__abc_21380_n3659_1), .Y(core__abc_21380_n3660) );
  OR2X2 OR2X2_145 ( .A(_abc_19068_n1214), .B(_abc_19068_n1215_1), .Y(_abc_19068_n1216_1) );
  OR2X2 OR2X2_1450 ( .A(core__abc_21380_n3317_bF_buf1), .B(core__abc_21380_n3660), .Y(core__abc_21380_n3661) );
  OR2X2 OR2X2_1451 ( .A(core__abc_21380_n3652), .B(core__abc_21380_n3661), .Y(core__abc_21380_n3662) );
  OR2X2 OR2X2_1452 ( .A(core__abc_21380_n3328_bF_buf2), .B(core_v3_reg_5_), .Y(core__abc_21380_n3663_1) );
  OR2X2 OR2X2_1453 ( .A(core__abc_21380_n3618), .B(core__abc_21380_n3551), .Y(core__abc_21380_n3666) );
  OR2X2 OR2X2_1454 ( .A(core__abc_21380_n3560), .B(core__abc_21380_n3666), .Y(core__abc_21380_n3667) );
  OR2X2 OR2X2_1455 ( .A(core__abc_21380_n3616), .B(core__abc_21380_n3549), .Y(core__abc_21380_n3669) );
  OR2X2 OR2X2_1456 ( .A(core__abc_21380_n3535_1), .B(core__abc_21380_n3675), .Y(core__abc_21380_n3676_1) );
  OR2X2 OR2X2_1457 ( .A(core__abc_21380_n3678), .B(core__abc_21380_n1949), .Y(core__abc_21380_n3679) );
  OR2X2 OR2X2_1458 ( .A(core__abc_21380_n3682), .B(core__abc_21380_n3683), .Y(core__abc_21380_n3684) );
  OR2X2 OR2X2_1459 ( .A(core__abc_21380_n3681_1), .B(core__abc_21380_n3685), .Y(core__abc_21380_n3686) );
  OR2X2 OR2X2_146 ( .A(_abc_19068_n1217), .B(_abc_19068_n1218_1), .Y(_abc_19068_n1219_1) );
  OR2X2 OR2X2_1460 ( .A(core__abc_21380_n3541), .B(core__abc_21380_n3019), .Y(core__abc_21380_n3688_1) );
  OR2X2 OR2X2_1461 ( .A(core__abc_21380_n3689), .B(core__abc_21380_n1383), .Y(core__abc_21380_n3691) );
  OR2X2 OR2X2_1462 ( .A(core__abc_21380_n3692), .B(core__abc_21380_n3690), .Y(core__abc_21380_n3693_1) );
  OR2X2 OR2X2_1463 ( .A(core__abc_21380_n3694), .B(core__abc_21380_n3687), .Y(core__abc_21380_n3695) );
  OR2X2 OR2X2_1464 ( .A(core__abc_21380_n3693_1), .B(core_v3_reg_54_), .Y(core__abc_21380_n3696) );
  OR2X2 OR2X2_1465 ( .A(core__abc_21380_n3686), .B(core__abc_21380_n3697), .Y(core__abc_21380_n3698) );
  OR2X2 OR2X2_1466 ( .A(core__abc_21380_n3699), .B(core__abc_21380_n3700), .Y(core__abc_21380_n3701) );
  OR2X2 OR2X2_1467 ( .A(core__abc_21380_n3703_1), .B(core__abc_21380_n3704), .Y(core__abc_21380_n3705) );
  OR2X2 OR2X2_1468 ( .A(core__abc_21380_n3713), .B(core__abc_21380_n3711), .Y(core__abc_21380_n3714) );
  OR2X2 OR2X2_1469 ( .A(core__abc_21380_n3710), .B(core__abc_21380_n3714), .Y(core__abc_21380_n3715) );
  OR2X2 OR2X2_147 ( .A(_abc_19068_n1216_1), .B(_abc_19068_n1219_1), .Y(_abc_19068_n1220) );
  OR2X2 OR2X2_1470 ( .A(core__abc_21380_n3718), .B(core__abc_21380_n3716_1), .Y(core__abc_21380_n3719) );
  OR2X2 OR2X2_1471 ( .A(core__abc_21380_n3706), .B(core__abc_21380_n3720_1), .Y(core__abc_21380_n3721) );
  OR2X2 OR2X2_1472 ( .A(core__abc_21380_n3705), .B(core__abc_21380_n3719), .Y(core__abc_21380_n3722) );
  OR2X2 OR2X2_1473 ( .A(core_v3_reg_6_), .B(core_mi_6_), .Y(core__abc_21380_n3727) );
  OR2X2 OR2X2_1474 ( .A(core__abc_21380_n3726), .B(core__abc_21380_n3731), .Y(core__abc_21380_n3732) );
  OR2X2 OR2X2_1475 ( .A(core__abc_21380_n3317_bF_buf0), .B(core__abc_21380_n3732), .Y(core__abc_21380_n3733) );
  OR2X2 OR2X2_1476 ( .A(core__abc_21380_n3724), .B(core__abc_21380_n3733), .Y(core__abc_21380_n3734) );
  OR2X2 OR2X2_1477 ( .A(core__abc_21380_n3328_bF_buf1), .B(core_v3_reg_6_), .Y(core__abc_21380_n3735) );
  OR2X2 OR2X2_1478 ( .A(core__abc_21380_n3703_1), .B(core__abc_21380_n3699), .Y(core__abc_21380_n3738) );
  OR2X2 OR2X2_1479 ( .A(core__abc_21380_n3680), .B(core__abc_21380_n1969), .Y(core__abc_21380_n3741) );
  OR2X2 OR2X2_148 ( .A(_abc_19068_n1220), .B(_abc_19068_n1213_1), .Y(_abc_19068_n1221_1) );
  OR2X2 OR2X2_1480 ( .A(core__abc_21380_n3685), .B(core__abc_21380_n1968), .Y(core__abc_21380_n3744) );
  OR2X2 OR2X2_1481 ( .A(core__abc_21380_n3743), .B(core__abc_21380_n3745_1), .Y(core__abc_21380_n3746) );
  OR2X2 OR2X2_1482 ( .A(core__abc_21380_n3692), .B(core__abc_21380_n1379), .Y(core__abc_21380_n3748) );
  OR2X2 OR2X2_1483 ( .A(core__abc_21380_n3750), .B(core__abc_21380_n3751), .Y(core__abc_21380_n3752_1) );
  OR2X2 OR2X2_1484 ( .A(core__abc_21380_n3755), .B(core__abc_21380_n3753), .Y(core__abc_21380_n3756_1) );
  OR2X2 OR2X2_1485 ( .A(core__abc_21380_n3746), .B(core__abc_21380_n3756_1), .Y(core__abc_21380_n3757) );
  OR2X2 OR2X2_1486 ( .A(core__abc_21380_n3744), .B(core__abc_21380_n1989), .Y(core__abc_21380_n3758) );
  OR2X2 OR2X2_1487 ( .A(core__abc_21380_n3742), .B(core__abc_21380_n1995_1), .Y(core__abc_21380_n3759) );
  OR2X2 OR2X2_1488 ( .A(core__abc_21380_n3760), .B(core__abc_21380_n3761), .Y(core__abc_21380_n3762) );
  OR2X2 OR2X2_1489 ( .A(core__abc_21380_n3765), .B(core__abc_21380_n3766), .Y(core__abc_21380_n3767_1) );
  OR2X2 OR2X2_149 ( .A(_abc_19068_n1221_1), .B(_abc_19068_n1208), .Y(_abc_19068_n1222_1) );
  OR2X2 OR2X2_1490 ( .A(core__abc_21380_n3711), .B(core__abc_21380_n2177), .Y(core__abc_21380_n3770) );
  OR2X2 OR2X2_1491 ( .A(core__abc_21380_n3713), .B(core__abc_21380_n3770), .Y(core__abc_21380_n3771) );
  OR2X2 OR2X2_1492 ( .A(core__abc_21380_n3771), .B(core__abc_21380_n2197), .Y(core__abc_21380_n3774) );
  OR2X2 OR2X2_1493 ( .A(core__abc_21380_n3775), .B(core__abc_21380_n3769), .Y(core__abc_21380_n3776) );
  OR2X2 OR2X2_1494 ( .A(core__abc_21380_n3777), .B(core_v3_reg_34_), .Y(core__abc_21380_n3778) );
  OR2X2 OR2X2_1495 ( .A(core__abc_21380_n3768), .B(core__abc_21380_n3780), .Y(core__abc_21380_n3781) );
  OR2X2 OR2X2_1496 ( .A(core__abc_21380_n3767_1), .B(core__abc_21380_n3779_1), .Y(core__abc_21380_n3782) );
  OR2X2 OR2X2_1497 ( .A(core_v3_reg_7_), .B(core_mi_7_), .Y(core__abc_21380_n3786) );
  OR2X2 OR2X2_1498 ( .A(core__abc_21380_n3785), .B(core__abc_21380_n3790), .Y(core__abc_21380_n3791) );
  OR2X2 OR2X2_1499 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n3791), .Y(core__abc_21380_n3792) );
  OR2X2 OR2X2_15 ( .A(_abc_19068_n928_1), .B(_abc_19068_n931_1), .Y(_abc_19068_n932) );
  OR2X2 OR2X2_150 ( .A(_abc_19068_n1225_1), .B(_abc_19068_n1226), .Y(_abc_19068_n1227_1) );
  OR2X2 OR2X2_1500 ( .A(core__abc_21380_n3784), .B(core__abc_21380_n3792), .Y(core__abc_21380_n3793) );
  OR2X2 OR2X2_1501 ( .A(core__abc_21380_n3328_bF_buf0), .B(core_v3_reg_7_), .Y(core__abc_21380_n3794) );
  OR2X2 OR2X2_1502 ( .A(core__abc_21380_n3801_1), .B(core__abc_21380_n1987), .Y(core__abc_21380_n3802) );
  OR2X2 OR2X2_1503 ( .A(core__abc_21380_n3800), .B(core__abc_21380_n3802), .Y(core__abc_21380_n3803) );
  OR2X2 OR2X2_1504 ( .A(core__abc_21380_n3799), .B(core__abc_21380_n3803), .Y(core__abc_21380_n3804) );
  OR2X2 OR2X2_1505 ( .A(core__abc_21380_n3806), .B(core__abc_21380_n3804), .Y(core__abc_21380_n3807) );
  OR2X2 OR2X2_1506 ( .A(core__abc_21380_n3287), .B(core__abc_21380_n3810), .Y(core__abc_21380_n3811) );
  OR2X2 OR2X2_1507 ( .A(core__abc_21380_n3813), .B(core__abc_21380_n3808), .Y(core__abc_21380_n3814_1) );
  OR2X2 OR2X2_1508 ( .A(core__abc_21380_n3819), .B(core__abc_21380_n3817), .Y(core__abc_21380_n3820) );
  OR2X2 OR2X2_1509 ( .A(core__abc_21380_n3821), .B(core__abc_21380_n3816), .Y(core__abc_21380_n3822) );
  OR2X2 OR2X2_151 ( .A(_abc_19068_n1228_1), .B(_abc_19068_n1229), .Y(_abc_19068_n1230_1) );
  OR2X2 OR2X2_1510 ( .A(core__abc_21380_n3820), .B(core_v3_reg_56_), .Y(core__abc_21380_n3823_1) );
  OR2X2 OR2X2_1511 ( .A(core__abc_21380_n3826), .B(core__abc_21380_n3827), .Y(core__abc_21380_n3828_1) );
  OR2X2 OR2X2_1512 ( .A(core__abc_21380_n3829), .B(core__abc_21380_n3698), .Y(core__abc_21380_n3830) );
  OR2X2 OR2X2_1513 ( .A(core__abc_21380_n3834_1), .B(core__abc_21380_n3829), .Y(core__abc_21380_n3835) );
  OR2X2 OR2X2_1514 ( .A(core__abc_21380_n3833), .B(core__abc_21380_n3835), .Y(core__abc_21380_n3836) );
  OR2X2 OR2X2_1515 ( .A(core__abc_21380_n3841), .B(core__abc_21380_n3839), .Y(core__abc_21380_n3842) );
  OR2X2 OR2X2_1516 ( .A(core__abc_21380_n3842), .B(core__abc_21380_n3845), .Y(core__abc_21380_n3846) );
  OR2X2 OR2X2_1517 ( .A(core__abc_21380_n3847), .B(core__abc_21380_n3837), .Y(core__abc_21380_n3848) );
  OR2X2 OR2X2_1518 ( .A(core__abc_21380_n3851), .B(core__abc_21380_n2220), .Y(core__abc_21380_n3854) );
  OR2X2 OR2X2_1519 ( .A(core__abc_21380_n3855), .B(core__abc_21380_n3850), .Y(core__abc_21380_n3856) );
  OR2X2 OR2X2_152 ( .A(_abc_19068_n1227_1), .B(_abc_19068_n1230_1), .Y(_abc_19068_n1231) );
  OR2X2 OR2X2_1520 ( .A(core__abc_21380_n3857_1), .B(core__abc_21380_n3858), .Y(core__abc_21380_n3859) );
  OR2X2 OR2X2_1521 ( .A(core__abc_21380_n3849), .B(core__abc_21380_n3859), .Y(core__abc_21380_n3860) );
  OR2X2 OR2X2_1522 ( .A(core__abc_21380_n3848), .B(core__abc_21380_n3862), .Y(core__abc_21380_n3863) );
  OR2X2 OR2X2_1523 ( .A(core_v3_reg_8_), .B(core_mi_8_), .Y(core__abc_21380_n3868) );
  OR2X2 OR2X2_1524 ( .A(core__abc_21380_n3867), .B(core__abc_21380_n3872), .Y(core__abc_21380_n3873) );
  OR2X2 OR2X2_1525 ( .A(core__abc_21380_n3317_bF_buf6), .B(core__abc_21380_n3873), .Y(core__abc_21380_n3874) );
  OR2X2 OR2X2_1526 ( .A(core__abc_21380_n3865), .B(core__abc_21380_n3874), .Y(core__abc_21380_n3875) );
  OR2X2 OR2X2_1527 ( .A(core__abc_21380_n3328_bF_buf7), .B(core_v3_reg_8_), .Y(core__abc_21380_n3876) );
  OR2X2 OR2X2_1528 ( .A(core__abc_21380_n3808), .B(core__abc_21380_n2003), .Y(core__abc_21380_n3884) );
  OR2X2 OR2X2_1529 ( .A(core__abc_21380_n3886_1), .B(core__abc_21380_n3888), .Y(core__abc_21380_n3889) );
  OR2X2 OR2X2_153 ( .A(_abc_19068_n1231), .B(_abc_19068_n1224_1), .Y(_abc_19068_n1232) );
  OR2X2 OR2X2_1530 ( .A(core__abc_21380_n3889), .B(core__abc_21380_n3883), .Y(core__abc_21380_n3890) );
  OR2X2 OR2X2_1531 ( .A(core__abc_21380_n3819), .B(core__abc_21380_n1415), .Y(core__abc_21380_n3892) );
  OR2X2 OR2X2_1532 ( .A(core__abc_21380_n3894), .B(core__abc_21380_n3895), .Y(core__abc_21380_n3896) );
  OR2X2 OR2X2_1533 ( .A(core__abc_21380_n3899), .B(core__abc_21380_n3897), .Y(core__abc_21380_n3900) );
  OR2X2 OR2X2_1534 ( .A(core__abc_21380_n3890), .B(core__abc_21380_n3900), .Y(core__abc_21380_n3901) );
  OR2X2 OR2X2_1535 ( .A(core__abc_21380_n3906), .B(core__abc_21380_n3907), .Y(core__abc_21380_n3908) );
  OR2X2 OR2X2_1536 ( .A(core__abc_21380_n3641), .B(core__abc_21380_n3912), .Y(core__abc_21380_n3913) );
  OR2X2 OR2X2_1537 ( .A(core__abc_21380_n3915), .B(core__abc_21380_n2216), .Y(core__abc_21380_n3916) );
  OR2X2 OR2X2_1538 ( .A(core__abc_21380_n3914_1), .B(core__abc_21380_n3916), .Y(core__abc_21380_n3917) );
  OR2X2 OR2X2_1539 ( .A(core__abc_21380_n3921), .B(core__abc_21380_n3922_1), .Y(core__abc_21380_n3923) );
  OR2X2 OR2X2_154 ( .A(_abc_19068_n1233_1), .B(_abc_19068_n1234), .Y(_abc_19068_n1235_1) );
  OR2X2 OR2X2_1540 ( .A(core__abc_21380_n3924), .B(core__abc_21380_n3909), .Y(core__abc_21380_n3925) );
  OR2X2 OR2X2_1541 ( .A(core__abc_21380_n3923), .B(core_v3_reg_36_), .Y(core__abc_21380_n3926) );
  OR2X2 OR2X2_1542 ( .A(core__abc_21380_n3908), .B(core__abc_21380_n3928), .Y(core__abc_21380_n3929) );
  OR2X2 OR2X2_1543 ( .A(core__abc_21380_n3930), .B(core__abc_21380_n3927_1), .Y(core__abc_21380_n3931) );
  OR2X2 OR2X2_1544 ( .A(core_v3_reg_9_), .B(core_mi_9_), .Y(core__abc_21380_n3935) );
  OR2X2 OR2X2_1545 ( .A(core__abc_21380_n3934), .B(core__abc_21380_n3939), .Y(core__abc_21380_n3940) );
  OR2X2 OR2X2_1546 ( .A(core__abc_21380_n3317_bF_buf5), .B(core__abc_21380_n3940), .Y(core__abc_21380_n3941) );
  OR2X2 OR2X2_1547 ( .A(core__abc_21380_n3933), .B(core__abc_21380_n3941), .Y(core__abc_21380_n3942_1) );
  OR2X2 OR2X2_1548 ( .A(core__abc_21380_n3328_bF_buf6), .B(core_v3_reg_9_), .Y(core__abc_21380_n3943) );
  OR2X2 OR2X2_1549 ( .A(core__abc_21380_n3883), .B(core__abc_21380_n2021), .Y(core__abc_21380_n3946) );
  OR2X2 OR2X2_155 ( .A(_abc_19068_n1235_1), .B(_abc_19068_n1236), .Y(_abc_19068_n1237_1) );
  OR2X2 OR2X2_1550 ( .A(core__abc_21380_n3888), .B(core__abc_21380_n3946), .Y(core__abc_21380_n3947) );
  OR2X2 OR2X2_1551 ( .A(core__abc_21380_n3950), .B(core__abc_21380_n3948_1), .Y(core__abc_21380_n3951) );
  OR2X2 OR2X2_1552 ( .A(core__abc_21380_n3956), .B(core__abc_21380_n1458), .Y(core__abc_21380_n3958) );
  OR2X2 OR2X2_1553 ( .A(core__abc_21380_n3959), .B(core__abc_21380_n3957), .Y(core__abc_21380_n3960) );
  OR2X2 OR2X2_1554 ( .A(core__abc_21380_n3961_1), .B(core__abc_21380_n3953), .Y(core__abc_21380_n3962) );
  OR2X2 OR2X2_1555 ( .A(core__abc_21380_n3960), .B(core_v3_reg_58_), .Y(core__abc_21380_n3963) );
  OR2X2 OR2X2_1556 ( .A(core__abc_21380_n3966), .B(core__abc_21380_n3967), .Y(core__abc_21380_n3968) );
  OR2X2 OR2X2_1557 ( .A(core__abc_21380_n3971), .B(core__abc_21380_n3902), .Y(core__abc_21380_n3972) );
  OR2X2 OR2X2_1558 ( .A(core__abc_21380_n3974_1), .B(core__abc_21380_n3975), .Y(core__abc_21380_n3976) );
  OR2X2 OR2X2_1559 ( .A(core__abc_21380_n3921), .B(core__abc_21380_n2232), .Y(core__abc_21380_n3979_1) );
  OR2X2 OR2X2_156 ( .A(_abc_19068_n1238), .B(_abc_19068_n1239_1), .Y(_abc_19068_n1240) );
  OR2X2 OR2X2_1560 ( .A(core__abc_21380_n3981), .B(core__abc_21380_n3982_1), .Y(core__abc_21380_n3983) );
  OR2X2 OR2X2_1561 ( .A(core__abc_21380_n3986_1), .B(core__abc_21380_n3984), .Y(core__abc_21380_n3987) );
  OR2X2 OR2X2_1562 ( .A(core__abc_21380_n3977), .B(core__abc_21380_n3988_1), .Y(core__abc_21380_n3989) );
  OR2X2 OR2X2_1563 ( .A(core__abc_21380_n3976), .B(core__abc_21380_n3987), .Y(core__abc_21380_n3990) );
  OR2X2 OR2X2_1564 ( .A(core_v3_reg_10_), .B(core_mi_10_), .Y(core__abc_21380_n3995_1) );
  OR2X2 OR2X2_1565 ( .A(core__abc_21380_n3994), .B(core__abc_21380_n3999), .Y(core__abc_21380_n4000_1) );
  OR2X2 OR2X2_1566 ( .A(core__abc_21380_n3317_bF_buf4), .B(core__abc_21380_n4000_1), .Y(core__abc_21380_n4001) );
  OR2X2 OR2X2_1567 ( .A(core__abc_21380_n3992_1), .B(core__abc_21380_n4001), .Y(core__abc_21380_n4002) );
  OR2X2 OR2X2_1568 ( .A(core__abc_21380_n3328_bF_buf5), .B(core_v3_reg_10_), .Y(core__abc_21380_n4003_1) );
  OR2X2 OR2X2_1569 ( .A(core__abc_21380_n3974_1), .B(core__abc_21380_n3966), .Y(core__abc_21380_n4006) );
  OR2X2 OR2X2_157 ( .A(_abc_19068_n910_1), .B(_abc_19068_n1240), .Y(_abc_19068_n1241_1) );
  OR2X2 OR2X2_1570 ( .A(core__abc_21380_n3948_1), .B(core__abc_21380_n2042), .Y(core__abc_21380_n4007) );
  OR2X2 OR2X2_1571 ( .A(core__abc_21380_n4009), .B(core__abc_21380_n4010), .Y(core__abc_21380_n4011) );
  OR2X2 OR2X2_1572 ( .A(core__abc_21380_n4013), .B(core__abc_21380_n1475), .Y(core__abc_21380_n4016_1) );
  OR2X2 OR2X2_1573 ( .A(core__abc_21380_n4019), .B(core__abc_21380_n4020), .Y(core__abc_21380_n4021) );
  OR2X2 OR2X2_1574 ( .A(core__abc_21380_n4011), .B(core__abc_21380_n4021), .Y(core__abc_21380_n4022) );
  OR2X2 OR2X2_1575 ( .A(core__abc_21380_n4006), .B(core__abc_21380_n4025), .Y(core__abc_21380_n4028) );
  OR2X2 OR2X2_1576 ( .A(core__abc_21380_n3919), .B(core__abc_21380_n4032), .Y(core__abc_21380_n4033) );
  OR2X2 OR2X2_1577 ( .A(core__abc_21380_n4035), .B(core__abc_21380_n4034_1), .Y(core__abc_21380_n4036) );
  OR2X2 OR2X2_1578 ( .A(core__abc_21380_n4039_1), .B(core__abc_21380_n4040), .Y(core__abc_21380_n4041) );
  OR2X2 OR2X2_1579 ( .A(core__abc_21380_n4042), .B(core_v3_reg_38_), .Y(core__abc_21380_n4043_1) );
  OR2X2 OR2X2_158 ( .A(_abc_19068_n1241_1), .B(_abc_19068_n1237_1), .Y(_abc_19068_n1242) );
  OR2X2 OR2X2_1580 ( .A(core__abc_21380_n4041), .B(core__abc_21380_n4044), .Y(core__abc_21380_n4045) );
  OR2X2 OR2X2_1581 ( .A(core__abc_21380_n4030), .B(core__abc_21380_n4047_1), .Y(core__abc_21380_n4048) );
  OR2X2 OR2X2_1582 ( .A(core__abc_21380_n4029), .B(core__abc_21380_n4046), .Y(core__abc_21380_n4049) );
  OR2X2 OR2X2_1583 ( .A(core_v3_reg_11_), .B(core_mi_11_), .Y(core__abc_21380_n4053) );
  OR2X2 OR2X2_1584 ( .A(core__abc_21380_n4052), .B(core__abc_21380_n4057_1), .Y(core__abc_21380_n4058) );
  OR2X2 OR2X2_1585 ( .A(core__abc_21380_n3317_bF_buf3), .B(core__abc_21380_n4058), .Y(core__abc_21380_n4059) );
  OR2X2 OR2X2_1586 ( .A(core__abc_21380_n4051), .B(core__abc_21380_n4059), .Y(core__abc_21380_n4060) );
  OR2X2 OR2X2_1587 ( .A(core__abc_21380_n3328_bF_buf4), .B(core_v3_reg_11_), .Y(core__abc_21380_n4061) );
  OR2X2 OR2X2_1588 ( .A(core__abc_21380_n3836), .B(core__abc_21380_n4067_1), .Y(core__abc_21380_n4068) );
  OR2X2 OR2X2_1589 ( .A(core__abc_21380_n3970), .B(core__abc_21380_n3902), .Y(core__abc_21380_n4069) );
  OR2X2 OR2X2_159 ( .A(_abc_19068_n1242), .B(_abc_19068_n1232), .Y(_abc_19068_n1243_1) );
  OR2X2 OR2X2_1590 ( .A(core__abc_21380_n4074), .B(core__abc_21380_n4023_1), .Y(core__abc_21380_n4075) );
  OR2X2 OR2X2_1591 ( .A(core__abc_21380_n4075), .B(core__abc_21380_n3968), .Y(core__abc_21380_n4076_1) );
  OR2X2 OR2X2_1592 ( .A(core__abc_21380_n4076_1), .B(core__abc_21380_n4069), .Y(core__abc_21380_n4077) );
  OR2X2 OR2X2_1593 ( .A(core__abc_21380_n4078), .B(core__abc_21380_n4074), .Y(core__abc_21380_n4079) );
  OR2X2 OR2X2_1594 ( .A(core__abc_21380_n4086), .B(core__abc_21380_n2061), .Y(core__abc_21380_n4087_1) );
  OR2X2 OR2X2_1595 ( .A(core__abc_21380_n4085), .B(core__abc_21380_n4087_1), .Y(core__abc_21380_n4088) );
  OR2X2 OR2X2_1596 ( .A(core__abc_21380_n4090), .B(core__abc_21380_n4088), .Y(core__abc_21380_n4091_1) );
  OR2X2 OR2X2_1597 ( .A(core__abc_21380_n3812), .B(core__abc_21380_n4094), .Y(core__abc_21380_n4095_1) );
  OR2X2 OR2X2_1598 ( .A(core__abc_21380_n4097), .B(core__abc_21380_n4092), .Y(core__abc_21380_n4098_1) );
  OR2X2 OR2X2_1599 ( .A(core__abc_21380_n4101), .B(core__abc_21380_n3049), .Y(core__abc_21380_n4102_1) );
  OR2X2 OR2X2_16 ( .A(_abc_19068_n934_1), .B(_abc_19068_n935), .Y(_abc_19068_n936_1) );
  OR2X2 OR2X2_160 ( .A(_abc_19068_n1245_1), .B(_abc_19068_n1246), .Y(_abc_19068_n1247_1) );
  OR2X2 OR2X2_1600 ( .A(core__abc_21380_n4105), .B(core__abc_21380_n4103), .Y(core__abc_21380_n4106_1) );
  OR2X2 OR2X2_1601 ( .A(core__abc_21380_n4107), .B(core__abc_21380_n4100), .Y(core__abc_21380_n4108) );
  OR2X2 OR2X2_1602 ( .A(core__abc_21380_n4106_1), .B(core_v3_reg_60_), .Y(core__abc_21380_n4109) );
  OR2X2 OR2X2_1603 ( .A(core__abc_21380_n4112), .B(core__abc_21380_n4113), .Y(core__abc_21380_n4114) );
  OR2X2 OR2X2_1604 ( .A(core__abc_21380_n4116), .B(core__abc_21380_n4117), .Y(core__abc_21380_n4118) );
  OR2X2 OR2X2_1605 ( .A(core__abc_21380_n4037), .B(core__abc_21380_n2275), .Y(core__abc_21380_n4120_1) );
  OR2X2 OR2X2_1606 ( .A(core__abc_21380_n4124_1), .B(core__abc_21380_n4122), .Y(core__abc_21380_n4125) );
  OR2X2 OR2X2_1607 ( .A(core__abc_21380_n4121), .B(core__abc_21380_n2295), .Y(core__abc_21380_n4129_1) );
  OR2X2 OR2X2_1608 ( .A(core__abc_21380_n4126), .B(core__abc_21380_n4131), .Y(core__abc_21380_n4132) );
  OR2X2 OR2X2_1609 ( .A(core__abc_21380_n4119), .B(core__abc_21380_n4132), .Y(core__abc_21380_n4133_1) );
  OR2X2 OR2X2_161 ( .A(_abc_19068_n906_1), .B(_abc_19068_n1185_1), .Y(_abc_19068_n1248) );
  OR2X2 OR2X2_1610 ( .A(core__abc_21380_n4130), .B(core__abc_21380_n4127), .Y(core__abc_21380_n4134) );
  OR2X2 OR2X2_1611 ( .A(core__abc_21380_n4125), .B(core_v3_reg_39_), .Y(core__abc_21380_n4135) );
  OR2X2 OR2X2_1612 ( .A(core__abc_21380_n4118), .B(core__abc_21380_n4136), .Y(core__abc_21380_n4137) );
  OR2X2 OR2X2_1613 ( .A(core_v3_reg_12_), .B(core_mi_12_), .Y(core__abc_21380_n4141_1) );
  OR2X2 OR2X2_1614 ( .A(core__abc_21380_n4140), .B(core__abc_21380_n4145_1), .Y(core__abc_21380_n4146) );
  OR2X2 OR2X2_1615 ( .A(core__abc_21380_n3317_bF_buf2), .B(core__abc_21380_n4146), .Y(core__abc_21380_n4147) );
  OR2X2 OR2X2_1616 ( .A(core__abc_21380_n4139), .B(core__abc_21380_n4147), .Y(core__abc_21380_n4148) );
  OR2X2 OR2X2_1617 ( .A(core__abc_21380_n3328_bF_buf3), .B(core_v3_reg_12_), .Y(core__abc_21380_n4149_1) );
  OR2X2 OR2X2_1618 ( .A(core__abc_21380_n4092), .B(core__abc_21380_n2077), .Y(core__abc_21380_n4156) );
  OR2X2 OR2X2_1619 ( .A(core__abc_21380_n4156), .B(core__abc_21380_n2101), .Y(core__abc_21380_n4157_1) );
  OR2X2 OR2X2_162 ( .A(_abc_19068_n1248), .B(_abc_19068_n1249_1), .Y(_abc_19068_n1250) );
  OR2X2 OR2X2_1620 ( .A(core__abc_21380_n4103), .B(core__abc_21380_n1488), .Y(core__abc_21380_n4162) );
  OR2X2 OR2X2_1621 ( .A(core__abc_21380_n4164), .B(core__abc_21380_n4165_1), .Y(core__abc_21380_n4166) );
  OR2X2 OR2X2_1622 ( .A(core__abc_21380_n4169), .B(core__abc_21380_n4167), .Y(core__abc_21380_n4170_1) );
  OR2X2 OR2X2_1623 ( .A(core__abc_21380_n4179), .B(core__abc_21380_n4180), .Y(core__abc_21380_n4181) );
  OR2X2 OR2X2_1624 ( .A(core__abc_21380_n4188), .B(core__abc_21380_n2290), .Y(core__abc_21380_n4189_1) );
  OR2X2 OR2X2_1625 ( .A(core__abc_21380_n4187), .B(core__abc_21380_n4189_1), .Y(core__abc_21380_n4190) );
  OR2X2 OR2X2_1626 ( .A(core__abc_21380_n4185), .B(core__abc_21380_n4190), .Y(core__abc_21380_n4191) );
  OR2X2 OR2X2_1627 ( .A(core__abc_21380_n4193), .B(core__abc_21380_n4191), .Y(core__abc_21380_n4194_1) );
  OR2X2 OR2X2_1628 ( .A(core__abc_21380_n4196), .B(core__abc_21380_n4197), .Y(core__abc_21380_n4198_1) );
  OR2X2 OR2X2_1629 ( .A(core__abc_21380_n4199), .B(core__abc_21380_n4182_1), .Y(core__abc_21380_n4200) );
  OR2X2 OR2X2_163 ( .A(_abc_19068_n1250), .B(_abc_19068_n1247_1), .Y(_abc_19068_n1251_1) );
  OR2X2 OR2X2_1630 ( .A(core__abc_21380_n4198_1), .B(core_v3_reg_40_), .Y(core__abc_21380_n4201) );
  OR2X2 OR2X2_1631 ( .A(core__abc_21380_n4181), .B(core__abc_21380_n4203_1), .Y(core__abc_21380_n4204) );
  OR2X2 OR2X2_1632 ( .A(core__abc_21380_n4205), .B(core__abc_21380_n4202), .Y(core__abc_21380_n4206_1) );
  OR2X2 OR2X2_1633 ( .A(core_v3_reg_13_), .B(core_mi_13_), .Y(core__abc_21380_n4211) );
  OR2X2 OR2X2_1634 ( .A(core__abc_21380_n4210_1), .B(core__abc_21380_n4215), .Y(core__abc_21380_n4216) );
  OR2X2 OR2X2_1635 ( .A(core__abc_21380_n3317_bF_buf1), .B(core__abc_21380_n4216), .Y(core__abc_21380_n4217) );
  OR2X2 OR2X2_1636 ( .A(core__abc_21380_n4208), .B(core__abc_21380_n4217), .Y(core__abc_21380_n4218_1) );
  OR2X2 OR2X2_1637 ( .A(core__abc_21380_n3328_bF_buf2), .B(core_v3_reg_13_), .Y(core__abc_21380_n4219) );
  OR2X2 OR2X2_1638 ( .A(core__abc_21380_n4096), .B(core__abc_21380_n4223), .Y(core__abc_21380_n4224_1) );
  OR2X2 OR2X2_1639 ( .A(core__abc_21380_n4226), .B(core__abc_21380_n2097), .Y(core__abc_21380_n4227) );
  OR2X2 OR2X2_164 ( .A(_abc_19068_n1253_1), .B(_abc_19068_n1254), .Y(_abc_19068_n1255_1) );
  OR2X2 OR2X2_1640 ( .A(core__abc_21380_n4230_1), .B(core__abc_21380_n4231), .Y(core__abc_21380_n4232) );
  OR2X2 OR2X2_1641 ( .A(core__abc_21380_n4229), .B(core__abc_21380_n4233), .Y(core__abc_21380_n4234) );
  OR2X2 OR2X2_1642 ( .A(core__abc_21380_n4237_1), .B(core__abc_21380_n3053), .Y(core__abc_21380_n4238) );
  OR2X2 OR2X2_1643 ( .A(core__abc_21380_n4240), .B(core__abc_21380_n4241), .Y(core__abc_21380_n4242) );
  OR2X2 OR2X2_1644 ( .A(core__abc_21380_n4243_1), .B(core__abc_21380_n4236), .Y(core__abc_21380_n4244) );
  OR2X2 OR2X2_1645 ( .A(core__abc_21380_n4242), .B(core_v3_reg_62_), .Y(core__abc_21380_n4245) );
  OR2X2 OR2X2_1646 ( .A(core__abc_21380_n4248), .B(core__abc_21380_n4249_1), .Y(core__abc_21380_n4250) );
  OR2X2 OR2X2_1647 ( .A(core__abc_21380_n4251), .B(core__abc_21380_n4175), .Y(core__abc_21380_n4252) );
  OR2X2 OR2X2_1648 ( .A(core__abc_21380_n4082_1), .B(core__abc_21380_n4254), .Y(core__abc_21380_n4255_1) );
  OR2X2 OR2X2_1649 ( .A(core__abc_21380_n4256), .B(core__abc_21380_n4250), .Y(core__abc_21380_n4258) );
  OR2X2 OR2X2_165 ( .A(_abc_19068_n1255_1), .B(_abc_19068_n1252), .Y(_abc_19068_n1256) );
  OR2X2 OR2X2_1650 ( .A(core__abc_21380_n4259), .B(core__abc_21380_n4257), .Y(core__abc_21380_n4260) );
  OR2X2 OR2X2_1651 ( .A(core__abc_21380_n4265), .B(core__abc_21380_n4266), .Y(core__abc_21380_n4267_1) );
  OR2X2 OR2X2_1652 ( .A(core__abc_21380_n4267_1), .B(core__abc_21380_n4262_1), .Y(core__abc_21380_n4268) );
  OR2X2 OR2X2_1653 ( .A(core__abc_21380_n4271), .B(core__abc_21380_n4269), .Y(core__abc_21380_n4272) );
  OR2X2 OR2X2_1654 ( .A(core__abc_21380_n4260), .B(core__abc_21380_n4272), .Y(core__abc_21380_n4273_1) );
  OR2X2 OR2X2_1655 ( .A(core__abc_21380_n4274), .B(core__abc_21380_n4275), .Y(core__abc_21380_n4276) );
  OR2X2 OR2X2_1656 ( .A(core_v3_reg_14_), .B(core_mi_14_), .Y(core__abc_21380_n4281) );
  OR2X2 OR2X2_1657 ( .A(core__abc_21380_n4280), .B(core__abc_21380_n4285), .Y(core__abc_21380_n4286) );
  OR2X2 OR2X2_1658 ( .A(core__abc_21380_n3317_bF_buf0), .B(core__abc_21380_n4286), .Y(core__abc_21380_n4287) );
  OR2X2 OR2X2_1659 ( .A(core__abc_21380_n4278_1), .B(core__abc_21380_n4287), .Y(core__abc_21380_n4288) );
  OR2X2 OR2X2_166 ( .A(_abc_19068_n1257_1), .B(_abc_19068_n1258), .Y(_abc_19068_n1259_1) );
  OR2X2 OR2X2_1660 ( .A(core__abc_21380_n3328_bF_buf1), .B(core_v3_reg_14_), .Y(core__abc_21380_n4289_1) );
  OR2X2 OR2X2_1661 ( .A(core__abc_21380_n4228), .B(core__abc_21380_n2119), .Y(core__abc_21380_n4295) );
  OR2X2 OR2X2_1662 ( .A(core__abc_21380_n4233), .B(core__abc_21380_n2115), .Y(core__abc_21380_n4298) );
  OR2X2 OR2X2_1663 ( .A(core__abc_21380_n4297), .B(core__abc_21380_n4299_1), .Y(core__abc_21380_n4300) );
  OR2X2 OR2X2_1664 ( .A(core__abc_21380_n4241), .B(core__abc_21380_n1524), .Y(core__abc_21380_n4302) );
  OR2X2 OR2X2_1665 ( .A(core__abc_21380_n4304_1), .B(core__abc_21380_n4305), .Y(core__abc_21380_n4306) );
  OR2X2 OR2X2_1666 ( .A(core__abc_21380_n4309_1), .B(core__abc_21380_n4307), .Y(core__abc_21380_n4310) );
  OR2X2 OR2X2_1667 ( .A(core__abc_21380_n4300), .B(core__abc_21380_n4311), .Y(core__abc_21380_n4312) );
  OR2X2 OR2X2_1668 ( .A(core__abc_21380_n4298), .B(core__abc_21380_n2139_1), .Y(core__abc_21380_n4313) );
  OR2X2 OR2X2_1669 ( .A(core__abc_21380_n4296), .B(core__abc_21380_n2140), .Y(core__abc_21380_n4314_1) );
  OR2X2 OR2X2_167 ( .A(_abc_19068_n1260), .B(_abc_19068_n1261_1), .Y(_abc_19068_n1262) );
  OR2X2 OR2X2_1670 ( .A(core__abc_21380_n4315), .B(core__abc_21380_n4310), .Y(core__abc_21380_n4316) );
  OR2X2 OR2X2_1671 ( .A(core__abc_21380_n4293), .B(core__abc_21380_n4317), .Y(core__abc_21380_n4320) );
  OR2X2 OR2X2_1672 ( .A(core__abc_21380_n4262_1), .B(core__abc_21380_n2327), .Y(core__abc_21380_n4323) );
  OR2X2 OR2X2_1673 ( .A(core__abc_21380_n4266), .B(core__abc_21380_n4323), .Y(core__abc_21380_n4324_1) );
  OR2X2 OR2X2_1674 ( .A(core__abc_21380_n4324_1), .B(core__abc_21380_n2347), .Y(core__abc_21380_n4327) );
  OR2X2 OR2X2_1675 ( .A(core__abc_21380_n4328), .B(core_v3_reg_42_), .Y(core__abc_21380_n4329_1) );
  OR2X2 OR2X2_1676 ( .A(core__abc_21380_n4331), .B(core__abc_21380_n4330), .Y(core__abc_21380_n4332) );
  OR2X2 OR2X2_1677 ( .A(core__abc_21380_n4322), .B(core__abc_21380_n4334_1), .Y(core__abc_21380_n4335) );
  OR2X2 OR2X2_1678 ( .A(core__abc_21380_n4321), .B(core__abc_21380_n4333), .Y(core__abc_21380_n4336) );
  OR2X2 OR2X2_1679 ( .A(core_v3_reg_15_), .B(core_mi_15_), .Y(core__abc_21380_n4340) );
  OR2X2 OR2X2_168 ( .A(_abc_19068_n1259_1), .B(_abc_19068_n1262), .Y(_abc_19068_n1263_1) );
  OR2X2 OR2X2_1680 ( .A(core__abc_21380_n4339_1), .B(core__abc_21380_n4344_1), .Y(core__abc_21380_n4345) );
  OR2X2 OR2X2_1681 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n4345), .Y(core__abc_21380_n4346) );
  OR2X2 OR2X2_1682 ( .A(core__abc_21380_n4338), .B(core__abc_21380_n4346), .Y(core__abc_21380_n4347) );
  OR2X2 OR2X2_1683 ( .A(core__abc_21380_n3328_bF_buf0), .B(core_v3_reg_15_), .Y(core__abc_21380_n4348) );
  OR2X2 OR2X2_1684 ( .A(core__abc_21380_n4300), .B(core__abc_21380_n4310), .Y(core__abc_21380_n4353) );
  OR2X2 OR2X2_1685 ( .A(core__abc_21380_n4315), .B(core__abc_21380_n4311), .Y(core__abc_21380_n4354) );
  OR2X2 OR2X2_1686 ( .A(core__abc_21380_n4360), .B(core__abc_21380_n4079), .Y(core__abc_21380_n4361_1) );
  OR2X2 OR2X2_1687 ( .A(core__abc_21380_n4366_1), .B(core__abc_21380_n4365), .Y(core__abc_21380_n4367) );
  OR2X2 OR2X2_1688 ( .A(core__abc_21380_n4364), .B(core__abc_21380_n4367), .Y(core__abc_21380_n4368) );
  OR2X2 OR2X2_1689 ( .A(core__abc_21380_n4368), .B(core__abc_21380_n4362), .Y(core__abc_21380_n4369) );
  OR2X2 OR2X2_169 ( .A(_abc_19068_n1263_1), .B(_abc_19068_n1256), .Y(_abc_19068_n1264) );
  OR2X2 OR2X2_1690 ( .A(core__abc_21380_n4369), .B(core__abc_21380_n4358), .Y(core__abc_21380_n4370) );
  OR2X2 OR2X2_1691 ( .A(core__abc_21380_n4379), .B(core__abc_21380_n2133), .Y(core__abc_21380_n4380) );
  OR2X2 OR2X2_1692 ( .A(core__abc_21380_n4378), .B(core__abc_21380_n4380), .Y(core__abc_21380_n4381_1) );
  OR2X2 OR2X2_1693 ( .A(core__abc_21380_n4377), .B(core__abc_21380_n4381_1), .Y(core__abc_21380_n4382) );
  OR2X2 OR2X2_1694 ( .A(core__abc_21380_n4376_1), .B(core__abc_21380_n4382), .Y(core__abc_21380_n4383) );
  OR2X2 OR2X2_1695 ( .A(core__abc_21380_n4375), .B(core__abc_21380_n4383), .Y(core__abc_21380_n4384) );
  OR2X2 OR2X2_1696 ( .A(core__abc_21380_n3287), .B(core__abc_21380_n4386_1), .Y(core__abc_21380_n4387) );
  OR2X2 OR2X2_1697 ( .A(core__abc_21380_n4390), .B(core__abc_21380_n4385), .Y(core__abc_21380_n4391) );
  OR2X2 OR2X2_1698 ( .A(core__abc_21380_n4395), .B(core__abc_21380_n4393), .Y(core__abc_21380_n4396) );
  OR2X2 OR2X2_1699 ( .A(core__abc_21380_n4397_1), .B(core_v3_reg_0_), .Y(core__abc_21380_n4398) );
  OR2X2 OR2X2_17 ( .A(_abc_19068_n936_1), .B(_abc_19068_n933_1), .Y(_abc_19068_n937_1) );
  OR2X2 OR2X2_170 ( .A(_abc_19068_n1264), .B(_abc_19068_n1251_1), .Y(_abc_19068_n1265_1) );
  OR2X2 OR2X2_1700 ( .A(core__abc_21380_n4396), .B(core__abc_21380_n1263), .Y(core__abc_21380_n4399) );
  OR2X2 OR2X2_1701 ( .A(core__abc_21380_n4403), .B(core__abc_21380_n4401), .Y(core__abc_21380_n4404) );
  OR2X2 OR2X2_1702 ( .A(core__abc_21380_n4317), .B(core__abc_21380_n4250), .Y(core__abc_21380_n4407_1) );
  OR2X2 OR2X2_1703 ( .A(core__abc_21380_n4407_1), .B(core__abc_21380_n4254), .Y(core__abc_21380_n4408) );
  OR2X2 OR2X2_1704 ( .A(core__abc_21380_n4068), .B(core__abc_21380_n4408), .Y(core__abc_21380_n4409) );
  OR2X2 OR2X2_1705 ( .A(core__abc_21380_n4408), .B(core__abc_21380_n4081), .Y(core__abc_21380_n4410) );
  OR2X2 OR2X2_1706 ( .A(core__abc_21380_n4407_1), .B(core__abc_21380_n4252), .Y(core__abc_21380_n4411) );
  OR2X2 OR2X2_1707 ( .A(core__abc_21380_n4406), .B(core__abc_21380_n4416), .Y(core__abc_21380_n4417_1) );
  OR2X2 OR2X2_1708 ( .A(core__abc_21380_n4418), .B(core__abc_21380_n2369_1), .Y(core__abc_21380_n4421) );
  OR2X2 OR2X2_1709 ( .A(core__abc_21380_n4422_1), .B(core_v3_reg_43_), .Y(core__abc_21380_n4423) );
  OR2X2 OR2X2_171 ( .A(_abc_19068_n1267_1), .B(_abc_19068_n1268), .Y(_abc_19068_n1269_1) );
  OR2X2 OR2X2_1710 ( .A(core__abc_21380_n4424), .B(core__abc_21380_n4425), .Y(core__abc_21380_n4426) );
  OR2X2 OR2X2_1711 ( .A(core__abc_21380_n4426), .B(core__abc_21380_n4417_1), .Y(core__abc_21380_n4427_1) );
  OR2X2 OR2X2_1712 ( .A(core__abc_21380_n4428), .B(core__abc_21380_n4430), .Y(core__abc_21380_n4431) );
  OR2X2 OR2X2_1713 ( .A(core_v3_reg_16_), .B(core_mi_16_), .Y(core__abc_21380_n4435) );
  OR2X2 OR2X2_1714 ( .A(core__abc_21380_n4434), .B(core__abc_21380_n4439), .Y(core__abc_21380_n4440) );
  OR2X2 OR2X2_1715 ( .A(core__abc_21380_n3317_bF_buf6), .B(core__abc_21380_n4440), .Y(core__abc_21380_n4441) );
  OR2X2 OR2X2_1716 ( .A(core__abc_21380_n4433), .B(core__abc_21380_n4441), .Y(core__abc_21380_n4442) );
  OR2X2 OR2X2_1717 ( .A(core__abc_21380_n3328_bF_buf7), .B(core_v3_reg_16_), .Y(core__abc_21380_n4443_1) );
  OR2X2 OR2X2_1718 ( .A(core__abc_21380_n4395), .B(core__abc_21380_n1562), .Y(core__abc_21380_n4462) );
  OR2X2 OR2X2_1719 ( .A(core__abc_21380_n4464_1), .B(core__abc_21380_n4465), .Y(core__abc_21380_n4466) );
  OR2X2 OR2X2_172 ( .A(_abc_19068_n1271_1), .B(_abc_19068_n1272), .Y(_abc_19068_n1273_1) );
  OR2X2 OR2X2_1720 ( .A(core__abc_21380_n4469_1), .B(core__abc_21380_n4467), .Y(core__abc_21380_n4470) );
  OR2X2 OR2X2_1721 ( .A(core__abc_21380_n4449), .B(core__abc_21380_n4477), .Y(core__abc_21380_n4478) );
  OR2X2 OR2X2_1722 ( .A(core__abc_21380_n4448_1), .B(core__abc_21380_n4479), .Y(core__abc_21380_n4480_1) );
  OR2X2 OR2X2_1723 ( .A(core__abc_21380_n4484), .B(core__abc_21380_n2364), .Y(core__abc_21380_n4485_1) );
  OR2X2 OR2X2_1724 ( .A(core__abc_21380_n4483), .B(core__abc_21380_n4485_1), .Y(core__abc_21380_n4486) );
  OR2X2 OR2X2_1725 ( .A(core__abc_21380_n4488), .B(core__abc_21380_n4489), .Y(core__abc_21380_n4490) );
  OR2X2 OR2X2_1726 ( .A(core__abc_21380_n4491_1), .B(core_v3_reg_44_), .Y(core__abc_21380_n4492) );
  OR2X2 OR2X2_1727 ( .A(core__abc_21380_n4490), .B(core__abc_21380_n4493), .Y(core__abc_21380_n4494) );
  OR2X2 OR2X2_1728 ( .A(core__abc_21380_n4482), .B(core__abc_21380_n4496_1), .Y(core__abc_21380_n4497) );
  OR2X2 OR2X2_1729 ( .A(core__abc_21380_n4481), .B(core__abc_21380_n4495), .Y(core__abc_21380_n4498) );
  OR2X2 OR2X2_173 ( .A(_abc_19068_n1273_1), .B(_abc_19068_n1270), .Y(_abc_19068_n1274) );
  OR2X2 OR2X2_1730 ( .A(core_v3_reg_17_), .B(core_mi_17_), .Y(core__abc_21380_n4502) );
  OR2X2 OR2X2_1731 ( .A(core__abc_21380_n4501_1), .B(core__abc_21380_n4506_1), .Y(core__abc_21380_n4507) );
  OR2X2 OR2X2_1732 ( .A(core__abc_21380_n3317_bF_buf5), .B(core__abc_21380_n4507), .Y(core__abc_21380_n4508) );
  OR2X2 OR2X2_1733 ( .A(core__abc_21380_n4500), .B(core__abc_21380_n4508), .Y(core__abc_21380_n4509) );
  OR2X2 OR2X2_1734 ( .A(core__abc_21380_n3328_bF_buf6), .B(core_v3_reg_17_), .Y(core__abc_21380_n4510) );
  OR2X2 OR2X2_1735 ( .A(core__abc_21380_n4475), .B(core__abc_21380_n4446), .Y(core__abc_21380_n4513) );
  OR2X2 OR2X2_1736 ( .A(core__abc_21380_n4517), .B(core__abc_21380_n4515), .Y(core__abc_21380_n4518) );
  OR2X2 OR2X2_1737 ( .A(core__abc_21380_n4455), .B(core__abc_21380_n2171), .Y(core__abc_21380_n4520) );
  OR2X2 OR2X2_1738 ( .A(core__abc_21380_n4458), .B(core__abc_21380_n4520), .Y(core__abc_21380_n4521) );
  OR2X2 OR2X2_1739 ( .A(core__abc_21380_n4523), .B(core__abc_21380_n4524), .Y(core__abc_21380_n4525) );
  OR2X2 OR2X2_174 ( .A(_abc_19068_n1274), .B(_abc_19068_n1269_1), .Y(_abc_19068_n1275_1) );
  OR2X2 OR2X2_1740 ( .A(core__abc_21380_n3060), .B(core__abc_21380_n4527_1), .Y(core__abc_21380_n4528) );
  OR2X2 OR2X2_1741 ( .A(core__abc_21380_n4529), .B(core__abc_21380_n1604), .Y(core__abc_21380_n4531) );
  OR2X2 OR2X2_1742 ( .A(core__abc_21380_n4532_1), .B(core__abc_21380_n4530), .Y(core__abc_21380_n4533) );
  OR2X2 OR2X2_1743 ( .A(core__abc_21380_n4534), .B(core__abc_21380_n1305), .Y(core__abc_21380_n4535) );
  OR2X2 OR2X2_1744 ( .A(core__abc_21380_n4533), .B(core_v3_reg_2_), .Y(core__abc_21380_n4536) );
  OR2X2 OR2X2_1745 ( .A(core__abc_21380_n4539), .B(core__abc_21380_n4540), .Y(core__abc_21380_n4541) );
  OR2X2 OR2X2_1746 ( .A(core__abc_21380_n4542_1), .B(core__abc_21380_n4544), .Y(core__abc_21380_n4545) );
  OR2X2 OR2X2_1747 ( .A(core__abc_21380_n4489), .B(core__abc_21380_n2383), .Y(core__abc_21380_n4546) );
  OR2X2 OR2X2_1748 ( .A(core__abc_21380_n4549), .B(core__abc_21380_n4547_1), .Y(core__abc_21380_n4550) );
  OR2X2 OR2X2_1749 ( .A(core__abc_21380_n4550), .B(core_v3_reg_45_), .Y(core__abc_21380_n4553) );
  OR2X2 OR2X2_175 ( .A(_abc_19068_n1277_1), .B(_abc_19068_n1278), .Y(_abc_19068_n1279_1) );
  OR2X2 OR2X2_1750 ( .A(core__abc_21380_n4555), .B(core__abc_21380_n4545), .Y(core__abc_21380_n4556) );
  OR2X2 OR2X2_1751 ( .A(core__abc_21380_n4554), .B(core__abc_21380_n4557), .Y(core__abc_21380_n4558) );
  OR2X2 OR2X2_1752 ( .A(core_v3_reg_18_), .B(core_mi_18_), .Y(core__abc_21380_n4563) );
  OR2X2 OR2X2_1753 ( .A(core__abc_21380_n4562), .B(core__abc_21380_n4567), .Y(core__abc_21380_n4568) );
  OR2X2 OR2X2_1754 ( .A(core__abc_21380_n3317_bF_buf4), .B(core__abc_21380_n4568), .Y(core__abc_21380_n4569) );
  OR2X2 OR2X2_1755 ( .A(core__abc_21380_n4560_1), .B(core__abc_21380_n4569), .Y(core__abc_21380_n4570) );
  OR2X2 OR2X2_1756 ( .A(core__abc_21380_n3328_bF_buf5), .B(core_v3_reg_18_), .Y(core__abc_21380_n4571_1) );
  OR2X2 OR2X2_1757 ( .A(core__abc_21380_n4576_1), .B(core__abc_21380_n4575), .Y(core__abc_21380_n4577) );
  OR2X2 OR2X2_1758 ( .A(core__abc_21380_n4579), .B(core__abc_21380_n4580), .Y(core__abc_21380_n4581) );
  OR2X2 OR2X2_1759 ( .A(core__abc_21380_n4584), .B(core__abc_21380_n4582_1), .Y(core__abc_21380_n4585) );
  OR2X2 OR2X2_176 ( .A(_abc_19068_n1280), .B(_abc_19068_n1281_1), .Y(_abc_19068_n1282) );
  OR2X2 OR2X2_1760 ( .A(core__abc_21380_n4524), .B(core__abc_21380_n2189), .Y(core__abc_21380_n4590) );
  OR2X2 OR2X2_1761 ( .A(core__abc_21380_n4590), .B(core__abc_21380_n2213_1), .Y(core__abc_21380_n4591) );
  OR2X2 OR2X2_1762 ( .A(core__abc_21380_n4595), .B(core__abc_21380_n1619), .Y(core__abc_21380_n4598) );
  OR2X2 OR2X2_1763 ( .A(core__abc_21380_n4601), .B(core__abc_21380_n4602), .Y(core__abc_21380_n4603_1) );
  OR2X2 OR2X2_1764 ( .A(core__abc_21380_n4607), .B(core__abc_21380_n4605), .Y(core__abc_21380_n4608_1) );
  OR2X2 OR2X2_1765 ( .A(core__abc_21380_n4589), .B(core__abc_21380_n4609), .Y(core__abc_21380_n4610) );
  OR2X2 OR2X2_1766 ( .A(core__abc_21380_n4588), .B(core__abc_21380_n4608_1), .Y(core__abc_21380_n4611) );
  OR2X2 OR2X2_1767 ( .A(core__abc_21380_n4614_1), .B(core__abc_21380_n4585), .Y(core__abc_21380_n4615) );
  OR2X2 OR2X2_1768 ( .A(core__abc_21380_n4616), .B(core__abc_21380_n4617), .Y(core__abc_21380_n4618) );
  OR2X2 OR2X2_1769 ( .A(core_v3_reg_19_), .B(core_mi_19_), .Y(core__abc_21380_n4623) );
  OR2X2 OR2X2_177 ( .A(_abc_19068_n1279_1), .B(_abc_19068_n1282), .Y(_abc_19068_n1283_1) );
  OR2X2 OR2X2_1770 ( .A(core__abc_21380_n4620), .B(core__abc_21380_n4625), .Y(core__abc_21380_n4626) );
  OR2X2 OR2X2_1771 ( .A(core__abc_21380_n3317_bF_buf3), .B(core__abc_21380_n4626), .Y(core__abc_21380_n4627) );
  OR2X2 OR2X2_1772 ( .A(core__abc_21380_n4619_1), .B(core__abc_21380_n4627), .Y(core__abc_21380_n4628) );
  OR2X2 OR2X2_1773 ( .A(core__abc_21380_n3328_bF_buf4), .B(core_v3_reg_19_), .Y(core__abc_21380_n4629_1) );
  OR2X2 OR2X2_1774 ( .A(core__abc_21380_n4634_1), .B(core__abc_21380_n2207), .Y(core__abc_21380_n4635) );
  OR2X2 OR2X2_1775 ( .A(core__abc_21380_n4633), .B(core__abc_21380_n4635), .Y(core__abc_21380_n4636) );
  OR2X2 OR2X2_1776 ( .A(core__abc_21380_n4638), .B(core__abc_21380_n4636), .Y(core__abc_21380_n4639_1) );
  OR2X2 OR2X2_1777 ( .A(core__abc_21380_n4641), .B(core__abc_21380_n4642), .Y(core__abc_21380_n4643) );
  OR2X2 OR2X2_1778 ( .A(core__abc_21380_n4645), .B(core__abc_21380_n3085), .Y(core__abc_21380_n4646) );
  OR2X2 OR2X2_1779 ( .A(core__abc_21380_n4649), .B(core__abc_21380_n4647), .Y(core__abc_21380_n4650_1) );
  OR2X2 OR2X2_178 ( .A(_abc_19068_n1283_1), .B(_abc_19068_n1276), .Y(_abc_19068_n1284) );
  OR2X2 OR2X2_1780 ( .A(core__abc_21380_n4651), .B(core__abc_21380_n1341), .Y(core__abc_21380_n4652) );
  OR2X2 OR2X2_1781 ( .A(core__abc_21380_n4650_1), .B(core_v3_reg_4_), .Y(core__abc_21380_n4653) );
  OR2X2 OR2X2_1782 ( .A(core__abc_21380_n4656), .B(core__abc_21380_n4657), .Y(core__abc_21380_n4658) );
  OR2X2 OR2X2_1783 ( .A(core__abc_21380_n4660_1), .B(core__abc_21380_n4607), .Y(core__abc_21380_n4661) );
  OR2X2 OR2X2_1784 ( .A(core__abc_21380_n4664), .B(core__abc_21380_n4662), .Y(core__abc_21380_n4665) );
  OR2X2 OR2X2_1785 ( .A(core__abc_21380_n4415), .B(core__abc_21380_n4668), .Y(core__abc_21380_n4669) );
  OR2X2 OR2X2_1786 ( .A(core__abc_21380_n4670), .B(core__abc_21380_n4658), .Y(core__abc_21380_n4672) );
  OR2X2 OR2X2_1787 ( .A(core__abc_21380_n4673), .B(core__abc_21380_n4671_1), .Y(core__abc_21380_n4674) );
  OR2X2 OR2X2_1788 ( .A(core__abc_21380_n4579), .B(core__abc_21380_n2419), .Y(core__abc_21380_n4676_1) );
  OR2X2 OR2X2_1789 ( .A(core__abc_21380_n4678), .B(core__abc_21380_n4679), .Y(core__abc_21380_n4680) );
  OR2X2 OR2X2_179 ( .A(_abc_19068_n1284), .B(_abc_19068_n1275_1), .Y(_abc_19068_n1285_1) );
  OR2X2 OR2X2_1790 ( .A(core__abc_21380_n4683), .B(core__abc_21380_n4681_1), .Y(core__abc_21380_n4684) );
  OR2X2 OR2X2_1791 ( .A(core__abc_21380_n4684), .B(core__abc_21380_n4674), .Y(core__abc_21380_n4685) );
  OR2X2 OR2X2_1792 ( .A(core__abc_21380_n4680), .B(core__abc_21380_n4675), .Y(core__abc_21380_n4688) );
  OR2X2 OR2X2_1793 ( .A(core__abc_21380_n4689), .B(core__abc_21380_n4686_1), .Y(core__abc_21380_n4690) );
  OR2X2 OR2X2_1794 ( .A(core_v3_reg_20_), .B(core_mi_20_), .Y(core__abc_21380_n4695) );
  OR2X2 OR2X2_1795 ( .A(core__abc_21380_n4694), .B(core__abc_21380_n4699), .Y(core__abc_21380_n4700) );
  OR2X2 OR2X2_1796 ( .A(core__abc_21380_n3317_bF_buf2), .B(core__abc_21380_n4700), .Y(core__abc_21380_n4701_1) );
  OR2X2 OR2X2_1797 ( .A(core__abc_21380_n4692), .B(core__abc_21380_n4701_1), .Y(core__abc_21380_n4702) );
  OR2X2 OR2X2_1798 ( .A(core__abc_21380_n3328_bF_buf3), .B(core_v3_reg_20_), .Y(core__abc_21380_n4703) );
  OR2X2 OR2X2_1799 ( .A(core__abc_21380_n4642), .B(core__abc_21380_n2228), .Y(core__abc_21380_n4706) );
  OR2X2 OR2X2_18 ( .A(_abc_19068_n932), .B(_abc_19068_n937_1), .Y(_abc_19068_n938) );
  OR2X2 OR2X2_180 ( .A(_abc_19068_n1248), .B(_abc_19068_n1287_1), .Y(_abc_19068_n1288) );
  OR2X2 OR2X2_1800 ( .A(core__abc_21380_n4708), .B(core__abc_21380_n4709), .Y(core__abc_21380_n4710) );
  OR2X2 OR2X2_1801 ( .A(core__abc_21380_n4647), .B(core__abc_21380_n1634), .Y(core__abc_21380_n4712_1) );
  OR2X2 OR2X2_1802 ( .A(core__abc_21380_n4714), .B(core__abc_21380_n4715), .Y(core__abc_21380_n4716) );
  OR2X2 OR2X2_1803 ( .A(core__abc_21380_n4719), .B(core__abc_21380_n4717_1), .Y(core__abc_21380_n4720) );
  OR2X2 OR2X2_1804 ( .A(core__abc_21380_n4722_1), .B(core__abc_21380_n4723), .Y(core__abc_21380_n4724) );
  OR2X2 OR2X2_1805 ( .A(core__abc_21380_n4726), .B(core__abc_21380_n4724), .Y(core__abc_21380_n4728) );
  OR2X2 OR2X2_1806 ( .A(core__abc_21380_n4729), .B(core__abc_21380_n4727_1), .Y(core__abc_21380_n4730) );
  OR2X2 OR2X2_1807 ( .A(core__abc_21380_n4731), .B(core__abc_21380_n3295), .Y(core__abc_21380_n4732_1) );
  OR2X2 OR2X2_1808 ( .A(core__abc_21380_n4730), .B(core__abc_21380_n3294), .Y(core__abc_21380_n4733) );
  OR2X2 OR2X2_1809 ( .A(core_v3_reg_21_), .B(core_mi_21_), .Y(core__abc_21380_n4738) );
  OR2X2 OR2X2_181 ( .A(_abc_19068_n1289_1), .B(_abc_19068_n1290), .Y(_abc_19068_n1291_1) );
  OR2X2 OR2X2_1810 ( .A(core__abc_21380_n4737_1), .B(core__abc_21380_n4742_1), .Y(core__abc_21380_n4743) );
  OR2X2 OR2X2_1811 ( .A(core__abc_21380_n3317_bF_buf1), .B(core__abc_21380_n4743), .Y(core__abc_21380_n4744) );
  OR2X2 OR2X2_1812 ( .A(core__abc_21380_n4735), .B(core__abc_21380_n4744), .Y(core__abc_21380_n4745) );
  OR2X2 OR2X2_1813 ( .A(core__abc_21380_n3328_bF_buf2), .B(core_v3_reg_21_), .Y(core__abc_21380_n4746) );
  OR2X2 OR2X2_1814 ( .A(core__abc_21380_n4724), .B(core__abc_21380_n4658), .Y(core__abc_21380_n4749) );
  OR2X2 OR2X2_1815 ( .A(core__abc_21380_n4670), .B(core__abc_21380_n4749), .Y(core__abc_21380_n4750) );
  OR2X2 OR2X2_1816 ( .A(core__abc_21380_n4752_1), .B(core__abc_21380_n4723), .Y(core__abc_21380_n4753) );
  OR2X2 OR2X2_1817 ( .A(core__abc_21380_n4755), .B(core__abc_21380_n2248), .Y(core__abc_21380_n4756) );
  OR2X2 OR2X2_1818 ( .A(core__abc_21380_n4759), .B(core__abc_21380_n4757_1), .Y(core__abc_21380_n4760) );
  OR2X2 OR2X2_1819 ( .A(core__abc_21380_n4762_1), .B(core__abc_21380_n4763), .Y(core__abc_21380_n4764) );
  OR2X2 OR2X2_182 ( .A(_abc_19068_n1288), .B(_abc_19068_n1291_1), .Y(_abc_19068_n1292) );
  OR2X2 OR2X2_1820 ( .A(core__abc_21380_n4766), .B(core__abc_21380_n3089), .Y(core__abc_21380_n4767_1) );
  OR2X2 OR2X2_1821 ( .A(core__abc_21380_n4769), .B(core__abc_21380_n4770), .Y(core__abc_21380_n4771) );
  OR2X2 OR2X2_1822 ( .A(core__abc_21380_n4772_1), .B(core__abc_21380_n1380), .Y(core__abc_21380_n4773) );
  OR2X2 OR2X2_1823 ( .A(core__abc_21380_n4771), .B(core_v3_reg_6_), .Y(core__abc_21380_n4774) );
  OR2X2 OR2X2_1824 ( .A(core__abc_21380_n4777_1), .B(core__abc_21380_n4778), .Y(core__abc_21380_n4779) );
  OR2X2 OR2X2_1825 ( .A(core__abc_21380_n4754), .B(core__abc_21380_n4779), .Y(core__abc_21380_n4781) );
  OR2X2 OR2X2_1826 ( .A(core__abc_21380_n4782), .B(core__abc_21380_n4780), .Y(core__abc_21380_n4783_1) );
  OR2X2 OR2X2_1827 ( .A(core__abc_21380_n4784), .B(core__abc_21380_n3349), .Y(core__abc_21380_n4785) );
  OR2X2 OR2X2_1828 ( .A(core__abc_21380_n4783_1), .B(core__abc_21380_n3348), .Y(core__abc_21380_n4786) );
  OR2X2 OR2X2_1829 ( .A(core_v3_reg_22_), .B(core_mi_22_), .Y(core__abc_21380_n4791) );
  OR2X2 OR2X2_183 ( .A(_abc_19068_n1294), .B(_abc_19068_n1295_1), .Y(_abc_19068_n1296) );
  OR2X2 OR2X2_1830 ( .A(core__abc_21380_n4790), .B(core__abc_21380_n4795), .Y(core__abc_21380_n4796) );
  OR2X2 OR2X2_1831 ( .A(core__abc_21380_n3317_bF_buf0), .B(core__abc_21380_n4796), .Y(core__abc_21380_n4797) );
  OR2X2 OR2X2_1832 ( .A(core__abc_21380_n4788_1), .B(core__abc_21380_n4797), .Y(core__abc_21380_n4798_1) );
  OR2X2 OR2X2_1833 ( .A(core__abc_21380_n3328_bF_buf1), .B(core_v3_reg_22_), .Y(core__abc_21380_n4799) );
  OR2X2 OR2X2_1834 ( .A(core__abc_21380_n4763), .B(core__abc_21380_n2267), .Y(core__abc_21380_n4805) );
  OR2X2 OR2X2_1835 ( .A(core__abc_21380_n4807), .B(core__abc_21380_n4808_1), .Y(core__abc_21380_n4809) );
  OR2X2 OR2X2_1836 ( .A(core__abc_21380_n4770), .B(core__abc_21380_n1670), .Y(core__abc_21380_n4810) );
  OR2X2 OR2X2_1837 ( .A(core__abc_21380_n4812), .B(core__abc_21380_n4813), .Y(core__abc_21380_n4814_1) );
  OR2X2 OR2X2_1838 ( .A(core__abc_21380_n4814_1), .B(core__abc_21380_n1399), .Y(core__abc_21380_n4816) );
  OR2X2 OR2X2_1839 ( .A(core__abc_21380_n4817), .B(core__abc_21380_n4815), .Y(core__abc_21380_n4818) );
  OR2X2 OR2X2_184 ( .A(_abc_19068_n1296), .B(_abc_19068_n1293_1), .Y(_abc_19068_n1297) );
  OR2X2 OR2X2_1840 ( .A(core__abc_21380_n4818), .B(core__abc_21380_n4809), .Y(core__abc_21380_n4819) );
  OR2X2 OR2X2_1841 ( .A(core__abc_21380_n4822), .B(core__abc_21380_n4824), .Y(core__abc_21380_n4825_1) );
  OR2X2 OR2X2_1842 ( .A(core__abc_21380_n4804), .B(core__abc_21380_n4826), .Y(core__abc_21380_n4827) );
  OR2X2 OR2X2_1843 ( .A(core__abc_21380_n4828), .B(core__abc_21380_n4829), .Y(core__abc_21380_n4830_1) );
  OR2X2 OR2X2_1844 ( .A(core__abc_21380_n4803_1), .B(core__abc_21380_n4830_1), .Y(core__abc_21380_n4831) );
  OR2X2 OR2X2_1845 ( .A(core__abc_21380_n4832), .B(core__abc_21380_n3420), .Y(core__abc_21380_n4833) );
  OR2X2 OR2X2_1846 ( .A(core__abc_21380_n4834), .B(core__abc_21380_n3419), .Y(core__abc_21380_n4835_1) );
  OR2X2 OR2X2_1847 ( .A(core_v3_reg_23_), .B(core_mi_23_), .Y(core__abc_21380_n4839) );
  OR2X2 OR2X2_1848 ( .A(core__abc_21380_n4838), .B(core__abc_21380_n4843), .Y(core__abc_21380_n4844) );
  OR2X2 OR2X2_1849 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n4844), .Y(core__abc_21380_n4845_1) );
  OR2X2 OR2X2_185 ( .A(_abc_19068_n1298_1), .B(_abc_19068_n1299), .Y(_abc_19068_n1300_1) );
  OR2X2 OR2X2_1850 ( .A(core__abc_21380_n4837), .B(core__abc_21380_n4845_1), .Y(core__abc_21380_n4846) );
  OR2X2 OR2X2_1851 ( .A(core__abc_21380_n3328_bF_buf0), .B(core_v3_reg_23_), .Y(core__abc_21380_n4847) );
  OR2X2 OR2X2_1852 ( .A(core__abc_21380_n4415), .B(core__abc_21380_n4855), .Y(core__abc_21380_n4856) );
  OR2X2 OR2X2_1853 ( .A(core__abc_21380_n4830_1), .B(core__abc_21380_n4779), .Y(core__abc_21380_n4857_1) );
  OR2X2 OR2X2_1854 ( .A(core__abc_21380_n4857_1), .B(core__abc_21380_n4749), .Y(core__abc_21380_n4858) );
  OR2X2 OR2X2_1855 ( .A(core__abc_21380_n4858), .B(core__abc_21380_n4666_1), .Y(core__abc_21380_n4859) );
  OR2X2 OR2X2_1856 ( .A(core__abc_21380_n4857_1), .B(core__abc_21380_n4753), .Y(core__abc_21380_n4860) );
  OR2X2 OR2X2_1857 ( .A(core__abc_21380_n4861), .B(core__abc_21380_n4828), .Y(core__abc_21380_n4862_1) );
  OR2X2 OR2X2_1858 ( .A(core__abc_21380_n4389), .B(core__abc_21380_n4871), .Y(core__abc_21380_n4872) );
  OR2X2 OR2X2_1859 ( .A(core__abc_21380_n4875), .B(core__abc_21380_n2286), .Y(core__abc_21380_n4876) );
  OR2X2 OR2X2_186 ( .A(_abc_19068_n1301), .B(_abc_19068_n1302_1), .Y(_abc_19068_n1303) );
  OR2X2 OR2X2_1860 ( .A(core__abc_21380_n4874), .B(core__abc_21380_n4876), .Y(core__abc_21380_n4877) );
  OR2X2 OR2X2_1861 ( .A(core__abc_21380_n4873_1), .B(core__abc_21380_n4877), .Y(core__abc_21380_n4878_1) );
  OR2X2 OR2X2_1862 ( .A(core__abc_21380_n4882), .B(core__abc_21380_n4878_1), .Y(core__abc_21380_n4883_1) );
  OR2X2 OR2X2_1863 ( .A(core__abc_21380_n4881), .B(core__abc_21380_n4884), .Y(core__abc_21380_n4885) );
  OR2X2 OR2X2_1864 ( .A(core__abc_21380_n3060), .B(core__abc_21380_n4889), .Y(core__abc_21380_n4890) );
  OR2X2 OR2X2_1865 ( .A(core__abc_21380_n4894), .B(core__abc_21380_n4892_1), .Y(core__abc_21380_n4895) );
  OR2X2 OR2X2_1866 ( .A(core__abc_21380_n4896_1), .B(core__abc_21380_n4887), .Y(core__abc_21380_n4897) );
  OR2X2 OR2X2_1867 ( .A(core__abc_21380_n4895), .B(core_v3_reg_8_), .Y(core__abc_21380_n4898_1) );
  OR2X2 OR2X2_1868 ( .A(core__abc_21380_n4901), .B(core__abc_21380_n4902_1), .Y(core__abc_21380_n4903) );
  OR2X2 OR2X2_1869 ( .A(core__abc_21380_n4905), .B(core__abc_21380_n4906), .Y(core__abc_21380_n4907) );
  OR2X2 OR2X2_187 ( .A(_abc_19068_n1300_1), .B(_abc_19068_n1303), .Y(_abc_19068_n1304_1) );
  OR2X2 OR2X2_1870 ( .A(core__abc_21380_n4908), .B(core__abc_21380_n3478), .Y(core__abc_21380_n4909) );
  OR2X2 OR2X2_1871 ( .A(core__abc_21380_n4907), .B(core__abc_21380_n3475), .Y(core__abc_21380_n4910) );
  OR2X2 OR2X2_1872 ( .A(core_v3_reg_24_), .B(core_mi_24_), .Y(core__abc_21380_n4915) );
  OR2X2 OR2X2_1873 ( .A(core__abc_21380_n4914), .B(core__abc_21380_n4919), .Y(core__abc_21380_n4920) );
  OR2X2 OR2X2_1874 ( .A(core__abc_21380_n3317_bF_buf6), .B(core__abc_21380_n4920), .Y(core__abc_21380_n4921) );
  OR2X2 OR2X2_1875 ( .A(core__abc_21380_n4912), .B(core__abc_21380_n4921), .Y(core__abc_21380_n4922) );
  OR2X2 OR2X2_1876 ( .A(core__abc_21380_n3328_bF_buf7), .B(core_v3_reg_24_), .Y(core__abc_21380_n4923) );
  OR2X2 OR2X2_1877 ( .A(core__abc_21380_n4884), .B(core__abc_21380_n2305), .Y(core__abc_21380_n4930) );
  OR2X2 OR2X2_1878 ( .A(core__abc_21380_n4932), .B(core__abc_21380_n4934), .Y(core__abc_21380_n4935) );
  OR2X2 OR2X2_1879 ( .A(core__abc_21380_n4935), .B(core__abc_21380_n4929), .Y(core__abc_21380_n4936) );
  OR2X2 OR2X2_188 ( .A(_abc_19068_n1304_1), .B(_abc_19068_n1297), .Y(_abc_19068_n1305) );
  OR2X2 OR2X2_1880 ( .A(core__abc_21380_n4894), .B(core__abc_21380_n1708), .Y(core__abc_21380_n4938) );
  OR2X2 OR2X2_1881 ( .A(core__abc_21380_n4940), .B(core__abc_21380_n4941), .Y(core__abc_21380_n4942) );
  OR2X2 OR2X2_1882 ( .A(core__abc_21380_n4945), .B(core__abc_21380_n4943), .Y(core__abc_21380_n4946) );
  OR2X2 OR2X2_1883 ( .A(core__abc_21380_n4936), .B(core__abc_21380_n4946), .Y(core__abc_21380_n4947) );
  OR2X2 OR2X2_1884 ( .A(core__abc_21380_n4928), .B(core__abc_21380_n4950), .Y(core__abc_21380_n4951) );
  OR2X2 OR2X2_1885 ( .A(core__abc_21380_n4952), .B(core__abc_21380_n4953), .Y(core__abc_21380_n4954) );
  OR2X2 OR2X2_1886 ( .A(core__abc_21380_n4956), .B(core__abc_21380_n3548_1), .Y(core__abc_21380_n4957) );
  OR2X2 OR2X2_1887 ( .A(core__abc_21380_n4955), .B(core__abc_21380_n3547), .Y(core__abc_21380_n4958) );
  OR2X2 OR2X2_1888 ( .A(core_v3_reg_25_), .B(core_mi_25_), .Y(core__abc_21380_n4962) );
  OR2X2 OR2X2_1889 ( .A(core__abc_21380_n4961), .B(core__abc_21380_n4966), .Y(core__abc_21380_n4967) );
  OR2X2 OR2X2_189 ( .A(_abc_19068_n1305), .B(_abc_19068_n1292), .Y(_abc_19068_n1306_1) );
  OR2X2 OR2X2_1890 ( .A(core__abc_21380_n3317_bF_buf5), .B(core__abc_21380_n4967), .Y(core__abc_21380_n4968) );
  OR2X2 OR2X2_1891 ( .A(core__abc_21380_n4960), .B(core__abc_21380_n4968), .Y(core__abc_21380_n4969) );
  OR2X2 OR2X2_1892 ( .A(core__abc_21380_n3328_bF_buf6), .B(core_v3_reg_25_), .Y(core__abc_21380_n4970) );
  OR2X2 OR2X2_1893 ( .A(core__abc_21380_n4929), .B(core__abc_21380_n2323), .Y(core__abc_21380_n4973) );
  OR2X2 OR2X2_1894 ( .A(core__abc_21380_n4934), .B(core__abc_21380_n4973), .Y(core__abc_21380_n4974) );
  OR2X2 OR2X2_1895 ( .A(core__abc_21380_n4977), .B(core__abc_21380_n4975), .Y(core__abc_21380_n4978) );
  OR2X2 OR2X2_1896 ( .A(core__abc_21380_n4981), .B(core__abc_21380_n3098), .Y(core__abc_21380_n4982) );
  OR2X2 OR2X2_1897 ( .A(core__abc_21380_n4984), .B(core__abc_21380_n4985), .Y(core__abc_21380_n4986) );
  OR2X2 OR2X2_1898 ( .A(core__abc_21380_n4987), .B(core__abc_21380_n4980), .Y(core__abc_21380_n4988) );
  OR2X2 OR2X2_1899 ( .A(core__abc_21380_n4986), .B(core_v3_reg_10_), .Y(core__abc_21380_n4989) );
  OR2X2 OR2X2_19 ( .A(_abc_19068_n940_1), .B(_abc_19068_n942_1), .Y(_abc_19068_n943_1) );
  OR2X2 OR2X2_190 ( .A(_abc_19068_n1308_1), .B(_abc_19068_n1309), .Y(_abc_19068_n1310_1) );
  OR2X2 OR2X2_1900 ( .A(core__abc_21380_n4992), .B(core__abc_21380_n4993), .Y(core__abc_21380_n4994) );
  OR2X2 OR2X2_1901 ( .A(core__abc_21380_n4995), .B(core__abc_21380_n4948), .Y(core__abc_21380_n4996) );
  OR2X2 OR2X2_1902 ( .A(core__abc_21380_n4866), .B(core__abc_21380_n4998), .Y(core__abc_21380_n4999) );
  OR2X2 OR2X2_1903 ( .A(core__abc_21380_n5000), .B(core__abc_21380_n4994), .Y(core__abc_21380_n5002) );
  OR2X2 OR2X2_1904 ( .A(core__abc_21380_n5003), .B(core__abc_21380_n5001), .Y(core__abc_21380_n5004) );
  OR2X2 OR2X2_1905 ( .A(core__abc_21380_n5004), .B(core__abc_21380_n3614), .Y(core__abc_21380_n5005) );
  OR2X2 OR2X2_1906 ( .A(core__abc_21380_n5006), .B(core__abc_21380_n3615), .Y(core__abc_21380_n5007) );
  OR2X2 OR2X2_1907 ( .A(core_v3_reg_26_), .B(core_mi_26_), .Y(core__abc_21380_n5011) );
  OR2X2 OR2X2_1908 ( .A(core__abc_21380_n5010), .B(core__abc_21380_n5015), .Y(core__abc_21380_n5016) );
  OR2X2 OR2X2_1909 ( .A(core__abc_21380_n3317_bF_buf4), .B(core__abc_21380_n5016), .Y(core__abc_21380_n5017) );
  OR2X2 OR2X2_191 ( .A(_abc_19068_n909_1), .B(_abc_19068_n1311), .Y(_abc_19068_n1312_1) );
  OR2X2 OR2X2_1910 ( .A(core__abc_21380_n5009), .B(core__abc_21380_n5017), .Y(core__abc_21380_n5018) );
  OR2X2 OR2X2_1911 ( .A(core__abc_21380_n3328_bF_buf5), .B(core_v3_reg_26_), .Y(core__abc_21380_n5019) );
  OR2X2 OR2X2_1912 ( .A(core__abc_21380_n4975), .B(core__abc_21380_n2341), .Y(core__abc_21380_n5025) );
  OR2X2 OR2X2_1913 ( .A(core__abc_21380_n4985), .B(core__abc_21380_n1744), .Y(core__abc_21380_n5033) );
  OR2X2 OR2X2_1914 ( .A(core__abc_21380_n5035), .B(core__abc_21380_n5036), .Y(core__abc_21380_n5037) );
  OR2X2 OR2X2_1915 ( .A(core__abc_21380_n5037), .B(core__abc_21380_n5032), .Y(core__abc_21380_n5040) );
  OR2X2 OR2X2_1916 ( .A(core__abc_21380_n5027), .B(core__abc_21380_n5029), .Y(core__abc_21380_n5043) );
  OR2X2 OR2X2_1917 ( .A(core__abc_21380_n5044), .B(core__abc_21380_n5038), .Y(core__abc_21380_n5045) );
  OR2X2 OR2X2_1918 ( .A(core__abc_21380_n5042), .B(core__abc_21380_n5046), .Y(core__abc_21380_n5047) );
  OR2X2 OR2X2_1919 ( .A(core__abc_21380_n5024), .B(core__abc_21380_n5047), .Y(core__abc_21380_n5048) );
  OR2X2 OR2X2_192 ( .A(_abc_19068_n1312_1), .B(_abc_19068_n1310_1), .Y(_abc_19068_n1313) );
  OR2X2 OR2X2_1920 ( .A(core__abc_21380_n5045), .B(core__abc_21380_n5043), .Y(core__abc_21380_n5050) );
  OR2X2 OR2X2_1921 ( .A(core__abc_21380_n5031), .B(core__abc_21380_n5041), .Y(core__abc_21380_n5051) );
  OR2X2 OR2X2_1922 ( .A(core__abc_21380_n5049), .B(core__abc_21380_n5052), .Y(core__abc_21380_n5053) );
  OR2X2 OR2X2_1923 ( .A(core__abc_21380_n5054), .B(core__abc_21380_n5022), .Y(core__abc_21380_n5055) );
  OR2X2 OR2X2_1924 ( .A(core__abc_21380_n5056), .B(core__abc_21380_n3697), .Y(core__abc_21380_n5057) );
  OR2X2 OR2X2_1925 ( .A(core_v3_reg_27_), .B(core_mi_27_), .Y(core__abc_21380_n5062) );
  OR2X2 OR2X2_1926 ( .A(core__abc_21380_n5061), .B(core__abc_21380_n5066), .Y(core__abc_21380_n5067) );
  OR2X2 OR2X2_1927 ( .A(core__abc_21380_n3317_bF_buf3), .B(core__abc_21380_n5067), .Y(core__abc_21380_n5068) );
  OR2X2 OR2X2_1928 ( .A(core__abc_21380_n5059), .B(core__abc_21380_n5068), .Y(core__abc_21380_n5069) );
  OR2X2 OR2X2_1929 ( .A(core__abc_21380_n3328_bF_buf4), .B(core_v3_reg_27_), .Y(core__abc_21380_n5070) );
  OR2X2 OR2X2_193 ( .A(_abc_19068_n1315), .B(_abc_19068_n1316_1), .Y(_abc_19068_n1317) );
  OR2X2 OR2X2_1930 ( .A(core__abc_21380_n5077), .B(core__abc_21380_n5042), .Y(core__abc_21380_n5078) );
  OR2X2 OR2X2_1931 ( .A(core__abc_21380_n5076), .B(core__abc_21380_n5078), .Y(core__abc_21380_n5079) );
  OR2X2 OR2X2_1932 ( .A(core__abc_21380_n5081), .B(core__abc_21380_n5079), .Y(core__abc_21380_n5082) );
  OR2X2 OR2X2_1933 ( .A(core__abc_21380_n5088), .B(core__abc_21380_n2360), .Y(core__abc_21380_n5089) );
  OR2X2 OR2X2_1934 ( .A(core__abc_21380_n5087), .B(core__abc_21380_n5089), .Y(core__abc_21380_n5090) );
  OR2X2 OR2X2_1935 ( .A(core__abc_21380_n5086), .B(core__abc_21380_n5090), .Y(core__abc_21380_n5091) );
  OR2X2 OR2X2_1936 ( .A(core__abc_21380_n4880), .B(core__abc_21380_n5093), .Y(core__abc_21380_n5094) );
  OR2X2 OR2X2_1937 ( .A(core__abc_21380_n5097), .B(core__abc_21380_n5092), .Y(core__abc_21380_n5098) );
  OR2X2 OR2X2_1938 ( .A(core__abc_21380_n4891), .B(core__abc_21380_n5102), .Y(core__abc_21380_n5103) );
  OR2X2 OR2X2_1939 ( .A(core__abc_21380_n5106), .B(core__abc_21380_n5107), .Y(core__abc_21380_n5108) );
  OR2X2 OR2X2_194 ( .A(_abc_19068_n1317), .B(_abc_19068_n1314_1), .Y(_abc_19068_n1318_1) );
  OR2X2 OR2X2_1940 ( .A(core__abc_21380_n5109), .B(core__abc_21380_n5100), .Y(core__abc_21380_n5110) );
  OR2X2 OR2X2_1941 ( .A(core__abc_21380_n5108), .B(core_v3_reg_12_), .Y(core__abc_21380_n5111) );
  OR2X2 OR2X2_1942 ( .A(core__abc_21380_n5114), .B(core__abc_21380_n5115), .Y(core__abc_21380_n5116) );
  OR2X2 OR2X2_1943 ( .A(core__abc_21380_n5117), .B(core__abc_21380_n5119), .Y(core__abc_21380_n5120) );
  OR2X2 OR2X2_1944 ( .A(core__abc_21380_n5120), .B(core__abc_21380_n3756_1), .Y(core__abc_21380_n5121) );
  OR2X2 OR2X2_1945 ( .A(core__abc_21380_n5122), .B(core__abc_21380_n3761), .Y(core__abc_21380_n5123) );
  OR2X2 OR2X2_1946 ( .A(core_v3_reg_28_), .B(core_mi_28_), .Y(core__abc_21380_n5128) );
  OR2X2 OR2X2_1947 ( .A(core__abc_21380_n5127), .B(core__abc_21380_n5132), .Y(core__abc_21380_n5133) );
  OR2X2 OR2X2_1948 ( .A(core__abc_21380_n3317_bF_buf2), .B(core__abc_21380_n5133), .Y(core__abc_21380_n5134) );
  OR2X2 OR2X2_1949 ( .A(core__abc_21380_n5125), .B(core__abc_21380_n5134), .Y(core__abc_21380_n5135) );
  OR2X2 OR2X2_195 ( .A(_abc_19068_n1319), .B(_abc_19068_n1320_1), .Y(_abc_19068_n1321) );
  OR2X2 OR2X2_1950 ( .A(core__abc_21380_n3328_bF_buf3), .B(core_v3_reg_28_), .Y(core__abc_21380_n5136) );
  OR2X2 OR2X2_1951 ( .A(core__abc_21380_n5143), .B(core__abc_21380_n5141), .Y(core__abc_21380_n5144) );
  OR2X2 OR2X2_1952 ( .A(core__abc_21380_n2399), .B(core__abc_21380_n2379), .Y(core__abc_21380_n5145) );
  OR2X2 OR2X2_1953 ( .A(core__abc_21380_n5092), .B(core__abc_21380_n5145), .Y(core__abc_21380_n5146) );
  OR2X2 OR2X2_1954 ( .A(core__abc_21380_n5147), .B(core__abc_21380_n5144), .Y(core__abc_21380_n5148) );
  OR2X2 OR2X2_1955 ( .A(core__abc_21380_n5106), .B(core__abc_21380_n1783), .Y(core__abc_21380_n5151) );
  OR2X2 OR2X2_1956 ( .A(core__abc_21380_n5153), .B(core__abc_21380_n5154), .Y(core__abc_21380_n5155) );
  OR2X2 OR2X2_1957 ( .A(core__abc_21380_n5155), .B(core__abc_21380_n5150), .Y(core__abc_21380_n5158) );
  OR2X2 OR2X2_1958 ( .A(core__abc_21380_n5161), .B(core__abc_21380_n5156), .Y(core__abc_21380_n5162) );
  OR2X2 OR2X2_1959 ( .A(core__abc_21380_n5163), .B(core__abc_21380_n5160), .Y(core__abc_21380_n5164) );
  OR2X2 OR2X2_196 ( .A(_abc_19068_n1322_1), .B(_abc_19068_n1323), .Y(_abc_19068_n1324_1) );
  OR2X2 OR2X2_1960 ( .A(core__abc_21380_n5164), .B(core__abc_21380_n5140), .Y(core__abc_21380_n5168) );
  OR2X2 OR2X2_1961 ( .A(core__abc_21380_n5162), .B(core__abc_21380_n5148), .Y(core__abc_21380_n5169) );
  OR2X2 OR2X2_1962 ( .A(core__abc_21380_n5159), .B(core__abc_21380_n5149), .Y(core__abc_21380_n5170) );
  OR2X2 OR2X2_1963 ( .A(core__abc_21380_n5176), .B(core__abc_21380_n3825), .Y(core__abc_21380_n5177) );
  OR2X2 OR2X2_1964 ( .A(core__abc_21380_n5178), .B(core__abc_21380_n3824), .Y(core__abc_21380_n5179) );
  OR2X2 OR2X2_1965 ( .A(core_v3_reg_29_), .B(core_mi_29_), .Y(core__abc_21380_n5184) );
  OR2X2 OR2X2_1966 ( .A(core__abc_21380_n5183), .B(core__abc_21380_n5188), .Y(core__abc_21380_n5189) );
  OR2X2 OR2X2_1967 ( .A(core__abc_21380_n3317_bF_buf1), .B(core__abc_21380_n5189), .Y(core__abc_21380_n5190) );
  OR2X2 OR2X2_1968 ( .A(core__abc_21380_n5181), .B(core__abc_21380_n5190), .Y(core__abc_21380_n5191) );
  OR2X2 OR2X2_1969 ( .A(core__abc_21380_n3328_bF_buf2), .B(core_v3_reg_29_), .Y(core__abc_21380_n5192) );
  OR2X2 OR2X2_197 ( .A(_abc_19068_n1321), .B(_abc_19068_n1324_1), .Y(_abc_19068_n1325) );
  OR2X2 OR2X2_1970 ( .A(core__abc_21380_n5096), .B(core__abc_21380_n5198), .Y(core__abc_21380_n5199) );
  OR2X2 OR2X2_1971 ( .A(core__abc_21380_n5141), .B(core__abc_21380_n2397), .Y(core__abc_21380_n5200) );
  OR2X2 OR2X2_1972 ( .A(core__abc_21380_n5143), .B(core__abc_21380_n5200), .Y(core__abc_21380_n5204) );
  OR2X2 OR2X2_1973 ( .A(core__abc_21380_n5203), .B(core__abc_21380_n5205), .Y(core__abc_21380_n5206) );
  OR2X2 OR2X2_1974 ( .A(core__abc_21380_n5104), .B(core__abc_21380_n5208), .Y(core__abc_21380_n5209) );
  OR2X2 OR2X2_1975 ( .A(core__abc_21380_n5210), .B(core__abc_21380_n1826), .Y(core__abc_21380_n5212) );
  OR2X2 OR2X2_1976 ( .A(core__abc_21380_n5213), .B(core__abc_21380_n5211), .Y(core__abc_21380_n5214) );
  OR2X2 OR2X2_1977 ( .A(core__abc_21380_n5215), .B(core_v3_reg_14_), .Y(core__abc_21380_n5216) );
  OR2X2 OR2X2_1978 ( .A(core__abc_21380_n5214), .B(core__abc_21380_n5217), .Y(core__abc_21380_n5218) );
  OR2X2 OR2X2_1979 ( .A(core__abc_21380_n5222), .B(core__abc_21380_n5220), .Y(core__abc_21380_n5223) );
  OR2X2 OR2X2_198 ( .A(_abc_19068_n1325), .B(_abc_19068_n1318_1), .Y(_abc_19068_n1326_1) );
  OR2X2 OR2X2_1980 ( .A(core__abc_21380_n5197), .B(core__abc_21380_n5223), .Y(core__abc_21380_n5225) );
  OR2X2 OR2X2_1981 ( .A(core__abc_21380_n5226), .B(core__abc_21380_n5224), .Y(core__abc_21380_n5227) );
  OR2X2 OR2X2_1982 ( .A(core__abc_21380_n5228), .B(core__abc_21380_n5195), .Y(core__abc_21380_n5229) );
  OR2X2 OR2X2_1983 ( .A(core__abc_21380_n5227), .B(core__abc_21380_n3900), .Y(core__abc_21380_n5230) );
  OR2X2 OR2X2_1984 ( .A(core_v3_reg_30_), .B(core_mi_30_), .Y(core__abc_21380_n5235) );
  OR2X2 OR2X2_1985 ( .A(core__abc_21380_n5234), .B(core__abc_21380_n5239), .Y(core__abc_21380_n5240) );
  OR2X2 OR2X2_1986 ( .A(core__abc_21380_n3317_bF_buf0), .B(core__abc_21380_n5240), .Y(core__abc_21380_n5241) );
  OR2X2 OR2X2_1987 ( .A(core__abc_21380_n5232), .B(core__abc_21380_n5241), .Y(core__abc_21380_n5242) );
  OR2X2 OR2X2_1988 ( .A(core__abc_21380_n3328_bF_buf1), .B(core_v3_reg_30_), .Y(core__abc_21380_n5243) );
  OR2X2 OR2X2_1989 ( .A(core__abc_21380_n5202), .B(core__abc_21380_n2416), .Y(core__abc_21380_n5250) );
  OR2X2 OR2X2_199 ( .A(_abc_19068_n1326_1), .B(_abc_19068_n1313), .Y(_abc_19068_n1327) );
  OR2X2 OR2X2_1990 ( .A(core__abc_21380_n5205), .B(core__abc_21380_n2415), .Y(core__abc_21380_n5253) );
  OR2X2 OR2X2_1991 ( .A(core__abc_21380_n5252), .B(core__abc_21380_n5254), .Y(core__abc_21380_n5255) );
  OR2X2 OR2X2_1992 ( .A(core__abc_21380_n5257), .B(core__abc_21380_n1846_1), .Y(core__abc_21380_n5259) );
  OR2X2 OR2X2_1993 ( .A(core__abc_21380_n5260), .B(core__abc_21380_n5258), .Y(core__abc_21380_n5261) );
  OR2X2 OR2X2_1994 ( .A(core__abc_21380_n5262), .B(core__abc_21380_n5265), .Y(core__abc_21380_n5266) );
  OR2X2 OR2X2_1995 ( .A(core__abc_21380_n5255), .B(core__abc_21380_n5266), .Y(core__abc_21380_n5267) );
  OR2X2 OR2X2_1996 ( .A(core__abc_21380_n5253), .B(core__abc_21380_n2435), .Y(core__abc_21380_n5268) );
  OR2X2 OR2X2_1997 ( .A(core__abc_21380_n5251), .B(core__abc_21380_n2434), .Y(core__abc_21380_n5269) );
  OR2X2 OR2X2_1998 ( .A(core__abc_21380_n5264), .B(core_v3_reg_15_), .Y(core__abc_21380_n5271) );
  OR2X2 OR2X2_1999 ( .A(core__abc_21380_n5270), .B(core__abc_21380_n5273), .Y(core__abc_21380_n5274) );
  OR2X2 OR2X2_2 ( .A(_abc_19068_n890), .B(_abc_19068_n882_1), .Y(_abc_19068_n891_1) );
  OR2X2 OR2X2_20 ( .A(_abc_19068_n944), .B(_abc_19068_n946_1), .Y(_abc_19068_n947) );
  OR2X2 OR2X2_200 ( .A(_abc_19068_n1330_1), .B(_abc_19068_n1331), .Y(_abc_19068_n1332_1) );
  OR2X2 OR2X2_2000 ( .A(core__abc_21380_n5248), .B(core__abc_21380_n5275), .Y(core__abc_21380_n5276) );
  OR2X2 OR2X2_2001 ( .A(core__abc_21380_n5255), .B(core__abc_21380_n5273), .Y(core__abc_21380_n5277) );
  OR2X2 OR2X2_2002 ( .A(core__abc_21380_n5270), .B(core__abc_21380_n5266), .Y(core__abc_21380_n5278) );
  OR2X2 OR2X2_2003 ( .A(core__abc_21380_n5247), .B(core__abc_21380_n5279), .Y(core__abc_21380_n5280) );
  OR2X2 OR2X2_2004 ( .A(core__abc_21380_n5281), .B(core__abc_21380_n3965_1), .Y(core__abc_21380_n5282) );
  OR2X2 OR2X2_2005 ( .A(core__abc_21380_n5283), .B(core__abc_21380_n3964), .Y(core__abc_21380_n5284) );
  OR2X2 OR2X2_2006 ( .A(core_v3_reg_31_), .B(core_mi_31_), .Y(core__abc_21380_n5288) );
  OR2X2 OR2X2_2007 ( .A(core__abc_21380_n5287), .B(core__abc_21380_n5292), .Y(core__abc_21380_n5293) );
  OR2X2 OR2X2_2008 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n5293), .Y(core__abc_21380_n5294) );
  OR2X2 OR2X2_2009 ( .A(core__abc_21380_n5286), .B(core__abc_21380_n5294), .Y(core__abc_21380_n5295) );
  OR2X2 OR2X2_201 ( .A(_abc_19068_n1332_1), .B(_abc_19068_n1329), .Y(_abc_19068_n1333) );
  OR2X2 OR2X2_2010 ( .A(core__abc_21380_n3328_bF_buf0), .B(core_v3_reg_31_), .Y(core__abc_21380_n5296) );
  OR2X2 OR2X2_2011 ( .A(core__abc_21380_n5279), .B(core__abc_21380_n5223), .Y(core__abc_21380_n5301) );
  OR2X2 OR2X2_2012 ( .A(core__abc_21380_n5301), .B(core__abc_21380_n5300), .Y(core__abc_21380_n5302) );
  OR2X2 OR2X2_2013 ( .A(core__abc_21380_n5302), .B(core__abc_21380_n5299), .Y(core__abc_21380_n5303) );
  OR2X2 OR2X2_2014 ( .A(core__abc_21380_n4856), .B(core__abc_21380_n5303), .Y(core__abc_21380_n5304) );
  OR2X2 OR2X2_2015 ( .A(core__abc_21380_n5303), .B(core__abc_21380_n4865), .Y(core__abc_21380_n5305) );
  OR2X2 OR2X2_2016 ( .A(core__abc_21380_n5047), .B(core__abc_21380_n4994), .Y(core__abc_21380_n5306) );
  OR2X2 OR2X2_2017 ( .A(core__abc_21380_n5306), .B(core__abc_21380_n4996), .Y(core__abc_21380_n5307) );
  OR2X2 OR2X2_2018 ( .A(core__abc_21380_n5302), .B(core__abc_21380_n5309), .Y(core__abc_21380_n5310) );
  OR2X2 OR2X2_2019 ( .A(core__abc_21380_n5301), .B(core__abc_21380_n5196), .Y(core__abc_21380_n5311) );
  OR2X2 OR2X2_202 ( .A(_abc_19068_n1334_1), .B(_abc_19068_n1038_1), .Y(_abc_19068_n1335) );
  OR2X2 OR2X2_2020 ( .A(core__abc_21380_n5313), .B(core__abc_21380_n5312), .Y(core__abc_21380_n5314) );
  OR2X2 OR2X2_2021 ( .A(core__abc_21380_n5322), .B(core__abc_21380_n5323), .Y(core__abc_21380_n5324) );
  OR2X2 OR2X2_2022 ( .A(core__abc_21380_n5325), .B(core__abc_21380_n5320), .Y(core__abc_21380_n5326) );
  OR2X2 OR2X2_2023 ( .A(core__abc_21380_n5324), .B(core_v3_reg_16_), .Y(core__abc_21380_n5327) );
  OR2X2 OR2X2_2024 ( .A(core__abc_21380_n5330), .B(core__abc_21380_n5331), .Y(core__abc_21380_n5332) );
  OR2X2 OR2X2_2025 ( .A(core__abc_21380_n5342), .B(core__abc_21380_n4862_1), .Y(core__abc_21380_n5343) );
  OR2X2 OR2X2_2026 ( .A(core__abc_21380_n5343), .B(core__abc_21380_n5340), .Y(core__abc_21380_n5344) );
  OR2X2 OR2X2_2027 ( .A(core__abc_21380_n5347), .B(core__abc_21380_n5160), .Y(core__abc_21380_n5348) );
  OR2X2 OR2X2_2028 ( .A(core__abc_21380_n5349), .B(core__abc_21380_n5314), .Y(core__abc_21380_n5350) );
  OR2X2 OR2X2_2029 ( .A(core__abc_21380_n5350), .B(core__abc_21380_n5346), .Y(core__abc_21380_n5351) );
  OR2X2 OR2X2_203 ( .A(_abc_19068_n1336_1), .B(_abc_19068_n1337), .Y(_abc_19068_n1338_1) );
  OR2X2 OR2X2_2030 ( .A(core__abc_21380_n5351), .B(core__abc_21380_n5345), .Y(core__abc_21380_n5352) );
  OR2X2 OR2X2_2031 ( .A(core__abc_21380_n5352), .B(core__abc_21380_n5339), .Y(core__abc_21380_n5353) );
  OR2X2 OR2X2_2032 ( .A(core__abc_21380_n5333), .B(core__abc_21380_n5355), .Y(core__abc_21380_n5356) );
  OR2X2 OR2X2_2033 ( .A(core__abc_21380_n5356), .B(core__abc_21380_n4021), .Y(core__abc_21380_n5357) );
  OR2X2 OR2X2_2034 ( .A(core__abc_21380_n5358), .B(core__abc_21380_n4073), .Y(core__abc_21380_n5359) );
  OR2X2 OR2X2_2035 ( .A(core_v3_reg_32_), .B(core_mi_32_), .Y(core__abc_21380_n5363) );
  OR2X2 OR2X2_2036 ( .A(core__abc_21380_n5362), .B(core__abc_21380_n5367), .Y(core__abc_21380_n5368) );
  OR2X2 OR2X2_2037 ( .A(core__abc_21380_n3317_bF_buf6), .B(core__abc_21380_n5368), .Y(core__abc_21380_n5369) );
  OR2X2 OR2X2_2038 ( .A(core__abc_21380_n5361), .B(core__abc_21380_n5369), .Y(core__abc_21380_n5370) );
  OR2X2 OR2X2_2039 ( .A(core__abc_21380_n3328_bF_buf7), .B(core_v3_reg_32_), .Y(core__abc_21380_n5371) );
  OR2X2 OR2X2_204 ( .A(_abc_19068_n1338_1), .B(_abc_19068_n1335), .Y(_abc_19068_n1339) );
  OR2X2 OR2X2_2040 ( .A(core__abc_21380_n5374), .B(core__abc_21380_n3168), .Y(core__abc_21380_n5375) );
  OR2X2 OR2X2_2041 ( .A(core__abc_21380_n5322), .B(core__abc_21380_n1859), .Y(core__abc_21380_n5378) );
  OR2X2 OR2X2_2042 ( .A(core__abc_21380_n5380), .B(core__abc_21380_n5381), .Y(core__abc_21380_n5382) );
  OR2X2 OR2X2_2043 ( .A(core__abc_21380_n5385), .B(core__abc_21380_n5383), .Y(core__abc_21380_n5386) );
  OR2X2 OR2X2_2044 ( .A(core__abc_21380_n5388), .B(core__abc_21380_n5389), .Y(core__abc_21380_n5390) );
  OR2X2 OR2X2_2045 ( .A(core__abc_21380_n5393), .B(core__abc_21380_n5390), .Y(core__abc_21380_n5395) );
  OR2X2 OR2X2_2046 ( .A(core__abc_21380_n5396), .B(core__abc_21380_n5394), .Y(core__abc_21380_n5397) );
  OR2X2 OR2X2_2047 ( .A(core__abc_21380_n5398), .B(core__abc_21380_n4111_1), .Y(core__abc_21380_n5399) );
  OR2X2 OR2X2_2048 ( .A(core__abc_21380_n5397), .B(core__abc_21380_n4110), .Y(core__abc_21380_n5400) );
  OR2X2 OR2X2_2049 ( .A(core_v3_reg_33_), .B(core_mi_33_), .Y(core__abc_21380_n5405) );
  OR2X2 OR2X2_205 ( .A(_abc_19068_n1340_1), .B(_abc_19068_n1341), .Y(_abc_19068_n1342_1) );
  OR2X2 OR2X2_2050 ( .A(core__abc_21380_n5404), .B(core__abc_21380_n5409), .Y(core__abc_21380_n5410) );
  OR2X2 OR2X2_2051 ( .A(core__abc_21380_n3317_bF_buf5), .B(core__abc_21380_n5410), .Y(core__abc_21380_n5411) );
  OR2X2 OR2X2_2052 ( .A(core__abc_21380_n5402), .B(core__abc_21380_n5411), .Y(core__abc_21380_n5412) );
  OR2X2 OR2X2_2053 ( .A(core__abc_21380_n3328_bF_buf6), .B(core_v3_reg_33_), .Y(core__abc_21380_n5413) );
  OR2X2 OR2X2_2054 ( .A(core__abc_21380_n5420), .B(core__abc_21380_n5388), .Y(core__abc_21380_n5421) );
  OR2X2 OR2X2_2055 ( .A(core__abc_21380_n5425), .B(core__abc_21380_n5424), .Y(core__abc_21380_n5426) );
  OR2X2 OR2X2_2056 ( .A(core__abc_21380_n3115), .B(core__abc_21380_n5429), .Y(core__abc_21380_n5430) );
  OR2X2 OR2X2_2057 ( .A(core__abc_21380_n5431), .B(core__abc_21380_n1900), .Y(core__abc_21380_n5433) );
  OR2X2 OR2X2_2058 ( .A(core__abc_21380_n5434), .B(core__abc_21380_n5432), .Y(core__abc_21380_n5435) );
  OR2X2 OR2X2_2059 ( .A(core__abc_21380_n5436), .B(core__abc_21380_n5428), .Y(core__abc_21380_n5437) );
  OR2X2 OR2X2_206 ( .A(_abc_19068_n1343), .B(_abc_19068_n1344_1), .Y(_abc_19068_n1345) );
  OR2X2 OR2X2_2060 ( .A(core__abc_21380_n5435), .B(core_v3_reg_18_), .Y(core__abc_21380_n5438) );
  OR2X2 OR2X2_2061 ( .A(core__abc_21380_n5441), .B(core__abc_21380_n5442), .Y(core__abc_21380_n5443) );
  OR2X2 OR2X2_2062 ( .A(core__abc_21380_n5423), .B(core__abc_21380_n5443), .Y(core__abc_21380_n5445) );
  OR2X2 OR2X2_2063 ( .A(core__abc_21380_n5446), .B(core__abc_21380_n5444), .Y(core__abc_21380_n5447) );
  OR2X2 OR2X2_2064 ( .A(core__abc_21380_n5447), .B(core__abc_21380_n4170_1), .Y(core__abc_21380_n5448) );
  OR2X2 OR2X2_2065 ( .A(core__abc_21380_n5449), .B(core__abc_21380_n4171), .Y(core__abc_21380_n5450) );
  OR2X2 OR2X2_2066 ( .A(core_v3_reg_34_), .B(core_mi_34_), .Y(core__abc_21380_n5454) );
  OR2X2 OR2X2_2067 ( .A(core__abc_21380_n5453), .B(core__abc_21380_n5458), .Y(core__abc_21380_n5459) );
  OR2X2 OR2X2_2068 ( .A(core__abc_21380_n3317_bF_buf4), .B(core__abc_21380_n5459), .Y(core__abc_21380_n5460) );
  OR2X2 OR2X2_2069 ( .A(core__abc_21380_n5452), .B(core__abc_21380_n5460), .Y(core__abc_21380_n5461) );
  OR2X2 OR2X2_207 ( .A(_abc_19068_n1342_1), .B(_abc_19068_n1345), .Y(_abc_19068_n1346_1) );
  OR2X2 OR2X2_2070 ( .A(core__abc_21380_n3328_bF_buf5), .B(core_v3_reg_34_), .Y(core__abc_21380_n5462) );
  OR2X2 OR2X2_2071 ( .A(core__abc_21380_n5424), .B(core__abc_21380_n1301), .Y(core__abc_21380_n5468) );
  OR2X2 OR2X2_2072 ( .A(core__abc_21380_n5470), .B(core__abc_21380_n5471), .Y(core__abc_21380_n5472) );
  OR2X2 OR2X2_2073 ( .A(core__abc_21380_n5475), .B(core__abc_21380_n1920), .Y(core__abc_21380_n5478) );
  OR2X2 OR2X2_2074 ( .A(core__abc_21380_n5481), .B(core__abc_21380_n5482), .Y(core__abc_21380_n5483) );
  OR2X2 OR2X2_2075 ( .A(core__abc_21380_n5485), .B(core__abc_21380_n5486), .Y(core__abc_21380_n5487) );
  OR2X2 OR2X2_2076 ( .A(core__abc_21380_n5467), .B(core__abc_21380_n5488), .Y(core__abc_21380_n5489) );
  OR2X2 OR2X2_2077 ( .A(core__abc_21380_n5466), .B(core__abc_21380_n5487), .Y(core__abc_21380_n5490) );
  OR2X2 OR2X2_2078 ( .A(core__abc_21380_n5491), .B(core__abc_21380_n4247), .Y(core__abc_21380_n5492) );
  OR2X2 OR2X2_2079 ( .A(core__abc_21380_n5493), .B(core__abc_21380_n4246), .Y(core__abc_21380_n5494) );
  OR2X2 OR2X2_208 ( .A(_abc_19068_n1346_1), .B(_abc_19068_n1339), .Y(_abc_19068_n1347) );
  OR2X2 OR2X2_2080 ( .A(core_v3_reg_35_), .B(core_mi_35_), .Y(core__abc_21380_n5498) );
  OR2X2 OR2X2_2081 ( .A(core__abc_21380_n5497), .B(core__abc_21380_n5502), .Y(core__abc_21380_n5503) );
  OR2X2 OR2X2_2082 ( .A(core__abc_21380_n3317_bF_buf3), .B(core__abc_21380_n5503), .Y(core__abc_21380_n5504) );
  OR2X2 OR2X2_2083 ( .A(core__abc_21380_n5496), .B(core__abc_21380_n5504), .Y(core__abc_21380_n5505) );
  OR2X2 OR2X2_2084 ( .A(core__abc_21380_n3328_bF_buf4), .B(core_v3_reg_35_), .Y(core__abc_21380_n5506) );
  OR2X2 OR2X2_2085 ( .A(core__abc_21380_n5487), .B(core__abc_21380_n5443), .Y(core__abc_21380_n5509) );
  OR2X2 OR2X2_2086 ( .A(core__abc_21380_n5486), .B(core__abc_21380_n5465), .Y(core__abc_21380_n5513) );
  OR2X2 OR2X2_2087 ( .A(core__abc_21380_n5511), .B(core__abc_21380_n5515), .Y(core__abc_21380_n5516) );
  OR2X2 OR2X2_2088 ( .A(core__abc_21380_n5518), .B(core__abc_21380_n5516), .Y(core__abc_21380_n5519) );
  OR2X2 OR2X2_2089 ( .A(core__abc_21380_n5521), .B(core__abc_21380_n5520), .Y(core__abc_21380_n5522) );
  OR2X2 OR2X2_209 ( .A(_abc_19068_n1347), .B(_abc_19068_n1333), .Y(_abc_19068_n1348_1) );
  OR2X2 OR2X2_2090 ( .A(core__abc_21380_n5525), .B(core__abc_21380_n3132), .Y(core__abc_21380_n5526) );
  OR2X2 OR2X2_2091 ( .A(core__abc_21380_n5529), .B(core__abc_21380_n5527), .Y(core__abc_21380_n5530) );
  OR2X2 OR2X2_2092 ( .A(core__abc_21380_n5531), .B(core__abc_21380_n5524), .Y(core__abc_21380_n5532) );
  OR2X2 OR2X2_2093 ( .A(core__abc_21380_n5530), .B(core_v3_reg_20_), .Y(core__abc_21380_n5533) );
  OR2X2 OR2X2_2094 ( .A(core__abc_21380_n5536), .B(core__abc_21380_n5537), .Y(core__abc_21380_n5538) );
  OR2X2 OR2X2_2095 ( .A(core__abc_21380_n5542), .B(core__abc_21380_n5540), .Y(core__abc_21380_n5543) );
  OR2X2 OR2X2_2096 ( .A(core__abc_21380_n5543), .B(core__abc_21380_n4310), .Y(core__abc_21380_n5544) );
  OR2X2 OR2X2_2097 ( .A(core__abc_21380_n5545), .B(core__abc_21380_n4311), .Y(core__abc_21380_n5546) );
  OR2X2 OR2X2_2098 ( .A(core_v3_reg_36_), .B(core_mi_36_), .Y(core__abc_21380_n5550) );
  OR2X2 OR2X2_2099 ( .A(core__abc_21380_n5549), .B(core__abc_21380_n5554), .Y(core__abc_21380_n5555) );
  OR2X2 OR2X2_21 ( .A(_abc_19068_n948_1), .B(_abc_19068_n949_1), .Y(_abc_19068_n950) );
  OR2X2 OR2X2_210 ( .A(_abc_19068_n1209_1), .B(_abc_19068_n1350_1), .Y(_abc_19068_n1351) );
  OR2X2 OR2X2_2100 ( .A(core__abc_21380_n3317_bF_buf2), .B(core__abc_21380_n5555), .Y(core__abc_21380_n5556) );
  OR2X2 OR2X2_2101 ( .A(core__abc_21380_n5548), .B(core__abc_21380_n5556), .Y(core__abc_21380_n5557) );
  OR2X2 OR2X2_2102 ( .A(core__abc_21380_n3328_bF_buf3), .B(core_v3_reg_36_), .Y(core__abc_21380_n5558) );
  OR2X2 OR2X2_2103 ( .A(core__abc_21380_n5540), .B(core__abc_21380_n5536), .Y(core__abc_21380_n5561) );
  OR2X2 OR2X2_2104 ( .A(core__abc_21380_n5520), .B(core__abc_21380_n1337), .Y(core__abc_21380_n5562) );
  OR2X2 OR2X2_2105 ( .A(core__abc_21380_n5564), .B(core__abc_21380_n5565), .Y(core__abc_21380_n5566) );
  OR2X2 OR2X2_2106 ( .A(core__abc_21380_n5527), .B(core__abc_21380_n1932), .Y(core__abc_21380_n5568) );
  OR2X2 OR2X2_2107 ( .A(core__abc_21380_n5570), .B(core__abc_21380_n5571), .Y(core__abc_21380_n5572) );
  OR2X2 OR2X2_2108 ( .A(core__abc_21380_n5572), .B(core_v3_reg_21_), .Y(core__abc_21380_n5575) );
  OR2X2 OR2X2_2109 ( .A(core__abc_21380_n5561), .B(core__abc_21380_n5582), .Y(core__abc_21380_n5583) );
  OR2X2 OR2X2_211 ( .A(_abc_19068_n1352_1), .B(_abc_19068_n1353), .Y(_abc_19068_n1354_1) );
  OR2X2 OR2X2_2110 ( .A(core__abc_21380_n5584), .B(core__abc_21380_n5585), .Y(core__abc_21380_n5586) );
  OR2X2 OR2X2_2111 ( .A(core__abc_21380_n5588), .B(core__abc_21380_n4402_1), .Y(core__abc_21380_n5589) );
  OR2X2 OR2X2_2112 ( .A(core__abc_21380_n5587), .B(core__abc_21380_n4400), .Y(core__abc_21380_n5590) );
  OR2X2 OR2X2_2113 ( .A(core_v3_reg_37_), .B(core_mi_37_), .Y(core__abc_21380_n5595) );
  OR2X2 OR2X2_2114 ( .A(core__abc_21380_n5594), .B(core__abc_21380_n5599), .Y(core__abc_21380_n5600) );
  OR2X2 OR2X2_2115 ( .A(core__abc_21380_n3317_bF_buf1), .B(core__abc_21380_n5600), .Y(core__abc_21380_n5601) );
  OR2X2 OR2X2_2116 ( .A(core__abc_21380_n5592), .B(core__abc_21380_n5601), .Y(core__abc_21380_n5602) );
  OR2X2 OR2X2_2117 ( .A(core__abc_21380_n3328_bF_buf2), .B(core_v3_reg_37_), .Y(core__abc_21380_n5603) );
  OR2X2 OR2X2_2118 ( .A(core__abc_21380_n5578), .B(core__abc_21380_n5536), .Y(core__abc_21380_n5606) );
  OR2X2 OR2X2_2119 ( .A(core__abc_21380_n5609), .B(core__abc_21380_n5607), .Y(core__abc_21380_n5610) );
  OR2X2 OR2X2_212 ( .A(_abc_19068_n1351), .B(_abc_19068_n1354_1), .Y(_abc_19068_n1355) );
  OR2X2 OR2X2_2120 ( .A(core__abc_21380_n5612), .B(core__abc_21380_n3183), .Y(core__abc_21380_n5613) );
  OR2X2 OR2X2_2121 ( .A(core__abc_21380_n5613), .B(core__abc_21380_n1378), .Y(core__abc_21380_n5616) );
  OR2X2 OR2X2_2122 ( .A(core__abc_21380_n5618), .B(core__abc_21380_n3136), .Y(core__abc_21380_n5619) );
  OR2X2 OR2X2_2123 ( .A(core__abc_21380_n5621), .B(core__abc_21380_n5622), .Y(core__abc_21380_n5623) );
  OR2X2 OR2X2_2124 ( .A(core__abc_21380_n5624), .B(core_v3_reg_22_), .Y(core__abc_21380_n5625) );
  OR2X2 OR2X2_2125 ( .A(core__abc_21380_n5623), .B(core__abc_21380_n5626), .Y(core__abc_21380_n5627) );
  OR2X2 OR2X2_2126 ( .A(core__abc_21380_n5632), .B(core__abc_21380_n5629), .Y(core__abc_21380_n5633) );
  OR2X2 OR2X2_2127 ( .A(core__abc_21380_n5634), .B(core__abc_21380_n5636), .Y(core__abc_21380_n5637) );
  OR2X2 OR2X2_2128 ( .A(core__abc_21380_n5637), .B(core__abc_21380_n4470), .Y(core__abc_21380_n5638) );
  OR2X2 OR2X2_2129 ( .A(core__abc_21380_n5639), .B(core__abc_21380_n4471), .Y(core__abc_21380_n5640) );
  OR2X2 OR2X2_213 ( .A(_abc_19068_n1357), .B(_abc_19068_n1358_1), .Y(_abc_19068_n1359) );
  OR2X2 OR2X2_2130 ( .A(core_v3_reg_38_), .B(core_mi_38_), .Y(core__abc_21380_n5645) );
  OR2X2 OR2X2_2131 ( .A(core__abc_21380_n5644), .B(core__abc_21380_n5649), .Y(core__abc_21380_n5650) );
  OR2X2 OR2X2_2132 ( .A(core__abc_21380_n3317_bF_buf0), .B(core__abc_21380_n5650), .Y(core__abc_21380_n5651) );
  OR2X2 OR2X2_2133 ( .A(core__abc_21380_n5642), .B(core__abc_21380_n5651), .Y(core__abc_21380_n5652) );
  OR2X2 OR2X2_2134 ( .A(core__abc_21380_n3328_bF_buf1), .B(core_v3_reg_38_), .Y(core__abc_21380_n5653) );
  OR2X2 OR2X2_2135 ( .A(core__abc_21380_n5636), .B(core__abc_21380_n5629), .Y(core__abc_21380_n5656) );
  OR2X2 OR2X2_2136 ( .A(core__abc_21380_n5658), .B(core__abc_21380_n1396), .Y(core__abc_21380_n5661) );
  OR2X2 OR2X2_2137 ( .A(core__abc_21380_n5622), .B(core__abc_21380_n1971), .Y(core__abc_21380_n5664) );
  OR2X2 OR2X2_2138 ( .A(core__abc_21380_n5666), .B(core__abc_21380_n5667), .Y(core__abc_21380_n5668) );
  OR2X2 OR2X2_2139 ( .A(core__abc_21380_n5668), .B(core__abc_21380_n5663), .Y(core__abc_21380_n5671) );
  OR2X2 OR2X2_214 ( .A(_abc_19068_n1359), .B(_abc_19068_n1356_1), .Y(_abc_19068_n1360_1) );
  OR2X2 OR2X2_2140 ( .A(core__abc_21380_n5672), .B(core__abc_21380_n5662), .Y(core__abc_21380_n5675) );
  OR2X2 OR2X2_2141 ( .A(core__abc_21380_n5656), .B(core__abc_21380_n5676), .Y(core__abc_21380_n5677) );
  OR2X2 OR2X2_2142 ( .A(core__abc_21380_n5680), .B(core__abc_21380_n5669), .Y(core__abc_21380_n5681) );
  OR2X2 OR2X2_2143 ( .A(core__abc_21380_n5682), .B(core__abc_21380_n5673), .Y(core__abc_21380_n5683) );
  OR2X2 OR2X2_2144 ( .A(core__abc_21380_n5678), .B(core__abc_21380_n5683), .Y(core__abc_21380_n5684) );
  OR2X2 OR2X2_2145 ( .A(core__abc_21380_n5685), .B(core__abc_21380_n4538), .Y(core__abc_21380_n5686) );
  OR2X2 OR2X2_2146 ( .A(core__abc_21380_n5687), .B(core__abc_21380_n4537_1), .Y(core__abc_21380_n5688) );
  OR2X2 OR2X2_2147 ( .A(core_v3_reg_39_), .B(core_mi_39_), .Y(core__abc_21380_n5692) );
  OR2X2 OR2X2_2148 ( .A(core__abc_21380_n5691), .B(core__abc_21380_n5696), .Y(core__abc_21380_n5697) );
  OR2X2 OR2X2_2149 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n5697), .Y(core__abc_21380_n5698) );
  OR2X2 OR2X2_215 ( .A(_abc_19068_n1361), .B(_abc_19068_n1362), .Y(_abc_19068_n1363_1) );
  OR2X2 OR2X2_2150 ( .A(core__abc_21380_n5690), .B(core__abc_21380_n5698), .Y(core__abc_21380_n5699) );
  OR2X2 OR2X2_2151 ( .A(core__abc_21380_n3328_bF_buf0), .B(core_v3_reg_39_), .Y(core__abc_21380_n5700) );
  OR2X2 OR2X2_2152 ( .A(core__abc_21380_n5707), .B(core__abc_21380_n5673), .Y(core__abc_21380_n5708) );
  OR2X2 OR2X2_2153 ( .A(core__abc_21380_n5706), .B(core__abc_21380_n5708), .Y(core__abc_21380_n5709) );
  OR2X2 OR2X2_2154 ( .A(core__abc_21380_n5709), .B(core__abc_21380_n5705), .Y(core__abc_21380_n5710) );
  OR2X2 OR2X2_2155 ( .A(core__abc_21380_n5712), .B(core__abc_21380_n5710), .Y(core__abc_21380_n5713) );
  OR2X2 OR2X2_2156 ( .A(core__abc_21380_n5715), .B(core__abc_21380_n5714), .Y(core__abc_21380_n5716) );
  OR2X2 OR2X2_2157 ( .A(core__abc_21380_n5720), .B(core__abc_21380_n5719), .Y(core__abc_21380_n5721) );
  OR2X2 OR2X2_2158 ( .A(core__abc_21380_n5722), .B(core__abc_21380_n5718), .Y(core__abc_21380_n5723) );
  OR2X2 OR2X2_2159 ( .A(core__abc_21380_n5721), .B(core_v3_reg_24_), .Y(core__abc_21380_n5724) );
  OR2X2 OR2X2_216 ( .A(_abc_19068_n1364), .B(_abc_19068_n1365_1), .Y(_abc_19068_n1366) );
  OR2X2 OR2X2_2160 ( .A(core__abc_21380_n5727), .B(core__abc_21380_n5728), .Y(core__abc_21380_n5729) );
  OR2X2 OR2X2_2161 ( .A(core__abc_21380_n5733), .B(core__abc_21380_n5731), .Y(core__abc_21380_n5734) );
  OR2X2 OR2X2_2162 ( .A(core__abc_21380_n5735), .B(core__abc_21380_n4604), .Y(core__abc_21380_n5736) );
  OR2X2 OR2X2_2163 ( .A(core__abc_21380_n5734), .B(core__abc_21380_n4603_1), .Y(core__abc_21380_n5737) );
  OR2X2 OR2X2_2164 ( .A(core_v3_reg_40_), .B(core_mi_40_), .Y(core__abc_21380_n5741) );
  OR2X2 OR2X2_2165 ( .A(core__abc_21380_n5740), .B(core__abc_21380_n5745), .Y(core__abc_21380_n5746) );
  OR2X2 OR2X2_2166 ( .A(core__abc_21380_n3317_bF_buf6), .B(core__abc_21380_n5746), .Y(core__abc_21380_n5747) );
  OR2X2 OR2X2_2167 ( .A(core__abc_21380_n5739), .B(core__abc_21380_n5747), .Y(core__abc_21380_n5748) );
  OR2X2 OR2X2_2168 ( .A(core__abc_21380_n3328_bF_buf7), .B(core_v3_reg_40_), .Y(core__abc_21380_n5749) );
  OR2X2 OR2X2_2169 ( .A(core__abc_21380_n5714), .B(core__abc_21380_n1411), .Y(core__abc_21380_n5755) );
  OR2X2 OR2X2_217 ( .A(_abc_19068_n1363_1), .B(_abc_19068_n1366), .Y(_abc_19068_n1367_1) );
  OR2X2 OR2X2_2170 ( .A(core__abc_21380_n5757), .B(core__abc_21380_n5758), .Y(core__abc_21380_n5759) );
  OR2X2 OR2X2_2171 ( .A(core__abc_21380_n5720), .B(core__abc_21380_n2009), .Y(core__abc_21380_n5762) );
  OR2X2 OR2X2_2172 ( .A(core__abc_21380_n5764), .B(core__abc_21380_n5765), .Y(core__abc_21380_n5766) );
  OR2X2 OR2X2_2173 ( .A(core__abc_21380_n5769), .B(core__abc_21380_n5767), .Y(core__abc_21380_n5770) );
  OR2X2 OR2X2_2174 ( .A(core__abc_21380_n5754), .B(core__abc_21380_n5776), .Y(core__abc_21380_n5777) );
  OR2X2 OR2X2_2175 ( .A(core__abc_21380_n5778), .B(core__abc_21380_n5779), .Y(core__abc_21380_n5780) );
  OR2X2 OR2X2_2176 ( .A(core__abc_21380_n5782), .B(core__abc_21380_n4655_1), .Y(core__abc_21380_n5783) );
  OR2X2 OR2X2_2177 ( .A(core__abc_21380_n5781), .B(core__abc_21380_n4654), .Y(core__abc_21380_n5784) );
  OR2X2 OR2X2_2178 ( .A(core_v3_reg_41_), .B(core_mi_41_), .Y(core__abc_21380_n5788) );
  OR2X2 OR2X2_2179 ( .A(core__abc_21380_n5787), .B(core__abc_21380_n5792), .Y(core__abc_21380_n5793) );
  OR2X2 OR2X2_218 ( .A(_abc_19068_n1367_1), .B(_abc_19068_n1360_1), .Y(_abc_19068_n1368) );
  OR2X2 OR2X2_2180 ( .A(core__abc_21380_n3317_bF_buf5), .B(core__abc_21380_n5793), .Y(core__abc_21380_n5794) );
  OR2X2 OR2X2_2181 ( .A(core__abc_21380_n5786), .B(core__abc_21380_n5794), .Y(core__abc_21380_n5795) );
  OR2X2 OR2X2_2182 ( .A(core__abc_21380_n3328_bF_buf6), .B(core_v3_reg_41_), .Y(core__abc_21380_n5796) );
  OR2X2 OR2X2_2183 ( .A(core__abc_21380_n5799), .B(core__abc_21380_n3200_1), .Y(core__abc_21380_n5800) );
  OR2X2 OR2X2_2184 ( .A(core__abc_21380_n5800), .B(core__abc_21380_n1451), .Y(core__abc_21380_n5803) );
  OR2X2 OR2X2_2185 ( .A(core__abc_21380_n3147), .B(core__abc_21380_n2048), .Y(core__abc_21380_n5806) );
  OR2X2 OR2X2_2186 ( .A(core__abc_21380_n5807), .B(core__abc_21380_n5805), .Y(core__abc_21380_n5808) );
  OR2X2 OR2X2_2187 ( .A(core__abc_21380_n5809), .B(core_v3_reg_26_), .Y(core__abc_21380_n5810) );
  OR2X2 OR2X2_2188 ( .A(core__abc_21380_n5813), .B(core__abc_21380_n5815), .Y(core__abc_21380_n5816) );
  OR2X2 OR2X2_2189 ( .A(core__abc_21380_n5818), .B(core__abc_21380_n5774), .Y(core__abc_21380_n5819) );
  OR2X2 OR2X2_219 ( .A(_abc_19068_n1368), .B(_abc_19068_n1355), .Y(_abc_19068_n1369_1) );
  OR2X2 OR2X2_2190 ( .A(core__abc_21380_n5819), .B(core__abc_21380_n5816), .Y(core__abc_21380_n5821) );
  OR2X2 OR2X2_2191 ( .A(core__abc_21380_n5822), .B(core__abc_21380_n5820), .Y(core__abc_21380_n5823) );
  OR2X2 OR2X2_2192 ( .A(core__abc_21380_n5823), .B(core__abc_21380_n4720), .Y(core__abc_21380_n5824) );
  OR2X2 OR2X2_2193 ( .A(core__abc_21380_n5825), .B(core__abc_21380_n4721), .Y(core__abc_21380_n5826) );
  OR2X2 OR2X2_2194 ( .A(core_v3_reg_42_), .B(core_mi_42_), .Y(core__abc_21380_n5831) );
  OR2X2 OR2X2_2195 ( .A(core__abc_21380_n5830), .B(core__abc_21380_n5835), .Y(core__abc_21380_n5836) );
  OR2X2 OR2X2_2196 ( .A(core__abc_21380_n3317_bF_buf4), .B(core__abc_21380_n5836), .Y(core__abc_21380_n5837) );
  OR2X2 OR2X2_2197 ( .A(core__abc_21380_n5828), .B(core__abc_21380_n5837), .Y(core__abc_21380_n5838) );
  OR2X2 OR2X2_2198 ( .A(core__abc_21380_n3328_bF_buf5), .B(core_v3_reg_42_), .Y(core__abc_21380_n5839) );
  OR2X2 OR2X2_2199 ( .A(core__abc_21380_n5844), .B(core__abc_21380_n1474), .Y(core__abc_21380_n5847) );
  OR2X2 OR2X2_22 ( .A(_abc_19068_n947), .B(_abc_19068_n950), .Y(_abc_19068_n951_1) );
  OR2X2 OR2X2_220 ( .A(_abc_19068_n1372), .B(_abc_19068_n1373_1), .Y(_abc_19068_n1374) );
  OR2X2 OR2X2_2200 ( .A(core__abc_21380_n3159), .B(core__abc_21380_n5849), .Y(core__abc_21380_n5850) );
  OR2X2 OR2X2_2201 ( .A(core__abc_21380_n3303), .B(core__abc_21380_n5848), .Y(core__abc_21380_n5851) );
  OR2X2 OR2X2_2202 ( .A(core__abc_21380_n5856), .B(core__abc_21380_n5854), .Y(core__abc_21380_n5857) );
  OR2X2 OR2X2_2203 ( .A(core__abc_21380_n5858), .B(core__abc_21380_n4776), .Y(core__abc_21380_n5859) );
  OR2X2 OR2X2_2204 ( .A(core__abc_21380_n5857), .B(core__abc_21380_n4775), .Y(core__abc_21380_n5860) );
  OR2X2 OR2X2_2205 ( .A(core_v3_reg_43_), .B(core_mi_43_), .Y(core__abc_21380_n5864) );
  OR2X2 OR2X2_2206 ( .A(core__abc_21380_n5863), .B(core__abc_21380_n5868), .Y(core__abc_21380_n5869) );
  OR2X2 OR2X2_2207 ( .A(core__abc_21380_n3317_bF_buf3), .B(core__abc_21380_n5869), .Y(core__abc_21380_n5870) );
  OR2X2 OR2X2_2208 ( .A(core__abc_21380_n5862), .B(core__abc_21380_n5870), .Y(core__abc_21380_n5871) );
  OR2X2 OR2X2_2209 ( .A(core__abc_21380_n3328_bF_buf4), .B(core_v3_reg_43_), .Y(core__abc_21380_n5872) );
  OR2X2 OR2X2_221 ( .A(_abc_19068_n1374), .B(_abc_19068_n1371_1), .Y(_abc_19068_n1375_1) );
  OR2X2 OR2X2_2210 ( .A(core__abc_21380_n5817), .B(core__abc_21380_n5774), .Y(core__abc_21380_n5875) );
  OR2X2 OR2X2_2211 ( .A(core__abc_21380_n5880), .B(core__abc_21380_n5842), .Y(core__abc_21380_n5881) );
  OR2X2 OR2X2_2212 ( .A(core__abc_21380_n5879), .B(core__abc_21380_n5883), .Y(core__abc_21380_n5884) );
  OR2X2 OR2X2_2213 ( .A(core__abc_21380_n5887), .B(core__abc_21380_n5884), .Y(core__abc_21380_n5888) );
  OR2X2 OR2X2_2214 ( .A(core__abc_21380_n5890), .B(core__abc_21380_n3204), .Y(core__abc_21380_n5891) );
  OR2X2 OR2X2_2215 ( .A(core__abc_21380_n5893), .B(core__abc_21380_n5894), .Y(core__abc_21380_n5895) );
  OR2X2 OR2X2_2216 ( .A(core__abc_21380_n5897), .B(core__abc_21380_n5898), .Y(core__abc_21380_n5899) );
  OR2X2 OR2X2_2217 ( .A(core__abc_21380_n5900), .B(core__abc_21380_n5902), .Y(core__abc_21380_n5903) );
  OR2X2 OR2X2_2218 ( .A(core__abc_21380_n5903), .B(core__abc_21380_n4818), .Y(core__abc_21380_n5904) );
  OR2X2 OR2X2_2219 ( .A(core__abc_21380_n5905), .B(core__abc_21380_n4824), .Y(core__abc_21380_n5906) );
  OR2X2 OR2X2_222 ( .A(_abc_19068_n1376), .B(_abc_19068_n1185_1), .Y(_abc_19068_n1377_1) );
  OR2X2 OR2X2_2220 ( .A(core_v3_reg_44_), .B(core_mi_44_), .Y(core__abc_21380_n5910) );
  OR2X2 OR2X2_2221 ( .A(core__abc_21380_n5909), .B(core__abc_21380_n5914), .Y(core__abc_21380_n5915) );
  OR2X2 OR2X2_2222 ( .A(core__abc_21380_n3317_bF_buf2), .B(core__abc_21380_n5915), .Y(core__abc_21380_n5916) );
  OR2X2 OR2X2_2223 ( .A(core__abc_21380_n5908), .B(core__abc_21380_n5916), .Y(core__abc_21380_n5917) );
  OR2X2 OR2X2_2224 ( .A(core__abc_21380_n3328_bF_buf3), .B(core_v3_reg_44_), .Y(core__abc_21380_n5918) );
  OR2X2 OR2X2_2225 ( .A(core__abc_21380_n5894), .B(core__abc_21380_n1482), .Y(core__abc_21380_n5921) );
  OR2X2 OR2X2_2226 ( .A(core__abc_21380_n5923), .B(core__abc_21380_n5924), .Y(core__abc_21380_n5925) );
  OR2X2 OR2X2_2227 ( .A(core__abc_21380_n3438), .B(core__abc_21380_n5925), .Y(core__abc_21380_n5926) );
  OR2X2 OR2X2_2228 ( .A(core__abc_21380_n3443), .B(core__abc_21380_n5927), .Y(core__abc_21380_n5928) );
  OR2X2 OR2X2_2229 ( .A(core__abc_21380_n5933), .B(core__abc_21380_n5930), .Y(core__abc_21380_n5935) );
  OR2X2 OR2X2_223 ( .A(_abc_19068_n1378), .B(_abc_19068_n1379_1), .Y(_abc_19068_n1380) );
  OR2X2 OR2X2_2230 ( .A(core__abc_21380_n5936), .B(core__abc_21380_n5934), .Y(core__abc_21380_n5937) );
  OR2X2 OR2X2_2231 ( .A(core__abc_21380_n5938), .B(core__abc_21380_n4900_1), .Y(core__abc_21380_n5939) );
  OR2X2 OR2X2_2232 ( .A(core__abc_21380_n5937), .B(core__abc_21380_n4899), .Y(core__abc_21380_n5940) );
  OR2X2 OR2X2_2233 ( .A(core_v3_reg_45_), .B(core_mi_45_), .Y(core__abc_21380_n5945) );
  OR2X2 OR2X2_2234 ( .A(core__abc_21380_n5944), .B(core__abc_21380_n5949), .Y(core__abc_21380_n5950) );
  OR2X2 OR2X2_2235 ( .A(core__abc_21380_n3317_bF_buf1), .B(core__abc_21380_n5950), .Y(core__abc_21380_n5951) );
  OR2X2 OR2X2_2236 ( .A(core__abc_21380_n5942), .B(core__abc_21380_n5951), .Y(core__abc_21380_n5952) );
  OR2X2 OR2X2_2237 ( .A(core__abc_21380_n3328_bF_buf2), .B(core_v3_reg_45_), .Y(core__abc_21380_n5953) );
  OR2X2 OR2X2_2238 ( .A(core__abc_21380_n5959), .B(core__abc_21380_n5958), .Y(core__abc_21380_n5960) );
  OR2X2 OR2X2_2239 ( .A(core__abc_21380_n5957), .B(core__abc_21380_n5960), .Y(core__abc_21380_n5961) );
  OR2X2 OR2X2_224 ( .A(_abc_19068_n1380), .B(_abc_19068_n1377_1), .Y(_abc_19068_n1381_1) );
  OR2X2 OR2X2_2240 ( .A(core__abc_21380_n5963), .B(core__abc_21380_n3209), .Y(core__abc_21380_n5964) );
  OR2X2 OR2X2_2241 ( .A(core__abc_21380_n5964), .B(core__abc_21380_n1523), .Y(core__abc_21380_n5967) );
  OR2X2 OR2X2_2242 ( .A(core__abc_21380_n5971), .B(core__abc_21380_n5969), .Y(core__abc_21380_n5972) );
  OR2X2 OR2X2_2243 ( .A(core__abc_21380_n5973), .B(core__abc_21380_n5975), .Y(core__abc_21380_n5976) );
  OR2X2 OR2X2_2244 ( .A(core__abc_21380_n5976), .B(core__abc_21380_n4946), .Y(core__abc_21380_n5977) );
  OR2X2 OR2X2_2245 ( .A(core__abc_21380_n5979), .B(core__abc_21380_n5978), .Y(core__abc_21380_n5980) );
  OR2X2 OR2X2_2246 ( .A(core_v3_reg_46_), .B(core_mi_46_), .Y(core__abc_21380_n5985) );
  OR2X2 OR2X2_2247 ( .A(core__abc_21380_n5984), .B(core__abc_21380_n5989), .Y(core__abc_21380_n5990) );
  OR2X2 OR2X2_2248 ( .A(core__abc_21380_n3317_bF_buf0), .B(core__abc_21380_n5990), .Y(core__abc_21380_n5991) );
  OR2X2 OR2X2_2249 ( .A(core__abc_21380_n5982), .B(core__abc_21380_n5991), .Y(core__abc_21380_n5992) );
  OR2X2 OR2X2_225 ( .A(_abc_19068_n1382), .B(_abc_19068_n1383_1), .Y(_abc_19068_n1384) );
  OR2X2 OR2X2_2250 ( .A(core__abc_21380_n3328_bF_buf1), .B(core_v3_reg_46_), .Y(core__abc_21380_n5993) );
  OR2X2 OR2X2_2251 ( .A(core__abc_21380_n5975), .B(core__abc_21380_n5969), .Y(core__abc_21380_n5996) );
  OR2X2 OR2X2_2252 ( .A(core__abc_21380_n5965), .B(core__abc_21380_n1521), .Y(core__abc_21380_n5997) );
  OR2X2 OR2X2_2253 ( .A(core__abc_21380_n5999), .B(core__abc_21380_n6000), .Y(core__abc_21380_n6001) );
  OR2X2 OR2X2_2254 ( .A(core__abc_21380_n6003), .B(core__abc_21380_n6004), .Y(core__abc_21380_n6005) );
  OR2X2 OR2X2_2255 ( .A(core__abc_21380_n5996), .B(core__abc_21380_n6005), .Y(core__abc_21380_n6006) );
  OR2X2 OR2X2_2256 ( .A(core__abc_21380_n3580), .B(core__abc_21380_n6001), .Y(core__abc_21380_n6008) );
  OR2X2 OR2X2_2257 ( .A(core__abc_21380_n3576), .B(core__abc_21380_n6002), .Y(core__abc_21380_n6009) );
  OR2X2 OR2X2_2258 ( .A(core__abc_21380_n6007), .B(core__abc_21380_n6010), .Y(core__abc_21380_n6011) );
  OR2X2 OR2X2_2259 ( .A(core__abc_21380_n6013), .B(core__abc_21380_n4991), .Y(core__abc_21380_n6014) );
  OR2X2 OR2X2_226 ( .A(_abc_19068_n1385_1), .B(_abc_19068_n1386), .Y(_abc_19068_n1387_1) );
  OR2X2 OR2X2_2260 ( .A(core__abc_21380_n6012), .B(core__abc_21380_n4990), .Y(core__abc_21380_n6015) );
  OR2X2 OR2X2_2261 ( .A(core_v3_reg_47_), .B(core_mi_47_), .Y(core__abc_21380_n6019) );
  OR2X2 OR2X2_2262 ( .A(core__abc_21380_n6018), .B(core__abc_21380_n6023), .Y(core__abc_21380_n6024) );
  OR2X2 OR2X2_2263 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n6024), .Y(core__abc_21380_n6025) );
  OR2X2 OR2X2_2264 ( .A(core__abc_21380_n6017), .B(core__abc_21380_n6025), .Y(core__abc_21380_n6026) );
  OR2X2 OR2X2_2265 ( .A(core__abc_21380_n3328_bF_buf0), .B(core_v3_reg_47_), .Y(core__abc_21380_n6027) );
  OR2X2 OR2X2_2266 ( .A(core__abc_21380_n6004), .B(core__abc_21380_n6038), .Y(core__abc_21380_n6039) );
  OR2X2 OR2X2_2267 ( .A(core__abc_21380_n6037), .B(core__abc_21380_n6041), .Y(core__abc_21380_n6042) );
  OR2X2 OR2X2_2268 ( .A(core__abc_21380_n6042), .B(core__abc_21380_n6036), .Y(core__abc_21380_n6043) );
  OR2X2 OR2X2_2269 ( .A(core__abc_21380_n6035), .B(core__abc_21380_n6043), .Y(core__abc_21380_n6044) );
  OR2X2 OR2X2_227 ( .A(_abc_19068_n1384), .B(_abc_19068_n1387_1), .Y(_abc_19068_n1388) );
  OR2X2 OR2X2_2270 ( .A(core__abc_21380_n6034), .B(core__abc_21380_n6044), .Y(core__abc_21380_n6045) );
  OR2X2 OR2X2_2271 ( .A(core__abc_21380_n6047), .B(core__abc_21380_n6046), .Y(core__abc_21380_n6048) );
  OR2X2 OR2X2_2272 ( .A(core__abc_21380_n6050), .B(core__abc_21380_n6051), .Y(core__abc_21380_n6052) );
  OR2X2 OR2X2_2273 ( .A(core__abc_21380_n5319), .B(core__abc_21380_n6055), .Y(core__abc_21380_n6056) );
  OR2X2 OR2X2_2274 ( .A(core__abc_21380_n5683), .B(core__abc_21380_n5633), .Y(core__abc_21380_n6059) );
  OR2X2 OR2X2_2275 ( .A(core__abc_21380_n6059), .B(core__abc_21380_n6058), .Y(core__abc_21380_n6060) );
  OR2X2 OR2X2_2276 ( .A(core__abc_21380_n6060), .B(core__abc_21380_n6057), .Y(core__abc_21380_n6061) );
  OR2X2 OR2X2_2277 ( .A(core__abc_21380_n6059), .B(core__abc_21380_n6062), .Y(core__abc_21380_n6063) );
  OR2X2 OR2X2_2278 ( .A(core__abc_21380_n6067), .B(core__abc_21380_n6066), .Y(core__abc_21380_n6068) );
  OR2X2 OR2X2_2279 ( .A(core__abc_21380_n6074), .B(core__abc_21380_n6054), .Y(core__abc_21380_n6075) );
  OR2X2 OR2X2_228 ( .A(_abc_19068_n1388), .B(_abc_19068_n1381_1), .Y(_abc_19068_n1389_1) );
  OR2X2 OR2X2_2280 ( .A(core__abc_21380_n6076), .B(core__abc_21380_n5041), .Y(core__abc_21380_n6077) );
  OR2X2 OR2X2_2281 ( .A(core__abc_21380_n6075), .B(core__abc_21380_n5045), .Y(core__abc_21380_n6078) );
  OR2X2 OR2X2_2282 ( .A(core_v3_reg_48_), .B(core_mi_48_), .Y(core__abc_21380_n6083) );
  OR2X2 OR2X2_2283 ( .A(core__abc_21380_n6082), .B(core__abc_21380_n6087), .Y(core__abc_21380_n6088) );
  OR2X2 OR2X2_2284 ( .A(core__abc_21380_n3317_bF_buf6), .B(core__abc_21380_n6088), .Y(core__abc_21380_n6089) );
  OR2X2 OR2X2_2285 ( .A(core__abc_21380_n6080), .B(core__abc_21380_n6089), .Y(core__abc_21380_n6090) );
  OR2X2 OR2X2_2286 ( .A(core__abc_21380_n3328_bF_buf7), .B(core_v3_reg_48_), .Y(core__abc_21380_n6091) );
  OR2X2 OR2X2_2287 ( .A(core__abc_21380_n6046), .B(core__abc_21380_n1556), .Y(core__abc_21380_n6098) );
  OR2X2 OR2X2_2288 ( .A(core__abc_21380_n6100), .B(core__abc_21380_n6101), .Y(core__abc_21380_n6102) );
  OR2X2 OR2X2_2289 ( .A(core__abc_21380_n6097), .B(core__abc_21380_n6108), .Y(core__abc_21380_n6109) );
  OR2X2 OR2X2_229 ( .A(_abc_19068_n1389_1), .B(_abc_19068_n1375_1), .Y(_abc_19068_n1390) );
  OR2X2 OR2X2_2290 ( .A(core__abc_21380_n6096), .B(core__abc_21380_n6110), .Y(core__abc_21380_n6111) );
  OR2X2 OR2X2_2291 ( .A(core__abc_21380_n6112), .B(core__abc_21380_n5113), .Y(core__abc_21380_n6113) );
  OR2X2 OR2X2_2292 ( .A(core__abc_21380_n6114), .B(core__abc_21380_n5112), .Y(core__abc_21380_n6115) );
  OR2X2 OR2X2_2293 ( .A(core_v3_reg_49_), .B(core_mi_49_), .Y(core__abc_21380_n6119) );
  OR2X2 OR2X2_2294 ( .A(core__abc_21380_n6118), .B(core__abc_21380_n6123), .Y(core__abc_21380_n6124) );
  OR2X2 OR2X2_2295 ( .A(core__abc_21380_n3317_bF_buf5), .B(core__abc_21380_n6124), .Y(core__abc_21380_n6125) );
  OR2X2 OR2X2_2296 ( .A(core__abc_21380_n6117), .B(core__abc_21380_n6125), .Y(core__abc_21380_n6126) );
  OR2X2 OR2X2_2297 ( .A(core__abc_21380_n3328_bF_buf6), .B(core_v3_reg_49_), .Y(core__abc_21380_n6127) );
  OR2X2 OR2X2_2298 ( .A(core__abc_21380_n6106), .B(core__abc_21380_n6094), .Y(core__abc_21380_n6130) );
  OR2X2 OR2X2_2299 ( .A(core__abc_21380_n6134), .B(core__abc_21380_n6132), .Y(core__abc_21380_n6135) );
  OR2X2 OR2X2_23 ( .A(_abc_19068_n951_1), .B(_abc_19068_n943_1), .Y(_abc_19068_n952_1) );
  OR2X2 OR2X2_230 ( .A(_abc_19068_n1392), .B(_abc_19068_n1393_1), .Y(_abc_19068_n1394) );
  OR2X2 OR2X2_2300 ( .A(core__abc_21380_n6137), .B(core__abc_21380_n3234), .Y(core__abc_21380_n6138) );
  OR2X2 OR2X2_2301 ( .A(core__abc_21380_n6138), .B(core__abc_21380_n1597), .Y(core__abc_21380_n6141) );
  OR2X2 OR2X2_2302 ( .A(core__abc_21380_n6143), .B(core__abc_21380_n6145), .Y(core__abc_21380_n6146) );
  OR2X2 OR2X2_2303 ( .A(core__abc_21380_n6147), .B(core__abc_21380_n6149), .Y(core__abc_21380_n6150) );
  OR2X2 OR2X2_2304 ( .A(core__abc_21380_n6150), .B(core__abc_21380_n5162), .Y(core__abc_21380_n6151) );
  OR2X2 OR2X2_2305 ( .A(core__abc_21380_n6152), .B(core__abc_21380_n5159), .Y(core__abc_21380_n6153) );
  OR2X2 OR2X2_2306 ( .A(core_v3_reg_50_), .B(core_mi_50_), .Y(core__abc_21380_n6158) );
  OR2X2 OR2X2_2307 ( .A(core__abc_21380_n6157), .B(core__abc_21380_n6162), .Y(core__abc_21380_n6163) );
  OR2X2 OR2X2_2308 ( .A(core__abc_21380_n3317_bF_buf4), .B(core__abc_21380_n6163), .Y(core__abc_21380_n6164) );
  OR2X2 OR2X2_2309 ( .A(core__abc_21380_n6155), .B(core__abc_21380_n6164), .Y(core__abc_21380_n6165) );
  OR2X2 OR2X2_231 ( .A(_abc_19068_n1395_1), .B(_abc_19068_n1396), .Y(_abc_19068_n1397_1) );
  OR2X2 OR2X2_2310 ( .A(core__abc_21380_n3328_bF_buf5), .B(core_v3_reg_50_), .Y(core__abc_21380_n6166) );
  OR2X2 OR2X2_2311 ( .A(core__abc_21380_n6149), .B(core__abc_21380_n6143), .Y(core__abc_21380_n6169) );
  OR2X2 OR2X2_2312 ( .A(core__abc_21380_n6170), .B(core__abc_21380_n1621), .Y(core__abc_21380_n6173) );
  OR2X2 OR2X2_2313 ( .A(core__abc_21380_n3862), .B(core__abc_21380_n6175), .Y(core__abc_21380_n6176) );
  OR2X2 OR2X2_2314 ( .A(core__abc_21380_n3859), .B(core__abc_21380_n6174), .Y(core__abc_21380_n6177) );
  OR2X2 OR2X2_2315 ( .A(core__abc_21380_n6169), .B(core__abc_21380_n6178), .Y(core__abc_21380_n6179) );
  OR2X2 OR2X2_2316 ( .A(core__abc_21380_n6181), .B(core__abc_21380_n6182), .Y(core__abc_21380_n6183) );
  OR2X2 OR2X2_2317 ( .A(core__abc_21380_n6180), .B(core__abc_21380_n6183), .Y(core__abc_21380_n6184) );
  OR2X2 OR2X2_2318 ( .A(core__abc_21380_n6186), .B(core__abc_21380_n5221), .Y(core__abc_21380_n6187) );
  OR2X2 OR2X2_2319 ( .A(core__abc_21380_n6185), .B(core__abc_21380_n5219), .Y(core__abc_21380_n6188) );
  OR2X2 OR2X2_232 ( .A(_abc_19068_n1394), .B(_abc_19068_n1397_1), .Y(_abc_19068_n1398) );
  OR2X2 OR2X2_2320 ( .A(core_v3_reg_51_), .B(core_mi_51_), .Y(core__abc_21380_n6192) );
  OR2X2 OR2X2_2321 ( .A(core__abc_21380_n6191), .B(core__abc_21380_n6196), .Y(core__abc_21380_n6197) );
  OR2X2 OR2X2_2322 ( .A(core__abc_21380_n3317_bF_buf3), .B(core__abc_21380_n6197), .Y(core__abc_21380_n6198) );
  OR2X2 OR2X2_2323 ( .A(core__abc_21380_n6190), .B(core__abc_21380_n6198), .Y(core__abc_21380_n6199) );
  OR2X2 OR2X2_2324 ( .A(core__abc_21380_n3328_bF_buf4), .B(core_v3_reg_51_), .Y(core__abc_21380_n6200) );
  OR2X2 OR2X2_2325 ( .A(core__abc_21380_n6181), .B(core__abc_21380_n6143), .Y(core__abc_21380_n6205) );
  OR2X2 OR2X2_2326 ( .A(core__abc_21380_n6204), .B(core__abc_21380_n6206), .Y(core__abc_21380_n6207) );
  OR2X2 OR2X2_2327 ( .A(core__abc_21380_n6209), .B(core__abc_21380_n6207), .Y(core__abc_21380_n6210) );
  OR2X2 OR2X2_2328 ( .A(core__abc_21380_n6212), .B(core__abc_21380_n3238), .Y(core__abc_21380_n6213) );
  OR2X2 OR2X2_2329 ( .A(core__abc_21380_n6215), .B(core__abc_21380_n6216), .Y(core__abc_21380_n6217) );
  OR2X2 OR2X2_233 ( .A(_abc_19068_n1399_1), .B(_abc_19068_n1400), .Y(_abc_19068_n1401_1) );
  OR2X2 OR2X2_2330 ( .A(core__abc_21380_n6219), .B(core__abc_21380_n6220), .Y(core__abc_21380_n6221) );
  OR2X2 OR2X2_2331 ( .A(core__abc_21380_n6222), .B(core__abc_21380_n6224), .Y(core__abc_21380_n6225) );
  OR2X2 OR2X2_2332 ( .A(core__abc_21380_n6225), .B(core__abc_21380_n5266), .Y(core__abc_21380_n6226) );
  OR2X2 OR2X2_2333 ( .A(core__abc_21380_n6227), .B(core__abc_21380_n5273), .Y(core__abc_21380_n6228) );
  OR2X2 OR2X2_2334 ( .A(core_v3_reg_52_), .B(core_mi_52_), .Y(core__abc_21380_n6232) );
  OR2X2 OR2X2_2335 ( .A(core__abc_21380_n6231), .B(core__abc_21380_n6236), .Y(core__abc_21380_n6237) );
  OR2X2 OR2X2_2336 ( .A(core__abc_21380_n3317_bF_buf2), .B(core__abc_21380_n6237), .Y(core__abc_21380_n6238) );
  OR2X2 OR2X2_2337 ( .A(core__abc_21380_n6230), .B(core__abc_21380_n6238), .Y(core__abc_21380_n6239) );
  OR2X2 OR2X2_2338 ( .A(core__abc_21380_n3328_bF_buf3), .B(core_v3_reg_52_), .Y(core__abc_21380_n6240) );
  OR2X2 OR2X2_2339 ( .A(core__abc_21380_n6224), .B(core__abc_21380_n6219), .Y(core__abc_21380_n6243) );
  OR2X2 OR2X2_234 ( .A(_abc_19068_n1402), .B(_abc_19068_n1403_1), .Y(_abc_19068_n1404) );
  OR2X2 OR2X2_2340 ( .A(core__abc_21380_n6216), .B(core__abc_21380_n1631), .Y(core__abc_21380_n6244) );
  OR2X2 OR2X2_2341 ( .A(core__abc_21380_n6246), .B(core__abc_21380_n6247), .Y(core__abc_21380_n6248) );
  OR2X2 OR2X2_2342 ( .A(core__abc_21380_n6250), .B(core__abc_21380_n6251), .Y(core__abc_21380_n6252) );
  OR2X2 OR2X2_2343 ( .A(core__abc_21380_n6243), .B(core__abc_21380_n6253), .Y(core__abc_21380_n6254) );
  OR2X2 OR2X2_2344 ( .A(core__abc_21380_n6255), .B(core__abc_21380_n6252), .Y(core__abc_21380_n6256) );
  OR2X2 OR2X2_2345 ( .A(core__abc_21380_n6257), .B(core__abc_21380_n5329), .Y(core__abc_21380_n6258) );
  OR2X2 OR2X2_2346 ( .A(core__abc_21380_n6259), .B(core__abc_21380_n5328), .Y(core__abc_21380_n6260) );
  OR2X2 OR2X2_2347 ( .A(core_v3_reg_53_), .B(core_mi_53_), .Y(core__abc_21380_n6265) );
  OR2X2 OR2X2_2348 ( .A(core__abc_21380_n6264), .B(core__abc_21380_n6269), .Y(core__abc_21380_n6270) );
  OR2X2 OR2X2_2349 ( .A(core__abc_21380_n3317_bF_buf1), .B(core__abc_21380_n6270), .Y(core__abc_21380_n6271) );
  OR2X2 OR2X2_235 ( .A(_abc_19068_n1401_1), .B(_abc_19068_n1404), .Y(_abc_19068_n1405_1) );
  OR2X2 OR2X2_2350 ( .A(core__abc_21380_n6262), .B(core__abc_21380_n6271), .Y(core__abc_21380_n6272) );
  OR2X2 OR2X2_2351 ( .A(core__abc_21380_n3328_bF_buf2), .B(core_v3_reg_53_), .Y(core__abc_21380_n6273) );
  OR2X2 OR2X2_2352 ( .A(core__abc_21380_n6251), .B(core__abc_21380_n6277), .Y(core__abc_21380_n6278) );
  OR2X2 OR2X2_2353 ( .A(core__abc_21380_n6252), .B(core__abc_21380_n6221), .Y(core__abc_21380_n6281) );
  OR2X2 OR2X2_2354 ( .A(core__abc_21380_n6283), .B(core__abc_21380_n6280), .Y(core__abc_21380_n6284) );
  OR2X2 OR2X2_2355 ( .A(core__abc_21380_n6286), .B(core__abc_21380_n3243), .Y(core__abc_21380_n6287) );
  OR2X2 OR2X2_2356 ( .A(core__abc_21380_n6287), .B(core__abc_21380_n1669), .Y(core__abc_21380_n6290) );
  OR2X2 OR2X2_2357 ( .A(core__abc_21380_n6294), .B(core__abc_21380_n6292), .Y(core__abc_21380_n6295) );
  OR2X2 OR2X2_2358 ( .A(core__abc_21380_n6296), .B(core__abc_21380_n6298), .Y(core__abc_21380_n6299) );
  OR2X2 OR2X2_2359 ( .A(core__abc_21380_n6299), .B(core__abc_21380_n5386), .Y(core__abc_21380_n6300) );
  OR2X2 OR2X2_236 ( .A(_abc_19068_n1406), .B(_abc_19068_n1407_1), .Y(_abc_19068_n1408) );
  OR2X2 OR2X2_2360 ( .A(core__abc_21380_n6301), .B(core__abc_21380_n5387), .Y(core__abc_21380_n6302) );
  OR2X2 OR2X2_2361 ( .A(core_v3_reg_54_), .B(core_mi_54_), .Y(core__abc_21380_n6307) );
  OR2X2 OR2X2_2362 ( .A(core__abc_21380_n6306), .B(core__abc_21380_n6311), .Y(core__abc_21380_n6312) );
  OR2X2 OR2X2_2363 ( .A(core__abc_21380_n3317_bF_buf0), .B(core__abc_21380_n6312), .Y(core__abc_21380_n6313) );
  OR2X2 OR2X2_2364 ( .A(core__abc_21380_n6304), .B(core__abc_21380_n6313), .Y(core__abc_21380_n6314) );
  OR2X2 OR2X2_2365 ( .A(core__abc_21380_n3328_bF_buf1), .B(core_v3_reg_54_), .Y(core__abc_21380_n6315) );
  OR2X2 OR2X2_2366 ( .A(core__abc_21380_n6298), .B(core__abc_21380_n6292), .Y(core__abc_21380_n6318) );
  OR2X2 OR2X2_2367 ( .A(core__abc_21380_n6288), .B(core__abc_21380_n1667), .Y(core__abc_21380_n6319) );
  OR2X2 OR2X2_2368 ( .A(core__abc_21380_n6319), .B(core__abc_21380_n1688), .Y(core__abc_21380_n6320) );
  OR2X2 OR2X2_2369 ( .A(core__abc_21380_n6324), .B(core__abc_21380_n6326), .Y(core__abc_21380_n6327) );
  OR2X2 OR2X2_237 ( .A(_abc_19068_n910_1), .B(_abc_19068_n1408), .Y(_abc_19068_n1409_1) );
  OR2X2 OR2X2_2370 ( .A(core__abc_21380_n6318), .B(core__abc_21380_n6327), .Y(core__abc_21380_n6328) );
  OR2X2 OR2X2_2371 ( .A(core__abc_21380_n4136), .B(core__abc_21380_n6325), .Y(core__abc_21380_n6330) );
  OR2X2 OR2X2_2372 ( .A(core__abc_21380_n4132), .B(core__abc_21380_n6323), .Y(core__abc_21380_n6331) );
  OR2X2 OR2X2_2373 ( .A(core__abc_21380_n6329), .B(core__abc_21380_n6332), .Y(core__abc_21380_n6333) );
  OR2X2 OR2X2_2374 ( .A(core__abc_21380_n6335), .B(core__abc_21380_n5440), .Y(core__abc_21380_n6336) );
  OR2X2 OR2X2_2375 ( .A(core__abc_21380_n6334), .B(core__abc_21380_n5439), .Y(core__abc_21380_n6337) );
  OR2X2 OR2X2_2376 ( .A(core_v3_reg_55_), .B(core_mi_55_), .Y(core__abc_21380_n6341) );
  OR2X2 OR2X2_2377 ( .A(core__abc_21380_n6340), .B(core__abc_21380_n6345), .Y(core__abc_21380_n6346) );
  OR2X2 OR2X2_2378 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n6346), .Y(core__abc_21380_n6347) );
  OR2X2 OR2X2_2379 ( .A(core__abc_21380_n6339), .B(core__abc_21380_n6347), .Y(core__abc_21380_n6348) );
  OR2X2 OR2X2_238 ( .A(_abc_19068_n1409_1), .B(_abc_19068_n1405_1), .Y(_abc_19068_n1410) );
  OR2X2 OR2X2_2380 ( .A(core__abc_21380_n3328_bF_buf0), .B(core_v3_reg_55_), .Y(core__abc_21380_n6349) );
  OR2X2 OR2X2_2381 ( .A(core__abc_21380_n6327), .B(core__abc_21380_n6295), .Y(core__abc_21380_n6353) );
  OR2X2 OR2X2_2382 ( .A(core__abc_21380_n6353), .B(core__abc_21380_n6281), .Y(core__abc_21380_n6354) );
  OR2X2 OR2X2_2383 ( .A(core__abc_21380_n6354), .B(core__abc_21380_n6352), .Y(core__abc_21380_n6355) );
  OR2X2 OR2X2_2384 ( .A(core__abc_21380_n6073), .B(core__abc_21380_n6355), .Y(core__abc_21380_n6356) );
  OR2X2 OR2X2_2385 ( .A(core__abc_21380_n6183), .B(core__abc_21380_n6146), .Y(core__abc_21380_n6357) );
  OR2X2 OR2X2_2386 ( .A(core__abc_21380_n6357), .B(core__abc_21380_n6131), .Y(core__abc_21380_n6358) );
  OR2X2 OR2X2_2387 ( .A(core__abc_21380_n6360), .B(core__abc_21380_n6354), .Y(core__abc_21380_n6361) );
  OR2X2 OR2X2_2388 ( .A(core__abc_21380_n6326), .B(core__abc_21380_n6364), .Y(core__abc_21380_n6365) );
  OR2X2 OR2X2_2389 ( .A(core__abc_21380_n6363), .B(core__abc_21380_n6367), .Y(core__abc_21380_n6368) );
  OR2X2 OR2X2_239 ( .A(_abc_19068_n1410), .B(_abc_19068_n1398), .Y(_abc_19068_n1411_1) );
  OR2X2 OR2X2_2390 ( .A(core__abc_21380_n6372), .B(core__abc_21380_n3248), .Y(core__abc_21380_n6373) );
  OR2X2 OR2X2_2391 ( .A(core__abc_21380_n3283), .B(core__abc_21380_n6376), .Y(core__abc_21380_n6377) );
  OR2X2 OR2X2_2392 ( .A(core__abc_21380_n6379), .B(core__abc_21380_n6374), .Y(core__abc_21380_n6380) );
  OR2X2 OR2X2_2393 ( .A(core__abc_21380_n6382), .B(core__abc_21380_n6383), .Y(core__abc_21380_n6384) );
  OR2X2 OR2X2_2394 ( .A(core__abc_21380_n6389), .B(core__abc_21380_n6368), .Y(core__abc_21380_n6390) );
  OR2X2 OR2X2_2395 ( .A(core__abc_21380_n6388), .B(core__abc_21380_n6390), .Y(core__abc_21380_n6391) );
  OR2X2 OR2X2_2396 ( .A(core__abc_21380_n6385), .B(core__abc_21380_n6393), .Y(core__abc_21380_n6394) );
  OR2X2 OR2X2_2397 ( .A(core__abc_21380_n6395), .B(core__abc_21380_n5484), .Y(core__abc_21380_n6396) );
  OR2X2 OR2X2_2398 ( .A(core__abc_21380_n6394), .B(core__abc_21380_n5483), .Y(core__abc_21380_n6397) );
  OR2X2 OR2X2_2399 ( .A(core_v3_reg_56_), .B(core_mi_56_), .Y(core__abc_21380_n6401) );
  OR2X2 OR2X2_24 ( .A(_abc_19068_n938), .B(_abc_19068_n952_1), .Y(_abc_19068_n953) );
  OR2X2 OR2X2_240 ( .A(_abc_19068_n1248), .B(_abc_19068_n1413_1), .Y(_abc_19068_n1414) );
  OR2X2 OR2X2_2400 ( .A(core__abc_21380_n6400), .B(core__abc_21380_n6405), .Y(core__abc_21380_n6406) );
  OR2X2 OR2X2_2401 ( .A(core__abc_21380_n3317_bF_buf6), .B(core__abc_21380_n6406), .Y(core__abc_21380_n6407) );
  OR2X2 OR2X2_2402 ( .A(core__abc_21380_n6399), .B(core__abc_21380_n6407), .Y(core__abc_21380_n6408) );
  OR2X2 OR2X2_2403 ( .A(core__abc_21380_n3328_bF_buf7), .B(core_v3_reg_56_), .Y(core__abc_21380_n6409) );
  OR2X2 OR2X2_2404 ( .A(core__abc_21380_n6374), .B(core__abc_21380_n1705), .Y(core__abc_21380_n6416) );
  OR2X2 OR2X2_2405 ( .A(core__abc_21380_n6418), .B(core__abc_21380_n6419), .Y(core__abc_21380_n6420) );
  OR2X2 OR2X2_2406 ( .A(core__abc_21380_n6415), .B(core__abc_21380_n6426), .Y(core__abc_21380_n6427) );
  OR2X2 OR2X2_2407 ( .A(core__abc_21380_n6414), .B(core__abc_21380_n6428), .Y(core__abc_21380_n6429) );
  OR2X2 OR2X2_2408 ( .A(core__abc_21380_n6430), .B(core__abc_21380_n5535), .Y(core__abc_21380_n6431) );
  OR2X2 OR2X2_2409 ( .A(core__abc_21380_n6432), .B(core__abc_21380_n5534), .Y(core__abc_21380_n6433) );
  OR2X2 OR2X2_241 ( .A(_abc_19068_n1415_1), .B(_abc_19068_n1416), .Y(_abc_19068_n1417_1) );
  OR2X2 OR2X2_2410 ( .A(core_v3_reg_57_), .B(core_mi_57_), .Y(core__abc_21380_n6437) );
  OR2X2 OR2X2_2411 ( .A(core__abc_21380_n6436), .B(core__abc_21380_n6441), .Y(core__abc_21380_n6442) );
  OR2X2 OR2X2_2412 ( .A(core__abc_21380_n3317_bF_buf5), .B(core__abc_21380_n6442), .Y(core__abc_21380_n6443) );
  OR2X2 OR2X2_2413 ( .A(core__abc_21380_n6435), .B(core__abc_21380_n6443), .Y(core__abc_21380_n6444) );
  OR2X2 OR2X2_2414 ( .A(core__abc_21380_n3328_bF_buf6), .B(core_v3_reg_57_), .Y(core__abc_21380_n6445) );
  OR2X2 OR2X2_2415 ( .A(core__abc_21380_n6424), .B(core__abc_21380_n6412), .Y(core__abc_21380_n6448) );
  OR2X2 OR2X2_2416 ( .A(core__abc_21380_n6452), .B(core__abc_21380_n6450), .Y(core__abc_21380_n6453) );
  OR2X2 OR2X2_2417 ( .A(core__abc_21380_n6378), .B(core__abc_21380_n6455), .Y(core__abc_21380_n6456) );
  OR2X2 OR2X2_2418 ( .A(core__abc_21380_n6459), .B(core__abc_21380_n6460), .Y(core__abc_21380_n6461) );
  OR2X2 OR2X2_2419 ( .A(core__abc_21380_n6464), .B(core__abc_21380_n6463), .Y(core__abc_21380_n6465) );
  OR2X2 OR2X2_242 ( .A(_abc_19068_n1414), .B(_abc_19068_n1417_1), .Y(_abc_19068_n1418) );
  OR2X2 OR2X2_2420 ( .A(core__abc_21380_n6466), .B(core__abc_21380_n6468), .Y(core__abc_21380_n6469) );
  OR2X2 OR2X2_2421 ( .A(core__abc_21380_n6470), .B(core__abc_21380_n5577), .Y(core__abc_21380_n6471) );
  OR2X2 OR2X2_2422 ( .A(core__abc_21380_n6469), .B(core__abc_21380_n5576), .Y(core__abc_21380_n6472) );
  OR2X2 OR2X2_2423 ( .A(core_v3_reg_58_), .B(core_mi_58_), .Y(core__abc_21380_n6477) );
  OR2X2 OR2X2_2424 ( .A(core__abc_21380_n6476), .B(core__abc_21380_n6481), .Y(core__abc_21380_n6482) );
  OR2X2 OR2X2_2425 ( .A(core__abc_21380_n3317_bF_buf4), .B(core__abc_21380_n6482), .Y(core__abc_21380_n6483) );
  OR2X2 OR2X2_2426 ( .A(core__abc_21380_n6474), .B(core__abc_21380_n6483), .Y(core__abc_21380_n6484) );
  OR2X2 OR2X2_2427 ( .A(core__abc_21380_n3328_bF_buf5), .B(core_v3_reg_58_), .Y(core__abc_21380_n6485) );
  OR2X2 OR2X2_2428 ( .A(core__abc_21380_n6468), .B(core__abc_21380_n6463), .Y(core__abc_21380_n6488) );
  OR2X2 OR2X2_2429 ( .A(core__abc_21380_n6459), .B(core__abc_21380_n1741), .Y(core__abc_21380_n6489) );
  OR2X2 OR2X2_243 ( .A(_abc_19068_n1420), .B(_abc_19068_n1421_1), .Y(_abc_19068_n1422) );
  OR2X2 OR2X2_2430 ( .A(core__abc_21380_n6491), .B(core__abc_21380_n6492), .Y(core__abc_21380_n6493) );
  OR2X2 OR2X2_2431 ( .A(core__abc_21380_n4430), .B(core__abc_21380_n6494), .Y(core__abc_21380_n6497) );
  OR2X2 OR2X2_2432 ( .A(core__abc_21380_n6488), .B(core__abc_21380_n6498), .Y(core__abc_21380_n6499) );
  OR2X2 OR2X2_2433 ( .A(core__abc_21380_n6501), .B(core__abc_21380_n6495), .Y(core__abc_21380_n6502) );
  OR2X2 OR2X2_2434 ( .A(core__abc_21380_n6500), .B(core__abc_21380_n6502), .Y(core__abc_21380_n6503) );
  OR2X2 OR2X2_2435 ( .A(core__abc_21380_n6505), .B(core__abc_21380_n5631), .Y(core__abc_21380_n6506) );
  OR2X2 OR2X2_2436 ( .A(core__abc_21380_n6504), .B(core__abc_21380_n5628), .Y(core__abc_21380_n6507) );
  OR2X2 OR2X2_2437 ( .A(core_v3_reg_59_), .B(core_mi_59_), .Y(core__abc_21380_n6511) );
  OR2X2 OR2X2_2438 ( .A(core__abc_21380_n6510), .B(core__abc_21380_n6515), .Y(core__abc_21380_n6516) );
  OR2X2 OR2X2_2439 ( .A(core__abc_21380_n3317_bF_buf3), .B(core__abc_21380_n6516), .Y(core__abc_21380_n6517) );
  OR2X2 OR2X2_244 ( .A(_abc_19068_n1422), .B(_abc_19068_n1419_1), .Y(_abc_19068_n1423_1) );
  OR2X2 OR2X2_2440 ( .A(core__abc_21380_n6509), .B(core__abc_21380_n6517), .Y(core__abc_21380_n6518) );
  OR2X2 OR2X2_2441 ( .A(core__abc_21380_n3328_bF_buf4), .B(core_v3_reg_59_), .Y(core__abc_21380_n6519) );
  OR2X2 OR2X2_2442 ( .A(core__abc_21380_n6527), .B(core__abc_21380_n6501), .Y(core__abc_21380_n6528) );
  OR2X2 OR2X2_2443 ( .A(core__abc_21380_n6525), .B(core__abc_21380_n6529), .Y(core__abc_21380_n6530) );
  OR2X2 OR2X2_2444 ( .A(core__abc_21380_n6524), .B(core__abc_21380_n6530), .Y(core__abc_21380_n6531) );
  OR2X2 OR2X2_2445 ( .A(core__abc_21380_n6532), .B(core__abc_21380_n3257), .Y(core__abc_21380_n6533) );
  OR2X2 OR2X2_2446 ( .A(core__abc_21380_n6535), .B(core__abc_21380_n6536), .Y(core__abc_21380_n6537) );
  OR2X2 OR2X2_2447 ( .A(core__abc_21380_n6538), .B(core__abc_21380_n6540), .Y(core__abc_21380_n6541) );
  OR2X2 OR2X2_2448 ( .A(core__abc_21380_n6502), .B(core__abc_21380_n6465), .Y(core__abc_21380_n6545) );
  OR2X2 OR2X2_2449 ( .A(core__abc_21380_n6545), .B(core__abc_21380_n6544), .Y(core__abc_21380_n6546) );
  OR2X2 OR2X2_245 ( .A(_abc_19068_n1424), .B(_abc_19068_n1425_1), .Y(_abc_19068_n1426) );
  OR2X2 OR2X2_2450 ( .A(core__abc_21380_n6371), .B(core__abc_21380_n6546), .Y(core__abc_21380_n6547) );
  OR2X2 OR2X2_2451 ( .A(core__abc_21380_n6545), .B(core__abc_21380_n6449), .Y(core__abc_21380_n6548) );
  OR2X2 OR2X2_2452 ( .A(core__abc_21380_n6551), .B(core__abc_21380_n6543), .Y(core__abc_21380_n6552) );
  OR2X2 OR2X2_2453 ( .A(core__abc_21380_n6553), .B(core__abc_21380_n5672), .Y(core__abc_21380_n6554) );
  OR2X2 OR2X2_2454 ( .A(core__abc_21380_n6552), .B(core__abc_21380_n5681), .Y(core__abc_21380_n6555) );
  OR2X2 OR2X2_2455 ( .A(core_v3_reg_60_), .B(core_mi_60_), .Y(core__abc_21380_n6560) );
  OR2X2 OR2X2_2456 ( .A(core__abc_21380_n6559), .B(core__abc_21380_n6564), .Y(core__abc_21380_n6565) );
  OR2X2 OR2X2_2457 ( .A(core__abc_21380_n3317_bF_buf2), .B(core__abc_21380_n6565), .Y(core__abc_21380_n6566) );
  OR2X2 OR2X2_2458 ( .A(core__abc_21380_n6557), .B(core__abc_21380_n6566), .Y(core__abc_21380_n6567) );
  OR2X2 OR2X2_2459 ( .A(core__abc_21380_n3328_bF_buf3), .B(core_v3_reg_60_), .Y(core__abc_21380_n6568) );
  OR2X2 OR2X2_246 ( .A(_abc_19068_n1427), .B(_abc_19068_n1428_1), .Y(_abc_19068_n1429) );
  OR2X2 OR2X2_2460 ( .A(core__abc_21380_n6543), .B(core__abc_21380_n6540), .Y(core__abc_21380_n6571) );
  OR2X2 OR2X2_2461 ( .A(core__abc_21380_n6536), .B(core__abc_21380_n1780), .Y(core__abc_21380_n6572) );
  OR2X2 OR2X2_2462 ( .A(core__abc_21380_n6574), .B(core__abc_21380_n6575), .Y(core__abc_21380_n6576) );
  OR2X2 OR2X2_2463 ( .A(core__abc_21380_n4554), .B(core__abc_21380_n6577), .Y(core__abc_21380_n6579) );
  OR2X2 OR2X2_2464 ( .A(core__abc_21380_n6580), .B(core__abc_21380_n6578), .Y(core__abc_21380_n6581) );
  OR2X2 OR2X2_2465 ( .A(core__abc_21380_n6571), .B(core__abc_21380_n6581), .Y(core__abc_21380_n6582) );
  OR2X2 OR2X2_2466 ( .A(core__abc_21380_n6583), .B(core__abc_21380_n6585), .Y(core__abc_21380_n6586) );
  OR2X2 OR2X2_2467 ( .A(core__abc_21380_n6588), .B(core__abc_21380_n5726), .Y(core__abc_21380_n6589) );
  OR2X2 OR2X2_2468 ( .A(core__abc_21380_n6587), .B(core__abc_21380_n5725), .Y(core__abc_21380_n6590) );
  OR2X2 OR2X2_2469 ( .A(core_v3_reg_61_), .B(core_mi_61_), .Y(core__abc_21380_n6595) );
  OR2X2 OR2X2_247 ( .A(_abc_19068_n1426), .B(_abc_19068_n1429), .Y(_abc_19068_n1430_1) );
  OR2X2 OR2X2_2470 ( .A(core__abc_21380_n6594), .B(core__abc_21380_n6599), .Y(core__abc_21380_n6600) );
  OR2X2 OR2X2_2471 ( .A(core__abc_21380_n3317_bF_buf1), .B(core__abc_21380_n6600), .Y(core__abc_21380_n6601) );
  OR2X2 OR2X2_2472 ( .A(core__abc_21380_n6592), .B(core__abc_21380_n6601), .Y(core__abc_21380_n6602) );
  OR2X2 OR2X2_2473 ( .A(core__abc_21380_n3328_bF_buf2), .B(core_v3_reg_61_), .Y(core__abc_21380_n6603) );
  OR2X2 OR2X2_2474 ( .A(core__abc_21380_n6608), .B(core__abc_21380_n6578), .Y(core__abc_21380_n6609) );
  OR2X2 OR2X2_2475 ( .A(core__abc_21380_n6607), .B(core__abc_21380_n6609), .Y(core__abc_21380_n6610) );
  OR2X2 OR2X2_2476 ( .A(core__abc_21380_n6611), .B(core__abc_21380_n3264), .Y(core__abc_21380_n6612) );
  OR2X2 OR2X2_2477 ( .A(core__abc_21380_n6612), .B(core__abc_21380_n1820), .Y(core__abc_21380_n6615) );
  OR2X2 OR2X2_2478 ( .A(core__abc_21380_n6617), .B(core__abc_21380_n6619), .Y(core__abc_21380_n6620) );
  OR2X2 OR2X2_2479 ( .A(core__abc_21380_n6610), .B(core__abc_21380_n6621), .Y(core__abc_21380_n6622) );
  OR2X2 OR2X2_248 ( .A(_abc_19068_n1430_1), .B(_abc_19068_n1423_1), .Y(_abc_19068_n1431) );
  OR2X2 OR2X2_2480 ( .A(core__abc_21380_n6581), .B(core__abc_21380_n6541), .Y(core__abc_21380_n6623) );
  OR2X2 OR2X2_2481 ( .A(core__abc_21380_n6550), .B(core__abc_21380_n6623), .Y(core__abc_21380_n6624) );
  OR2X2 OR2X2_2482 ( .A(core__abc_21380_n6627), .B(core__abc_21380_n6620), .Y(core__abc_21380_n6628) );
  OR2X2 OR2X2_2483 ( .A(core__abc_21380_n6630), .B(core__abc_21380_n5770), .Y(core__abc_21380_n6631) );
  OR2X2 OR2X2_2484 ( .A(core__abc_21380_n6629), .B(core__abc_21380_n5771), .Y(core__abc_21380_n6632) );
  OR2X2 OR2X2_2485 ( .A(core_v3_reg_62_), .B(core_mi_62_), .Y(core__abc_21380_n6637) );
  OR2X2 OR2X2_2486 ( .A(core__abc_21380_n6636), .B(core__abc_21380_n6641), .Y(core__abc_21380_n6642) );
  OR2X2 OR2X2_2487 ( .A(core__abc_21380_n3317_bF_buf0), .B(core__abc_21380_n6642), .Y(core__abc_21380_n6643) );
  OR2X2 OR2X2_2488 ( .A(core__abc_21380_n6634), .B(core__abc_21380_n6643), .Y(core__abc_21380_n6644) );
  OR2X2 OR2X2_2489 ( .A(core__abc_21380_n3328_bF_buf1), .B(core_v3_reg_62_), .Y(core__abc_21380_n6645) );
  OR2X2 OR2X2_249 ( .A(_abc_19068_n1431), .B(_abc_19068_n1418), .Y(_abc_19068_n1432_1) );
  OR2X2 OR2X2_2490 ( .A(core__abc_21380_n6648), .B(core__abc_21380_n6617), .Y(core__abc_21380_n6649) );
  OR2X2 OR2X2_2491 ( .A(core__abc_21380_n6613), .B(core__abc_21380_n1818), .Y(core__abc_21380_n6650) );
  OR2X2 OR2X2_2492 ( .A(core__abc_21380_n6650), .B(core__abc_21380_n1839), .Y(core__abc_21380_n6651) );
  OR2X2 OR2X2_2493 ( .A(core__abc_21380_n6649), .B(core__abc_21380_n6660), .Y(core__abc_21380_n6661) );
  OR2X2 OR2X2_2494 ( .A(core__abc_21380_n6655), .B(core__abc_21380_n6658), .Y(core__abc_21380_n6664) );
  OR2X2 OR2X2_2495 ( .A(core__abc_21380_n6663), .B(core__abc_21380_n6664), .Y(core__abc_21380_n6665) );
  OR2X2 OR2X2_2496 ( .A(core__abc_21380_n6667), .B(core__abc_21380_n5812), .Y(core__abc_21380_n6668) );
  OR2X2 OR2X2_2497 ( .A(core__abc_21380_n6666), .B(core__abc_21380_n5811), .Y(core__abc_21380_n6669) );
  OR2X2 OR2X2_2498 ( .A(core_v3_reg_63_), .B(core_mi_63_), .Y(core__abc_21380_n6673) );
  OR2X2 OR2X2_2499 ( .A(core__abc_21380_n6672), .B(core__abc_21380_n6677), .Y(core__abc_21380_n6678) );
  OR2X2 OR2X2_25 ( .A(_abc_19068_n955_1), .B(_abc_19068_n956), .Y(_abc_19068_n957_1) );
  OR2X2 OR2X2_250 ( .A(_abc_19068_n1434_1), .B(_abc_19068_n1435), .Y(_abc_19068_n1436_1) );
  OR2X2 OR2X2_2500 ( .A(core__abc_21380_n3317_bF_buf7), .B(core__abc_21380_n6678), .Y(core__abc_21380_n6679) );
  OR2X2 OR2X2_2501 ( .A(core__abc_21380_n6671), .B(core__abc_21380_n6679), .Y(core__abc_21380_n6680) );
  OR2X2 OR2X2_2502 ( .A(core__abc_21380_n3328_bF_buf0), .B(core_v3_reg_63_), .Y(core__abc_21380_n6681) );
  OR2X2 OR2X2_2503 ( .A(core__abc_21380_n6654), .B(core__abc_21380_n6684), .Y(core__abc_21380_n6685) );
  OR2X2 OR2X2_2504 ( .A(core__abc_21380_n6688), .B(core__abc_21380_n5261), .Y(core__abc_21380_n6689) );
  OR2X2 OR2X2_2505 ( .A(core__abc_21380_n6690), .B(core__abc_21380_n6686), .Y(core__abc_21380_n6691) );
  OR2X2 OR2X2_2506 ( .A(core__abc_21380_n6691), .B(core__abc_21380_n5264), .Y(core__abc_21380_n6692) );
  OR2X2 OR2X2_2507 ( .A(core__abc_21380_n6616), .B(core__abc_21380_n1577), .Y(core__abc_21380_n6694) );
  OR2X2 OR2X2_2508 ( .A(core__abc_21380_n6618), .B(core_v1_reg_17_), .Y(core__abc_21380_n6695) );
  OR2X2 OR2X2_2509 ( .A(core__abc_21380_n6698), .B(core__abc_21380_n6699), .Y(core__abc_21380_n6700) );
  OR2X2 OR2X2_251 ( .A(_abc_19068_n1438_1), .B(_abc_19068_n1439), .Y(_abc_19068_n1440_1) );
  OR2X2 OR2X2_2510 ( .A(core__abc_21380_n6705), .B(core__abc_21380_n6704), .Y(core__abc_21380_n6706) );
  OR2X2 OR2X2_2511 ( .A(core__abc_21380_n6539), .B(core__abc_21380_n1537), .Y(core__abc_21380_n6713) );
  OR2X2 OR2X2_2512 ( .A(core__abc_21380_n6537), .B(core_v1_reg_15_), .Y(core__abc_21380_n6714) );
  OR2X2 OR2X2_2513 ( .A(core__abc_21380_n6717), .B(core__abc_21380_n6718), .Y(core__abc_21380_n6719) );
  OR2X2 OR2X2_2514 ( .A(core__abc_21380_n6493), .B(core_v1_reg_14_), .Y(core__abc_21380_n6725) );
  OR2X2 OR2X2_2515 ( .A(core__abc_21380_n6726), .B(core__abc_21380_n5037), .Y(core__abc_21380_n6727) );
  OR2X2 OR2X2_2516 ( .A(core__abc_21380_n6462), .B(core__abc_21380_n1501), .Y(core__abc_21380_n6731) );
  OR2X2 OR2X2_2517 ( .A(core__abc_21380_n6461), .B(core_v1_reg_13_), .Y(core__abc_21380_n6732) );
  OR2X2 OR2X2_2518 ( .A(core__abc_21380_n6735), .B(core__abc_21380_n6736), .Y(core__abc_21380_n6737) );
  OR2X2 OR2X2_2519 ( .A(core__abc_21380_n6741), .B(core__abc_21380_n6740), .Y(core__abc_21380_n6742) );
  OR2X2 OR2X2_252 ( .A(_abc_19068_n1440_1), .B(_abc_19068_n1437), .Y(_abc_19068_n1441) );
  OR2X2 OR2X2_2520 ( .A(core__abc_21380_n6381), .B(core__abc_21380_n6748), .Y(core__abc_21380_n6749) );
  OR2X2 OR2X2_2521 ( .A(core__abc_21380_n6380), .B(core_v1_reg_11_), .Y(core__abc_21380_n6750) );
  OR2X2 OR2X2_2522 ( .A(core__abc_21380_n6728), .B(core__abc_21380_n6759), .Y(core__abc_21380_n6760) );
  OR2X2 OR2X2_2523 ( .A(core__abc_21380_n6758), .B(core__abc_21380_n6762), .Y(core__abc_21380_n6763) );
  OR2X2 OR2X2_2524 ( .A(core__abc_21380_n6770), .B(core__abc_21380_n6771), .Y(core__abc_21380_n6772) );
  OR2X2 OR2X2_2525 ( .A(core__abc_21380_n6769), .B(core__abc_21380_n6774), .Y(core__abc_21380_n6775) );
  OR2X2 OR2X2_2526 ( .A(core__abc_21380_n6775), .B(core__abc_21380_n6764), .Y(core__abc_21380_n6776) );
  OR2X2 OR2X2_2527 ( .A(core__abc_21380_n6753), .B(core__abc_21380_n6778), .Y(core__abc_21380_n6779) );
  OR2X2 OR2X2_2528 ( .A(core__abc_21380_n6323), .B(core__abc_21380_n6784), .Y(core__abc_21380_n6785) );
  OR2X2 OR2X2_2529 ( .A(core__abc_21380_n6788), .B(core__abc_21380_n4814_1), .Y(core__abc_21380_n6789) );
  OR2X2 OR2X2_253 ( .A(_abc_19068_n1441), .B(_abc_19068_n1436_1), .Y(_abc_19068_n1442_1) );
  OR2X2 OR2X2_2530 ( .A(core__abc_21380_n6791), .B(core__abc_21380_n6786), .Y(core__abc_21380_n6792) );
  OR2X2 OR2X2_2531 ( .A(core__abc_21380_n6792), .B(core__abc_21380_n6790), .Y(core__abc_21380_n6793) );
  OR2X2 OR2X2_2532 ( .A(core__abc_21380_n6291), .B(core__abc_21380_n1431), .Y(core__abc_21380_n6795) );
  OR2X2 OR2X2_2533 ( .A(core__abc_21380_n6293), .B(core_v1_reg_9_), .Y(core__abc_21380_n6796) );
  OR2X2 OR2X2_2534 ( .A(core__abc_21380_n6799), .B(core__abc_21380_n6800), .Y(core__abc_21380_n6801) );
  OR2X2 OR2X2_2535 ( .A(core__abc_21380_n6806), .B(core__abc_21380_n6805), .Y(core__abc_21380_n6807) );
  OR2X2 OR2X2_2536 ( .A(core__abc_21380_n6218), .B(core__abc_21380_n1393), .Y(core__abc_21380_n6814) );
  OR2X2 OR2X2_2537 ( .A(core__abc_21380_n6217), .B(core_v1_reg_7_), .Y(core__abc_21380_n6815) );
  OR2X2 OR2X2_2538 ( .A(core__abc_21380_n6818), .B(core__abc_21380_n6819), .Y(core__abc_21380_n6820) );
  OR2X2 OR2X2_2539 ( .A(core__abc_21380_n6824), .B(core__abc_21380_n6825), .Y(core__abc_21380_n6826) );
  OR2X2 OR2X2_254 ( .A(_abc_19068_n1444_1), .B(_abc_19068_n1445), .Y(_abc_19068_n1446_1) );
  OR2X2 OR2X2_2540 ( .A(core__abc_21380_n6826), .B(core__abc_21380_n4599), .Y(core__abc_21380_n6829) );
  OR2X2 OR2X2_2541 ( .A(core__abc_21380_n6142), .B(core__abc_21380_n1356), .Y(core__abc_21380_n6831) );
  OR2X2 OR2X2_2542 ( .A(core__abc_21380_n6144), .B(core_v1_reg_5_), .Y(core__abc_21380_n6832) );
  OR2X2 OR2X2_2543 ( .A(core__abc_21380_n6835), .B(core__abc_21380_n6836), .Y(core__abc_21380_n6837) );
  OR2X2 OR2X2_2544 ( .A(core__abc_21380_n6842), .B(core__abc_21380_n6841), .Y(core__abc_21380_n6843) );
  OR2X2 OR2X2_2545 ( .A(core__abc_21380_n6049), .B(core__abc_21380_n1319), .Y(core__abc_21380_n6846) );
  OR2X2 OR2X2_2546 ( .A(core__abc_21380_n6048), .B(core_v1_reg_3_), .Y(core__abc_21380_n6847) );
  OR2X2 OR2X2_2547 ( .A(core__abc_21380_n6853), .B(core__abc_21380_n6845), .Y(core__abc_21380_n6854) );
  OR2X2 OR2X2_2548 ( .A(core__abc_21380_n6858), .B(core__abc_21380_n6856), .Y(core__abc_21380_n6859) );
  OR2X2 OR2X2_2549 ( .A(core__abc_21380_n6855), .B(core__abc_21380_n6860), .Y(core__abc_21380_n6861) );
  OR2X2 OR2X2_255 ( .A(_abc_19068_n1447), .B(_abc_19068_n1448_1), .Y(_abc_19068_n1449) );
  OR2X2 OR2X2_2550 ( .A(core__abc_21380_n6868), .B(core__abc_21380_n6869), .Y(core__abc_21380_n6870) );
  OR2X2 OR2X2_2551 ( .A(core__abc_21380_n6867), .B(core__abc_21380_n6872), .Y(core__abc_21380_n6873) );
  OR2X2 OR2X2_2552 ( .A(core__abc_21380_n6873), .B(core__abc_21380_n6862), .Y(core__abc_21380_n6874) );
  OR2X2 OR2X2_2553 ( .A(core__abc_21380_n6876), .B(core__abc_21380_n6875), .Y(core__abc_21380_n6877) );
  OR2X2 OR2X2_2554 ( .A(core__abc_21380_n6877), .B(core__abc_21380_n4308), .Y(core__abc_21380_n6880) );
  OR2X2 OR2X2_2555 ( .A(core__abc_21380_n5968), .B(core__abc_21380_n1289), .Y(core__abc_21380_n6882) );
  OR2X2 OR2X2_2556 ( .A(core__abc_21380_n5970), .B(core_v1_reg_1_), .Y(core__abc_21380_n6883) );
  OR2X2 OR2X2_2557 ( .A(core__abc_21380_n6886), .B(core__abc_21380_n6887), .Y(core__abc_21380_n6888) );
  OR2X2 OR2X2_2558 ( .A(core__abc_21380_n6893), .B(core__abc_21380_n6892), .Y(core__abc_21380_n6894) );
  OR2X2 OR2X2_2559 ( .A(core__abc_21380_n5896), .B(core__abc_21380_n2432), .Y(core__abc_21380_n6899) );
  OR2X2 OR2X2_256 ( .A(_abc_19068_n1446_1), .B(_abc_19068_n1449), .Y(_abc_19068_n1450_1) );
  OR2X2 OR2X2_2560 ( .A(core__abc_21380_n5895), .B(core_v1_reg_63_), .Y(core__abc_21380_n6900) );
  OR2X2 OR2X2_2561 ( .A(core__abc_21380_n6905), .B(core__abc_21380_n6895), .Y(core__abc_21380_n6906) );
  OR2X2 OR2X2_2562 ( .A(core__abc_21380_n6878), .B(core__abc_21380_n6886), .Y(core__abc_21380_n6909) );
  OR2X2 OR2X2_2563 ( .A(core__abc_21380_n6908), .B(core__abc_21380_n6910), .Y(core__abc_21380_n6911) );
  OR2X2 OR2X2_2564 ( .A(core__abc_21380_n6903), .B(core__abc_21380_n6914), .Y(core__abc_21380_n6915) );
  OR2X2 OR2X2_2565 ( .A(core__abc_21380_n5848), .B(core__abc_21380_n2413), .Y(core__abc_21380_n6919) );
  OR2X2 OR2X2_2566 ( .A(core__abc_21380_n5804), .B(core__abc_21380_n2395_1), .Y(core__abc_21380_n6924) );
  OR2X2 OR2X2_2567 ( .A(core__abc_21380_n5814), .B(core_v1_reg_61_), .Y(core__abc_21380_n6925) );
  OR2X2 OR2X2_2568 ( .A(core__abc_21380_n6922), .B(core__abc_21380_n4018_1), .Y(core__abc_21380_n6930) );
  OR2X2 OR2X2_2569 ( .A(core__abc_21380_n6931), .B(core__abc_21380_n6923), .Y(core__abc_21380_n6932) );
  OR2X2 OR2X2_257 ( .A(_abc_19068_n1450_1), .B(_abc_19068_n1443), .Y(_abc_19068_n1451) );
  OR2X2 OR2X2_2570 ( .A(core__abc_21380_n6935), .B(core__abc_21380_n6934), .Y(core__abc_21380_n6936) );
  OR2X2 OR2X2_2571 ( .A(core__abc_21380_n5717), .B(core__abc_21380_n2357), .Y(core__abc_21380_n6941) );
  OR2X2 OR2X2_2572 ( .A(core__abc_21380_n5716), .B(core_v1_reg_59_), .Y(core__abc_21380_n6942) );
  OR2X2 OR2X2_2573 ( .A(core__abc_21380_n6940), .B(core__abc_21380_n6946), .Y(core__abc_21380_n6947) );
  OR2X2 OR2X2_2574 ( .A(core__abc_21380_n6928), .B(core__abc_21380_n6952), .Y(core__abc_21380_n6953) );
  OR2X2 OR2X2_2575 ( .A(core__abc_21380_n6956), .B(core__abc_21380_n6933), .Y(core__abc_21380_n6957) );
  OR2X2 OR2X2_2576 ( .A(core__abc_21380_n6958), .B(core__abc_21380_n6959), .Y(core__abc_21380_n6960) );
  OR2X2 OR2X2_2577 ( .A(core__abc_21380_n5617), .B(core__abc_21380_n2321), .Y(core__abc_21380_n6965) );
  OR2X2 OR2X2_2578 ( .A(core__abc_21380_n5630), .B(core_v1_reg_57_), .Y(core__abc_21380_n6966) );
  OR2X2 OR2X2_2579 ( .A(core__abc_21380_n6970), .B(core__abc_21380_n6961), .Y(core__abc_21380_n6971) );
  OR2X2 OR2X2_258 ( .A(_abc_19068_n1451), .B(_abc_19068_n1442_1), .Y(_abc_19068_n1452_1) );
  OR2X2 OR2X2_2580 ( .A(core__abc_21380_n6969), .B(core__abc_21380_n6974), .Y(core__abc_21380_n6975) );
  OR2X2 OR2X2_2581 ( .A(core__abc_21380_n6979), .B(core__abc_21380_n6978), .Y(core__abc_21380_n6980) );
  OR2X2 OR2X2_2582 ( .A(core__abc_21380_n6982), .B(core__abc_21380_n6983), .Y(core__abc_21380_n6984) );
  OR2X2 OR2X2_2583 ( .A(core__abc_21380_n5523), .B(core__abc_21380_n2283), .Y(core__abc_21380_n6986) );
  OR2X2 OR2X2_2584 ( .A(core__abc_21380_n5522), .B(core_v1_reg_55_), .Y(core__abc_21380_n6987) );
  OR2X2 OR2X2_2585 ( .A(core__abc_21380_n6992), .B(core__abc_21380_n6991), .Y(core__abc_21380_n6993) );
  OR2X2 OR2X2_2586 ( .A(core__abc_21380_n6993), .B(core__abc_21380_n3471), .Y(core__abc_21380_n6994) );
  OR2X2 OR2X2_2587 ( .A(core__abc_21380_n5427), .B(core__abc_21380_n2247_1), .Y(core__abc_21380_n6999) );
  OR2X2 OR2X2_2588 ( .A(core__abc_21380_n5426), .B(core_v1_reg_53_), .Y(core__abc_21380_n7000) );
  OR2X2 OR2X2_2589 ( .A(core__abc_21380_n5376), .B(core__abc_21380_n7004), .Y(core__abc_21380_n7005) );
  OR2X2 OR2X2_259 ( .A(_abc_19068_n1248), .B(_abc_19068_n1454_1), .Y(_abc_19068_n1455) );
  OR2X2 OR2X2_2590 ( .A(core__abc_21380_n5375), .B(core_v1_reg_52_), .Y(core__abc_21380_n7006) );
  OR2X2 OR2X2_2591 ( .A(core__abc_21380_n7010), .B(core__abc_21380_n7011), .Y(core__abc_21380_n7012) );
  OR2X2 OR2X2_2592 ( .A(core__abc_21380_n7018), .B(core__abc_21380_n7009), .Y(core__abc_21380_n7019) );
  OR2X2 OR2X2_2593 ( .A(core__abc_21380_n7024), .B(core__abc_21380_n7003), .Y(core__abc_21380_n7025) );
  OR2X2 OR2X2_2594 ( .A(core__abc_21380_n7026), .B(core__abc_21380_n6995), .Y(core__abc_21380_n7027) );
  OR2X2 OR2X2_2595 ( .A(core__abc_21380_n6990), .B(core__abc_21380_n7028), .Y(core__abc_21380_n7029) );
  OR2X2 OR2X2_2596 ( .A(core__abc_21380_n7031), .B(core__abc_21380_n6990), .Y(core__abc_21380_n7032) );
  OR2X2 OR2X2_2597 ( .A(core__abc_21380_n7033), .B(core__abc_21380_n6982), .Y(core__abc_21380_n7034) );
  OR2X2 OR2X2_2598 ( .A(core__abc_21380_n7035), .B(core__abc_21380_n6971), .Y(core__abc_21380_n7036) );
  OR2X2 OR2X2_2599 ( .A(core__abc_21380_n6945), .B(core__abc_21380_n7039), .Y(core__abc_21380_n7040) );
  OR2X2 OR2X2_26 ( .A(_abc_19068_n958_1), .B(_abc_19068_n959), .Y(_abc_19068_n960_1) );
  OR2X2 OR2X2_260 ( .A(_abc_19068_n1456_1), .B(_abc_19068_n1457), .Y(_abc_19068_n1458_1) );
  OR2X2 OR2X2_2600 ( .A(core__abc_21380_n7044), .B(core__abc_21380_n6957), .Y(core__abc_21380_n7045) );
  OR2X2 OR2X2_2601 ( .A(core__abc_21380_n7046), .B(core__abc_21380_n6911), .Y(core__abc_21380_n7047) );
  OR2X2 OR2X2_2602 ( .A(core__abc_21380_n6850), .B(core__abc_21380_n7050), .Y(core__abc_21380_n7051) );
  OR2X2 OR2X2_2603 ( .A(core__abc_21380_n6874), .B(core__abc_21380_n7056), .Y(core__abc_21380_n7057) );
  OR2X2 OR2X2_2604 ( .A(core__abc_21380_n6776), .B(core__abc_21380_n7058), .Y(core__abc_21380_n7059) );
  OR2X2 OR2X2_2605 ( .A(core__abc_21380_n3290), .B(core__abc_21380_n7061), .Y(core__abc_21380_n7062) );
  OR2X2 OR2X2_2606 ( .A(core__abc_21380_n3289), .B(core_v1_reg_19_), .Y(core__abc_21380_n7063) );
  OR2X2 OR2X2_2607 ( .A(core__abc_21380_n7066), .B(core__abc_21380_n7067), .Y(core__abc_21380_n7068) );
  OR2X2 OR2X2_2608 ( .A(core__abc_21380_n7069), .B(core__abc_21380_n7071), .Y(core__abc_21380_n7072) );
  OR2X2 OR2X2_2609 ( .A(core__abc_21380_n7075), .B(core__abc_21380_n3311), .Y(core__abc_21380_n7076) );
  OR2X2 OR2X2_261 ( .A(_abc_19068_n1455), .B(_abc_19068_n1458_1), .Y(_abc_19068_n1459) );
  OR2X2 OR2X2_2610 ( .A(core__abc_21380_n7079), .B(core_v2_reg_0_), .Y(core__abc_21380_n7080) );
  OR2X2 OR2X2_2611 ( .A(core__abc_21380_n1264_1), .B(core_long), .Y(core__abc_21380_n7081) );
  OR2X2 OR2X2_2612 ( .A(core__abc_21380_n7078), .B(core__abc_21380_n7083), .Y(core__abc_21380_n7084) );
  OR2X2 OR2X2_2613 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n7084), .Y(core__abc_21380_n7085) );
  OR2X2 OR2X2_2614 ( .A(core__abc_21380_n7074), .B(core__abc_21380_n7085), .Y(core__abc_21380_n7086) );
  OR2X2 OR2X2_2615 ( .A(core__abc_21380_n7087_bF_buf7), .B(core_v2_reg_0_), .Y(core__abc_21380_n7088) );
  OR2X2 OR2X2_2616 ( .A(core__abc_21380_n7092), .B(core__abc_21380_n7091), .Y(core__abc_21380_n7093) );
  OR2X2 OR2X2_2617 ( .A(core__abc_21380_n7094), .B(core__abc_21380_n7096), .Y(core__abc_21380_n7097) );
  OR2X2 OR2X2_2618 ( .A(core__abc_21380_n7100), .B(core__abc_21380_n7097), .Y(core__abc_21380_n7102) );
  OR2X2 OR2X2_2619 ( .A(core__abc_21380_n7103), .B(core__abc_21380_n7101), .Y(core__abc_21380_n7104) );
  OR2X2 OR2X2_262 ( .A(_abc_19068_n1461), .B(_abc_19068_n1462_1), .Y(_abc_19068_n1463) );
  OR2X2 OR2X2_2620 ( .A(core__abc_21380_n7107), .B(core__abc_21380_n7108), .Y(core__abc_21380_n7109) );
  OR2X2 OR2X2_2621 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n7109), .Y(core__abc_21380_n7110) );
  OR2X2 OR2X2_2622 ( .A(core__abc_21380_n7106), .B(core__abc_21380_n7110), .Y(core__abc_21380_n7111) );
  OR2X2 OR2X2_2623 ( .A(core__abc_21380_n7087_bF_buf6), .B(core_v2_reg_1_), .Y(core__abc_21380_n7112) );
  OR2X2 OR2X2_2624 ( .A(core__abc_21380_n7118), .B(core__abc_21380_n7094), .Y(core__abc_21380_n7119) );
  OR2X2 OR2X2_2625 ( .A(core__abc_21380_n7117), .B(core__abc_21380_n7119), .Y(core__abc_21380_n7120) );
  OR2X2 OR2X2_2626 ( .A(core__abc_21380_n3410), .B(core__abc_21380_n1647), .Y(core__abc_21380_n7122) );
  OR2X2 OR2X2_2627 ( .A(core__abc_21380_n3409), .B(core_v1_reg_21_), .Y(core__abc_21380_n7123) );
  OR2X2 OR2X2_2628 ( .A(core__abc_21380_n7126), .B(core__abc_21380_n7127), .Y(core__abc_21380_n7128) );
  OR2X2 OR2X2_2629 ( .A(core__abc_21380_n7129), .B(core__abc_21380_n7131), .Y(core__abc_21380_n7132) );
  OR2X2 OR2X2_263 ( .A(_abc_19068_n1463), .B(_abc_19068_n1460_1), .Y(_abc_19068_n1464_1) );
  OR2X2 OR2X2_2630 ( .A(core__abc_21380_n7135), .B(core__abc_21380_n7136), .Y(core__abc_21380_n7137) );
  OR2X2 OR2X2_2631 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n7137), .Y(core__abc_21380_n7138) );
  OR2X2 OR2X2_2632 ( .A(core__abc_21380_n7134), .B(core__abc_21380_n7138), .Y(core__abc_21380_n7139) );
  OR2X2 OR2X2_2633 ( .A(core__abc_21380_n7087_bF_buf5), .B(core_v2_reg_2_), .Y(core__abc_21380_n7140) );
  OR2X2 OR2X2_2634 ( .A(core__abc_21380_n7131), .B(core__abc_21380_n7126), .Y(core__abc_21380_n7143) );
  OR2X2 OR2X2_2635 ( .A(core__abc_21380_n7146), .B(core__abc_21380_n7145), .Y(core__abc_21380_n7147) );
  OR2X2 OR2X2_2636 ( .A(core__abc_21380_n7155), .B(core__abc_21380_n7156), .Y(core__abc_21380_n7157) );
  OR2X2 OR2X2_2637 ( .A(core__abc_21380_n7160), .B(core__abc_21380_n7161), .Y(core__abc_21380_n7162) );
  OR2X2 OR2X2_2638 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n7162), .Y(core__abc_21380_n7163) );
  OR2X2 OR2X2_2639 ( .A(core__abc_21380_n7159), .B(core__abc_21380_n7163), .Y(core__abc_21380_n7164) );
  OR2X2 OR2X2_264 ( .A(_abc_19068_n1465), .B(_abc_19068_n1466_1), .Y(_abc_19068_n1467) );
  OR2X2 OR2X2_2640 ( .A(core__abc_21380_n7087_bF_buf4), .B(core_v2_reg_3_), .Y(core__abc_21380_n7165) );
  OR2X2 OR2X2_2641 ( .A(core__abc_21380_n7168), .B(core__abc_21380_n7149), .Y(core__abc_21380_n7169) );
  OR2X2 OR2X2_2642 ( .A(core__abc_21380_n7171), .B(core__abc_21380_n7169), .Y(core__abc_21380_n7172) );
  OR2X2 OR2X2_2643 ( .A(core__abc_21380_n7174), .B(core__abc_21380_n7172), .Y(core__abc_21380_n7175) );
  OR2X2 OR2X2_2644 ( .A(core__abc_21380_n3538), .B(core__abc_21380_n1683), .Y(core__abc_21380_n7176) );
  OR2X2 OR2X2_2645 ( .A(core__abc_21380_n3537), .B(core_v1_reg_23_), .Y(core__abc_21380_n7177) );
  OR2X2 OR2X2_2646 ( .A(core__abc_21380_n7180), .B(core__abc_21380_n7181), .Y(core__abc_21380_n7182) );
  OR2X2 OR2X2_2647 ( .A(core__abc_21380_n7175), .B(core__abc_21380_n7183), .Y(core__abc_21380_n7186) );
  OR2X2 OR2X2_2648 ( .A(core__abc_21380_n1342), .B(core_long), .Y(core__abc_21380_n7190) );
  OR2X2 OR2X2_2649 ( .A(core__abc_21380_n7079), .B(core_v2_reg_4_), .Y(core__abc_21380_n7191) );
  OR2X2 OR2X2_265 ( .A(_abc_19068_n1468_1), .B(_abc_19068_n1469), .Y(_abc_19068_n1470_1) );
  OR2X2 OR2X2_2650 ( .A(core__abc_21380_n7189), .B(core__abc_21380_n7193), .Y(core__abc_21380_n7194) );
  OR2X2 OR2X2_2651 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n7194), .Y(core__abc_21380_n7195) );
  OR2X2 OR2X2_2652 ( .A(core__abc_21380_n7188), .B(core__abc_21380_n7195), .Y(core__abc_21380_n7196) );
  OR2X2 OR2X2_2653 ( .A(core__abc_21380_n7087_bF_buf3), .B(core_v2_reg_4_), .Y(core__abc_21380_n7197) );
  OR2X2 OR2X2_2654 ( .A(core__abc_21380_n7205), .B(core__abc_21380_n7204), .Y(core__abc_21380_n7206) );
  OR2X2 OR2X2_2655 ( .A(core__abc_21380_n7214), .B(core__abc_21380_n7215), .Y(core__abc_21380_n7216) );
  OR2X2 OR2X2_2656 ( .A(core__abc_21380_n7219), .B(core__abc_21380_n7220), .Y(core__abc_21380_n7221) );
  OR2X2 OR2X2_2657 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n7221), .Y(core__abc_21380_n7222) );
  OR2X2 OR2X2_2658 ( .A(core__abc_21380_n7217), .B(core__abc_21380_n7222), .Y(core__abc_21380_n7223) );
  OR2X2 OR2X2_2659 ( .A(core__abc_21380_n7087_bF_buf2), .B(core_v2_reg_5_), .Y(core__abc_21380_n7224) );
  OR2X2 OR2X2_266 ( .A(_abc_19068_n1467), .B(_abc_19068_n1470_1), .Y(_abc_19068_n1471) );
  OR2X2 OR2X2_2660 ( .A(core__abc_21380_n7227), .B(core__abc_21380_n1721), .Y(core__abc_21380_n7228) );
  OR2X2 OR2X2_2661 ( .A(core__abc_21380_n3686), .B(core_v1_reg_25_), .Y(core__abc_21380_n7229) );
  OR2X2 OR2X2_2662 ( .A(core__abc_21380_n7232), .B(core__abc_21380_n7233), .Y(core__abc_21380_n7234) );
  OR2X2 OR2X2_2663 ( .A(core__abc_21380_n7236), .B(core__abc_21380_n7210), .Y(core__abc_21380_n7237) );
  OR2X2 OR2X2_2664 ( .A(core__abc_21380_n7237), .B(core__abc_21380_n7234), .Y(core__abc_21380_n7239) );
  OR2X2 OR2X2_2665 ( .A(core__abc_21380_n7240), .B(core__abc_21380_n7238), .Y(core__abc_21380_n7241) );
  OR2X2 OR2X2_2666 ( .A(core__abc_21380_n7245), .B(core__abc_21380_n7246), .Y(core__abc_21380_n7247) );
  OR2X2 OR2X2_2667 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n7247), .Y(core__abc_21380_n7248) );
  OR2X2 OR2X2_2668 ( .A(core__abc_21380_n7243), .B(core__abc_21380_n7248), .Y(core__abc_21380_n7249) );
  OR2X2 OR2X2_2669 ( .A(core__abc_21380_n7087_bF_buf1), .B(core_v2_reg_6_), .Y(core__abc_21380_n7250) );
  OR2X2 OR2X2_267 ( .A(_abc_19068_n1471), .B(_abc_19068_n1464_1), .Y(_abc_19068_n1472_1) );
  OR2X2 OR2X2_2670 ( .A(core__abc_21380_n7257), .B(core__abc_21380_n7258), .Y(core__abc_21380_n7259) );
  OR2X2 OR2X2_2671 ( .A(core__abc_21380_n7261), .B(core__abc_21380_n7262), .Y(core__abc_21380_n7263) );
  OR2X2 OR2X2_2672 ( .A(core__abc_21380_n7254), .B(core__abc_21380_n7263), .Y(core__abc_21380_n7266) );
  OR2X2 OR2X2_2673 ( .A(core__abc_21380_n7269), .B(core__abc_21380_n7270), .Y(core__abc_21380_n7271) );
  OR2X2 OR2X2_2674 ( .A(core__abc_21380_n7076_bF_buf5), .B(core__abc_21380_n7271), .Y(core__abc_21380_n7272) );
  OR2X2 OR2X2_2675 ( .A(core__abc_21380_n7268), .B(core__abc_21380_n7272), .Y(core__abc_21380_n7273) );
  OR2X2 OR2X2_2676 ( .A(core__abc_21380_n7087_bF_buf0), .B(core_v2_reg_7_), .Y(core__abc_21380_n7274) );
  OR2X2 OR2X2_2677 ( .A(core__abc_21380_n7263), .B(core__abc_21380_n7234), .Y(core__abc_21380_n7278) );
  OR2X2 OR2X2_2678 ( .A(core__abc_21380_n7235), .B(core__abc_21380_n7210), .Y(core__abc_21380_n7285) );
  OR2X2 OR2X2_2679 ( .A(core__abc_21380_n7278), .B(core__abc_21380_n7285), .Y(core__abc_21380_n7286) );
  OR2X2 OR2X2_268 ( .A(_abc_19068_n1472_1), .B(_abc_19068_n1459), .Y(_abc_19068_n1473) );
  OR2X2 OR2X2_2680 ( .A(core__abc_21380_n7288), .B(core__abc_21380_n7261), .Y(core__abc_21380_n7289) );
  OR2X2 OR2X2_2681 ( .A(core__abc_21380_n7282), .B(core__abc_21380_n7293), .Y(core__abc_21380_n7294) );
  OR2X2 OR2X2_2682 ( .A(core__abc_21380_n3815), .B(core__abc_21380_n1758), .Y(core__abc_21380_n7295) );
  OR2X2 OR2X2_2683 ( .A(core__abc_21380_n3814_1), .B(core_v1_reg_27_), .Y(core__abc_21380_n7296) );
  OR2X2 OR2X2_2684 ( .A(core__abc_21380_n7299), .B(core__abc_21380_n7300), .Y(core__abc_21380_n7301) );
  OR2X2 OR2X2_2685 ( .A(core__abc_21380_n7305), .B(core__abc_21380_n7303), .Y(core__abc_21380_n7306) );
  OR2X2 OR2X2_2686 ( .A(core__abc_21380_n7309), .B(core__abc_21380_n7310), .Y(core__abc_21380_n7311) );
  OR2X2 OR2X2_2687 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n7311), .Y(core__abc_21380_n7312) );
  OR2X2 OR2X2_2688 ( .A(core__abc_21380_n7308), .B(core__abc_21380_n7312), .Y(core__abc_21380_n7313) );
  OR2X2 OR2X2_2689 ( .A(core__abc_21380_n7087_bF_buf7), .B(core_v2_reg_8_), .Y(core__abc_21380_n7314) );
  OR2X2 OR2X2_269 ( .A(_abc_19068_n1209_1), .B(_abc_19068_n1475), .Y(_abc_19068_n1476_1) );
  OR2X2 OR2X2_2690 ( .A(core__abc_21380_n3890), .B(core__abc_21380_n1778), .Y(core__abc_21380_n7322) );
  OR2X2 OR2X2_2691 ( .A(core__abc_21380_n7319), .B(core__abc_21380_n7330), .Y(core__abc_21380_n7333) );
  OR2X2 OR2X2_2692 ( .A(core__abc_21380_n7337), .B(core__abc_21380_n7338), .Y(core__abc_21380_n7339) );
  OR2X2 OR2X2_2693 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n7339), .Y(core__abc_21380_n7340) );
  OR2X2 OR2X2_2694 ( .A(core__abc_21380_n7335), .B(core__abc_21380_n7340), .Y(core__abc_21380_n7341) );
  OR2X2 OR2X2_2695 ( .A(core__abc_21380_n7087_bF_buf6), .B(core_v2_reg_9_), .Y(core__abc_21380_n7342) );
  OR2X2 OR2X2_2696 ( .A(core__abc_21380_n7327), .B(core__abc_21380_n7317), .Y(core__abc_21380_n7345) );
  OR2X2 OR2X2_2697 ( .A(core__abc_21380_n7349), .B(core__abc_21380_n7347), .Y(core__abc_21380_n7350) );
  OR2X2 OR2X2_2698 ( .A(core__abc_21380_n3952_1), .B(core__abc_21380_n1796), .Y(core__abc_21380_n7352) );
  OR2X2 OR2X2_2699 ( .A(core__abc_21380_n3951), .B(core_v1_reg_29_), .Y(core__abc_21380_n7353) );
  OR2X2 OR2X2_27 ( .A(_abc_19068_n957_1), .B(_abc_19068_n960_1), .Y(_abc_19068_n961_1) );
  OR2X2 OR2X2_270 ( .A(_abc_19068_n1477), .B(_abc_19068_n1478_1), .Y(_abc_19068_n1479) );
  OR2X2 OR2X2_2700 ( .A(core__abc_21380_n7356), .B(core__abc_21380_n7357), .Y(core__abc_21380_n7358) );
  OR2X2 OR2X2_2701 ( .A(core__abc_21380_n7359), .B(core__abc_21380_n7361), .Y(core__abc_21380_n7362) );
  OR2X2 OR2X2_2702 ( .A(core__abc_21380_n7365), .B(core__abc_21380_n7366), .Y(core__abc_21380_n7367) );
  OR2X2 OR2X2_2703 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n7367), .Y(core__abc_21380_n7368) );
  OR2X2 OR2X2_2704 ( .A(core__abc_21380_n7364), .B(core__abc_21380_n7368), .Y(core__abc_21380_n7369) );
  OR2X2 OR2X2_2705 ( .A(core__abc_21380_n7087_bF_buf5), .B(core_v2_reg_10_), .Y(core__abc_21380_n7370) );
  OR2X2 OR2X2_2706 ( .A(core__abc_21380_n7361), .B(core__abc_21380_n7356), .Y(core__abc_21380_n7373) );
  OR2X2 OR2X2_2707 ( .A(core__abc_21380_n7376), .B(core__abc_21380_n7375), .Y(core__abc_21380_n7377) );
  OR2X2 OR2X2_2708 ( .A(core__abc_21380_n7380), .B(core__abc_21380_n7378), .Y(core__abc_21380_n7381) );
  OR2X2 OR2X2_2709 ( .A(core__abc_21380_n7382), .B(core__abc_21380_n7384), .Y(core__abc_21380_n7385) );
  OR2X2 OR2X2_271 ( .A(_abc_19068_n1476_1), .B(_abc_19068_n1479), .Y(_abc_19068_n1480_1) );
  OR2X2 OR2X2_2710 ( .A(core__abc_21380_n7388), .B(core__abc_21380_n7389), .Y(core__abc_21380_n7390) );
  OR2X2 OR2X2_2711 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n7390), .Y(core__abc_21380_n7391) );
  OR2X2 OR2X2_2712 ( .A(core__abc_21380_n7387), .B(core__abc_21380_n7391), .Y(core__abc_21380_n7392) );
  OR2X2 OR2X2_2713 ( .A(core__abc_21380_n7087_bF_buf4), .B(core_v2_reg_11_), .Y(core__abc_21380_n7393) );
  OR2X2 OR2X2_2714 ( .A(core__abc_21380_n7398), .B(core__abc_21380_n7378), .Y(core__abc_21380_n7399) );
  OR2X2 OR2X2_2715 ( .A(core__abc_21380_n7399), .B(core__abc_21380_n7397), .Y(core__abc_21380_n7400) );
  OR2X2 OR2X2_2716 ( .A(core__abc_21380_n7402), .B(core__abc_21380_n7400), .Y(core__abc_21380_n7403) );
  OR2X2 OR2X2_2717 ( .A(core__abc_21380_n4099), .B(core__abc_21380_n1834), .Y(core__abc_21380_n7405) );
  OR2X2 OR2X2_2718 ( .A(core__abc_21380_n4098_1), .B(core_v1_reg_31_), .Y(core__abc_21380_n7406) );
  OR2X2 OR2X2_2719 ( .A(core__abc_21380_n7409), .B(core__abc_21380_n7410), .Y(core__abc_21380_n7411) );
  OR2X2 OR2X2_272 ( .A(_abc_19068_n1482_1), .B(_abc_19068_n1483), .Y(_abc_19068_n1484_1) );
  OR2X2 OR2X2_2720 ( .A(core__abc_21380_n7412), .B(core__abc_21380_n7414), .Y(core__abc_21380_n7415) );
  OR2X2 OR2X2_2721 ( .A(core__abc_21380_n7419), .B(core__abc_21380_n7420), .Y(core__abc_21380_n7421) );
  OR2X2 OR2X2_2722 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n7421), .Y(core__abc_21380_n7422) );
  OR2X2 OR2X2_2723 ( .A(core__abc_21380_n7417), .B(core__abc_21380_n7422), .Y(core__abc_21380_n7423) );
  OR2X2 OR2X2_2724 ( .A(core__abc_21380_n7087_bF_buf3), .B(core_v2_reg_12_), .Y(core__abc_21380_n7424) );
  OR2X2 OR2X2_2725 ( .A(core__abc_21380_n7427), .B(core__abc_21380_n7428), .Y(core__abc_21380_n7429) );
  OR2X2 OR2X2_2726 ( .A(core__abc_21380_n7429), .B(core__abc_21380_n3434), .Y(core__abc_21380_n7430) );
  OR2X2 OR2X2_2727 ( .A(core__abc_21380_n7437), .B(core__abc_21380_n7434), .Y(core__abc_21380_n7439) );
  OR2X2 OR2X2_2728 ( .A(core__abc_21380_n7440), .B(core__abc_21380_n7438), .Y(core__abc_21380_n7441) );
  OR2X2 OR2X2_2729 ( .A(core__abc_21380_n7445), .B(core__abc_21380_n7446), .Y(core__abc_21380_n7447) );
  OR2X2 OR2X2_273 ( .A(_abc_19068_n1484_1), .B(_abc_19068_n1481), .Y(_abc_19068_n1485) );
  OR2X2 OR2X2_2730 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n7447), .Y(core__abc_21380_n7448) );
  OR2X2 OR2X2_2731 ( .A(core__abc_21380_n7443), .B(core__abc_21380_n7448), .Y(core__abc_21380_n7449) );
  OR2X2 OR2X2_2732 ( .A(core__abc_21380_n7087_bF_buf2), .B(core_v2_reg_13_), .Y(core__abc_21380_n7450) );
  OR2X2 OR2X2_2733 ( .A(core__abc_21380_n7456), .B(core__abc_21380_n7455), .Y(core__abc_21380_n7457) );
  OR2X2 OR2X2_2734 ( .A(core__abc_21380_n7454), .B(core__abc_21380_n7457), .Y(core__abc_21380_n7458) );
  OR2X2 OR2X2_2735 ( .A(core__abc_21380_n4235), .B(core_v1_reg_33_), .Y(core__abc_21380_n7460) );
  OR2X2 OR2X2_2736 ( .A(core__abc_21380_n4234), .B(core__abc_21380_n1872), .Y(core__abc_21380_n7461) );
  OR2X2 OR2X2_2737 ( .A(core__abc_21380_n7464), .B(core__abc_21380_n7465), .Y(core__abc_21380_n7466) );
  OR2X2 OR2X2_2738 ( .A(core__abc_21380_n7467), .B(core__abc_21380_n7469), .Y(core__abc_21380_n7470) );
  OR2X2 OR2X2_2739 ( .A(core__abc_21380_n7474), .B(core__abc_21380_n7475), .Y(core__abc_21380_n7476) );
  OR2X2 OR2X2_274 ( .A(_abc_19068_n1486_1), .B(_abc_19068_n1487), .Y(_abc_19068_n1488_1) );
  OR2X2 OR2X2_2740 ( .A(core__abc_21380_n7076_bF_buf5), .B(core__abc_21380_n7476), .Y(core__abc_21380_n7477) );
  OR2X2 OR2X2_2741 ( .A(core__abc_21380_n7472), .B(core__abc_21380_n7477), .Y(core__abc_21380_n7478) );
  OR2X2 OR2X2_2742 ( .A(core__abc_21380_n7087_bF_buf1), .B(core_v2_reg_14_), .Y(core__abc_21380_n7479) );
  OR2X2 OR2X2_2743 ( .A(core__abc_21380_n7469), .B(core__abc_21380_n7465), .Y(core__abc_21380_n7482) );
  OR2X2 OR2X2_2744 ( .A(core__abc_21380_n7484), .B(core__abc_21380_n7485), .Y(core__abc_21380_n7486) );
  OR2X2 OR2X2_2745 ( .A(core__abc_21380_n7488), .B(core__abc_21380_n7489), .Y(core__abc_21380_n7490) );
  OR2X2 OR2X2_2746 ( .A(core__abc_21380_n7491), .B(core__abc_21380_n7493), .Y(core__abc_21380_n7494) );
  OR2X2 OR2X2_2747 ( .A(core__abc_21380_n7497), .B(core__abc_21380_n7498), .Y(core__abc_21380_n7499) );
  OR2X2 OR2X2_2748 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n7499), .Y(core__abc_21380_n7500) );
  OR2X2 OR2X2_2749 ( .A(core__abc_21380_n7496), .B(core__abc_21380_n7500), .Y(core__abc_21380_n7501) );
  OR2X2 OR2X2_275 ( .A(_abc_19068_n1489), .B(_abc_19068_n1490_1), .Y(_abc_19068_n1491) );
  OR2X2 OR2X2_2750 ( .A(core__abc_21380_n7087_bF_buf0), .B(core_v2_reg_15_), .Y(core__abc_21380_n7502) );
  OR2X2 OR2X2_2751 ( .A(core__abc_21380_n7510), .B(core__abc_21380_n7488), .Y(core__abc_21380_n7511) );
  OR2X2 OR2X2_2752 ( .A(core__abc_21380_n7508), .B(core__abc_21380_n7511), .Y(core__abc_21380_n7512) );
  OR2X2 OR2X2_2753 ( .A(core__abc_21380_n7512), .B(core__abc_21380_n7507), .Y(core__abc_21380_n7513) );
  OR2X2 OR2X2_2754 ( .A(core__abc_21380_n7515), .B(core__abc_21380_n7513), .Y(core__abc_21380_n7516) );
  OR2X2 OR2X2_2755 ( .A(core__abc_21380_n4392_1), .B(core__abc_21380_n1908), .Y(core__abc_21380_n7517) );
  OR2X2 OR2X2_2756 ( .A(core__abc_21380_n4391), .B(core_v1_reg_35_), .Y(core__abc_21380_n7518) );
  OR2X2 OR2X2_2757 ( .A(core__abc_21380_n7522), .B(core__abc_21380_n7520), .Y(core__abc_21380_n7523) );
  OR2X2 OR2X2_2758 ( .A(core__abc_21380_n7527), .B(core__abc_21380_n7292), .Y(core__abc_21380_n7528) );
  OR2X2 OR2X2_2759 ( .A(core__abc_21380_n7525), .B(core__abc_21380_n7534), .Y(core__abc_21380_n7535) );
  OR2X2 OR2X2_276 ( .A(_abc_19068_n1488_1), .B(_abc_19068_n1491), .Y(_abc_19068_n1492) );
  OR2X2 OR2X2_2760 ( .A(core__abc_21380_n7539), .B(core__abc_21380_n7540), .Y(core__abc_21380_n7541) );
  OR2X2 OR2X2_2761 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n7541), .Y(core__abc_21380_n7542) );
  OR2X2 OR2X2_2762 ( .A(core__abc_21380_n7537), .B(core__abc_21380_n7542), .Y(core__abc_21380_n7543) );
  OR2X2 OR2X2_2763 ( .A(core__abc_21380_n7087_bF_buf7), .B(core_v2_reg_16_), .Y(core__abc_21380_n7544) );
  OR2X2 OR2X2_2764 ( .A(core__abc_21380_n7551), .B(core__abc_21380_n7552), .Y(core__abc_21380_n7553) );
  OR2X2 OR2X2_2765 ( .A(core__abc_21380_n7550), .B(core__abc_21380_n7559), .Y(core__abc_21380_n7560) );
  OR2X2 OR2X2_2766 ( .A(core__abc_21380_n7549), .B(core__abc_21380_n7561), .Y(core__abc_21380_n7562) );
  OR2X2 OR2X2_2767 ( .A(core__abc_21380_n7565), .B(core__abc_21380_n7566), .Y(core__abc_21380_n7567) );
  OR2X2 OR2X2_2768 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n7567), .Y(core__abc_21380_n7568) );
  OR2X2 OR2X2_2769 ( .A(core__abc_21380_n7564), .B(core__abc_21380_n7568), .Y(core__abc_21380_n7569) );
  OR2X2 OR2X2_277 ( .A(_abc_19068_n1492), .B(_abc_19068_n1485), .Y(_abc_19068_n1493_1) );
  OR2X2 OR2X2_2770 ( .A(core__abc_21380_n7087_bF_buf6), .B(core_v2_reg_17_), .Y(core__abc_21380_n7570) );
  OR2X2 OR2X2_2771 ( .A(core__abc_21380_n7555), .B(core__abc_21380_n7522), .Y(core__abc_21380_n7573) );
  OR2X2 OR2X2_2772 ( .A(core__abc_21380_n7576), .B(core__abc_21380_n7574), .Y(core__abc_21380_n7577) );
  OR2X2 OR2X2_2773 ( .A(core__abc_21380_n4526), .B(core__abc_21380_n1948), .Y(core__abc_21380_n7579) );
  OR2X2 OR2X2_2774 ( .A(core__abc_21380_n4525), .B(core_v1_reg_37_), .Y(core__abc_21380_n7580) );
  OR2X2 OR2X2_2775 ( .A(core__abc_21380_n7582), .B(core__abc_21380_n7584), .Y(core__abc_21380_n7585) );
  OR2X2 OR2X2_2776 ( .A(core__abc_21380_n7586), .B(core__abc_21380_n7588), .Y(core__abc_21380_n7589) );
  OR2X2 OR2X2_2777 ( .A(core__abc_21380_n7593), .B(core__abc_21380_n7594), .Y(core__abc_21380_n7595) );
  OR2X2 OR2X2_2778 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n7595), .Y(core__abc_21380_n7596) );
  OR2X2 OR2X2_2779 ( .A(core__abc_21380_n7591), .B(core__abc_21380_n7596), .Y(core__abc_21380_n7597) );
  OR2X2 OR2X2_278 ( .A(_abc_19068_n1493_1), .B(_abc_19068_n1480_1), .Y(_abc_19068_n1494) );
  OR2X2 OR2X2_2780 ( .A(core__abc_21380_n7087_bF_buf5), .B(core_v2_reg_18_), .Y(core__abc_21380_n7598) );
  OR2X2 OR2X2_2781 ( .A(core__abc_21380_n7588), .B(core__abc_21380_n7584), .Y(core__abc_21380_n7601) );
  OR2X2 OR2X2_2782 ( .A(core__abc_21380_n7602), .B(core__abc_21380_n7603), .Y(core__abc_21380_n7604) );
  OR2X2 OR2X2_2783 ( .A(core__abc_21380_n3855), .B(core__abc_21380_n7605), .Y(core__abc_21380_n7608) );
  OR2X2 OR2X2_2784 ( .A(core__abc_21380_n7601), .B(core__abc_21380_n7609), .Y(core__abc_21380_n7610) );
  OR2X2 OR2X2_2785 ( .A(core__abc_21380_n7611), .B(core__abc_21380_n7612), .Y(core__abc_21380_n7613) );
  OR2X2 OR2X2_2786 ( .A(core__abc_21380_n7616), .B(core__abc_21380_n7617), .Y(core__abc_21380_n7618) );
  OR2X2 OR2X2_2787 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n7618), .Y(core__abc_21380_n7619) );
  OR2X2 OR2X2_2788 ( .A(core__abc_21380_n7615), .B(core__abc_21380_n7619), .Y(core__abc_21380_n7620) );
  OR2X2 OR2X2_2789 ( .A(core__abc_21380_n7087_bF_buf4), .B(core_v2_reg_19_), .Y(core__abc_21380_n7621) );
  OR2X2 OR2X2_279 ( .A(_abc_19068_n1496), .B(_abc_19068_n1497_1), .Y(_abc_19068_n1498) );
  OR2X2 OR2X2_2790 ( .A(core__abc_21380_n7606), .B(core__abc_21380_n7584), .Y(core__abc_21380_n7626) );
  OR2X2 OR2X2_2791 ( .A(core__abc_21380_n7625), .B(core__abc_21380_n7627), .Y(core__abc_21380_n7628) );
  OR2X2 OR2X2_2792 ( .A(core__abc_21380_n7533), .B(core__abc_21380_n7631), .Y(core__abc_21380_n7632) );
  OR2X2 OR2X2_2793 ( .A(core__abc_21380_n4644_1), .B(core__abc_21380_n1984), .Y(core__abc_21380_n7634) );
  OR2X2 OR2X2_2794 ( .A(core__abc_21380_n4643), .B(core_v1_reg_39_), .Y(core__abc_21380_n7635) );
  OR2X2 OR2X2_2795 ( .A(core__abc_21380_n7638), .B(core__abc_21380_n7639), .Y(core__abc_21380_n7640) );
  OR2X2 OR2X2_2796 ( .A(core__abc_21380_n7633), .B(core__abc_21380_n7640), .Y(core__abc_21380_n7642) );
  OR2X2 OR2X2_2797 ( .A(core__abc_21380_n7643), .B(core__abc_21380_n7641), .Y(core__abc_21380_n7644) );
  OR2X2 OR2X2_2798 ( .A(core__abc_21380_n7647), .B(core__abc_21380_n7648), .Y(core__abc_21380_n7649) );
  OR2X2 OR2X2_2799 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n7649), .Y(core__abc_21380_n7650) );
  OR2X2 OR2X2_28 ( .A(_abc_19068_n963_1), .B(_abc_19068_n964_1), .Y(_abc_19068_n965) );
  OR2X2 OR2X2_280 ( .A(_abc_19068_n1500), .B(_abc_19068_n1501_1), .Y(_abc_19068_n1502) );
  OR2X2 OR2X2_2800 ( .A(core__abc_21380_n7646), .B(core__abc_21380_n7650), .Y(core__abc_21380_n7651) );
  OR2X2 OR2X2_2801 ( .A(core__abc_21380_n7087_bF_buf3), .B(core_v2_reg_20_), .Y(core__abc_21380_n7652) );
  OR2X2 OR2X2_2802 ( .A(core__abc_21380_n7656), .B(core__abc_21380_n7655), .Y(core__abc_21380_n7657) );
  OR2X2 OR2X2_2803 ( .A(core__abc_21380_n7659), .B(core__abc_21380_n7660), .Y(core__abc_21380_n7661) );
  OR2X2 OR2X2_2804 ( .A(core__abc_21380_n7663), .B(core__abc_21380_n7661), .Y(core__abc_21380_n7666) );
  OR2X2 OR2X2_2805 ( .A(core__abc_21380_n7670), .B(core__abc_21380_n7671), .Y(core__abc_21380_n7672) );
  OR2X2 OR2X2_2806 ( .A(core__abc_21380_n7076_bF_buf5), .B(core__abc_21380_n7672), .Y(core__abc_21380_n7673) );
  OR2X2 OR2X2_2807 ( .A(core__abc_21380_n7668), .B(core__abc_21380_n7673), .Y(core__abc_21380_n7674) );
  OR2X2 OR2X2_2808 ( .A(core__abc_21380_n7087_bF_buf2), .B(core_v2_reg_21_), .Y(core__abc_21380_n7675) );
  OR2X2 OR2X2_2809 ( .A(core__abc_21380_n7680), .B(core__abc_21380_n7659), .Y(core__abc_21380_n7681) );
  OR2X2 OR2X2_281 ( .A(_abc_19068_n1502), .B(_abc_19068_n1499_1), .Y(_abc_19068_n1503_1) );
  OR2X2 OR2X2_2810 ( .A(core__abc_21380_n7679), .B(core__abc_21380_n7681), .Y(core__abc_21380_n7682) );
  OR2X2 OR2X2_2811 ( .A(core__abc_21380_n4765), .B(core__abc_21380_n2023), .Y(core__abc_21380_n7684) );
  OR2X2 OR2X2_2812 ( .A(core__abc_21380_n4764), .B(core_v1_reg_41_), .Y(core__abc_21380_n7685) );
  OR2X2 OR2X2_2813 ( .A(core__abc_21380_n7688), .B(core__abc_21380_n7689), .Y(core__abc_21380_n7690) );
  OR2X2 OR2X2_2814 ( .A(core__abc_21380_n7691), .B(core__abc_21380_n7693), .Y(core__abc_21380_n7694) );
  OR2X2 OR2X2_2815 ( .A(core__abc_21380_n7698), .B(core__abc_21380_n7699), .Y(core__abc_21380_n7700) );
  OR2X2 OR2X2_2816 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n7700), .Y(core__abc_21380_n7701) );
  OR2X2 OR2X2_2817 ( .A(core__abc_21380_n7696), .B(core__abc_21380_n7701), .Y(core__abc_21380_n7702) );
  OR2X2 OR2X2_2818 ( .A(core__abc_21380_n7087_bF_buf1), .B(core_v2_reg_22_), .Y(core__abc_21380_n7703) );
  OR2X2 OR2X2_2819 ( .A(core__abc_21380_n7693), .B(core__abc_21380_n7688), .Y(core__abc_21380_n7706) );
  OR2X2 OR2X2_282 ( .A(_abc_19068_n1503_1), .B(_abc_19068_n1498), .Y(_abc_19068_n1504) );
  OR2X2 OR2X2_2820 ( .A(core__abc_21380_n7708), .B(core__abc_21380_n7707), .Y(core__abc_21380_n7709) );
  OR2X2 OR2X2_2821 ( .A(core__abc_21380_n7706), .B(core__abc_21380_n7716), .Y(core__abc_21380_n7717) );
  OR2X2 OR2X2_2822 ( .A(core__abc_21380_n7718), .B(core__abc_21380_n7715), .Y(core__abc_21380_n7719) );
  OR2X2 OR2X2_2823 ( .A(core__abc_21380_n7723), .B(core__abc_21380_n7724), .Y(core__abc_21380_n7725) );
  OR2X2 OR2X2_2824 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n7725), .Y(core__abc_21380_n7726) );
  OR2X2 OR2X2_2825 ( .A(core__abc_21380_n7722), .B(core__abc_21380_n7726), .Y(core__abc_21380_n7727) );
  OR2X2 OR2X2_2826 ( .A(core__abc_21380_n7087_bF_buf0), .B(core_v2_reg_23_), .Y(core__abc_21380_n7728) );
  OR2X2 OR2X2_2827 ( .A(core__abc_21380_n7661), .B(core__abc_21380_n7640), .Y(core__abc_21380_n7731) );
  OR2X2 OR2X2_2828 ( .A(core__abc_21380_n7733), .B(core__abc_21380_n7731), .Y(core__abc_21380_n7734) );
  OR2X2 OR2X2_2829 ( .A(core__abc_21380_n7737), .B(core__abc_21380_n7533), .Y(core__abc_21380_n7738) );
  OR2X2 OR2X2_283 ( .A(_abc_19068_n1506), .B(_abc_19068_n1507_1), .Y(_abc_19068_n1508) );
  OR2X2 OR2X2_2830 ( .A(core__abc_21380_n7741), .B(core__abc_21380_n7711), .Y(core__abc_21380_n7742) );
  OR2X2 OR2X2_2831 ( .A(core__abc_21380_n7740), .B(core__abc_21380_n7742), .Y(core__abc_21380_n7743) );
  OR2X2 OR2X2_2832 ( .A(core__abc_21380_n7739), .B(core__abc_21380_n7743), .Y(core__abc_21380_n7744) );
  OR2X2 OR2X2_2833 ( .A(core__abc_21380_n4886), .B(core__abc_21380_n2058), .Y(core__abc_21380_n7747) );
  OR2X2 OR2X2_2834 ( .A(core__abc_21380_n4885), .B(core_v1_reg_43_), .Y(core__abc_21380_n7748) );
  OR2X2 OR2X2_2835 ( .A(core__abc_21380_n7752), .B(core__abc_21380_n7750), .Y(core__abc_21380_n7753) );
  OR2X2 OR2X2_2836 ( .A(core__abc_21380_n7746), .B(core__abc_21380_n7753), .Y(core__abc_21380_n7755) );
  OR2X2 OR2X2_2837 ( .A(core__abc_21380_n7756), .B(core__abc_21380_n7754), .Y(core__abc_21380_n7757) );
  OR2X2 OR2X2_2838 ( .A(core__abc_21380_n7760), .B(core__abc_21380_n7761), .Y(core__abc_21380_n7762) );
  OR2X2 OR2X2_2839 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n7762), .Y(core__abc_21380_n7763) );
  OR2X2 OR2X2_284 ( .A(_abc_19068_n1509_1), .B(_abc_19068_n1510), .Y(_abc_19068_n1511_1) );
  OR2X2 OR2X2_2840 ( .A(core__abc_21380_n7759), .B(core__abc_21380_n7763), .Y(core__abc_21380_n7764) );
  OR2X2 OR2X2_2841 ( .A(core__abc_21380_n7087_bF_buf7), .B(core_v2_reg_24_), .Y(core__abc_21380_n7765) );
  OR2X2 OR2X2_2842 ( .A(core__abc_21380_n4936), .B(core__abc_21380_n2079), .Y(core__abc_21380_n7772) );
  OR2X2 OR2X2_2843 ( .A(core__abc_21380_n7769), .B(core__abc_21380_n7779), .Y(core__abc_21380_n7780) );
  OR2X2 OR2X2_2844 ( .A(core__abc_21380_n7781), .B(core__abc_21380_n7782), .Y(core__abc_21380_n7783) );
  OR2X2 OR2X2_2845 ( .A(core__abc_21380_n7788), .B(core__abc_21380_n7789), .Y(core__abc_21380_n7790) );
  OR2X2 OR2X2_2846 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n7790), .Y(core__abc_21380_n7791) );
  OR2X2 OR2X2_2847 ( .A(core__abc_21380_n7786), .B(core__abc_21380_n7791), .Y(core__abc_21380_n7792) );
  OR2X2 OR2X2_2848 ( .A(core__abc_21380_n7087_bF_buf6), .B(core_v2_reg_25_), .Y(core__abc_21380_n7793) );
  OR2X2 OR2X2_2849 ( .A(core__abc_21380_n4979), .B(core__abc_21380_n2096), .Y(core__abc_21380_n7796) );
  OR2X2 OR2X2_285 ( .A(_abc_19068_n1508), .B(_abc_19068_n1511_1), .Y(_abc_19068_n1512) );
  OR2X2 OR2X2_2850 ( .A(core__abc_21380_n4978), .B(core_v1_reg_45_), .Y(core__abc_21380_n7797) );
  OR2X2 OR2X2_2851 ( .A(core__abc_21380_n7799), .B(core__abc_21380_n7801), .Y(core__abc_21380_n7802) );
  OR2X2 OR2X2_2852 ( .A(core__abc_21380_n7782), .B(core__abc_21380_n7753), .Y(core__abc_21380_n7803) );
  OR2X2 OR2X2_2853 ( .A(core__abc_21380_n7746), .B(core__abc_21380_n7803), .Y(core__abc_21380_n7804) );
  OR2X2 OR2X2_2854 ( .A(core__abc_21380_n7805), .B(core__abc_21380_n7777), .Y(core__abc_21380_n7806) );
  OR2X2 OR2X2_2855 ( .A(core__abc_21380_n7807), .B(core__abc_21380_n7802), .Y(core__abc_21380_n7809) );
  OR2X2 OR2X2_2856 ( .A(core__abc_21380_n7810), .B(core__abc_21380_n7808), .Y(core__abc_21380_n7811) );
  OR2X2 OR2X2_2857 ( .A(core__abc_21380_n7815), .B(core__abc_21380_n7816), .Y(core__abc_21380_n7817) );
  OR2X2 OR2X2_2858 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n7817), .Y(core__abc_21380_n7818) );
  OR2X2 OR2X2_2859 ( .A(core__abc_21380_n7813), .B(core__abc_21380_n7818), .Y(core__abc_21380_n7819) );
  OR2X2 OR2X2_286 ( .A(_abc_19068_n1512), .B(_abc_19068_n1505_1), .Y(_abc_19068_n1513_1) );
  OR2X2 OR2X2_2860 ( .A(core__abc_21380_n7087_bF_buf5), .B(core_v2_reg_26_), .Y(core__abc_21380_n7820) );
  OR2X2 OR2X2_2861 ( .A(core__abc_21380_n7826), .B(core__abc_21380_n7825), .Y(core__abc_21380_n7827) );
  OR2X2 OR2X2_2862 ( .A(core__abc_21380_n7838), .B(core__abc_21380_n7836), .Y(core__abc_21380_n7839) );
  OR2X2 OR2X2_2863 ( .A(core__abc_21380_n7843), .B(core__abc_21380_n7844), .Y(core__abc_21380_n7845) );
  OR2X2 OR2X2_2864 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n7845), .Y(core__abc_21380_n7846) );
  OR2X2 OR2X2_2865 ( .A(core__abc_21380_n7841), .B(core__abc_21380_n7846), .Y(core__abc_21380_n7847) );
  OR2X2 OR2X2_2866 ( .A(core__abc_21380_n7087_bF_buf4), .B(core_v2_reg_27_), .Y(core__abc_21380_n7848) );
  OR2X2 OR2X2_2867 ( .A(core__abc_21380_n7851), .B(core__abc_21380_n7744), .Y(core__abc_21380_n7852) );
  OR2X2 OR2X2_2868 ( .A(core__abc_21380_n7835), .B(core__abc_21380_n7802), .Y(core__abc_21380_n7853) );
  OR2X2 OR2X2_2869 ( .A(core__abc_21380_n7853), .B(core__abc_21380_n7803), .Y(core__abc_21380_n7854) );
  OR2X2 OR2X2_287 ( .A(_abc_19068_n1513_1), .B(_abc_19068_n1504), .Y(_abc_19068_n1514) );
  OR2X2 OR2X2_2870 ( .A(core__abc_21380_n7853), .B(core__abc_21380_n7806), .Y(core__abc_21380_n7857) );
  OR2X2 OR2X2_2871 ( .A(core__abc_21380_n7858), .B(core__abc_21380_n7829), .Y(core__abc_21380_n7859) );
  OR2X2 OR2X2_2872 ( .A(core__abc_21380_n7856), .B(core__abc_21380_n7862), .Y(core__abc_21380_n7863) );
  OR2X2 OR2X2_2873 ( .A(core__abc_21380_n5099), .B(core__abc_21380_n2136), .Y(core__abc_21380_n7864) );
  OR2X2 OR2X2_2874 ( .A(core__abc_21380_n5098), .B(core_v1_reg_47_), .Y(core__abc_21380_n7865) );
  OR2X2 OR2X2_2875 ( .A(core__abc_21380_n7869), .B(core__abc_21380_n7867), .Y(core__abc_21380_n7870) );
  OR2X2 OR2X2_2876 ( .A(core__abc_21380_n7746), .B(core__abc_21380_n7854), .Y(core__abc_21380_n7873) );
  OR2X2 OR2X2_2877 ( .A(core__abc_21380_n7872), .B(core__abc_21380_n7875), .Y(core__abc_21380_n7876) );
  OR2X2 OR2X2_2878 ( .A(core__abc_21380_n7879), .B(core__abc_21380_n7880), .Y(core__abc_21380_n7881) );
  OR2X2 OR2X2_2879 ( .A(core__abc_21380_n7076_bF_buf5), .B(core__abc_21380_n7881), .Y(core__abc_21380_n7882) );
  OR2X2 OR2X2_288 ( .A(_abc_19068_n1516), .B(_abc_19068_n1517_1), .Y(_abc_19068_n1518) );
  OR2X2 OR2X2_2880 ( .A(core__abc_21380_n7878), .B(core__abc_21380_n7882), .Y(core__abc_21380_n7883) );
  OR2X2 OR2X2_2881 ( .A(core__abc_21380_n7087_bF_buf3), .B(core_v2_reg_28_), .Y(core__abc_21380_n7884) );
  OR2X2 OR2X2_2882 ( .A(core__abc_21380_n7872), .B(core__abc_21380_n7869), .Y(core__abc_21380_n7887) );
  OR2X2 OR2X2_2883 ( .A(core__abc_21380_n7889), .B(core__abc_21380_n7890), .Y(core__abc_21380_n7891) );
  OR2X2 OR2X2_2884 ( .A(core__abc_21380_n7892), .B(core__abc_21380_n7894), .Y(core__abc_21380_n7895) );
  OR2X2 OR2X2_2885 ( .A(core__abc_21380_n7887), .B(core__abc_21380_n7895), .Y(core__abc_21380_n7896) );
  OR2X2 OR2X2_2886 ( .A(core__abc_21380_n7897), .B(core__abc_21380_n7898), .Y(core__abc_21380_n7899) );
  OR2X2 OR2X2_2887 ( .A(core__abc_21380_n7904), .B(core__abc_21380_n7905), .Y(core__abc_21380_n7906) );
  OR2X2 OR2X2_2888 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n7906), .Y(core__abc_21380_n7907) );
  OR2X2 OR2X2_2889 ( .A(core__abc_21380_n7902), .B(core__abc_21380_n7907), .Y(core__abc_21380_n7908) );
  OR2X2 OR2X2_289 ( .A(_abc_19068_n1520), .B(_abc_19068_n1521_1), .Y(_abc_19068_n1522) );
  OR2X2 OR2X2_2890 ( .A(core__abc_21380_n7087_bF_buf2), .B(core_v2_reg_29_), .Y(core__abc_21380_n7909) );
  OR2X2 OR2X2_2891 ( .A(core__abc_21380_n7874), .B(core__abc_21380_n7913), .Y(core__abc_21380_n7914) );
  OR2X2 OR2X2_2892 ( .A(core__abc_21380_n7915), .B(core__abc_21380_n7894), .Y(core__abc_21380_n7916) );
  OR2X2 OR2X2_2893 ( .A(core__abc_21380_n5207), .B(core__abc_21380_n2173), .Y(core__abc_21380_n7919) );
  OR2X2 OR2X2_2894 ( .A(core__abc_21380_n5206), .B(core_v1_reg_49_), .Y(core__abc_21380_n7920) );
  OR2X2 OR2X2_2895 ( .A(core__abc_21380_n7923), .B(core__abc_21380_n7924), .Y(core__abc_21380_n7925) );
  OR2X2 OR2X2_2896 ( .A(core__abc_21380_n7927), .B(core__abc_21380_n7916), .Y(core__abc_21380_n7928) );
  OR2X2 OR2X2_2897 ( .A(core__abc_21380_n7930), .B(core__abc_21380_n7926), .Y(core__abc_21380_n7931) );
  OR2X2 OR2X2_2898 ( .A(core__abc_21380_n7935), .B(core__abc_21380_n7936), .Y(core__abc_21380_n7937) );
  OR2X2 OR2X2_2899 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n7937), .Y(core__abc_21380_n7938) );
  OR2X2 OR2X2_29 ( .A(_abc_19068_n965), .B(_abc_19068_n962), .Y(_abc_19068_n966_1) );
  OR2X2 OR2X2_290 ( .A(_abc_19068_n1522), .B(_abc_19068_n1519_1), .Y(_abc_19068_n1523_1) );
  OR2X2 OR2X2_2900 ( .A(core__abc_21380_n7933), .B(core__abc_21380_n7938), .Y(core__abc_21380_n7939) );
  OR2X2 OR2X2_2901 ( .A(core__abc_21380_n7087_bF_buf1), .B(core_v2_reg_30_), .Y(core__abc_21380_n7940) );
  OR2X2 OR2X2_2902 ( .A(core__abc_21380_n7918), .B(core__abc_21380_n7925), .Y(core__abc_21380_n7944) );
  OR2X2 OR2X2_2903 ( .A(core__abc_21380_n7946), .B(core__abc_21380_n7947), .Y(core__abc_21380_n7948) );
  OR2X2 OR2X2_2904 ( .A(core__abc_21380_n4682), .B(core__abc_21380_n7949), .Y(core__abc_21380_n7950) );
  OR2X2 OR2X2_2905 ( .A(core__abc_21380_n4680), .B(core__abc_21380_n7948), .Y(core__abc_21380_n7951) );
  OR2X2 OR2X2_2906 ( .A(core__abc_21380_n7945), .B(core__abc_21380_n7953), .Y(core__abc_21380_n7956) );
  OR2X2 OR2X2_2907 ( .A(core__abc_21380_n7959), .B(core__abc_21380_n7960), .Y(core__abc_21380_n7961) );
  OR2X2 OR2X2_2908 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n7961), .Y(core__abc_21380_n7962) );
  OR2X2 OR2X2_2909 ( .A(core__abc_21380_n7958), .B(core__abc_21380_n7962), .Y(core__abc_21380_n7963) );
  OR2X2 OR2X2_291 ( .A(_abc_19068_n1523_1), .B(_abc_19068_n1518), .Y(_abc_19068_n1524) );
  OR2X2 OR2X2_2910 ( .A(core__abc_21380_n7087_bF_buf0), .B(core_v2_reg_31_), .Y(core__abc_21380_n7964) );
  OR2X2 OR2X2_2911 ( .A(core__abc_21380_n7970), .B(core__abc_21380_n7013), .Y(core__abc_21380_n7971) );
  OR2X2 OR2X2_2912 ( .A(core__abc_21380_n7973), .B(core__abc_21380_n7968), .Y(core__abc_21380_n7974) );
  OR2X2 OR2X2_2913 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n3163_1_bF_buf1), .Y(core__abc_21380_n7976) );
  OR2X2 OR2X2_2914 ( .A(core__abc_21380_n7977), .B(core__abc_21380_n7975), .Y(core__abc_21380_n7978) );
  OR2X2 OR2X2_2915 ( .A(core__abc_21380_n7017), .B(core__abc_21380_n7013), .Y(core__abc_21380_n7981) );
  OR2X2 OR2X2_2916 ( .A(core__abc_21380_n7983), .B(core__abc_21380_n7984), .Y(core__abc_21380_n7985) );
  OR2X2 OR2X2_2917 ( .A(core__abc_21380_n7986), .B(core__abc_21380_n7987), .Y(core__abc_21380_n7988) );
  OR2X2 OR2X2_2918 ( .A(core__abc_21380_n7019), .B(core__abc_21380_n7023), .Y(core__abc_21380_n7992) );
  OR2X2 OR2X2_2919 ( .A(core__abc_21380_n7994), .B(core__abc_21380_n7996), .Y(core__abc_21380_n7997) );
  OR2X2 OR2X2_292 ( .A(_abc_19068_n1526), .B(_abc_19068_n1527_1), .Y(_abc_19068_n1528) );
  OR2X2 OR2X2_2920 ( .A(core__abc_21380_n7998), .B(core__abc_21380_n7990), .Y(core__abc_21380_n7999) );
  OR2X2 OR2X2_2921 ( .A(core__abc_21380_n7025), .B(core__abc_21380_n6998), .Y(core__abc_21380_n8002) );
  OR2X2 OR2X2_2922 ( .A(core__abc_21380_n8005), .B(core__abc_21380_n8006), .Y(core__abc_21380_n8007) );
  OR2X2 OR2X2_2923 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n8007), .Y(core__abc_21380_n8008) );
  OR2X2 OR2X2_2924 ( .A(core__abc_21380_n8004), .B(core__abc_21380_n8008), .Y(core__abc_21380_n8009) );
  OR2X2 OR2X2_2925 ( .A(core__abc_21380_n7087_bF_buf4), .B(core_v2_reg_35_), .Y(core__abc_21380_n8010) );
  OR2X2 OR2X2_2926 ( .A(core__abc_21380_n7027), .B(core__abc_21380_n7030), .Y(core__abc_21380_n8014) );
  OR2X2 OR2X2_2927 ( .A(core__abc_21380_n8017), .B(core__abc_21380_n8018), .Y(core__abc_21380_n8019) );
  OR2X2 OR2X2_2928 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n8019), .Y(core__abc_21380_n8020) );
  OR2X2 OR2X2_2929 ( .A(core__abc_21380_n8016), .B(core__abc_21380_n8020), .Y(core__abc_21380_n8021) );
  OR2X2 OR2X2_293 ( .A(_abc_19068_n1529_1), .B(_abc_19068_n1530), .Y(_abc_19068_n1531_1) );
  OR2X2 OR2X2_2930 ( .A(core__abc_21380_n7087_bF_buf3), .B(core_v2_reg_36_), .Y(core__abc_21380_n8022) );
  OR2X2 OR2X2_2931 ( .A(core__abc_21380_n7032), .B(core__abc_21380_n6985), .Y(core__abc_21380_n8026) );
  OR2X2 OR2X2_2932 ( .A(core__abc_21380_n8030), .B(core__abc_21380_n8031), .Y(core__abc_21380_n8032) );
  OR2X2 OR2X2_2933 ( .A(core__abc_21380_n7076_bF_buf5), .B(core__abc_21380_n8032), .Y(core__abc_21380_n8033) );
  OR2X2 OR2X2_2934 ( .A(core__abc_21380_n8028), .B(core__abc_21380_n8033), .Y(core__abc_21380_n8034) );
  OR2X2 OR2X2_2935 ( .A(core__abc_21380_n7087_bF_buf2), .B(core_v2_reg_37_), .Y(core__abc_21380_n8035) );
  OR2X2 OR2X2_2936 ( .A(core__abc_21380_n7034), .B(core__abc_21380_n6976), .Y(core__abc_21380_n8040) );
  OR2X2 OR2X2_2937 ( .A(core__abc_21380_n8044), .B(core__abc_21380_n8045), .Y(core__abc_21380_n8046) );
  OR2X2 OR2X2_2938 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n8046), .Y(core__abc_21380_n8047) );
  OR2X2 OR2X2_2939 ( .A(core__abc_21380_n8042), .B(core__abc_21380_n8047), .Y(core__abc_21380_n8048) );
  OR2X2 OR2X2_294 ( .A(_abc_19068_n1528), .B(_abc_19068_n1531_1), .Y(_abc_19068_n1532) );
  OR2X2 OR2X2_2940 ( .A(core__abc_21380_n7087_bF_buf1), .B(core_v2_reg_38_), .Y(core__abc_21380_n8049) );
  OR2X2 OR2X2_2941 ( .A(core__abc_21380_n8038), .B(core__abc_21380_n6969), .Y(core__abc_21380_n8052) );
  OR2X2 OR2X2_2942 ( .A(core__abc_21380_n8052), .B(core__abc_21380_n6973), .Y(core__abc_21380_n8053) );
  OR2X2 OR2X2_2943 ( .A(core__abc_21380_n8055), .B(core__abc_21380_n8054), .Y(core__abc_21380_n8056) );
  OR2X2 OR2X2_2944 ( .A(core__abc_21380_n8059), .B(core__abc_21380_n8060), .Y(core__abc_21380_n8061) );
  OR2X2 OR2X2_2945 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n8061), .Y(core__abc_21380_n8062) );
  OR2X2 OR2X2_2946 ( .A(core__abc_21380_n8058), .B(core__abc_21380_n8062), .Y(core__abc_21380_n8063) );
  OR2X2 OR2X2_2947 ( .A(core__abc_21380_n7087_bF_buf0), .B(core_v2_reg_39_), .Y(core__abc_21380_n8064) );
  OR2X2 OR2X2_2948 ( .A(core__abc_21380_n8068), .B(core__abc_21380_n8069), .Y(core__abc_21380_n8070) );
  OR2X2 OR2X2_2949 ( .A(core__abc_21380_n8074), .B(core__abc_21380_n8075), .Y(core__abc_21380_n8076) );
  OR2X2 OR2X2_295 ( .A(_abc_19068_n1532), .B(_abc_19068_n1525_1), .Y(_abc_19068_n1533_1) );
  OR2X2 OR2X2_2950 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n8076), .Y(core__abc_21380_n8077) );
  OR2X2 OR2X2_2951 ( .A(core__abc_21380_n8072), .B(core__abc_21380_n8077), .Y(core__abc_21380_n8078) );
  OR2X2 OR2X2_2952 ( .A(core__abc_21380_n7087_bF_buf7), .B(core_v2_reg_40_), .Y(core__abc_21380_n8079) );
  OR2X2 OR2X2_2953 ( .A(core__abc_21380_n8069), .B(core__abc_21380_n6945), .Y(core__abc_21380_n8083) );
  OR2X2 OR2X2_2954 ( .A(core__abc_21380_n8085), .B(core__abc_21380_n8086), .Y(core__abc_21380_n8087) );
  OR2X2 OR2X2_2955 ( .A(core__abc_21380_n8091), .B(core__abc_21380_n8092), .Y(core__abc_21380_n8093) );
  OR2X2 OR2X2_2956 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n8093), .Y(core__abc_21380_n8094) );
  OR2X2 OR2X2_2957 ( .A(core__abc_21380_n8089), .B(core__abc_21380_n8094), .Y(core__abc_21380_n8095) );
  OR2X2 OR2X2_2958 ( .A(core__abc_21380_n7087_bF_buf6), .B(core_v2_reg_41_), .Y(core__abc_21380_n8096) );
  OR2X2 OR2X2_2959 ( .A(core__abc_21380_n8099), .B(core__abc_21380_n6949), .Y(core__abc_21380_n8100) );
  OR2X2 OR2X2_296 ( .A(_abc_19068_n1533_1), .B(_abc_19068_n1524), .Y(_abc_19068_n1534) );
  OR2X2 OR2X2_2960 ( .A(core__abc_21380_n8100), .B(core__abc_21380_n6954), .Y(core__abc_21380_n8103) );
  OR2X2 OR2X2_2961 ( .A(core__abc_21380_n8107), .B(core__abc_21380_n8108), .Y(core__abc_21380_n8109) );
  OR2X2 OR2X2_2962 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n8109), .Y(core__abc_21380_n8110) );
  OR2X2 OR2X2_2963 ( .A(core__abc_21380_n8105), .B(core__abc_21380_n8110), .Y(core__abc_21380_n8111) );
  OR2X2 OR2X2_2964 ( .A(core__abc_21380_n7087_bF_buf5), .B(core_v2_reg_42_), .Y(core__abc_21380_n8112) );
  OR2X2 OR2X2_2965 ( .A(core__abc_21380_n8116), .B(core__abc_21380_n8115), .Y(core__abc_21380_n8119) );
  OR2X2 OR2X2_2966 ( .A(core__abc_21380_n8122), .B(core__abc_21380_n8123), .Y(core__abc_21380_n8124) );
  OR2X2 OR2X2_2967 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n8124), .Y(core__abc_21380_n8125) );
  OR2X2 OR2X2_2968 ( .A(core__abc_21380_n8121), .B(core__abc_21380_n8125), .Y(core__abc_21380_n8126) );
  OR2X2 OR2X2_2969 ( .A(core__abc_21380_n7087_bF_buf4), .B(core_v2_reg_43_), .Y(core__abc_21380_n8127) );
  OR2X2 OR2X2_297 ( .A(_abc_19068_n1209_1), .B(_abc_19068_n1536), .Y(_abc_19068_n1537_1) );
  OR2X2 OR2X2_2970 ( .A(core__abc_21380_n8132), .B(core__abc_21380_n8130), .Y(core__abc_21380_n8133) );
  OR2X2 OR2X2_2971 ( .A(core__abc_21380_n8136), .B(core__abc_21380_n8137), .Y(core__abc_21380_n8138) );
  OR2X2 OR2X2_2972 ( .A(core__abc_21380_n7076_bF_buf5), .B(core__abc_21380_n8138), .Y(core__abc_21380_n8139) );
  OR2X2 OR2X2_2973 ( .A(core__abc_21380_n8135), .B(core__abc_21380_n8139), .Y(core__abc_21380_n8140) );
  OR2X2 OR2X2_2974 ( .A(core__abc_21380_n7087_bF_buf3), .B(core_v2_reg_44_), .Y(core__abc_21380_n8141) );
  OR2X2 OR2X2_2975 ( .A(core__abc_21380_n8130), .B(core__abc_21380_n6903), .Y(core__abc_21380_n8145) );
  OR2X2 OR2X2_2976 ( .A(core__abc_21380_n8145), .B(core__abc_21380_n8144), .Y(core__abc_21380_n8148) );
  OR2X2 OR2X2_2977 ( .A(core__abc_21380_n8153), .B(core__abc_21380_n8154), .Y(core__abc_21380_n8155) );
  OR2X2 OR2X2_2978 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n8155), .Y(core__abc_21380_n8156) );
  OR2X2 OR2X2_2979 ( .A(core__abc_21380_n8151), .B(core__abc_21380_n8156), .Y(core__abc_21380_n8157) );
  OR2X2 OR2X2_298 ( .A(_abc_19068_n1538), .B(_abc_19068_n1539_1), .Y(_abc_19068_n1540) );
  OR2X2 OR2X2_2980 ( .A(core__abc_21380_n7087_bF_buf2), .B(core_v2_reg_45_), .Y(core__abc_21380_n8158) );
  OR2X2 OR2X2_2981 ( .A(core__abc_21380_n8161), .B(core__abc_21380_n6907), .Y(core__abc_21380_n8162) );
  OR2X2 OR2X2_2982 ( .A(core__abc_21380_n8162), .B(core__abc_21380_n6889), .Y(core__abc_21380_n8165) );
  OR2X2 OR2X2_2983 ( .A(core__abc_21380_n8169), .B(core__abc_21380_n8170), .Y(core__abc_21380_n8171) );
  OR2X2 OR2X2_2984 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n8171), .Y(core__abc_21380_n8172) );
  OR2X2 OR2X2_2985 ( .A(core__abc_21380_n8167), .B(core__abc_21380_n8172), .Y(core__abc_21380_n8173) );
  OR2X2 OR2X2_2986 ( .A(core__abc_21380_n7087_bF_buf1), .B(core_v2_reg_46_), .Y(core__abc_21380_n8174) );
  OR2X2 OR2X2_2987 ( .A(core__abc_21380_n8163), .B(core__abc_21380_n6886), .Y(core__abc_21380_n8178) );
  OR2X2 OR2X2_2988 ( .A(core__abc_21380_n8180), .B(core__abc_21380_n8181), .Y(core__abc_21380_n8182) );
  OR2X2 OR2X2_2989 ( .A(core__abc_21380_n8185), .B(core__abc_21380_n8186), .Y(core__abc_21380_n8187) );
  OR2X2 OR2X2_299 ( .A(_abc_19068_n1537_1), .B(_abc_19068_n1540), .Y(_abc_19068_n1541_1) );
  OR2X2 OR2X2_2990 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n8187), .Y(core__abc_21380_n8188) );
  OR2X2 OR2X2_2991 ( .A(core__abc_21380_n8184), .B(core__abc_21380_n8188), .Y(core__abc_21380_n8189) );
  OR2X2 OR2X2_2992 ( .A(core__abc_21380_n7087_bF_buf0), .B(core_v2_reg_47_), .Y(core__abc_21380_n8190) );
  OR2X2 OR2X2_2993 ( .A(core__abc_21380_n8194), .B(core__abc_21380_n8195), .Y(core__abc_21380_n8196) );
  OR2X2 OR2X2_2994 ( .A(core__abc_21380_n8200), .B(core__abc_21380_n8201), .Y(core__abc_21380_n8202) );
  OR2X2 OR2X2_2995 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n8202), .Y(core__abc_21380_n8203) );
  OR2X2 OR2X2_2996 ( .A(core__abc_21380_n8198), .B(core__abc_21380_n8203), .Y(core__abc_21380_n8204) );
  OR2X2 OR2X2_2997 ( .A(core__abc_21380_n7087_bF_buf7), .B(core_v2_reg_48_), .Y(core__abc_21380_n8205) );
  OR2X2 OR2X2_2998 ( .A(core__abc_21380_n8195), .B(core__abc_21380_n6850), .Y(core__abc_21380_n8209) );
  OR2X2 OR2X2_2999 ( .A(core__abc_21380_n8212), .B(core__abc_21380_n8210), .Y(core__abc_21380_n8213) );
  OR2X2 OR2X2_3 ( .A(_abc_19068_n899_bF_buf4), .B(_abc_19068_n902_bF_buf4), .Y(_abc_19068_n903_1) );
  OR2X2 OR2X2_30 ( .A(_abc_19068_n961_1), .B(_abc_19068_n966_1), .Y(_abc_19068_n967_1) );
  OR2X2 OR2X2_300 ( .A(_abc_19068_n1543_1), .B(_abc_19068_n1544), .Y(_abc_19068_n1545_1) );
  OR2X2 OR2X2_3000 ( .A(core__abc_21380_n8215), .B(core__abc_21380_n8216), .Y(core__abc_21380_n8217) );
  OR2X2 OR2X2_3001 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n8217), .Y(core__abc_21380_n8218) );
  OR2X2 OR2X2_3002 ( .A(core__abc_21380_n8214), .B(core__abc_21380_n8218), .Y(core__abc_21380_n8219) );
  OR2X2 OR2X2_3003 ( .A(core__abc_21380_n7087_bF_buf6), .B(core_v2_reg_49_), .Y(core__abc_21380_n8220) );
  OR2X2 OR2X2_3004 ( .A(core__abc_21380_n8223), .B(core__abc_21380_n6851), .Y(core__abc_21380_n8224) );
  OR2X2 OR2X2_3005 ( .A(core__abc_21380_n8226), .B(core__abc_21380_n8227), .Y(core__abc_21380_n8228) );
  OR2X2 OR2X2_3006 ( .A(core__abc_21380_n8231), .B(core__abc_21380_n8232), .Y(core__abc_21380_n8233) );
  OR2X2 OR2X2_3007 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n8233), .Y(core__abc_21380_n8234) );
  OR2X2 OR2X2_3008 ( .A(core__abc_21380_n8230), .B(core__abc_21380_n8234), .Y(core__abc_21380_n8235) );
  OR2X2 OR2X2_3009 ( .A(core__abc_21380_n7087_bF_buf5), .B(core_v2_reg_50_), .Y(core__abc_21380_n8236) );
  OR2X2 OR2X2_301 ( .A(_abc_19068_n1545_1), .B(_abc_19068_n1542), .Y(_abc_19068_n1546) );
  OR2X2 OR2X2_3010 ( .A(core__abc_21380_n8226), .B(core__abc_21380_n6835), .Y(core__abc_21380_n8240) );
  OR2X2 OR2X2_3011 ( .A(core__abc_21380_n8242), .B(core__abc_21380_n8243), .Y(core__abc_21380_n8244) );
  OR2X2 OR2X2_3012 ( .A(core__abc_21380_n8248), .B(core__abc_21380_n8249), .Y(core__abc_21380_n8250) );
  OR2X2 OR2X2_3013 ( .A(core__abc_21380_n7076_bF_buf5), .B(core__abc_21380_n8250), .Y(core__abc_21380_n8251) );
  OR2X2 OR2X2_3014 ( .A(core__abc_21380_n8246), .B(core__abc_21380_n8251), .Y(core__abc_21380_n8252) );
  OR2X2 OR2X2_3015 ( .A(core__abc_21380_n7087_bF_buf4), .B(core_v2_reg_51_), .Y(core__abc_21380_n8253) );
  OR2X2 OR2X2_3016 ( .A(core__abc_21380_n8256), .B(core__abc_21380_n6861), .Y(core__abc_21380_n8257) );
  OR2X2 OR2X2_3017 ( .A(core__abc_21380_n8257), .B(core__abc_21380_n6821), .Y(core__abc_21380_n8260) );
  OR2X2 OR2X2_3018 ( .A(core__abc_21380_n8264), .B(core__abc_21380_n8265), .Y(core__abc_21380_n8266) );
  OR2X2 OR2X2_3019 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n8266), .Y(core__abc_21380_n8267) );
  OR2X2 OR2X2_302 ( .A(_abc_19068_n1547_1), .B(_abc_19068_n1548), .Y(_abc_19068_n1549_1) );
  OR2X2 OR2X2_3020 ( .A(core__abc_21380_n8262), .B(core__abc_21380_n8267), .Y(core__abc_21380_n8268) );
  OR2X2 OR2X2_3021 ( .A(core__abc_21380_n7087_bF_buf3), .B(core_v2_reg_52_), .Y(core__abc_21380_n8269) );
  OR2X2 OR2X2_3022 ( .A(core__abc_21380_n8275), .B(core__abc_21380_n8276), .Y(core__abc_21380_n8277) );
  OR2X2 OR2X2_3023 ( .A(core__abc_21380_n8280), .B(core__abc_21380_n8281), .Y(core__abc_21380_n8282) );
  OR2X2 OR2X2_3024 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n8282), .Y(core__abc_21380_n8283) );
  OR2X2 OR2X2_3025 ( .A(core__abc_21380_n8278), .B(core__abc_21380_n8283), .Y(core__abc_21380_n8284) );
  OR2X2 OR2X2_3026 ( .A(core__abc_21380_n7087_bF_buf2), .B(core_v2_reg_53_), .Y(core__abc_21380_n8285) );
  OR2X2 OR2X2_3027 ( .A(core__abc_21380_n8288), .B(core__abc_21380_n6811), .Y(core__abc_21380_n8289) );
  OR2X2 OR2X2_3028 ( .A(core__abc_21380_n8289), .B(core__abc_21380_n6801), .Y(core__abc_21380_n8291) );
  OR2X2 OR2X2_3029 ( .A(core__abc_21380_n8292), .B(core__abc_21380_n8290), .Y(core__abc_21380_n8293) );
  OR2X2 OR2X2_303 ( .A(_abc_19068_n1550), .B(_abc_19068_n1551_1), .Y(_abc_19068_n1552) );
  OR2X2 OR2X2_3030 ( .A(core__abc_21380_n8297), .B(core__abc_21380_n8298), .Y(core__abc_21380_n8299) );
  OR2X2 OR2X2_3031 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n8299), .Y(core__abc_21380_n8300) );
  OR2X2 OR2X2_3032 ( .A(core__abc_21380_n8295), .B(core__abc_21380_n8300), .Y(core__abc_21380_n8301) );
  OR2X2 OR2X2_3033 ( .A(core__abc_21380_n7087_bF_buf1), .B(core_v2_reg_54_), .Y(core__abc_21380_n8302) );
  OR2X2 OR2X2_3034 ( .A(core__abc_21380_n8306), .B(core__abc_21380_n8305), .Y(core__abc_21380_n8309) );
  OR2X2 OR2X2_3035 ( .A(core__abc_21380_n8312), .B(core__abc_21380_n8313), .Y(core__abc_21380_n8314) );
  OR2X2 OR2X2_3036 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n8314), .Y(core__abc_21380_n8315) );
  OR2X2 OR2X2_3037 ( .A(core__abc_21380_n8311), .B(core__abc_21380_n8315), .Y(core__abc_21380_n8316) );
  OR2X2 OR2X2_3038 ( .A(core__abc_21380_n7087_bF_buf0), .B(core_v2_reg_55_), .Y(core__abc_21380_n8317) );
  OR2X2 OR2X2_3039 ( .A(core__abc_21380_n8322), .B(core__abc_21380_n8320), .Y(core__abc_21380_n8323) );
  OR2X2 OR2X2_304 ( .A(_abc_19068_n1549_1), .B(_abc_19068_n1552), .Y(_abc_19068_n1553_1) );
  OR2X2 OR2X2_3040 ( .A(core__abc_21380_n8326), .B(core__abc_21380_n8327), .Y(core__abc_21380_n8328) );
  OR2X2 OR2X2_3041 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n8328), .Y(core__abc_21380_n8329) );
  OR2X2 OR2X2_3042 ( .A(core__abc_21380_n8325), .B(core__abc_21380_n8329), .Y(core__abc_21380_n8330) );
  OR2X2 OR2X2_3043 ( .A(core__abc_21380_n7087_bF_buf7), .B(core_v2_reg_56_), .Y(core__abc_21380_n8331) );
  OR2X2 OR2X2_3044 ( .A(core__abc_21380_n8338), .B(core__abc_21380_n8339), .Y(core__abc_21380_n8340) );
  OR2X2 OR2X2_3045 ( .A(core__abc_21380_n8342), .B(core__abc_21380_n8343), .Y(core__abc_21380_n8344) );
  OR2X2 OR2X2_3046 ( .A(core__abc_21380_n7076_bF_buf6), .B(core__abc_21380_n8344), .Y(core__abc_21380_n8345) );
  OR2X2 OR2X2_3047 ( .A(core__abc_21380_n8341), .B(core__abc_21380_n8345), .Y(core__abc_21380_n8346) );
  OR2X2 OR2X2_3048 ( .A(core__abc_21380_n7087_bF_buf6), .B(core_v2_reg_57_), .Y(core__abc_21380_n8347) );
  OR2X2 OR2X2_3049 ( .A(core__abc_21380_n8350), .B(core__abc_21380_n6743), .Y(core__abc_21380_n8351) );
  OR2X2 OR2X2_305 ( .A(_abc_19068_n1553_1), .B(_abc_19068_n1546), .Y(_abc_19068_n1554) );
  OR2X2 OR2X2_3050 ( .A(core__abc_21380_n8351), .B(core__abc_21380_n6737), .Y(core__abc_21380_n8353) );
  OR2X2 OR2X2_3051 ( .A(core__abc_21380_n8354), .B(core__abc_21380_n8352), .Y(core__abc_21380_n8355) );
  OR2X2 OR2X2_3052 ( .A(core__abc_21380_n8359), .B(core__abc_21380_n8360), .Y(core__abc_21380_n8361) );
  OR2X2 OR2X2_3053 ( .A(core__abc_21380_n7076_bF_buf5), .B(core__abc_21380_n8361), .Y(core__abc_21380_n8362) );
  OR2X2 OR2X2_3054 ( .A(core__abc_21380_n8357), .B(core__abc_21380_n8362), .Y(core__abc_21380_n8363) );
  OR2X2 OR2X2_3055 ( .A(core__abc_21380_n7087_bF_buf5), .B(core_v2_reg_58_), .Y(core__abc_21380_n8364) );
  OR2X2 OR2X2_3056 ( .A(core__abc_21380_n8368), .B(core__abc_21380_n8367), .Y(core__abc_21380_n8371) );
  OR2X2 OR2X2_3057 ( .A(core__abc_21380_n8375), .B(core__abc_21380_n8376), .Y(core__abc_21380_n8377) );
  OR2X2 OR2X2_3058 ( .A(core__abc_21380_n7076_bF_buf4), .B(core__abc_21380_n8377), .Y(core__abc_21380_n8378) );
  OR2X2 OR2X2_3059 ( .A(core__abc_21380_n8373), .B(core__abc_21380_n8378), .Y(core__abc_21380_n8379) );
  OR2X2 OR2X2_306 ( .A(_abc_19068_n1554), .B(_abc_19068_n1541_1), .Y(_abc_19068_n1555_1) );
  OR2X2 OR2X2_3060 ( .A(core__abc_21380_n7087_bF_buf4), .B(core_v2_reg_59_), .Y(core__abc_21380_n8380) );
  OR2X2 OR2X2_3061 ( .A(core__abc_21380_n8383), .B(core__abc_21380_n6763), .Y(core__abc_21380_n8384) );
  OR2X2 OR2X2_3062 ( .A(core__abc_21380_n8386), .B(core__abc_21380_n8387), .Y(core__abc_21380_n8388) );
  OR2X2 OR2X2_3063 ( .A(core__abc_21380_n8391), .B(core__abc_21380_n8392), .Y(core__abc_21380_n8393) );
  OR2X2 OR2X2_3064 ( .A(core__abc_21380_n7076_bF_buf3), .B(core__abc_21380_n8393), .Y(core__abc_21380_n8394) );
  OR2X2 OR2X2_3065 ( .A(core__abc_21380_n8390), .B(core__abc_21380_n8394), .Y(core__abc_21380_n8395) );
  OR2X2 OR2X2_3066 ( .A(core__abc_21380_n7087_bF_buf3), .B(core_v2_reg_60_), .Y(core__abc_21380_n8396) );
  OR2X2 OR2X2_3067 ( .A(core__abc_21380_n8403), .B(core__abc_21380_n8404), .Y(core__abc_21380_n8405) );
  OR2X2 OR2X2_3068 ( .A(core__abc_21380_n8408), .B(core__abc_21380_n8409), .Y(core__abc_21380_n8410) );
  OR2X2 OR2X2_3069 ( .A(core__abc_21380_n7076_bF_buf2), .B(core__abc_21380_n8410), .Y(core__abc_21380_n8411) );
  OR2X2 OR2X2_307 ( .A(_abc_19068_n1557), .B(_abc_19068_n1558_1), .Y(_abc_19068_n1559) );
  OR2X2 OR2X2_3070 ( .A(core__abc_21380_n8406), .B(core__abc_21380_n8411), .Y(core__abc_21380_n8412) );
  OR2X2 OR2X2_3071 ( .A(core__abc_21380_n7087_bF_buf2), .B(core_v2_reg_61_), .Y(core__abc_21380_n8413) );
  OR2X2 OR2X2_3072 ( .A(core__abc_21380_n8416), .B(core__abc_21380_n6710), .Y(core__abc_21380_n8417) );
  OR2X2 OR2X2_3073 ( .A(core__abc_21380_n8417), .B(core__abc_21380_n6700), .Y(core__abc_21380_n8419) );
  OR2X2 OR2X2_3074 ( .A(core__abc_21380_n8420), .B(core__abc_21380_n8418), .Y(core__abc_21380_n8421) );
  OR2X2 OR2X2_3075 ( .A(core__abc_21380_n8425), .B(core__abc_21380_n8426), .Y(core__abc_21380_n8427) );
  OR2X2 OR2X2_3076 ( .A(core__abc_21380_n7076_bF_buf1), .B(core__abc_21380_n8427), .Y(core__abc_21380_n8428) );
  OR2X2 OR2X2_3077 ( .A(core__abc_21380_n8423), .B(core__abc_21380_n8428), .Y(core__abc_21380_n8429) );
  OR2X2 OR2X2_3078 ( .A(core__abc_21380_n7087_bF_buf1), .B(core_v2_reg_62_), .Y(core__abc_21380_n8430) );
  OR2X2 OR2X2_3079 ( .A(core__abc_21380_n8434), .B(core__abc_21380_n8433), .Y(core__abc_21380_n8437) );
  OR2X2 OR2X2_308 ( .A(_abc_19068_n1560), .B(_abc_19068_n1561_1), .Y(_abc_19068_n1562) );
  OR2X2 OR2X2_3080 ( .A(core__abc_21380_n8440), .B(core__abc_21380_n8441), .Y(core__abc_21380_n8442) );
  OR2X2 OR2X2_3081 ( .A(core__abc_21380_n7076_bF_buf0), .B(core__abc_21380_n8442), .Y(core__abc_21380_n8443) );
  OR2X2 OR2X2_3082 ( .A(core__abc_21380_n8439), .B(core__abc_21380_n8443), .Y(core__abc_21380_n8444) );
  OR2X2 OR2X2_3083 ( .A(core__abc_21380_n7087_bF_buf0), .B(core_v2_reg_63_), .Y(core__abc_21380_n8445) );
  OR2X2 OR2X2_3084 ( .A(core__abc_21380_n7487), .B(core__abc_21380_n7973), .Y(core__abc_21380_n8448) );
  OR2X2 OR2X2_3085 ( .A(core__abc_21380_n7486), .B(core__abc_21380_n8449), .Y(core__abc_21380_n8450) );
  OR2X2 OR2X2_3086 ( .A(core__abc_21380_n3313_bF_buf0), .B(core__abc_21380_n3166), .Y(core__abc_21380_n8453) );
  OR2X2 OR2X2_3087 ( .A(core__abc_21380_n8457), .B(core__abc_21380_n3319), .Y(core__abc_21380_n8458) );
  OR2X2 OR2X2_3088 ( .A(core__abc_21380_n8458), .B(core__abc_21380_n8455_bF_buf7), .Y(core__abc_21380_n8459) );
  OR2X2 OR2X2_3089 ( .A(core__abc_21380_n8451), .B(core__abc_21380_n8459), .Y(core__abc_21380_n8460) );
  OR2X2 OR2X2_309 ( .A(_abc_19068_n1559), .B(_abc_19068_n1562), .Y(_abc_19068_n1563_1) );
  OR2X2 OR2X2_3090 ( .A(core__abc_21380_n8454_bF_buf6), .B(core_v1_reg_0_), .Y(core__abc_21380_n8461) );
  OR2X2 OR2X2_3091 ( .A(core__abc_21380_n7521), .B(core__abc_21380_n7982), .Y(core__abc_21380_n8464) );
  OR2X2 OR2X2_3092 ( .A(core__abc_21380_n7519), .B(core__abc_21380_n8465), .Y(core__abc_21380_n8466) );
  OR2X2 OR2X2_3093 ( .A(core__abc_21380_n8470), .B(core__abc_21380_n8471), .Y(core__abc_21380_n8472) );
  OR2X2 OR2X2_3094 ( .A(core__abc_21380_n8469), .B(core__abc_21380_n8473), .Y(core__abc_21380_n8474) );
  OR2X2 OR2X2_3095 ( .A(core__abc_21380_n8474), .B(core__abc_21380_n8455_bF_buf6), .Y(core__abc_21380_n8475) );
  OR2X2 OR2X2_3096 ( .A(core__abc_21380_n8468), .B(core__abc_21380_n8475), .Y(core__abc_21380_n8476) );
  OR2X2 OR2X2_3097 ( .A(core__abc_21380_n8454_bF_buf5), .B(core_v1_reg_1_), .Y(core__abc_21380_n8477) );
  OR2X2 OR2X2_3098 ( .A(core__abc_21380_n7553), .B(core__abc_21380_n8481), .Y(core__abc_21380_n8482) );
  OR2X2 OR2X2_3099 ( .A(core__abc_21380_n7554), .B(core__abc_21380_n7994), .Y(core__abc_21380_n8483) );
  OR2X2 OR2X2_31 ( .A(_abc_19068_n968), .B(_abc_19068_n969_1), .Y(_abc_19068_n970_1) );
  OR2X2 OR2X2_310 ( .A(_abc_19068_n1564), .B(_abc_19068_n1565_1), .Y(_abc_19068_n1566) );
  OR2X2 OR2X2_3100 ( .A(core__abc_21380_n7079), .B(core_key_66_), .Y(core__abc_21380_n8486) );
  OR2X2 OR2X2_3101 ( .A(core__abc_21380_n8487), .B(core_long), .Y(core__abc_21380_n8488) );
  OR2X2 OR2X2_3102 ( .A(core__abc_21380_n8485), .B(core__abc_21380_n8490), .Y(core__abc_21380_n8491) );
  OR2X2 OR2X2_3103 ( .A(core__abc_21380_n8491), .B(core__abc_21380_n8455_bF_buf5), .Y(core__abc_21380_n8492) );
  OR2X2 OR2X2_3104 ( .A(core__abc_21380_n8484), .B(core__abc_21380_n8492), .Y(core__abc_21380_n8493) );
  OR2X2 OR2X2_3105 ( .A(core__abc_21380_n8454_bF_buf4), .B(core_v1_reg_2_), .Y(core__abc_21380_n8494) );
  OR2X2 OR2X2_3106 ( .A(core__abc_21380_n7583), .B(core__abc_21380_n8003), .Y(core__abc_21380_n8497) );
  OR2X2 OR2X2_3107 ( .A(core__abc_21380_n7581), .B(core__abc_21380_n8498), .Y(core__abc_21380_n8499) );
  OR2X2 OR2X2_3108 ( .A(core__abc_21380_n7079), .B(core_key_67_), .Y(core__abc_21380_n8503) );
  OR2X2 OR2X2_3109 ( .A(core__abc_21380_n8504), .B(core_long), .Y(core__abc_21380_n8505) );
  OR2X2 OR2X2_311 ( .A(_abc_19068_n1567_1), .B(_abc_19068_n1568), .Y(_abc_19068_n1569_1) );
  OR2X2 OR2X2_3110 ( .A(core__abc_21380_n8502), .B(core__abc_21380_n8507), .Y(core__abc_21380_n8508) );
  OR2X2 OR2X2_3111 ( .A(core__abc_21380_n8508), .B(core__abc_21380_n8455_bF_buf4), .Y(core__abc_21380_n8509) );
  OR2X2 OR2X2_3112 ( .A(core__abc_21380_n8501), .B(core__abc_21380_n8509), .Y(core__abc_21380_n8510) );
  OR2X2 OR2X2_3113 ( .A(core__abc_21380_n8454_bF_buf3), .B(core_v1_reg_3_), .Y(core__abc_21380_n8511) );
  OR2X2 OR2X2_3114 ( .A(core__abc_21380_n7604), .B(core__abc_21380_n8515), .Y(core__abc_21380_n8516) );
  OR2X2 OR2X2_3115 ( .A(core__abc_21380_n7605), .B(core__abc_21380_n8016), .Y(core__abc_21380_n8517) );
  OR2X2 OR2X2_3116 ( .A(core__abc_21380_n8455_bF_buf3), .B(core__abc_21380_n8520), .Y(core__abc_21380_n8521) );
  OR2X2 OR2X2_3117 ( .A(core__abc_21380_n8521), .B(core__abc_21380_n8519), .Y(core__abc_21380_n8522) );
  OR2X2 OR2X2_3118 ( .A(core__abc_21380_n8518), .B(core__abc_21380_n8522), .Y(core__abc_21380_n8523) );
  OR2X2 OR2X2_3119 ( .A(core__abc_21380_n8454_bF_buf2), .B(core_v1_reg_4_), .Y(core__abc_21380_n8524) );
  OR2X2 OR2X2_312 ( .A(_abc_19068_n1566), .B(_abc_19068_n1569_1), .Y(_abc_19068_n1570) );
  OR2X2 OR2X2_3120 ( .A(core__abc_21380_n7637), .B(core__abc_21380_n8027), .Y(core__abc_21380_n8527) );
  OR2X2 OR2X2_3121 ( .A(core__abc_21380_n7636), .B(core__abc_21380_n8528), .Y(core__abc_21380_n8529) );
  OR2X2 OR2X2_3122 ( .A(core__abc_21380_n7079), .B(core_key_69_), .Y(core__abc_21380_n8533) );
  OR2X2 OR2X2_3123 ( .A(core__abc_21380_n3653), .B(core_long), .Y(core__abc_21380_n8534) );
  OR2X2 OR2X2_3124 ( .A(core__abc_21380_n8532), .B(core__abc_21380_n8536), .Y(core__abc_21380_n8537) );
  OR2X2 OR2X2_3125 ( .A(core__abc_21380_n8537), .B(core__abc_21380_n8455_bF_buf2), .Y(core__abc_21380_n8538) );
  OR2X2 OR2X2_3126 ( .A(core__abc_21380_n8531), .B(core__abc_21380_n8538), .Y(core__abc_21380_n8539) );
  OR2X2 OR2X2_3127 ( .A(core__abc_21380_n8454_bF_buf1), .B(core_v1_reg_5_), .Y(core__abc_21380_n8540) );
  OR2X2 OR2X2_3128 ( .A(core__abc_21380_n8544), .B(core__abc_21380_n7657), .Y(core__abc_21380_n8545) );
  OR2X2 OR2X2_3129 ( .A(core__abc_21380_n7658), .B(core__abc_21380_n8042), .Y(core__abc_21380_n8546) );
  OR2X2 OR2X2_313 ( .A(_abc_19068_n1571_1), .B(_abc_19068_n1572), .Y(_abc_19068_n1573_1) );
  OR2X2 OR2X2_3130 ( .A(core__abc_21380_n8549), .B(core__abc_21380_n8550), .Y(core__abc_21380_n8551) );
  OR2X2 OR2X2_3131 ( .A(core__abc_21380_n8455_bF_buf1), .B(core__abc_21380_n8552), .Y(core__abc_21380_n8553) );
  OR2X2 OR2X2_3132 ( .A(core__abc_21380_n8553), .B(core__abc_21380_n8548), .Y(core__abc_21380_n8554) );
  OR2X2 OR2X2_3133 ( .A(core__abc_21380_n8547), .B(core__abc_21380_n8554), .Y(core__abc_21380_n8555) );
  OR2X2 OR2X2_3134 ( .A(core__abc_21380_n8454_bF_buf0), .B(core_v1_reg_6_), .Y(core__abc_21380_n8556) );
  OR2X2 OR2X2_3135 ( .A(core__abc_21380_n8057), .B(core__abc_21380_n7687), .Y(core__abc_21380_n8559) );
  OR2X2 OR2X2_3136 ( .A(core__abc_21380_n8560), .B(core__abc_21380_n7686), .Y(core__abc_21380_n8561) );
  OR2X2 OR2X2_3137 ( .A(core_key_71_), .B(core_long), .Y(core__abc_21380_n8567) );
  OR2X2 OR2X2_3138 ( .A(core__abc_21380_n8564), .B(core__abc_21380_n8569), .Y(core__abc_21380_n8570) );
  OR2X2 OR2X2_3139 ( .A(core__abc_21380_n8570), .B(core__abc_21380_n8455_bF_buf0), .Y(core__abc_21380_n8571) );
  OR2X2 OR2X2_314 ( .A(_abc_19068_n910_1), .B(_abc_19068_n1573_1), .Y(_abc_19068_n1574) );
  OR2X2 OR2X2_3140 ( .A(core__abc_21380_n8563), .B(core__abc_21380_n8571), .Y(core__abc_21380_n8572) );
  OR2X2 OR2X2_3141 ( .A(core__abc_21380_n8454_bF_buf7), .B(core_v1_reg_7_), .Y(core__abc_21380_n8573) );
  OR2X2 OR2X2_3142 ( .A(core__abc_21380_n8576), .B(core__abc_21380_n7709), .Y(core__abc_21380_n8577) );
  OR2X2 OR2X2_3143 ( .A(core__abc_21380_n8072), .B(core__abc_21380_n7710), .Y(core__abc_21380_n8578) );
  OR2X2 OR2X2_3144 ( .A(core__abc_21380_n8580), .B(core__abc_21380_n3867), .Y(core__abc_21380_n8581) );
  OR2X2 OR2X2_3145 ( .A(core__abc_21380_n8581), .B(core__abc_21380_n8455_bF_buf7), .Y(core__abc_21380_n8582) );
  OR2X2 OR2X2_3146 ( .A(core__abc_21380_n8579), .B(core__abc_21380_n8582), .Y(core__abc_21380_n8583) );
  OR2X2 OR2X2_3147 ( .A(core__abc_21380_n8454_bF_buf6), .B(core_v1_reg_8_), .Y(core__abc_21380_n8584) );
  OR2X2 OR2X2_3148 ( .A(core__abc_21380_n8088), .B(core__abc_21380_n7751), .Y(core__abc_21380_n8587) );
  OR2X2 OR2X2_3149 ( .A(core__abc_21380_n8087), .B(core__abc_21380_n7749), .Y(core__abc_21380_n8588) );
  OR2X2 OR2X2_315 ( .A(_abc_19068_n1574), .B(_abc_19068_n1570), .Y(_abc_19068_n1575) );
  OR2X2 OR2X2_3150 ( .A(core__abc_21380_n8591), .B(core__abc_21380_n8593), .Y(core__abc_21380_n8594) );
  OR2X2 OR2X2_3151 ( .A(core__abc_21380_n8594), .B(core__abc_21380_n8455_bF_buf6), .Y(core__abc_21380_n8595) );
  OR2X2 OR2X2_3152 ( .A(core__abc_21380_n8590), .B(core__abc_21380_n8595), .Y(core__abc_21380_n8596) );
  OR2X2 OR2X2_3153 ( .A(core__abc_21380_n8454_bF_buf5), .B(core_v1_reg_9_), .Y(core__abc_21380_n8597) );
  OR2X2 OR2X2_3154 ( .A(core__abc_21380_n8600), .B(core__abc_21380_n7776), .Y(core__abc_21380_n8601) );
  OR2X2 OR2X2_3155 ( .A(core__abc_21380_n8104), .B(core__abc_21380_n7773), .Y(core__abc_21380_n8602) );
  OR2X2 OR2X2_3156 ( .A(core__abc_21380_n8605), .B(core__abc_21380_n3994), .Y(core__abc_21380_n8606) );
  OR2X2 OR2X2_3157 ( .A(core__abc_21380_n8606), .B(core__abc_21380_n8455_bF_buf5), .Y(core__abc_21380_n8607) );
  OR2X2 OR2X2_3158 ( .A(core__abc_21380_n8604), .B(core__abc_21380_n8607), .Y(core__abc_21380_n8608) );
  OR2X2 OR2X2_3159 ( .A(core__abc_21380_n8454_bF_buf4), .B(core_v1_reg_10_), .Y(core__abc_21380_n8609) );
  OR2X2 OR2X2_316 ( .A(_abc_19068_n1575), .B(_abc_19068_n1563_1), .Y(_abc_19068_n1576) );
  OR2X2 OR2X2_3160 ( .A(core__abc_21380_n8120), .B(core__abc_21380_n7800), .Y(core__abc_21380_n8612) );
  OR2X2 OR2X2_3161 ( .A(core__abc_21380_n8613), .B(core__abc_21380_n7798), .Y(core__abc_21380_n8614) );
  OR2X2 OR2X2_3162 ( .A(core__abc_21380_n8617), .B(core__abc_21380_n8619), .Y(core__abc_21380_n8620) );
  OR2X2 OR2X2_3163 ( .A(core__abc_21380_n8620), .B(core__abc_21380_n8455_bF_buf4), .Y(core__abc_21380_n8621) );
  OR2X2 OR2X2_3164 ( .A(core__abc_21380_n8616), .B(core__abc_21380_n8621), .Y(core__abc_21380_n8622) );
  OR2X2 OR2X2_3165 ( .A(core__abc_21380_n8454_bF_buf3), .B(core_v1_reg_11_), .Y(core__abc_21380_n8623) );
  OR2X2 OR2X2_3166 ( .A(core__abc_21380_n8133), .B(core__abc_21380_n7827), .Y(core__abc_21380_n8626) );
  OR2X2 OR2X2_3167 ( .A(core__abc_21380_n8134), .B(core__abc_21380_n7828), .Y(core__abc_21380_n8627) );
  OR2X2 OR2X2_3168 ( .A(core__abc_21380_n8630), .B(core__abc_21380_n4140), .Y(core__abc_21380_n8631) );
  OR2X2 OR2X2_3169 ( .A(core__abc_21380_n8631), .B(core__abc_21380_n8455_bF_buf3), .Y(core__abc_21380_n8632) );
  OR2X2 OR2X2_317 ( .A(_abc_19068_n1248), .B(_abc_19068_n1578), .Y(_abc_19068_n1579) );
  OR2X2 OR2X2_3170 ( .A(core__abc_21380_n8629), .B(core__abc_21380_n8632), .Y(core__abc_21380_n8633) );
  OR2X2 OR2X2_3171 ( .A(core__abc_21380_n8454_bF_buf2), .B(core_v1_reg_12_), .Y(core__abc_21380_n8634) );
  OR2X2 OR2X2_3172 ( .A(core__abc_21380_n8150), .B(core__abc_21380_n7868), .Y(core__abc_21380_n8637) );
  OR2X2 OR2X2_3173 ( .A(core__abc_21380_n8149), .B(core__abc_21380_n7866), .Y(core__abc_21380_n8638) );
  OR2X2 OR2X2_3174 ( .A(core__abc_21380_n8641), .B(core__abc_21380_n4210_1), .Y(core__abc_21380_n8642) );
  OR2X2 OR2X2_3175 ( .A(core__abc_21380_n8642), .B(core__abc_21380_n8455_bF_buf2), .Y(core__abc_21380_n8643) );
  OR2X2 OR2X2_3176 ( .A(core__abc_21380_n8640), .B(core__abc_21380_n8643), .Y(core__abc_21380_n8644) );
  OR2X2 OR2X2_3177 ( .A(core__abc_21380_n8454_bF_buf1), .B(core_v1_reg_13_), .Y(core__abc_21380_n8645) );
  OR2X2 OR2X2_3178 ( .A(core__abc_21380_n8648), .B(core__abc_21380_n7891), .Y(core__abc_21380_n8649) );
  OR2X2 OR2X2_3179 ( .A(core__abc_21380_n8166), .B(core__abc_21380_n7893), .Y(core__abc_21380_n8650) );
  OR2X2 OR2X2_318 ( .A(_abc_19068_n1580_1), .B(_abc_19068_n1581), .Y(_abc_19068_n1582) );
  OR2X2 OR2X2_3180 ( .A(core__abc_21380_n8653), .B(core__abc_21380_n4280), .Y(core__abc_21380_n8654) );
  OR2X2 OR2X2_3181 ( .A(core__abc_21380_n8654), .B(core__abc_21380_n8455_bF_buf1), .Y(core__abc_21380_n8655) );
  OR2X2 OR2X2_3182 ( .A(core__abc_21380_n8652), .B(core__abc_21380_n8655), .Y(core__abc_21380_n8656) );
  OR2X2 OR2X2_3183 ( .A(core__abc_21380_n8454_bF_buf0), .B(core_v1_reg_14_), .Y(core__abc_21380_n8657) );
  OR2X2 OR2X2_3184 ( .A(core__abc_21380_n8183), .B(core__abc_21380_n7922), .Y(core__abc_21380_n8660) );
  OR2X2 OR2X2_3185 ( .A(core__abc_21380_n8182), .B(core__abc_21380_n7921), .Y(core__abc_21380_n8661) );
  OR2X2 OR2X2_3186 ( .A(core__abc_21380_n8664), .B(core__abc_21380_n4339_1), .Y(core__abc_21380_n8665) );
  OR2X2 OR2X2_3187 ( .A(core__abc_21380_n8665), .B(core__abc_21380_n8455_bF_buf0), .Y(core__abc_21380_n8666) );
  OR2X2 OR2X2_3188 ( .A(core__abc_21380_n8663), .B(core__abc_21380_n8666), .Y(core__abc_21380_n8667) );
  OR2X2 OR2X2_3189 ( .A(core__abc_21380_n8454_bF_buf7), .B(core_v1_reg_15_), .Y(core__abc_21380_n8668) );
  OR2X2 OR2X2_319 ( .A(_abc_19068_n1579), .B(_abc_19068_n1582), .Y(_abc_19068_n1583_1) );
  OR2X2 OR2X2_3190 ( .A(core__abc_21380_n8196), .B(core__abc_21380_n7948), .Y(core__abc_21380_n8671) );
  OR2X2 OR2X2_3191 ( .A(core__abc_21380_n8197), .B(core__abc_21380_n7949), .Y(core__abc_21380_n8672) );
  OR2X2 OR2X2_3192 ( .A(core__abc_21380_n8675), .B(core__abc_21380_n4434), .Y(core__abc_21380_n8676) );
  OR2X2 OR2X2_3193 ( .A(core__abc_21380_n8676), .B(core__abc_21380_n8455_bF_buf7), .Y(core__abc_21380_n8677) );
  OR2X2 OR2X2_3194 ( .A(core__abc_21380_n8674), .B(core__abc_21380_n8677), .Y(core__abc_21380_n8678) );
  OR2X2 OR2X2_3195 ( .A(core__abc_21380_n8454_bF_buf6), .B(core_v1_reg_16_), .Y(core__abc_21380_n8679) );
  OR2X2 OR2X2_3196 ( .A(core__abc_21380_n8213), .B(core__abc_21380_n7012), .Y(core__abc_21380_n8682) );
  OR2X2 OR2X2_3197 ( .A(core__abc_21380_n8683), .B(core__abc_21380_n7969), .Y(core__abc_21380_n8684) );
  OR2X2 OR2X2_3198 ( .A(core__abc_21380_n8687), .B(core__abc_21380_n4501_1), .Y(core__abc_21380_n8688) );
  OR2X2 OR2X2_3199 ( .A(core__abc_21380_n8688), .B(core__abc_21380_n8455_bF_buf6), .Y(core__abc_21380_n8689) );
  OR2X2 OR2X2_32 ( .A(_abc_19068_n971), .B(_abc_19068_n972_1), .Y(_abc_19068_n973_1) );
  OR2X2 OR2X2_320 ( .A(_abc_19068_n1585), .B(_abc_19068_n1586), .Y(_abc_19068_n1587_1) );
  OR2X2 OR2X2_3200 ( .A(core__abc_21380_n8686), .B(core__abc_21380_n8689), .Y(core__abc_21380_n8690) );
  OR2X2 OR2X2_3201 ( .A(core__abc_21380_n8454_bF_buf5), .B(core_v1_reg_17_), .Y(core__abc_21380_n8691) );
  OR2X2 OR2X2_3202 ( .A(core__abc_21380_n8229), .B(core__abc_21380_n7008), .Y(core__abc_21380_n8694) );
  OR2X2 OR2X2_3203 ( .A(core__abc_21380_n8228), .B(core__abc_21380_n7007), .Y(core__abc_21380_n8695) );
  OR2X2 OR2X2_3204 ( .A(core__abc_21380_n8698), .B(core__abc_21380_n4562), .Y(core__abc_21380_n8699) );
  OR2X2 OR2X2_3205 ( .A(core__abc_21380_n8699), .B(core__abc_21380_n8455_bF_buf5), .Y(core__abc_21380_n8700) );
  OR2X2 OR2X2_3206 ( .A(core__abc_21380_n8697), .B(core__abc_21380_n8700), .Y(core__abc_21380_n8701) );
  OR2X2 OR2X2_3207 ( .A(core__abc_21380_n8454_bF_buf4), .B(core_v1_reg_18_), .Y(core__abc_21380_n8702) );
  OR2X2 OR2X2_3208 ( .A(core__abc_21380_n8245), .B(core__abc_21380_n7002), .Y(core__abc_21380_n8705) );
  OR2X2 OR2X2_3209 ( .A(core__abc_21380_n8244), .B(core__abc_21380_n7001), .Y(core__abc_21380_n8706) );
  OR2X2 OR2X2_321 ( .A(_abc_19068_n1587_1), .B(_abc_19068_n1584), .Y(_abc_19068_n1588) );
  OR2X2 OR2X2_3210 ( .A(core__abc_21380_n8709), .B(core__abc_21380_n4620), .Y(core__abc_21380_n8710) );
  OR2X2 OR2X2_3211 ( .A(core__abc_21380_n8710), .B(core__abc_21380_n8455_bF_buf4), .Y(core__abc_21380_n8711) );
  OR2X2 OR2X2_3212 ( .A(core__abc_21380_n8708), .B(core__abc_21380_n8711), .Y(core__abc_21380_n8712) );
  OR2X2 OR2X2_3213 ( .A(core__abc_21380_n8454_bF_buf3), .B(core_v1_reg_19_), .Y(core__abc_21380_n8713) );
  OR2X2 OR2X2_3214 ( .A(core__abc_21380_n8716), .B(core__abc_21380_n6993), .Y(core__abc_21380_n8717) );
  OR2X2 OR2X2_3215 ( .A(core__abc_21380_n8261), .B(core__abc_21380_n8718), .Y(core__abc_21380_n8719) );
  OR2X2 OR2X2_3216 ( .A(core__abc_21380_n8722), .B(core__abc_21380_n8723), .Y(core__abc_21380_n8724) );
  OR2X2 OR2X2_3217 ( .A(core__abc_21380_n8724), .B(core__abc_21380_n8455_bF_buf3), .Y(core__abc_21380_n8725) );
  OR2X2 OR2X2_3218 ( .A(core__abc_21380_n8721), .B(core__abc_21380_n8725), .Y(core__abc_21380_n8726) );
  OR2X2 OR2X2_3219 ( .A(core__abc_21380_n8454_bF_buf2), .B(core_v1_reg_20_), .Y(core__abc_21380_n8727) );
  OR2X2 OR2X2_322 ( .A(_abc_19068_n1589_1), .B(_abc_19068_n1590), .Y(_abc_19068_n1591) );
  OR2X2 OR2X2_3220 ( .A(core__abc_21380_n8277), .B(core__abc_21380_n6989), .Y(core__abc_21380_n8730) );
  OR2X2 OR2X2_3221 ( .A(core__abc_21380_n8731), .B(core__abc_21380_n6988), .Y(core__abc_21380_n8732) );
  OR2X2 OR2X2_3222 ( .A(core__abc_21380_n8735), .B(core__abc_21380_n4737_1), .Y(core__abc_21380_n8736) );
  OR2X2 OR2X2_3223 ( .A(core__abc_21380_n8736), .B(core__abc_21380_n8455_bF_buf2), .Y(core__abc_21380_n8737) );
  OR2X2 OR2X2_3224 ( .A(core__abc_21380_n8734), .B(core__abc_21380_n8737), .Y(core__abc_21380_n8738) );
  OR2X2 OR2X2_3225 ( .A(core__abc_21380_n8454_bF_buf1), .B(core_v1_reg_21_), .Y(core__abc_21380_n8739) );
  OR2X2 OR2X2_3226 ( .A(core__abc_21380_n8293), .B(core__abc_21380_n6980), .Y(core__abc_21380_n8742) );
  OR2X2 OR2X2_3227 ( .A(core__abc_21380_n8294), .B(core__abc_21380_n6981), .Y(core__abc_21380_n8743) );
  OR2X2 OR2X2_3228 ( .A(core__abc_21380_n8746), .B(core__abc_21380_n4790), .Y(core__abc_21380_n8747) );
  OR2X2 OR2X2_3229 ( .A(core__abc_21380_n8747), .B(core__abc_21380_n8455_bF_buf1), .Y(core__abc_21380_n8748) );
  OR2X2 OR2X2_323 ( .A(_abc_19068_n1592), .B(_abc_19068_n1593), .Y(_abc_19068_n1594) );
  OR2X2 OR2X2_3230 ( .A(core__abc_21380_n8745), .B(core__abc_21380_n8748), .Y(core__abc_21380_n8749) );
  OR2X2 OR2X2_3231 ( .A(core__abc_21380_n8454_bF_buf0), .B(core_v1_reg_22_), .Y(core__abc_21380_n8750) );
  OR2X2 OR2X2_3232 ( .A(core__abc_21380_n8310), .B(core__abc_21380_n6968), .Y(core__abc_21380_n8753) );
  OR2X2 OR2X2_3233 ( .A(core__abc_21380_n8754), .B(core__abc_21380_n6967), .Y(core__abc_21380_n8755) );
  OR2X2 OR2X2_3234 ( .A(core__abc_21380_n8758), .B(core__abc_21380_n4838), .Y(core__abc_21380_n8759) );
  OR2X2 OR2X2_3235 ( .A(core__abc_21380_n8759), .B(core__abc_21380_n8455_bF_buf0), .Y(core__abc_21380_n8760) );
  OR2X2 OR2X2_3236 ( .A(core__abc_21380_n8757), .B(core__abc_21380_n8760), .Y(core__abc_21380_n8761) );
  OR2X2 OR2X2_3237 ( .A(core__abc_21380_n8454_bF_buf7), .B(core_v1_reg_23_), .Y(core__abc_21380_n8762) );
  OR2X2 OR2X2_3238 ( .A(core__abc_21380_n8324), .B(core__abc_21380_n6960), .Y(core__abc_21380_n8765) );
  OR2X2 OR2X2_3239 ( .A(core__abc_21380_n8323), .B(core__abc_21380_n6962), .Y(core__abc_21380_n8766) );
  OR2X2 OR2X2_324 ( .A(_abc_19068_n1591), .B(_abc_19068_n1594), .Y(_abc_19068_n1595) );
  OR2X2 OR2X2_3240 ( .A(core__abc_21380_n8769), .B(core__abc_21380_n8770), .Y(core__abc_21380_n8771) );
  OR2X2 OR2X2_3241 ( .A(core__abc_21380_n8771), .B(core__abc_21380_n8455_bF_buf7), .Y(core__abc_21380_n8772) );
  OR2X2 OR2X2_3242 ( .A(core__abc_21380_n8768), .B(core__abc_21380_n8772), .Y(core__abc_21380_n8773) );
  OR2X2 OR2X2_3243 ( .A(core__abc_21380_n8454_bF_buf6), .B(core_v1_reg_24_), .Y(core__abc_21380_n8774) );
  OR2X2 OR2X2_3244 ( .A(core__abc_21380_n8340), .B(core__abc_21380_n6944), .Y(core__abc_21380_n8777) );
  OR2X2 OR2X2_3245 ( .A(core__abc_21380_n8778), .B(core__abc_21380_n6943), .Y(core__abc_21380_n8779) );
  OR2X2 OR2X2_3246 ( .A(core__abc_21380_n8782), .B(core__abc_21380_n8784), .Y(core__abc_21380_n8785) );
  OR2X2 OR2X2_3247 ( .A(core__abc_21380_n8785), .B(core__abc_21380_n8455_bF_buf6), .Y(core__abc_21380_n8786) );
  OR2X2 OR2X2_3248 ( .A(core__abc_21380_n8781), .B(core__abc_21380_n8786), .Y(core__abc_21380_n8787) );
  OR2X2 OR2X2_3249 ( .A(core__abc_21380_n8454_bF_buf5), .B(core_v1_reg_25_), .Y(core__abc_21380_n8788) );
  OR2X2 OR2X2_325 ( .A(_abc_19068_n1595), .B(_abc_19068_n1588), .Y(_abc_19068_n1596) );
  OR2X2 OR2X2_3250 ( .A(core__abc_21380_n8355), .B(core__abc_21380_n6936), .Y(core__abc_21380_n8791) );
  OR2X2 OR2X2_3251 ( .A(core__abc_21380_n8356), .B(core__abc_21380_n6937), .Y(core__abc_21380_n8792) );
  OR2X2 OR2X2_3252 ( .A(core__abc_21380_n8795), .B(core__abc_21380_n8797), .Y(core__abc_21380_n8798) );
  OR2X2 OR2X2_3253 ( .A(core__abc_21380_n8798), .B(core__abc_21380_n8455_bF_buf5), .Y(core__abc_21380_n8799) );
  OR2X2 OR2X2_3254 ( .A(core__abc_21380_n8794), .B(core__abc_21380_n8799), .Y(core__abc_21380_n8800) );
  OR2X2 OR2X2_3255 ( .A(core__abc_21380_n8454_bF_buf4), .B(core_v1_reg_26_), .Y(core__abc_21380_n8801) );
  OR2X2 OR2X2_3256 ( .A(core__abc_21380_n8372), .B(core__abc_21380_n6927), .Y(core__abc_21380_n8804) );
  OR2X2 OR2X2_3257 ( .A(core__abc_21380_n8805), .B(core__abc_21380_n6926), .Y(core__abc_21380_n8806) );
  OR2X2 OR2X2_3258 ( .A(core__abc_21380_n8809), .B(core__abc_21380_n5061), .Y(core__abc_21380_n8810) );
  OR2X2 OR2X2_3259 ( .A(core__abc_21380_n8810), .B(core__abc_21380_n8455_bF_buf4), .Y(core__abc_21380_n8811) );
  OR2X2 OR2X2_326 ( .A(_abc_19068_n1596), .B(_abc_19068_n1583_1), .Y(_abc_19068_n1597) );
  OR2X2 OR2X2_3260 ( .A(core__abc_21380_n8808), .B(core__abc_21380_n8811), .Y(core__abc_21380_n8812) );
  OR2X2 OR2X2_3261 ( .A(core__abc_21380_n8454_bF_buf3), .B(core_v1_reg_27_), .Y(core__abc_21380_n8813) );
  OR2X2 OR2X2_3262 ( .A(core__abc_21380_n8389), .B(core__abc_21380_n8816), .Y(core__abc_21380_n8817) );
  OR2X2 OR2X2_3263 ( .A(core__abc_21380_n8388), .B(core__abc_21380_n6922), .Y(core__abc_21380_n8818) );
  OR2X2 OR2X2_3264 ( .A(core__abc_21380_n8821), .B(core__abc_21380_n8822), .Y(core__abc_21380_n8823) );
  OR2X2 OR2X2_3265 ( .A(core__abc_21380_n8823), .B(core__abc_21380_n8455_bF_buf3), .Y(core__abc_21380_n8824) );
  OR2X2 OR2X2_3266 ( .A(core__abc_21380_n8820), .B(core__abc_21380_n8824), .Y(core__abc_21380_n8825) );
  OR2X2 OR2X2_3267 ( .A(core__abc_21380_n8454_bF_buf2), .B(core_v1_reg_28_), .Y(core__abc_21380_n8826) );
  OR2X2 OR2X2_3268 ( .A(core__abc_21380_n8405), .B(core__abc_21380_n6902), .Y(core__abc_21380_n8829) );
  OR2X2 OR2X2_3269 ( .A(core__abc_21380_n8830), .B(core__abc_21380_n6901), .Y(core__abc_21380_n8831) );
  OR2X2 OR2X2_327 ( .A(_abc_19068_n1599), .B(_abc_19068_n1600), .Y(_abc_19068_n1601) );
  OR2X2 OR2X2_3270 ( .A(core__abc_21380_n8834), .B(core__abc_21380_n5183), .Y(core__abc_21380_n8835) );
  OR2X2 OR2X2_3271 ( .A(core__abc_21380_n8835), .B(core__abc_21380_n8455_bF_buf2), .Y(core__abc_21380_n8836) );
  OR2X2 OR2X2_3272 ( .A(core__abc_21380_n8833), .B(core__abc_21380_n8836), .Y(core__abc_21380_n8837) );
  OR2X2 OR2X2_3273 ( .A(core__abc_21380_n8454_bF_buf1), .B(core_v1_reg_29_), .Y(core__abc_21380_n8838) );
  OR2X2 OR2X2_3274 ( .A(core__abc_21380_n8421), .B(core__abc_21380_n6894), .Y(core__abc_21380_n8841) );
  OR2X2 OR2X2_3275 ( .A(core__abc_21380_n8422), .B(core__abc_21380_n6896), .Y(core__abc_21380_n8842) );
  OR2X2 OR2X2_3276 ( .A(core__abc_21380_n8845), .B(core__abc_21380_n5234), .Y(core__abc_21380_n8846) );
  OR2X2 OR2X2_3277 ( .A(core__abc_21380_n8846), .B(core__abc_21380_n8455_bF_buf1), .Y(core__abc_21380_n8847) );
  OR2X2 OR2X2_3278 ( .A(core__abc_21380_n8844), .B(core__abc_21380_n8847), .Y(core__abc_21380_n8848) );
  OR2X2 OR2X2_3279 ( .A(core__abc_21380_n8454_bF_buf0), .B(core_v1_reg_30_), .Y(core__abc_21380_n8849) );
  OR2X2 OR2X2_328 ( .A(_abc_19068_n1603), .B(_abc_19068_n1604), .Y(_abc_19068_n1605) );
  OR2X2 OR2X2_3280 ( .A(core__abc_21380_n8438), .B(core__abc_21380_n6885), .Y(core__abc_21380_n8852) );
  OR2X2 OR2X2_3281 ( .A(core__abc_21380_n8853), .B(core__abc_21380_n6884), .Y(core__abc_21380_n8854) );
  OR2X2 OR2X2_3282 ( .A(core__abc_21380_n8857), .B(core__abc_21380_n5287), .Y(core__abc_21380_n8858) );
  OR2X2 OR2X2_3283 ( .A(core__abc_21380_n8858), .B(core__abc_21380_n8455_bF_buf0), .Y(core__abc_21380_n8859) );
  OR2X2 OR2X2_3284 ( .A(core__abc_21380_n8856), .B(core__abc_21380_n8859), .Y(core__abc_21380_n8860) );
  OR2X2 OR2X2_3285 ( .A(core__abc_21380_n8454_bF_buf7), .B(core_v1_reg_31_), .Y(core__abc_21380_n8861) );
  OR2X2 OR2X2_3286 ( .A(core__abc_21380_n7073), .B(core__abc_21380_n6877), .Y(core__abc_21380_n8864) );
  OR2X2 OR2X2_3287 ( .A(core__abc_21380_n7072), .B(core__abc_21380_n8865), .Y(core__abc_21380_n8866) );
  OR2X2 OR2X2_3288 ( .A(core__abc_21380_n8869), .B(core__abc_21380_n8871), .Y(core__abc_21380_n8872) );
  OR2X2 OR2X2_3289 ( .A(core__abc_21380_n8872), .B(core__abc_21380_n8455_bF_buf7), .Y(core__abc_21380_n8873) );
  OR2X2 OR2X2_329 ( .A(_abc_19068_n1605), .B(_abc_19068_n1602), .Y(_abc_19068_n1606) );
  OR2X2 OR2X2_3290 ( .A(core__abc_21380_n8868), .B(core__abc_21380_n8873), .Y(core__abc_21380_n8874) );
  OR2X2 OR2X2_3291 ( .A(core__abc_21380_n8454_bF_buf6), .B(core_v1_reg_32_), .Y(core__abc_21380_n8875) );
  OR2X2 OR2X2_3292 ( .A(core__abc_21380_n7105), .B(core__abc_21380_n6849), .Y(core__abc_21380_n8878) );
  OR2X2 OR2X2_3293 ( .A(core__abc_21380_n7104), .B(core__abc_21380_n6848), .Y(core__abc_21380_n8879) );
  OR2X2 OR2X2_3294 ( .A(core__abc_21380_n8882), .B(core__abc_21380_n8883), .Y(core__abc_21380_n8884) );
  OR2X2 OR2X2_3295 ( .A(core__abc_21380_n8884), .B(core__abc_21380_n8455_bF_buf6), .Y(core__abc_21380_n8885) );
  OR2X2 OR2X2_3296 ( .A(core__abc_21380_n8881), .B(core__abc_21380_n8885), .Y(core__abc_21380_n8886) );
  OR2X2 OR2X2_3297 ( .A(core__abc_21380_n8454_bF_buf5), .B(core_v1_reg_33_), .Y(core__abc_21380_n8887) );
  OR2X2 OR2X2_3298 ( .A(core__abc_21380_n7132), .B(core__abc_21380_n6843), .Y(core__abc_21380_n8890) );
  OR2X2 OR2X2_3299 ( .A(core__abc_21380_n7133), .B(core__abc_21380_n6844), .Y(core__abc_21380_n8891) );
  OR2X2 OR2X2_33 ( .A(_abc_19068_n974), .B(_abc_19068_n975_1), .Y(_abc_19068_n976_1) );
  OR2X2 OR2X2_330 ( .A(_abc_19068_n1606), .B(_abc_19068_n1601), .Y(_abc_19068_n1607) );
  OR2X2 OR2X2_3300 ( .A(core__abc_21380_n8894), .B(core__abc_21380_n5453), .Y(core__abc_21380_n8895) );
  OR2X2 OR2X2_3301 ( .A(core__abc_21380_n8895), .B(core__abc_21380_n8455_bF_buf5), .Y(core__abc_21380_n8896) );
  OR2X2 OR2X2_3302 ( .A(core__abc_21380_n8893), .B(core__abc_21380_n8896), .Y(core__abc_21380_n8897) );
  OR2X2 OR2X2_3303 ( .A(core__abc_21380_n8454_bF_buf4), .B(core_v1_reg_34_), .Y(core__abc_21380_n8898) );
  OR2X2 OR2X2_3304 ( .A(core__abc_21380_n7158), .B(core__abc_21380_n6834), .Y(core__abc_21380_n8901) );
  OR2X2 OR2X2_3305 ( .A(core__abc_21380_n7157), .B(core__abc_21380_n6833), .Y(core__abc_21380_n8902) );
  OR2X2 OR2X2_3306 ( .A(core__abc_21380_n8905), .B(core__abc_21380_n5497), .Y(core__abc_21380_n8906) );
  OR2X2 OR2X2_3307 ( .A(core__abc_21380_n8906), .B(core__abc_21380_n8455_bF_buf4), .Y(core__abc_21380_n8907) );
  OR2X2 OR2X2_3308 ( .A(core__abc_21380_n8904), .B(core__abc_21380_n8907), .Y(core__abc_21380_n8908) );
  OR2X2 OR2X2_3309 ( .A(core__abc_21380_n8454_bF_buf3), .B(core_v1_reg_35_), .Y(core__abc_21380_n8909) );
  OR2X2 OR2X2_331 ( .A(_abc_19068_n1609), .B(_abc_19068_n1610), .Y(_abc_19068_n1611) );
  OR2X2 OR2X2_3310 ( .A(core__abc_21380_n7187), .B(core__abc_21380_n6826), .Y(core__abc_21380_n8912) );
  OR2X2 OR2X2_3311 ( .A(core__abc_21380_n8914), .B(core__abc_21380_n8913), .Y(core__abc_21380_n8915) );
  OR2X2 OR2X2_3312 ( .A(core__abc_21380_n8918), .B(core__abc_21380_n5549), .Y(core__abc_21380_n8919) );
  OR2X2 OR2X2_3313 ( .A(core__abc_21380_n8919), .B(core__abc_21380_n8455_bF_buf3), .Y(core__abc_21380_n8920) );
  OR2X2 OR2X2_3314 ( .A(core__abc_21380_n8917), .B(core__abc_21380_n8920), .Y(core__abc_21380_n8921) );
  OR2X2 OR2X2_3315 ( .A(core__abc_21380_n8454_bF_buf2), .B(core_v1_reg_36_), .Y(core__abc_21380_n8922) );
  OR2X2 OR2X2_3316 ( .A(core__abc_21380_n7216), .B(core__abc_21380_n6817), .Y(core__abc_21380_n8925) );
  OR2X2 OR2X2_3317 ( .A(core__abc_21380_n8926), .B(core__abc_21380_n6816), .Y(core__abc_21380_n8927) );
  OR2X2 OR2X2_3318 ( .A(core__abc_21380_n8930), .B(core__abc_21380_n5594), .Y(core__abc_21380_n8931) );
  OR2X2 OR2X2_3319 ( .A(core__abc_21380_n8931), .B(core__abc_21380_n8455_bF_buf2), .Y(core__abc_21380_n8932) );
  OR2X2 OR2X2_332 ( .A(_abc_19068_n1612), .B(_abc_19068_n1613), .Y(_abc_19068_n1614) );
  OR2X2 OR2X2_3320 ( .A(core__abc_21380_n8929), .B(core__abc_21380_n8932), .Y(core__abc_21380_n8933) );
  OR2X2 OR2X2_3321 ( .A(core__abc_21380_n8454_bF_buf1), .B(core_v1_reg_37_), .Y(core__abc_21380_n8934) );
  OR2X2 OR2X2_3322 ( .A(core__abc_21380_n7241), .B(core__abc_21380_n6807), .Y(core__abc_21380_n8937) );
  OR2X2 OR2X2_3323 ( .A(core__abc_21380_n7242), .B(core__abc_21380_n6808), .Y(core__abc_21380_n8938) );
  OR2X2 OR2X2_3324 ( .A(core__abc_21380_n8941), .B(core__abc_21380_n5644), .Y(core__abc_21380_n8942) );
  OR2X2 OR2X2_3325 ( .A(core__abc_21380_n8942), .B(core__abc_21380_n8455_bF_buf1), .Y(core__abc_21380_n8943) );
  OR2X2 OR2X2_3326 ( .A(core__abc_21380_n8940), .B(core__abc_21380_n8943), .Y(core__abc_21380_n8944) );
  OR2X2 OR2X2_3327 ( .A(core__abc_21380_n8454_bF_buf0), .B(core_v1_reg_38_), .Y(core__abc_21380_n8945) );
  OR2X2 OR2X2_3328 ( .A(core__abc_21380_n7267), .B(core__abc_21380_n6798), .Y(core__abc_21380_n8948) );
  OR2X2 OR2X2_3329 ( .A(core__abc_21380_n8949), .B(core__abc_21380_n6797), .Y(core__abc_21380_n8950) );
  OR2X2 OR2X2_333 ( .A(_abc_19068_n1611), .B(_abc_19068_n1614), .Y(_abc_19068_n1615) );
  OR2X2 OR2X2_3330 ( .A(core__abc_21380_n8953), .B(core__abc_21380_n5691), .Y(core__abc_21380_n8954) );
  OR2X2 OR2X2_3331 ( .A(core__abc_21380_n8954), .B(core__abc_21380_n8455_bF_buf0), .Y(core__abc_21380_n8955) );
  OR2X2 OR2X2_3332 ( .A(core__abc_21380_n8952), .B(core__abc_21380_n8955), .Y(core__abc_21380_n8956) );
  OR2X2 OR2X2_3333 ( .A(core__abc_21380_n8454_bF_buf7), .B(core_v1_reg_39_), .Y(core__abc_21380_n8957) );
  OR2X2 OR2X2_3334 ( .A(core__abc_21380_n7307), .B(core__abc_21380_n6792), .Y(core__abc_21380_n8960) );
  OR2X2 OR2X2_3335 ( .A(core__abc_21380_n7306), .B(core__abc_21380_n6788), .Y(core__abc_21380_n8961) );
  OR2X2 OR2X2_3336 ( .A(core__abc_21380_n8964), .B(core__abc_21380_n5740), .Y(core__abc_21380_n8965) );
  OR2X2 OR2X2_3337 ( .A(core__abc_21380_n8965), .B(core__abc_21380_n8455_bF_buf7), .Y(core__abc_21380_n8966) );
  OR2X2 OR2X2_3338 ( .A(core__abc_21380_n8963), .B(core__abc_21380_n8966), .Y(core__abc_21380_n8967) );
  OR2X2 OR2X2_3339 ( .A(core__abc_21380_n8454_bF_buf6), .B(core_v1_reg_40_), .Y(core__abc_21380_n8968) );
  OR2X2 OR2X2_334 ( .A(_abc_19068_n1615), .B(_abc_19068_n1608), .Y(_abc_19068_n1616) );
  OR2X2 OR2X2_3340 ( .A(core__abc_21380_n7334), .B(core__abc_21380_n6752), .Y(core__abc_21380_n8971) );
  OR2X2 OR2X2_3341 ( .A(core__abc_21380_n8972), .B(core__abc_21380_n6751), .Y(core__abc_21380_n8973) );
  OR2X2 OR2X2_3342 ( .A(core__abc_21380_n8976), .B(core__abc_21380_n8978), .Y(core__abc_21380_n8979) );
  OR2X2 OR2X2_3343 ( .A(core__abc_21380_n8979), .B(core__abc_21380_n8455_bF_buf6), .Y(core__abc_21380_n8980) );
  OR2X2 OR2X2_3344 ( .A(core__abc_21380_n8975), .B(core__abc_21380_n8980), .Y(core__abc_21380_n8981) );
  OR2X2 OR2X2_3345 ( .A(core__abc_21380_n8454_bF_buf5), .B(core_v1_reg_41_), .Y(core__abc_21380_n8982) );
  OR2X2 OR2X2_3346 ( .A(core__abc_21380_n7362), .B(core__abc_21380_n6742), .Y(core__abc_21380_n8985) );
  OR2X2 OR2X2_3347 ( .A(core__abc_21380_n7363), .B(core__abc_21380_n6745), .Y(core__abc_21380_n8986) );
  OR2X2 OR2X2_3348 ( .A(core__abc_21380_n8989), .B(core__abc_21380_n8990), .Y(core__abc_21380_n8991) );
  OR2X2 OR2X2_3349 ( .A(core__abc_21380_n8991), .B(core__abc_21380_n8455_bF_buf5), .Y(core__abc_21380_n8992) );
  OR2X2 OR2X2_335 ( .A(_abc_19068_n1616), .B(_abc_19068_n1607), .Y(_abc_19068_n1617) );
  OR2X2 OR2X2_3350 ( .A(core__abc_21380_n8988), .B(core__abc_21380_n8992), .Y(core__abc_21380_n8993) );
  OR2X2 OR2X2_3351 ( .A(core__abc_21380_n8454_bF_buf4), .B(core_v1_reg_42_), .Y(core__abc_21380_n8994) );
  OR2X2 OR2X2_3352 ( .A(core__abc_21380_n7386), .B(core__abc_21380_n6734), .Y(core__abc_21380_n8997) );
  OR2X2 OR2X2_3353 ( .A(core__abc_21380_n7385), .B(core__abc_21380_n6733), .Y(core__abc_21380_n8998) );
  OR2X2 OR2X2_3354 ( .A(core__abc_21380_n9001), .B(core__abc_21380_n5863), .Y(core__abc_21380_n9002) );
  OR2X2 OR2X2_3355 ( .A(core__abc_21380_n9002), .B(core__abc_21380_n8455_bF_buf4), .Y(core__abc_21380_n9003) );
  OR2X2 OR2X2_3356 ( .A(core__abc_21380_n9000), .B(core__abc_21380_n9003), .Y(core__abc_21380_n9004) );
  OR2X2 OR2X2_3357 ( .A(core__abc_21380_n8454_bF_buf3), .B(core_v1_reg_43_), .Y(core__abc_21380_n9005) );
  OR2X2 OR2X2_3358 ( .A(core__abc_21380_n9008), .B(core__abc_21380_n6723), .Y(core__abc_21380_n9009) );
  OR2X2 OR2X2_3359 ( .A(core__abc_21380_n7416), .B(core__abc_21380_n9009), .Y(core__abc_21380_n9010) );
  OR2X2 OR2X2_336 ( .A(_abc_19068_n1621), .B(_abc_19068_n1619), .Y(_abc_19068_n1622) );
  OR2X2 OR2X2_3360 ( .A(core__abc_21380_n7415), .B(core__abc_21380_n6726), .Y(core__abc_21380_n9011) );
  OR2X2 OR2X2_3361 ( .A(core__abc_21380_n9014), .B(core__abc_21380_n9016), .Y(core__abc_21380_n9017) );
  OR2X2 OR2X2_3362 ( .A(core__abc_21380_n9017), .B(core__abc_21380_n8455_bF_buf3), .Y(core__abc_21380_n9018) );
  OR2X2 OR2X2_3363 ( .A(core__abc_21380_n9013), .B(core__abc_21380_n9018), .Y(core__abc_21380_n9019) );
  OR2X2 OR2X2_3364 ( .A(core__abc_21380_n8454_bF_buf2), .B(core_v1_reg_44_), .Y(core__abc_21380_n9020) );
  OR2X2 OR2X2_3365 ( .A(core__abc_21380_n7442), .B(core__abc_21380_n6716), .Y(core__abc_21380_n9023) );
  OR2X2 OR2X2_3366 ( .A(core__abc_21380_n7441), .B(core__abc_21380_n6715), .Y(core__abc_21380_n9024) );
  OR2X2 OR2X2_3367 ( .A(core__abc_21380_n9027), .B(core__abc_21380_n5944), .Y(core__abc_21380_n9028) );
  OR2X2 OR2X2_3368 ( .A(core__abc_21380_n9028), .B(core__abc_21380_n8455_bF_buf2), .Y(core__abc_21380_n9029) );
  OR2X2 OR2X2_3369 ( .A(core__abc_21380_n9026), .B(core__abc_21380_n9029), .Y(core__abc_21380_n9030) );
  OR2X2 OR2X2_337 ( .A(_abc_19068_n1625), .B(_abc_19068_n1624), .Y(_abc_19068_n1626) );
  OR2X2 OR2X2_3370 ( .A(core__abc_21380_n8454_bF_buf1), .B(core_v1_reg_45_), .Y(core__abc_21380_n9031) );
  OR2X2 OR2X2_3371 ( .A(core__abc_21380_n7470), .B(core__abc_21380_n6706), .Y(core__abc_21380_n9034) );
  OR2X2 OR2X2_3372 ( .A(core__abc_21380_n7471), .B(core__abc_21380_n6707), .Y(core__abc_21380_n9035) );
  OR2X2 OR2X2_3373 ( .A(core__abc_21380_n9038), .B(core__abc_21380_n5984), .Y(core__abc_21380_n9039) );
  OR2X2 OR2X2_3374 ( .A(core__abc_21380_n9039), .B(core__abc_21380_n8455_bF_buf1), .Y(core__abc_21380_n9040) );
  OR2X2 OR2X2_3375 ( .A(core__abc_21380_n9037), .B(core__abc_21380_n9040), .Y(core__abc_21380_n9041) );
  OR2X2 OR2X2_3376 ( .A(core__abc_21380_n8454_bF_buf0), .B(core_v1_reg_46_), .Y(core__abc_21380_n9042) );
  OR2X2 OR2X2_3377 ( .A(core__abc_21380_n7495), .B(core__abc_21380_n6697), .Y(core__abc_21380_n9045) );
  OR2X2 OR2X2_3378 ( .A(core__abc_21380_n7494), .B(core__abc_21380_n6696), .Y(core__abc_21380_n9046) );
  OR2X2 OR2X2_3379 ( .A(core__abc_21380_n9049), .B(core__abc_21380_n6018), .Y(core__abc_21380_n9050) );
  OR2X2 OR2X2_338 ( .A(_abc_19068_n1629), .B(_abc_19068_n1628), .Y(_abc_19068_n1630) );
  OR2X2 OR2X2_3380 ( .A(core__abc_21380_n9050), .B(core__abc_21380_n8455_bF_buf0), .Y(core__abc_21380_n9051) );
  OR2X2 OR2X2_3381 ( .A(core__abc_21380_n9048), .B(core__abc_21380_n9051), .Y(core__abc_21380_n9052) );
  OR2X2 OR2X2_3382 ( .A(core__abc_21380_n8454_bF_buf7), .B(core_v1_reg_47_), .Y(core__abc_21380_n9053) );
  OR2X2 OR2X2_3383 ( .A(core__abc_21380_n7536), .B(core__abc_21380_n6691), .Y(core__abc_21380_n9056) );
  OR2X2 OR2X2_3384 ( .A(core__abc_21380_n7535), .B(core__abc_21380_n6688), .Y(core__abc_21380_n9057) );
  OR2X2 OR2X2_3385 ( .A(core__abc_21380_n9060), .B(core__abc_21380_n6082), .Y(core__abc_21380_n9061) );
  OR2X2 OR2X2_3386 ( .A(core__abc_21380_n9061), .B(core__abc_21380_n8455_bF_buf7), .Y(core__abc_21380_n9062) );
  OR2X2 OR2X2_3387 ( .A(core__abc_21380_n9059), .B(core__abc_21380_n9062), .Y(core__abc_21380_n9063) );
  OR2X2 OR2X2_3388 ( .A(core__abc_21380_n8454_bF_buf6), .B(core_v1_reg_48_), .Y(core__abc_21380_n9064) );
  OR2X2 OR2X2_3389 ( .A(core__abc_21380_n7563), .B(core__abc_21380_n7065), .Y(core__abc_21380_n9067) );
  OR2X2 OR2X2_339 ( .A(_abc_19068_n1633), .B(_abc_19068_n1632), .Y(_abc_19068_n1634) );
  OR2X2 OR2X2_3390 ( .A(core__abc_21380_n9068), .B(core__abc_21380_n7064), .Y(core__abc_21380_n9069) );
  OR2X2 OR2X2_3391 ( .A(core__abc_21380_n9072), .B(core__abc_21380_n9074), .Y(core__abc_21380_n9075) );
  OR2X2 OR2X2_3392 ( .A(core__abc_21380_n9075), .B(core__abc_21380_n8455_bF_buf6), .Y(core__abc_21380_n9076) );
  OR2X2 OR2X2_3393 ( .A(core__abc_21380_n9071), .B(core__abc_21380_n9076), .Y(core__abc_21380_n9077) );
  OR2X2 OR2X2_3394 ( .A(core__abc_21380_n8454_bF_buf5), .B(core_v1_reg_49_), .Y(core__abc_21380_n9078) );
  OR2X2 OR2X2_3395 ( .A(core__abc_21380_n7590), .B(core__abc_21380_n7093), .Y(core__abc_21380_n9081) );
  OR2X2 OR2X2_3396 ( .A(core__abc_21380_n7589), .B(core__abc_21380_n7095), .Y(core__abc_21380_n9082) );
  OR2X2 OR2X2_3397 ( .A(core__abc_21380_n9085), .B(core__abc_21380_n6157), .Y(core__abc_21380_n9086) );
  OR2X2 OR2X2_3398 ( .A(core__abc_21380_n9086), .B(core__abc_21380_n8455_bF_buf5), .Y(core__abc_21380_n9087) );
  OR2X2 OR2X2_3399 ( .A(core__abc_21380_n9084), .B(core__abc_21380_n9087), .Y(core__abc_21380_n9088) );
  OR2X2 OR2X2_34 ( .A(_abc_19068_n973_1), .B(_abc_19068_n976_1), .Y(_abc_19068_n977) );
  OR2X2 OR2X2_340 ( .A(_abc_19068_n1637), .B(_abc_19068_n1636), .Y(_abc_19068_n1638) );
  OR2X2 OR2X2_3400 ( .A(core__abc_21380_n8454_bF_buf4), .B(core_v1_reg_50_), .Y(core__abc_21380_n9089) );
  OR2X2 OR2X2_3401 ( .A(core__abc_21380_n7614), .B(core__abc_21380_n7125), .Y(core__abc_21380_n9092) );
  OR2X2 OR2X2_3402 ( .A(core__abc_21380_n9093), .B(core__abc_21380_n7124), .Y(core__abc_21380_n9094) );
  OR2X2 OR2X2_3403 ( .A(core__abc_21380_n9097), .B(core__abc_21380_n9099), .Y(core__abc_21380_n9100) );
  OR2X2 OR2X2_3404 ( .A(core__abc_21380_n9100), .B(core__abc_21380_n8455_bF_buf4), .Y(core__abc_21380_n9101) );
  OR2X2 OR2X2_3405 ( .A(core__abc_21380_n9096), .B(core__abc_21380_n9101), .Y(core__abc_21380_n9102) );
  OR2X2 OR2X2_3406 ( .A(core__abc_21380_n8454_bF_buf3), .B(core_v1_reg_51_), .Y(core__abc_21380_n9103) );
  OR2X2 OR2X2_3407 ( .A(core__abc_21380_n7644), .B(core__abc_21380_n7147), .Y(core__abc_21380_n9106) );
  OR2X2 OR2X2_3408 ( .A(core__abc_21380_n7645), .B(core__abc_21380_n7148), .Y(core__abc_21380_n9107) );
  OR2X2 OR2X2_3409 ( .A(core__abc_21380_n9110), .B(core__abc_21380_n6231), .Y(core__abc_21380_n9111) );
  OR2X2 OR2X2_341 ( .A(_abc_19068_n1641), .B(_abc_19068_n1640), .Y(_abc_19068_n1642) );
  OR2X2 OR2X2_3410 ( .A(core__abc_21380_n9111), .B(core__abc_21380_n8455_bF_buf3), .Y(core__abc_21380_n9112) );
  OR2X2 OR2X2_3411 ( .A(core__abc_21380_n9109), .B(core__abc_21380_n9112), .Y(core__abc_21380_n9113) );
  OR2X2 OR2X2_3412 ( .A(core__abc_21380_n8454_bF_buf2), .B(core_v1_reg_52_), .Y(core__abc_21380_n9114) );
  OR2X2 OR2X2_3413 ( .A(core__abc_21380_n7667), .B(core__abc_21380_n7179), .Y(core__abc_21380_n9117) );
  OR2X2 OR2X2_3414 ( .A(core__abc_21380_n9118), .B(core__abc_21380_n7178), .Y(core__abc_21380_n9119) );
  OR2X2 OR2X2_3415 ( .A(core__abc_21380_n9122), .B(core__abc_21380_n6264), .Y(core__abc_21380_n9123) );
  OR2X2 OR2X2_3416 ( .A(core__abc_21380_n9123), .B(core__abc_21380_n8455_bF_buf2), .Y(core__abc_21380_n9124) );
  OR2X2 OR2X2_3417 ( .A(core__abc_21380_n9121), .B(core__abc_21380_n9124), .Y(core__abc_21380_n9125) );
  OR2X2 OR2X2_3418 ( .A(core__abc_21380_n8454_bF_buf1), .B(core_v1_reg_53_), .Y(core__abc_21380_n9126) );
  OR2X2 OR2X2_3419 ( .A(core__abc_21380_n7694), .B(core__abc_21380_n7206), .Y(core__abc_21380_n9129) );
  OR2X2 OR2X2_342 ( .A(_abc_19068_n1645), .B(_abc_19068_n1644), .Y(_abc_19068_n1646) );
  OR2X2 OR2X2_3420 ( .A(core__abc_21380_n7695), .B(core__abc_21380_n7207), .Y(core__abc_21380_n9130) );
  OR2X2 OR2X2_3421 ( .A(core__abc_21380_n9133), .B(core__abc_21380_n6306), .Y(core__abc_21380_n9134) );
  OR2X2 OR2X2_3422 ( .A(core__abc_21380_n9134), .B(core__abc_21380_n8455_bF_buf1), .Y(core__abc_21380_n9135) );
  OR2X2 OR2X2_3423 ( .A(core__abc_21380_n9132), .B(core__abc_21380_n9135), .Y(core__abc_21380_n9136) );
  OR2X2 OR2X2_3424 ( .A(core__abc_21380_n8454_bF_buf0), .B(core_v1_reg_54_), .Y(core__abc_21380_n9137) );
  OR2X2 OR2X2_3425 ( .A(core__abc_21380_n7721), .B(core__abc_21380_n7231), .Y(core__abc_21380_n9140) );
  OR2X2 OR2X2_3426 ( .A(core__abc_21380_n7720), .B(core__abc_21380_n7230), .Y(core__abc_21380_n9141) );
  OR2X2 OR2X2_3427 ( .A(core__abc_21380_n9144), .B(core__abc_21380_n6340), .Y(core__abc_21380_n9145) );
  OR2X2 OR2X2_3428 ( .A(core__abc_21380_n9145), .B(core__abc_21380_n8455_bF_buf0), .Y(core__abc_21380_n9146) );
  OR2X2 OR2X2_3429 ( .A(core__abc_21380_n9143), .B(core__abc_21380_n9146), .Y(core__abc_21380_n9147) );
  OR2X2 OR2X2_343 ( .A(_abc_19068_n1649), .B(_abc_19068_n1648), .Y(_abc_19068_n1650) );
  OR2X2 OR2X2_3430 ( .A(core__abc_21380_n8454_bF_buf7), .B(core_v1_reg_55_), .Y(core__abc_21380_n9148) );
  OR2X2 OR2X2_3431 ( .A(core__abc_21380_n7757), .B(core__abc_21380_n7259), .Y(core__abc_21380_n9151) );
  OR2X2 OR2X2_3432 ( .A(core__abc_21380_n7758), .B(core__abc_21380_n7260), .Y(core__abc_21380_n9152) );
  OR2X2 OR2X2_3433 ( .A(core__abc_21380_n9155), .B(core__abc_21380_n6400), .Y(core__abc_21380_n9156) );
  OR2X2 OR2X2_3434 ( .A(core__abc_21380_n9156), .B(core__abc_21380_n8455_bF_buf7), .Y(core__abc_21380_n9157) );
  OR2X2 OR2X2_3435 ( .A(core__abc_21380_n9154), .B(core__abc_21380_n9157), .Y(core__abc_21380_n9158) );
  OR2X2 OR2X2_3436 ( .A(core__abc_21380_n8454_bF_buf6), .B(core_v1_reg_56_), .Y(core__abc_21380_n9159) );
  OR2X2 OR2X2_3437 ( .A(core__abc_21380_n7785), .B(core__abc_21380_n7298), .Y(core__abc_21380_n9162) );
  OR2X2 OR2X2_3438 ( .A(core__abc_21380_n7784), .B(core__abc_21380_n7297), .Y(core__abc_21380_n9163) );
  OR2X2 OR2X2_3439 ( .A(core__abc_21380_n9166), .B(core__abc_21380_n6436), .Y(core__abc_21380_n9167) );
  OR2X2 OR2X2_344 ( .A(_abc_19068_n1653), .B(_abc_19068_n1652), .Y(_abc_19068_n1654) );
  OR2X2 OR2X2_3440 ( .A(core__abc_21380_n9167), .B(core__abc_21380_n8455_bF_buf6), .Y(core__abc_21380_n9168) );
  OR2X2 OR2X2_3441 ( .A(core__abc_21380_n9165), .B(core__abc_21380_n9168), .Y(core__abc_21380_n9169) );
  OR2X2 OR2X2_3442 ( .A(core__abc_21380_n8454_bF_buf5), .B(core_v1_reg_57_), .Y(core__abc_21380_n9170) );
  OR2X2 OR2X2_3443 ( .A(core__abc_21380_n7811), .B(core__abc_21380_n7326), .Y(core__abc_21380_n9173) );
  OR2X2 OR2X2_3444 ( .A(core__abc_21380_n7812), .B(core__abc_21380_n7323), .Y(core__abc_21380_n9174) );
  OR2X2 OR2X2_3445 ( .A(core__abc_21380_n9177), .B(core__abc_21380_n6476), .Y(core__abc_21380_n9178) );
  OR2X2 OR2X2_3446 ( .A(core__abc_21380_n9178), .B(core__abc_21380_n8455_bF_buf5), .Y(core__abc_21380_n9179) );
  OR2X2 OR2X2_3447 ( .A(core__abc_21380_n9176), .B(core__abc_21380_n9179), .Y(core__abc_21380_n9180) );
  OR2X2 OR2X2_3448 ( .A(core__abc_21380_n8454_bF_buf4), .B(core_v1_reg_58_), .Y(core__abc_21380_n9181) );
  OR2X2 OR2X2_3449 ( .A(core__abc_21380_n7840), .B(core__abc_21380_n7355), .Y(core__abc_21380_n9184) );
  OR2X2 OR2X2_345 ( .A(_abc_19068_n1657), .B(_abc_19068_n1656), .Y(_abc_19068_n1658) );
  OR2X2 OR2X2_3450 ( .A(core__abc_21380_n7839), .B(core__abc_21380_n7354), .Y(core__abc_21380_n9185) );
  OR2X2 OR2X2_3451 ( .A(core__abc_21380_n9188), .B(core__abc_21380_n6510), .Y(core__abc_21380_n9189) );
  OR2X2 OR2X2_3452 ( .A(core__abc_21380_n9189), .B(core__abc_21380_n8455_bF_buf4), .Y(core__abc_21380_n9190) );
  OR2X2 OR2X2_3453 ( .A(core__abc_21380_n9187), .B(core__abc_21380_n9190), .Y(core__abc_21380_n9191) );
  OR2X2 OR2X2_3454 ( .A(core__abc_21380_n8454_bF_buf3), .B(core_v1_reg_59_), .Y(core__abc_21380_n9192) );
  OR2X2 OR2X2_3455 ( .A(core__abc_21380_n7877), .B(core__abc_21380_n7377), .Y(core__abc_21380_n9195) );
  OR2X2 OR2X2_3456 ( .A(core__abc_21380_n7876), .B(core__abc_21380_n7379), .Y(core__abc_21380_n9196) );
  OR2X2 OR2X2_3457 ( .A(core__abc_21380_n9199), .B(core__abc_21380_n9200), .Y(core__abc_21380_n9201) );
  OR2X2 OR2X2_3458 ( .A(core__abc_21380_n9201), .B(core__abc_21380_n8455_bF_buf3), .Y(core__abc_21380_n9202) );
  OR2X2 OR2X2_3459 ( .A(core__abc_21380_n9198), .B(core__abc_21380_n9202), .Y(core__abc_21380_n9203) );
  OR2X2 OR2X2_346 ( .A(_abc_19068_n1661), .B(_abc_19068_n1660), .Y(_abc_19068_n1662) );
  OR2X2 OR2X2_3460 ( .A(core__abc_21380_n8454_bF_buf2), .B(core_v1_reg_60_), .Y(core__abc_21380_n9204) );
  OR2X2 OR2X2_3461 ( .A(core__abc_21380_n7901), .B(core__abc_21380_n7408), .Y(core__abc_21380_n9207) );
  OR2X2 OR2X2_3462 ( .A(core__abc_21380_n7900), .B(core__abc_21380_n7407), .Y(core__abc_21380_n9208) );
  OR2X2 OR2X2_3463 ( .A(core__abc_21380_n9211), .B(core__abc_21380_n6594), .Y(core__abc_21380_n9212) );
  OR2X2 OR2X2_3464 ( .A(core__abc_21380_n9212), .B(core__abc_21380_n8455_bF_buf2), .Y(core__abc_21380_n9213) );
  OR2X2 OR2X2_3465 ( .A(core__abc_21380_n9210), .B(core__abc_21380_n9213), .Y(core__abc_21380_n9214) );
  OR2X2 OR2X2_3466 ( .A(core__abc_21380_n8454_bF_buf1), .B(core_v1_reg_61_), .Y(core__abc_21380_n9215) );
  OR2X2 OR2X2_3467 ( .A(core__abc_21380_n7931), .B(core__abc_21380_n7429), .Y(core__abc_21380_n9218) );
  OR2X2 OR2X2_3468 ( .A(core__abc_21380_n7932), .B(core__abc_21380_n9219), .Y(core__abc_21380_n9220) );
  OR2X2 OR2X2_3469 ( .A(core__abc_21380_n9223), .B(core__abc_21380_n6636), .Y(core__abc_21380_n9224) );
  OR2X2 OR2X2_347 ( .A(_abc_19068_n1665), .B(_abc_19068_n1664), .Y(_abc_19068_n1666) );
  OR2X2 OR2X2_3470 ( .A(core__abc_21380_n9224), .B(core__abc_21380_n8455_bF_buf1), .Y(core__abc_21380_n9225) );
  OR2X2 OR2X2_3471 ( .A(core__abc_21380_n9222), .B(core__abc_21380_n9225), .Y(core__abc_21380_n9226) );
  OR2X2 OR2X2_3472 ( .A(core__abc_21380_n8454_bF_buf0), .B(core_v1_reg_62_), .Y(core__abc_21380_n9227) );
  OR2X2 OR2X2_3473 ( .A(core__abc_21380_n7930), .B(core__abc_21380_n7923), .Y(core__abc_21380_n9231) );
  OR2X2 OR2X2_3474 ( .A(core__abc_21380_n9232), .B(core__abc_21380_n7954), .Y(core__abc_21380_n9233) );
  OR2X2 OR2X2_3475 ( .A(core__abc_21380_n9230), .B(core__abc_21380_n9234), .Y(core__abc_21380_n9235) );
  OR2X2 OR2X2_3476 ( .A(core__abc_21380_n9237), .B(core__abc_21380_n6672), .Y(core__abc_21380_n9238) );
  OR2X2 OR2X2_3477 ( .A(core__abc_21380_n9238), .B(core__abc_21380_n8455_bF_buf0), .Y(core__abc_21380_n9239) );
  OR2X2 OR2X2_3478 ( .A(core__abc_21380_n9236), .B(core__abc_21380_n9239), .Y(core__abc_21380_n9240) );
  OR2X2 OR2X2_3479 ( .A(core__abc_21380_n8454_bF_buf7), .B(core_v1_reg_63_), .Y(core__abc_21380_n9241) );
  OR2X2 OR2X2_348 ( .A(_abc_19068_n1669), .B(_abc_19068_n1668), .Y(_abc_19068_n1670) );
  OR2X2 OR2X2_3480 ( .A(core__abc_21380_n3167_1_bF_buf12), .B(core__abc_21380_n3312), .Y(core__abc_21380_n9244) );
  OR2X2 OR2X2_3481 ( .A(core_v0_reg_0_), .B(core_mi_reg_0_), .Y(core__abc_21380_n9251) );
  OR2X2 OR2X2_3482 ( .A(core__abc_21380_n9253), .B(core__abc_21380_n7078), .Y(core__abc_21380_n9254) );
  OR2X2 OR2X2_3483 ( .A(core__abc_21380_n9246_bF_buf7), .B(core__abc_21380_n9254), .Y(core__abc_21380_n9255) );
  OR2X2 OR2X2_3484 ( .A(core__abc_21380_n3305), .B(core__abc_21380_n9255), .Y(core__abc_21380_n9256) );
  OR2X2 OR2X2_3485 ( .A(core__abc_21380_n9245_bF_buf6), .B(core_v0_reg_0_), .Y(core__abc_21380_n9257) );
  OR2X2 OR2X2_3486 ( .A(core__abc_21380_n9262), .B(core__abc_21380_n9263), .Y(core__abc_21380_n9264) );
  OR2X2 OR2X2_3487 ( .A(core__abc_21380_n9265), .B(core__abc_21380_n7107), .Y(core__abc_21380_n9266) );
  OR2X2 OR2X2_3488 ( .A(core__abc_21380_n9246_bF_buf6), .B(core__abc_21380_n9266), .Y(core__abc_21380_n9267) );
  OR2X2 OR2X2_3489 ( .A(core__abc_21380_n9260), .B(core__abc_21380_n9267), .Y(core__abc_21380_n9268) );
  OR2X2 OR2X2_349 ( .A(_abc_19068_n1673), .B(_abc_19068_n1672), .Y(_abc_19068_n1674) );
  OR2X2 OR2X2_3490 ( .A(core__abc_21380_n9245_bF_buf5), .B(core_v0_reg_1_), .Y(core__abc_21380_n9269) );
  OR2X2 OR2X2_3491 ( .A(core__abc_21380_n9276), .B(core__abc_21380_n9277), .Y(core__abc_21380_n9278) );
  OR2X2 OR2X2_3492 ( .A(core__abc_21380_n9279), .B(core__abc_21380_n9274), .Y(core__abc_21380_n9280) );
  OR2X2 OR2X2_3493 ( .A(core__abc_21380_n9246_bF_buf5), .B(core__abc_21380_n9280), .Y(core__abc_21380_n9281) );
  OR2X2 OR2X2_3494 ( .A(core__abc_21380_n9272), .B(core__abc_21380_n9281), .Y(core__abc_21380_n9282) );
  OR2X2 OR2X2_3495 ( .A(core__abc_21380_n9245_bF_buf4), .B(core_v0_reg_2_), .Y(core__abc_21380_n9283) );
  OR2X2 OR2X2_3496 ( .A(core__abc_21380_n9288), .B(core__abc_21380_n9289), .Y(core__abc_21380_n9290) );
  OR2X2 OR2X2_3497 ( .A(core__abc_21380_n9291), .B(core__abc_21380_n7160), .Y(core__abc_21380_n9292) );
  OR2X2 OR2X2_3498 ( .A(core__abc_21380_n9246_bF_buf4), .B(core__abc_21380_n9292), .Y(core__abc_21380_n9293) );
  OR2X2 OR2X2_3499 ( .A(core__abc_21380_n9286), .B(core__abc_21380_n9293), .Y(core__abc_21380_n9294) );
  OR2X2 OR2X2_35 ( .A(_abc_19068_n977), .B(_abc_19068_n970_1), .Y(_abc_19068_n978_1) );
  OR2X2 OR2X2_350 ( .A(_abc_19068_n1677), .B(_abc_19068_n1676), .Y(_abc_19068_n1678) );
  OR2X2 OR2X2_3500 ( .A(core__abc_21380_n9245_bF_buf3), .B(core_v0_reg_3_), .Y(core__abc_21380_n9295) );
  OR2X2 OR2X2_3501 ( .A(core_v0_reg_4_), .B(core_mi_reg_4_), .Y(core__abc_21380_n9303) );
  OR2X2 OR2X2_3502 ( .A(core__abc_21380_n9305), .B(core__abc_21380_n9300), .Y(core__abc_21380_n9306) );
  OR2X2 OR2X2_3503 ( .A(core__abc_21380_n9246_bF_buf3), .B(core__abc_21380_n9306), .Y(core__abc_21380_n9307) );
  OR2X2 OR2X2_3504 ( .A(core__abc_21380_n9298), .B(core__abc_21380_n9307), .Y(core__abc_21380_n9308) );
  OR2X2 OR2X2_3505 ( .A(core__abc_21380_n9245_bF_buf2), .B(core_v0_reg_4_), .Y(core__abc_21380_n9309) );
  OR2X2 OR2X2_3506 ( .A(core__abc_21380_n9314), .B(core__abc_21380_n9315), .Y(core__abc_21380_n9316) );
  OR2X2 OR2X2_3507 ( .A(core__abc_21380_n9317), .B(core__abc_21380_n7219), .Y(core__abc_21380_n9318) );
  OR2X2 OR2X2_3508 ( .A(core__abc_21380_n9246_bF_buf2), .B(core__abc_21380_n9318), .Y(core__abc_21380_n9319) );
  OR2X2 OR2X2_3509 ( .A(core__abc_21380_n9312), .B(core__abc_21380_n9319), .Y(core__abc_21380_n9320) );
  OR2X2 OR2X2_351 ( .A(_abc_19068_n1681), .B(_abc_19068_n1680), .Y(_abc_19068_n1682) );
  OR2X2 OR2X2_3510 ( .A(core__abc_21380_n9245_bF_buf1), .B(core_v0_reg_5_), .Y(core__abc_21380_n9321) );
  OR2X2 OR2X2_3511 ( .A(core__abc_21380_n9326), .B(core__abc_21380_n9327), .Y(core__abc_21380_n9328) );
  OR2X2 OR2X2_3512 ( .A(core__abc_21380_n9329), .B(core__abc_21380_n7245), .Y(core__abc_21380_n9330) );
  OR2X2 OR2X2_3513 ( .A(core__abc_21380_n9246_bF_buf1), .B(core__abc_21380_n9330), .Y(core__abc_21380_n9331) );
  OR2X2 OR2X2_3514 ( .A(core__abc_21380_n9324), .B(core__abc_21380_n9331), .Y(core__abc_21380_n9332) );
  OR2X2 OR2X2_3515 ( .A(core__abc_21380_n9245_bF_buf0), .B(core_v0_reg_6_), .Y(core__abc_21380_n9333) );
  OR2X2 OR2X2_3516 ( .A(core__abc_21380_n9338), .B(core__abc_21380_n9339), .Y(core__abc_21380_n9340) );
  OR2X2 OR2X2_3517 ( .A(core__abc_21380_n9341), .B(core__abc_21380_n7269), .Y(core__abc_21380_n9342) );
  OR2X2 OR2X2_3518 ( .A(core__abc_21380_n9246_bF_buf0), .B(core__abc_21380_n9342), .Y(core__abc_21380_n9343) );
  OR2X2 OR2X2_3519 ( .A(core__abc_21380_n9336), .B(core__abc_21380_n9343), .Y(core__abc_21380_n9344) );
  OR2X2 OR2X2_352 ( .A(_abc_19068_n1685), .B(_abc_19068_n1684), .Y(_abc_19068_n1686) );
  OR2X2 OR2X2_3520 ( .A(core__abc_21380_n9245_bF_buf7), .B(core_v0_reg_7_), .Y(core__abc_21380_n9345) );
  OR2X2 OR2X2_3521 ( .A(core_v0_reg_8_), .B(core_mi_reg_8_), .Y(core__abc_21380_n9353) );
  OR2X2 OR2X2_3522 ( .A(core__abc_21380_n9355), .B(core__abc_21380_n9350), .Y(core__abc_21380_n9356) );
  OR2X2 OR2X2_3523 ( .A(core__abc_21380_n9246_bF_buf7), .B(core__abc_21380_n9356), .Y(core__abc_21380_n9357) );
  OR2X2 OR2X2_3524 ( .A(core__abc_21380_n9348), .B(core__abc_21380_n9357), .Y(core__abc_21380_n9358) );
  OR2X2 OR2X2_3525 ( .A(core__abc_21380_n9245_bF_buf6), .B(core_v0_reg_8_), .Y(core__abc_21380_n9359) );
  OR2X2 OR2X2_3526 ( .A(core__abc_21380_n9365), .B(core__abc_21380_n9366), .Y(core__abc_21380_n9367) );
  OR2X2 OR2X2_3527 ( .A(core__abc_21380_n9368), .B(core__abc_21380_n9363), .Y(core__abc_21380_n9369) );
  OR2X2 OR2X2_3528 ( .A(core__abc_21380_n9246_bF_buf6), .B(core__abc_21380_n9369), .Y(core__abc_21380_n9370) );
  OR2X2 OR2X2_3529 ( .A(core__abc_21380_n9362), .B(core__abc_21380_n9370), .Y(core__abc_21380_n9371) );
  OR2X2 OR2X2_353 ( .A(_abc_19068_n1689), .B(_abc_19068_n1688), .Y(_abc_19068_n1690) );
  OR2X2 OR2X2_3530 ( .A(core__abc_21380_n9245_bF_buf5), .B(core_v0_reg_9_), .Y(core__abc_21380_n9372) );
  OR2X2 OR2X2_3531 ( .A(core_v0_reg_10_), .B(core_mi_reg_10_), .Y(core__abc_21380_n9380) );
  OR2X2 OR2X2_3532 ( .A(core__abc_21380_n9382), .B(core__abc_21380_n9377), .Y(core__abc_21380_n9383) );
  OR2X2 OR2X2_3533 ( .A(core__abc_21380_n9246_bF_buf5), .B(core__abc_21380_n9383), .Y(core__abc_21380_n9384) );
  OR2X2 OR2X2_3534 ( .A(core__abc_21380_n9375), .B(core__abc_21380_n9384), .Y(core__abc_21380_n9385) );
  OR2X2 OR2X2_3535 ( .A(core__abc_21380_n9245_bF_buf4), .B(core_v0_reg_10_), .Y(core__abc_21380_n9386) );
  OR2X2 OR2X2_3536 ( .A(core__abc_21380_n9391), .B(core__abc_21380_n9393), .Y(core__abc_21380_n9394) );
  OR2X2 OR2X2_3537 ( .A(core__abc_21380_n9395), .B(core__abc_21380_n7388), .Y(core__abc_21380_n9396) );
  OR2X2 OR2X2_3538 ( .A(core__abc_21380_n9246_bF_buf4), .B(core__abc_21380_n9396), .Y(core__abc_21380_n9397) );
  OR2X2 OR2X2_3539 ( .A(core__abc_21380_n9389), .B(core__abc_21380_n9397), .Y(core__abc_21380_n9398) );
  OR2X2 OR2X2_354 ( .A(_abc_19068_n1693), .B(_abc_19068_n1692), .Y(_abc_19068_n1694) );
  OR2X2 OR2X2_3540 ( .A(core__abc_21380_n9245_bF_buf3), .B(core_v0_reg_11_), .Y(core__abc_21380_n9399) );
  OR2X2 OR2X2_3541 ( .A(core__abc_21380_n9405), .B(core__abc_21380_n9406), .Y(core__abc_21380_n9407) );
  OR2X2 OR2X2_3542 ( .A(core__abc_21380_n9408), .B(core__abc_21380_n9403), .Y(core__abc_21380_n9409) );
  OR2X2 OR2X2_3543 ( .A(core__abc_21380_n9246_bF_buf3), .B(core__abc_21380_n9409), .Y(core__abc_21380_n9410) );
  OR2X2 OR2X2_3544 ( .A(core__abc_21380_n9402), .B(core__abc_21380_n9410), .Y(core__abc_21380_n9411) );
  OR2X2 OR2X2_3545 ( .A(core__abc_21380_n9245_bF_buf2), .B(core_v0_reg_12_), .Y(core__abc_21380_n9412) );
  OR2X2 OR2X2_3546 ( .A(core__abc_21380_n9417), .B(core__abc_21380_n9418), .Y(core__abc_21380_n9419) );
  OR2X2 OR2X2_3547 ( .A(core__abc_21380_n9420), .B(core__abc_21380_n7445), .Y(core__abc_21380_n9421) );
  OR2X2 OR2X2_3548 ( .A(core__abc_21380_n9246_bF_buf2), .B(core__abc_21380_n9421), .Y(core__abc_21380_n9422) );
  OR2X2 OR2X2_3549 ( .A(core__abc_21380_n9415), .B(core__abc_21380_n9422), .Y(core__abc_21380_n9423) );
  OR2X2 OR2X2_355 ( .A(_abc_19068_n1697), .B(_abc_19068_n1696), .Y(_abc_19068_n1698) );
  OR2X2 OR2X2_3550 ( .A(core__abc_21380_n9245_bF_buf1), .B(core_v0_reg_13_), .Y(core__abc_21380_n9424) );
  OR2X2 OR2X2_3551 ( .A(core__abc_21380_n9429), .B(core__abc_21380_n9430), .Y(core__abc_21380_n9431) );
  OR2X2 OR2X2_3552 ( .A(core__abc_21380_n9432), .B(core__abc_21380_n7474), .Y(core__abc_21380_n9433) );
  OR2X2 OR2X2_3553 ( .A(core__abc_21380_n9246_bF_buf1), .B(core__abc_21380_n9433), .Y(core__abc_21380_n9434) );
  OR2X2 OR2X2_3554 ( .A(core__abc_21380_n9427), .B(core__abc_21380_n9434), .Y(core__abc_21380_n9435) );
  OR2X2 OR2X2_3555 ( .A(core__abc_21380_n9245_bF_buf0), .B(core_v0_reg_14_), .Y(core__abc_21380_n9436) );
  OR2X2 OR2X2_3556 ( .A(core__abc_21380_n9441), .B(core__abc_21380_n9442), .Y(core__abc_21380_n9443) );
  OR2X2 OR2X2_3557 ( .A(core__abc_21380_n9444), .B(core__abc_21380_n7497), .Y(core__abc_21380_n9445) );
  OR2X2 OR2X2_3558 ( .A(core__abc_21380_n9246_bF_buf0), .B(core__abc_21380_n9445), .Y(core__abc_21380_n9446) );
  OR2X2 OR2X2_3559 ( .A(core__abc_21380_n9439), .B(core__abc_21380_n9446), .Y(core__abc_21380_n9447) );
  OR2X2 OR2X2_356 ( .A(_abc_19068_n1701), .B(_abc_19068_n1700), .Y(_abc_19068_n1702) );
  OR2X2 OR2X2_3560 ( .A(core__abc_21380_n9245_bF_buf7), .B(core_v0_reg_15_), .Y(core__abc_21380_n9448) );
  OR2X2 OR2X2_3561 ( .A(core__abc_21380_n9453), .B(core__abc_21380_n9454), .Y(core__abc_21380_n9455) );
  OR2X2 OR2X2_3562 ( .A(core__abc_21380_n9456), .B(core__abc_21380_n7539), .Y(core__abc_21380_n9457) );
  OR2X2 OR2X2_3563 ( .A(core__abc_21380_n9246_bF_buf7), .B(core__abc_21380_n9457), .Y(core__abc_21380_n9458) );
  OR2X2 OR2X2_3564 ( .A(core__abc_21380_n9451), .B(core__abc_21380_n9458), .Y(core__abc_21380_n9459) );
  OR2X2 OR2X2_3565 ( .A(core__abc_21380_n9245_bF_buf6), .B(core_v0_reg_16_), .Y(core__abc_21380_n9460) );
  OR2X2 OR2X2_3566 ( .A(core__abc_21380_n9467), .B(core__abc_21380_n9468), .Y(core__abc_21380_n9469) );
  OR2X2 OR2X2_3567 ( .A(core__abc_21380_n9470), .B(core__abc_21380_n9465), .Y(core__abc_21380_n9471) );
  OR2X2 OR2X2_3568 ( .A(core__abc_21380_n9246_bF_buf6), .B(core__abc_21380_n9471), .Y(core__abc_21380_n9472) );
  OR2X2 OR2X2_3569 ( .A(core__abc_21380_n9463), .B(core__abc_21380_n9472), .Y(core__abc_21380_n9473) );
  OR2X2 OR2X2_357 ( .A(_abc_19068_n1705), .B(_abc_19068_n1704), .Y(_abc_19068_n1706) );
  OR2X2 OR2X2_3570 ( .A(core__abc_21380_n9245_bF_buf5), .B(core_v0_reg_17_), .Y(core__abc_21380_n9474) );
  OR2X2 OR2X2_3571 ( .A(core__abc_21380_n9480), .B(core__abc_21380_n9482), .Y(core__abc_21380_n9483) );
  OR2X2 OR2X2_3572 ( .A(core__abc_21380_n9484), .B(core__abc_21380_n9478), .Y(core__abc_21380_n9485) );
  OR2X2 OR2X2_3573 ( .A(core__abc_21380_n9246_bF_buf5), .B(core__abc_21380_n9485), .Y(core__abc_21380_n9486) );
  OR2X2 OR2X2_3574 ( .A(core__abc_21380_n9477), .B(core__abc_21380_n9486), .Y(core__abc_21380_n9487) );
  OR2X2 OR2X2_3575 ( .A(core__abc_21380_n9245_bF_buf4), .B(core_v0_reg_18_), .Y(core__abc_21380_n9488) );
  OR2X2 OR2X2_3576 ( .A(core__abc_21380_n9492), .B(core__abc_21380_n9494), .Y(core__abc_21380_n9495) );
  OR2X2 OR2X2_3577 ( .A(core__abc_21380_n9496), .B(core__abc_21380_n7616), .Y(core__abc_21380_n9497) );
  OR2X2 OR2X2_3578 ( .A(core__abc_21380_n9246_bF_buf4), .B(core__abc_21380_n9497), .Y(core__abc_21380_n9498) );
  OR2X2 OR2X2_3579 ( .A(core__abc_21380_n4617), .B(core__abc_21380_n9498), .Y(core__abc_21380_n9499) );
  OR2X2 OR2X2_358 ( .A(_abc_19068_n1709), .B(_abc_19068_n1708), .Y(_abc_19068_n1710) );
  OR2X2 OR2X2_3580 ( .A(core__abc_21380_n9245_bF_buf3), .B(core_v0_reg_19_), .Y(core__abc_21380_n9500) );
  OR2X2 OR2X2_3581 ( .A(core__abc_21380_n9507), .B(core__abc_21380_n9508), .Y(core__abc_21380_n9509) );
  OR2X2 OR2X2_3582 ( .A(core__abc_21380_n9510), .B(core__abc_21380_n9505), .Y(core__abc_21380_n9511) );
  OR2X2 OR2X2_3583 ( .A(core__abc_21380_n9246_bF_buf3), .B(core__abc_21380_n9511), .Y(core__abc_21380_n9512) );
  OR2X2 OR2X2_3584 ( .A(core__abc_21380_n9503), .B(core__abc_21380_n9512), .Y(core__abc_21380_n9513) );
  OR2X2 OR2X2_3585 ( .A(core__abc_21380_n9245_bF_buf2), .B(core_v0_reg_20_), .Y(core__abc_21380_n9514) );
  OR2X2 OR2X2_3586 ( .A(core__abc_21380_n9519), .B(core__abc_21380_n9520), .Y(core__abc_21380_n9521) );
  OR2X2 OR2X2_3587 ( .A(core__abc_21380_n9522), .B(core__abc_21380_n7670), .Y(core__abc_21380_n9523) );
  OR2X2 OR2X2_3588 ( .A(core__abc_21380_n9246_bF_buf2), .B(core__abc_21380_n9523), .Y(core__abc_21380_n9524) );
  OR2X2 OR2X2_3589 ( .A(core__abc_21380_n9517), .B(core__abc_21380_n9524), .Y(core__abc_21380_n9525) );
  OR2X2 OR2X2_359 ( .A(_abc_19068_n1713), .B(_abc_19068_n1712), .Y(_abc_19068_n1714) );
  OR2X2 OR2X2_3590 ( .A(core__abc_21380_n9245_bF_buf1), .B(core_v0_reg_21_), .Y(core__abc_21380_n9526) );
  OR2X2 OR2X2_3591 ( .A(core__abc_21380_n9531), .B(core__abc_21380_n9532), .Y(core__abc_21380_n9533) );
  OR2X2 OR2X2_3592 ( .A(core__abc_21380_n9534), .B(core__abc_21380_n7698), .Y(core__abc_21380_n9535) );
  OR2X2 OR2X2_3593 ( .A(core__abc_21380_n9246_bF_buf1), .B(core__abc_21380_n9535), .Y(core__abc_21380_n9536) );
  OR2X2 OR2X2_3594 ( .A(core__abc_21380_n9529), .B(core__abc_21380_n9536), .Y(core__abc_21380_n9537) );
  OR2X2 OR2X2_3595 ( .A(core__abc_21380_n9245_bF_buf0), .B(core_v0_reg_22_), .Y(core__abc_21380_n9538) );
  OR2X2 OR2X2_3596 ( .A(core__abc_21380_n9543), .B(core__abc_21380_n9544), .Y(core__abc_21380_n9545) );
  OR2X2 OR2X2_3597 ( .A(core__abc_21380_n9546), .B(core__abc_21380_n7723), .Y(core__abc_21380_n9547) );
  OR2X2 OR2X2_3598 ( .A(core__abc_21380_n9246_bF_buf0), .B(core__abc_21380_n9547), .Y(core__abc_21380_n9548) );
  OR2X2 OR2X2_3599 ( .A(core__abc_21380_n9541), .B(core__abc_21380_n9548), .Y(core__abc_21380_n9549) );
  OR2X2 OR2X2_36 ( .A(_abc_19068_n967_1), .B(_abc_19068_n978_1), .Y(_abc_19068_n979_1) );
  OR2X2 OR2X2_360 ( .A(_abc_19068_n1717), .B(_abc_19068_n1716), .Y(_abc_19068_n1718) );
  OR2X2 OR2X2_3600 ( .A(core__abc_21380_n9245_bF_buf7), .B(core_v0_reg_23_), .Y(core__abc_21380_n9550) );
  OR2X2 OR2X2_3601 ( .A(core__abc_21380_n9555), .B(core__abc_21380_n9556), .Y(core__abc_21380_n9557) );
  OR2X2 OR2X2_3602 ( .A(core__abc_21380_n9558), .B(core__abc_21380_n7760), .Y(core__abc_21380_n9559) );
  OR2X2 OR2X2_3603 ( .A(core__abc_21380_n9246_bF_buf7), .B(core__abc_21380_n9559), .Y(core__abc_21380_n9560) );
  OR2X2 OR2X2_3604 ( .A(core__abc_21380_n9553), .B(core__abc_21380_n9560), .Y(core__abc_21380_n9561) );
  OR2X2 OR2X2_3605 ( .A(core__abc_21380_n9245_bF_buf6), .B(core_v0_reg_24_), .Y(core__abc_21380_n9562) );
  OR2X2 OR2X2_3606 ( .A(core__abc_21380_n9568), .B(core__abc_21380_n9569), .Y(core__abc_21380_n9570) );
  OR2X2 OR2X2_3607 ( .A(core__abc_21380_n9571), .B(core__abc_21380_n9566), .Y(core__abc_21380_n9572) );
  OR2X2 OR2X2_3608 ( .A(core__abc_21380_n9246_bF_buf6), .B(core__abc_21380_n9572), .Y(core__abc_21380_n9573) );
  OR2X2 OR2X2_3609 ( .A(core__abc_21380_n9565), .B(core__abc_21380_n9573), .Y(core__abc_21380_n9574) );
  OR2X2 OR2X2_361 ( .A(_abc_19068_n1721), .B(_abc_19068_n1720), .Y(_abc_19068_n1722) );
  OR2X2 OR2X2_3610 ( .A(core__abc_21380_n9245_bF_buf5), .B(core_v0_reg_25_), .Y(core__abc_21380_n9575) );
  OR2X2 OR2X2_3611 ( .A(core_v0_reg_26_), .B(core_mi_reg_26_), .Y(core__abc_21380_n9582) );
  OR2X2 OR2X2_3612 ( .A(core__abc_21380_n9584), .B(core__abc_21380_n9579), .Y(core__abc_21380_n9585) );
  OR2X2 OR2X2_3613 ( .A(core__abc_21380_n9246_bF_buf5), .B(core__abc_21380_n9585), .Y(core__abc_21380_n9586) );
  OR2X2 OR2X2_3614 ( .A(core__abc_21380_n9578), .B(core__abc_21380_n9586), .Y(core__abc_21380_n9587) );
  OR2X2 OR2X2_3615 ( .A(core__abc_21380_n9245_bF_buf4), .B(core_v0_reg_26_), .Y(core__abc_21380_n9588) );
  OR2X2 OR2X2_3616 ( .A(core__abc_21380_n9594), .B(core__abc_21380_n9595), .Y(core__abc_21380_n9596) );
  OR2X2 OR2X2_3617 ( .A(core__abc_21380_n9597), .B(core__abc_21380_n9592), .Y(core__abc_21380_n9598) );
  OR2X2 OR2X2_3618 ( .A(core__abc_21380_n9246_bF_buf4), .B(core__abc_21380_n9598), .Y(core__abc_21380_n9599) );
  OR2X2 OR2X2_3619 ( .A(core__abc_21380_n9591), .B(core__abc_21380_n9599), .Y(core__abc_21380_n9600) );
  OR2X2 OR2X2_362 ( .A(_abc_19068_n1725), .B(_abc_19068_n1724), .Y(_abc_19068_n1726) );
  OR2X2 OR2X2_3620 ( .A(core__abc_21380_n9245_bF_buf3), .B(core_v0_reg_27_), .Y(core__abc_21380_n9601) );
  OR2X2 OR2X2_3621 ( .A(core__abc_21380_n9608), .B(core__abc_21380_n9609), .Y(core__abc_21380_n9610) );
  OR2X2 OR2X2_3622 ( .A(core__abc_21380_n9611), .B(core__abc_21380_n9606), .Y(core__abc_21380_n9612) );
  OR2X2 OR2X2_3623 ( .A(core__abc_21380_n9246_bF_buf3), .B(core__abc_21380_n9612), .Y(core__abc_21380_n9613) );
  OR2X2 OR2X2_3624 ( .A(core__abc_21380_n9604), .B(core__abc_21380_n9613), .Y(core__abc_21380_n9614) );
  OR2X2 OR2X2_3625 ( .A(core__abc_21380_n9245_bF_buf2), .B(core_v0_reg_28_), .Y(core__abc_21380_n9615) );
  OR2X2 OR2X2_3626 ( .A(core__abc_21380_n9620), .B(core__abc_21380_n9621), .Y(core__abc_21380_n9622) );
  OR2X2 OR2X2_3627 ( .A(core__abc_21380_n9623), .B(core__abc_21380_n7904), .Y(core__abc_21380_n9624) );
  OR2X2 OR2X2_3628 ( .A(core__abc_21380_n9246_bF_buf2), .B(core__abc_21380_n9624), .Y(core__abc_21380_n9625) );
  OR2X2 OR2X2_3629 ( .A(core__abc_21380_n9618), .B(core__abc_21380_n9625), .Y(core__abc_21380_n9626) );
  OR2X2 OR2X2_363 ( .A(_abc_19068_n1729), .B(_abc_19068_n1728), .Y(_abc_19068_n1730) );
  OR2X2 OR2X2_3630 ( .A(core__abc_21380_n9245_bF_buf1), .B(core_v0_reg_29_), .Y(core__abc_21380_n9627) );
  OR2X2 OR2X2_3631 ( .A(core__abc_21380_n9632), .B(core__abc_21380_n9633), .Y(core__abc_21380_n9634) );
  OR2X2 OR2X2_3632 ( .A(core__abc_21380_n9635), .B(core__abc_21380_n7935), .Y(core__abc_21380_n9636) );
  OR2X2 OR2X2_3633 ( .A(core__abc_21380_n9246_bF_buf1), .B(core__abc_21380_n9636), .Y(core__abc_21380_n9637) );
  OR2X2 OR2X2_3634 ( .A(core__abc_21380_n9630), .B(core__abc_21380_n9637), .Y(core__abc_21380_n9638) );
  OR2X2 OR2X2_3635 ( .A(core__abc_21380_n9245_bF_buf0), .B(core_v0_reg_30_), .Y(core__abc_21380_n9639) );
  OR2X2 OR2X2_3636 ( .A(core__abc_21380_n9644), .B(core__abc_21380_n9645), .Y(core__abc_21380_n9646) );
  OR2X2 OR2X2_3637 ( .A(core__abc_21380_n9647), .B(core__abc_21380_n7959), .Y(core__abc_21380_n9648) );
  OR2X2 OR2X2_3638 ( .A(core__abc_21380_n9246_bF_buf0), .B(core__abc_21380_n9648), .Y(core__abc_21380_n9649) );
  OR2X2 OR2X2_3639 ( .A(core__abc_21380_n9642), .B(core__abc_21380_n9649), .Y(core__abc_21380_n9650) );
  OR2X2 OR2X2_364 ( .A(_abc_19068_n1733), .B(_abc_19068_n1732), .Y(_abc_19068_n1734) );
  OR2X2 OR2X2_3640 ( .A(core__abc_21380_n9245_bF_buf7), .B(core_v0_reg_31_), .Y(core__abc_21380_n9651) );
  OR2X2 OR2X2_3641 ( .A(core__abc_21380_n9656), .B(core__abc_21380_n9657), .Y(core__abc_21380_n9658) );
  OR2X2 OR2X2_3642 ( .A(core__abc_21380_n9659), .B(core__abc_21380_n7968), .Y(core__abc_21380_n9660) );
  OR2X2 OR2X2_3643 ( .A(core__abc_21380_n9246_bF_buf7), .B(core__abc_21380_n9660), .Y(core__abc_21380_n9661) );
  OR2X2 OR2X2_3644 ( .A(core__abc_21380_n9654), .B(core__abc_21380_n9661), .Y(core__abc_21380_n9662) );
  OR2X2 OR2X2_3645 ( .A(core__abc_21380_n9245_bF_buf6), .B(core_v0_reg_32_), .Y(core__abc_21380_n9663) );
  OR2X2 OR2X2_3646 ( .A(core__abc_21380_n9668), .B(core__abc_21380_n9669), .Y(core__abc_21380_n9670) );
  OR2X2 OR2X2_3647 ( .A(core__abc_21380_n9671), .B(core__abc_21380_n7984), .Y(core__abc_21380_n9672) );
  OR2X2 OR2X2_3648 ( .A(core__abc_21380_n9246_bF_buf6), .B(core__abc_21380_n9672), .Y(core__abc_21380_n9673) );
  OR2X2 OR2X2_3649 ( .A(core__abc_21380_n9666), .B(core__abc_21380_n9673), .Y(core__abc_21380_n9674) );
  OR2X2 OR2X2_365 ( .A(_abc_19068_n1737), .B(_abc_19068_n1736), .Y(_abc_19068_n1738) );
  OR2X2 OR2X2_3650 ( .A(core__abc_21380_n9245_bF_buf5), .B(core_v0_reg_33_), .Y(core__abc_21380_n9675) );
  OR2X2 OR2X2_3651 ( .A(core__abc_21380_n9680), .B(core__abc_21380_n9681), .Y(core__abc_21380_n9682) );
  OR2X2 OR2X2_3652 ( .A(core__abc_21380_n9683), .B(core__abc_21380_n7996), .Y(core__abc_21380_n9684) );
  OR2X2 OR2X2_3653 ( .A(core__abc_21380_n9246_bF_buf5), .B(core__abc_21380_n9684), .Y(core__abc_21380_n9685) );
  OR2X2 OR2X2_3654 ( .A(core__abc_21380_n9678), .B(core__abc_21380_n9685), .Y(core__abc_21380_n9686) );
  OR2X2 OR2X2_3655 ( .A(core__abc_21380_n9245_bF_buf4), .B(core_v0_reg_34_), .Y(core__abc_21380_n9687) );
  OR2X2 OR2X2_3656 ( .A(core__abc_21380_n9692), .B(core__abc_21380_n9693), .Y(core__abc_21380_n9694) );
  OR2X2 OR2X2_3657 ( .A(core__abc_21380_n9695), .B(core__abc_21380_n8005), .Y(core__abc_21380_n9696) );
  OR2X2 OR2X2_3658 ( .A(core__abc_21380_n9246_bF_buf4), .B(core__abc_21380_n9696), .Y(core__abc_21380_n9697) );
  OR2X2 OR2X2_3659 ( .A(core__abc_21380_n9690), .B(core__abc_21380_n9697), .Y(core__abc_21380_n9698) );
  OR2X2 OR2X2_366 ( .A(_abc_19068_n1741), .B(_abc_19068_n1740), .Y(_abc_19068_n1742) );
  OR2X2 OR2X2_3660 ( .A(core__abc_21380_n9245_bF_buf3), .B(core_v0_reg_35_), .Y(core__abc_21380_n9699) );
  OR2X2 OR2X2_3661 ( .A(core__abc_21380_n9704), .B(core__abc_21380_n9705), .Y(core__abc_21380_n9706) );
  OR2X2 OR2X2_3662 ( .A(core__abc_21380_n9707), .B(core__abc_21380_n8017), .Y(core__abc_21380_n9708) );
  OR2X2 OR2X2_3663 ( .A(core__abc_21380_n9246_bF_buf3), .B(core__abc_21380_n9708), .Y(core__abc_21380_n9709) );
  OR2X2 OR2X2_3664 ( .A(core__abc_21380_n9702), .B(core__abc_21380_n9709), .Y(core__abc_21380_n9710) );
  OR2X2 OR2X2_3665 ( .A(core__abc_21380_n9245_bF_buf2), .B(core_v0_reg_36_), .Y(core__abc_21380_n9711) );
  OR2X2 OR2X2_3666 ( .A(core__abc_21380_n9716), .B(core__abc_21380_n9717), .Y(core__abc_21380_n9718) );
  OR2X2 OR2X2_3667 ( .A(core__abc_21380_n9719), .B(core__abc_21380_n8030), .Y(core__abc_21380_n9720) );
  OR2X2 OR2X2_3668 ( .A(core__abc_21380_n9246_bF_buf2), .B(core__abc_21380_n9720), .Y(core__abc_21380_n9721) );
  OR2X2 OR2X2_3669 ( .A(core__abc_21380_n9714), .B(core__abc_21380_n9721), .Y(core__abc_21380_n9722) );
  OR2X2 OR2X2_367 ( .A(_abc_19068_n1745), .B(_abc_19068_n1744), .Y(_abc_19068_n1746) );
  OR2X2 OR2X2_3670 ( .A(core__abc_21380_n9245_bF_buf1), .B(core_v0_reg_37_), .Y(core__abc_21380_n9723) );
  OR2X2 OR2X2_3671 ( .A(core__abc_21380_n9728), .B(core__abc_21380_n9729), .Y(core__abc_21380_n9730) );
  OR2X2 OR2X2_3672 ( .A(core__abc_21380_n9731), .B(core__abc_21380_n8044), .Y(core__abc_21380_n9732) );
  OR2X2 OR2X2_3673 ( .A(core__abc_21380_n9246_bF_buf1), .B(core__abc_21380_n9732), .Y(core__abc_21380_n9733) );
  OR2X2 OR2X2_3674 ( .A(core__abc_21380_n9726), .B(core__abc_21380_n9733), .Y(core__abc_21380_n9734) );
  OR2X2 OR2X2_3675 ( .A(core__abc_21380_n9245_bF_buf0), .B(core_v0_reg_38_), .Y(core__abc_21380_n9735) );
  OR2X2 OR2X2_3676 ( .A(core__abc_21380_n9740), .B(core__abc_21380_n9741), .Y(core__abc_21380_n9742) );
  OR2X2 OR2X2_3677 ( .A(core__abc_21380_n9743), .B(core__abc_21380_n8059), .Y(core__abc_21380_n9744) );
  OR2X2 OR2X2_3678 ( .A(core__abc_21380_n9246_bF_buf0), .B(core__abc_21380_n9744), .Y(core__abc_21380_n9745) );
  OR2X2 OR2X2_3679 ( .A(core__abc_21380_n9738), .B(core__abc_21380_n9745), .Y(core__abc_21380_n9746) );
  OR2X2 OR2X2_368 ( .A(_abc_19068_n1749), .B(_abc_19068_n1748), .Y(_abc_19068_n1750) );
  OR2X2 OR2X2_3680 ( .A(core__abc_21380_n9245_bF_buf7), .B(core_v0_reg_39_), .Y(core__abc_21380_n9747) );
  OR2X2 OR2X2_3681 ( .A(core__abc_21380_n9752), .B(core__abc_21380_n9753), .Y(core__abc_21380_n9754) );
  OR2X2 OR2X2_3682 ( .A(core__abc_21380_n9755), .B(core__abc_21380_n8074), .Y(core__abc_21380_n9756) );
  OR2X2 OR2X2_3683 ( .A(core__abc_21380_n9246_bF_buf7), .B(core__abc_21380_n9756), .Y(core__abc_21380_n9757) );
  OR2X2 OR2X2_3684 ( .A(core__abc_21380_n9750), .B(core__abc_21380_n9757), .Y(core__abc_21380_n9758) );
  OR2X2 OR2X2_3685 ( .A(core__abc_21380_n9245_bF_buf6), .B(core_v0_reg_40_), .Y(core__abc_21380_n9759) );
  OR2X2 OR2X2_3686 ( .A(core__abc_21380_n9765), .B(core__abc_21380_n9766), .Y(core__abc_21380_n9767) );
  OR2X2 OR2X2_3687 ( .A(core__abc_21380_n9768), .B(core__abc_21380_n9763), .Y(core__abc_21380_n9769) );
  OR2X2 OR2X2_3688 ( .A(core__abc_21380_n9246_bF_buf6), .B(core__abc_21380_n9769), .Y(core__abc_21380_n9770) );
  OR2X2 OR2X2_3689 ( .A(core__abc_21380_n9762), .B(core__abc_21380_n9770), .Y(core__abc_21380_n9771) );
  OR2X2 OR2X2_369 ( .A(_abc_19068_n1753), .B(_abc_19068_n1752), .Y(_abc_19068_n1754) );
  OR2X2 OR2X2_3690 ( .A(core__abc_21380_n9245_bF_buf5), .B(core_v0_reg_41_), .Y(core__abc_21380_n9772) );
  OR2X2 OR2X2_3691 ( .A(core__abc_21380_n9777), .B(core__abc_21380_n9778), .Y(core__abc_21380_n9779) );
  OR2X2 OR2X2_3692 ( .A(core__abc_21380_n9780), .B(core__abc_21380_n8107), .Y(core__abc_21380_n9781) );
  OR2X2 OR2X2_3693 ( .A(core__abc_21380_n9246_bF_buf5), .B(core__abc_21380_n9781), .Y(core__abc_21380_n9782) );
  OR2X2 OR2X2_3694 ( .A(core__abc_21380_n9775), .B(core__abc_21380_n9782), .Y(core__abc_21380_n9783) );
  OR2X2 OR2X2_3695 ( .A(core__abc_21380_n9245_bF_buf4), .B(core_v0_reg_42_), .Y(core__abc_21380_n9784) );
  OR2X2 OR2X2_3696 ( .A(core__abc_21380_n9791), .B(core__abc_21380_n9792), .Y(core__abc_21380_n9793) );
  OR2X2 OR2X2_3697 ( .A(core__abc_21380_n9794), .B(core__abc_21380_n9789), .Y(core__abc_21380_n9795) );
  OR2X2 OR2X2_3698 ( .A(core__abc_21380_n9246_bF_buf4), .B(core__abc_21380_n9795), .Y(core__abc_21380_n9796) );
  OR2X2 OR2X2_3699 ( .A(core__abc_21380_n9787), .B(core__abc_21380_n9796), .Y(core__abc_21380_n9797) );
  OR2X2 OR2X2_37 ( .A(_abc_19068_n982_1), .B(_abc_19068_n983), .Y(_abc_19068_n984_1) );
  OR2X2 OR2X2_370 ( .A(_abc_19068_n1757), .B(_abc_19068_n1756), .Y(_abc_19068_n1758) );
  OR2X2 OR2X2_3700 ( .A(core__abc_21380_n9245_bF_buf3), .B(core_v0_reg_43_), .Y(core__abc_21380_n9798) );
  OR2X2 OR2X2_3701 ( .A(core__abc_21380_n9803), .B(core__abc_21380_n9804), .Y(core__abc_21380_n9805) );
  OR2X2 OR2X2_3702 ( .A(core__abc_21380_n9806), .B(core__abc_21380_n8136), .Y(core__abc_21380_n9807) );
  OR2X2 OR2X2_3703 ( .A(core__abc_21380_n9246_bF_buf3), .B(core__abc_21380_n9807), .Y(core__abc_21380_n9808) );
  OR2X2 OR2X2_3704 ( .A(core__abc_21380_n9801), .B(core__abc_21380_n9808), .Y(core__abc_21380_n9809) );
  OR2X2 OR2X2_3705 ( .A(core__abc_21380_n9245_bF_buf2), .B(core_v0_reg_44_), .Y(core__abc_21380_n9810) );
  OR2X2 OR2X2_3706 ( .A(core__abc_21380_n9815), .B(core__abc_21380_n9816), .Y(core__abc_21380_n9817) );
  OR2X2 OR2X2_3707 ( .A(core__abc_21380_n9818), .B(core__abc_21380_n8153), .Y(core__abc_21380_n9819) );
  OR2X2 OR2X2_3708 ( .A(core__abc_21380_n9246_bF_buf2), .B(core__abc_21380_n9819), .Y(core__abc_21380_n9820) );
  OR2X2 OR2X2_3709 ( .A(core__abc_21380_n9813), .B(core__abc_21380_n9820), .Y(core__abc_21380_n9821) );
  OR2X2 OR2X2_371 ( .A(_abc_19068_n1761), .B(_abc_19068_n1760), .Y(_abc_19068_n1762) );
  OR2X2 OR2X2_3710 ( .A(core__abc_21380_n9245_bF_buf1), .B(core_v0_reg_45_), .Y(core__abc_21380_n9822) );
  OR2X2 OR2X2_3711 ( .A(core__abc_21380_n9827), .B(core__abc_21380_n9828), .Y(core__abc_21380_n9829) );
  OR2X2 OR2X2_3712 ( .A(core__abc_21380_n9830), .B(core__abc_21380_n8169), .Y(core__abc_21380_n9831) );
  OR2X2 OR2X2_3713 ( .A(core__abc_21380_n9246_bF_buf1), .B(core__abc_21380_n9831), .Y(core__abc_21380_n9832) );
  OR2X2 OR2X2_3714 ( .A(core__abc_21380_n9825), .B(core__abc_21380_n9832), .Y(core__abc_21380_n9833) );
  OR2X2 OR2X2_3715 ( .A(core__abc_21380_n9245_bF_buf0), .B(core_v0_reg_46_), .Y(core__abc_21380_n9834) );
  OR2X2 OR2X2_3716 ( .A(core__abc_21380_n9839), .B(core__abc_21380_n9840), .Y(core__abc_21380_n9841) );
  OR2X2 OR2X2_3717 ( .A(core__abc_21380_n9842), .B(core__abc_21380_n8185), .Y(core__abc_21380_n9843) );
  OR2X2 OR2X2_3718 ( .A(core__abc_21380_n9246_bF_buf0), .B(core__abc_21380_n9843), .Y(core__abc_21380_n9844) );
  OR2X2 OR2X2_3719 ( .A(core__abc_21380_n9837), .B(core__abc_21380_n9844), .Y(core__abc_21380_n9845) );
  OR2X2 OR2X2_372 ( .A(_abc_19068_n1765), .B(_abc_19068_n1764), .Y(_abc_19068_n1766) );
  OR2X2 OR2X2_3720 ( .A(core__abc_21380_n9245_bF_buf7), .B(core_v0_reg_47_), .Y(core__abc_21380_n9846) );
  OR2X2 OR2X2_3721 ( .A(core__abc_21380_n9851), .B(core__abc_21380_n9852), .Y(core__abc_21380_n9853) );
  OR2X2 OR2X2_3722 ( .A(core__abc_21380_n9854), .B(core__abc_21380_n8200), .Y(core__abc_21380_n9855) );
  OR2X2 OR2X2_3723 ( .A(core__abc_21380_n9246_bF_buf7), .B(core__abc_21380_n9855), .Y(core__abc_21380_n9856) );
  OR2X2 OR2X2_3724 ( .A(core__abc_21380_n9849), .B(core__abc_21380_n9856), .Y(core__abc_21380_n9857) );
  OR2X2 OR2X2_3725 ( .A(core__abc_21380_n9245_bF_buf6), .B(core_v0_reg_48_), .Y(core__abc_21380_n9858) );
  OR2X2 OR2X2_3726 ( .A(core__abc_21380_n9865), .B(core__abc_21380_n9866), .Y(core__abc_21380_n9867) );
  OR2X2 OR2X2_3727 ( .A(core__abc_21380_n9868), .B(core__abc_21380_n9863), .Y(core__abc_21380_n9869) );
  OR2X2 OR2X2_3728 ( .A(core__abc_21380_n9246_bF_buf6), .B(core__abc_21380_n9869), .Y(core__abc_21380_n9870) );
  OR2X2 OR2X2_3729 ( .A(core__abc_21380_n9861), .B(core__abc_21380_n9870), .Y(core__abc_21380_n9871) );
  OR2X2 OR2X2_373 ( .A(_abc_19068_n1769), .B(_abc_19068_n1768), .Y(_abc_19068_n1770) );
  OR2X2 OR2X2_3730 ( .A(core__abc_21380_n9245_bF_buf5), .B(core_v0_reg_49_), .Y(core__abc_21380_n9872) );
  OR2X2 OR2X2_3731 ( .A(core__abc_21380_n9879), .B(core__abc_21380_n9880), .Y(core__abc_21380_n9881) );
  OR2X2 OR2X2_3732 ( .A(core__abc_21380_n9882), .B(core__abc_21380_n9877), .Y(core__abc_21380_n9883) );
  OR2X2 OR2X2_3733 ( .A(core__abc_21380_n9246_bF_buf5), .B(core__abc_21380_n9883), .Y(core__abc_21380_n9884) );
  OR2X2 OR2X2_3734 ( .A(core__abc_21380_n9875), .B(core__abc_21380_n9884), .Y(core__abc_21380_n9885) );
  OR2X2 OR2X2_3735 ( .A(core__abc_21380_n9245_bF_buf4), .B(core_v0_reg_50_), .Y(core__abc_21380_n9886) );
  OR2X2 OR2X2_3736 ( .A(core__abc_21380_n9891), .B(core__abc_21380_n9892), .Y(core__abc_21380_n9893) );
  OR2X2 OR2X2_3737 ( .A(core__abc_21380_n9894), .B(core__abc_21380_n8248), .Y(core__abc_21380_n9895) );
  OR2X2 OR2X2_3738 ( .A(core__abc_21380_n9246_bF_buf4), .B(core__abc_21380_n9895), .Y(core__abc_21380_n9896) );
  OR2X2 OR2X2_3739 ( .A(core__abc_21380_n9889), .B(core__abc_21380_n9896), .Y(core__abc_21380_n9897) );
  OR2X2 OR2X2_374 ( .A(_abc_19068_n1773), .B(_abc_19068_n1772), .Y(_abc_19068_n1774) );
  OR2X2 OR2X2_3740 ( .A(core__abc_21380_n9245_bF_buf3), .B(core_v0_reg_51_), .Y(core__abc_21380_n9898) );
  OR2X2 OR2X2_3741 ( .A(core_v0_reg_52_), .B(core_mi_reg_52_), .Y(core__abc_21380_n9905) );
  OR2X2 OR2X2_3742 ( .A(core__abc_21380_n9907), .B(core__abc_21380_n9902), .Y(core__abc_21380_n9908) );
  OR2X2 OR2X2_3743 ( .A(core__abc_21380_n9246_bF_buf3), .B(core__abc_21380_n9908), .Y(core__abc_21380_n9909) );
  OR2X2 OR2X2_3744 ( .A(core__abc_21380_n9901), .B(core__abc_21380_n9909), .Y(core__abc_21380_n9910) );
  OR2X2 OR2X2_3745 ( .A(core__abc_21380_n9245_bF_buf2), .B(core_v0_reg_52_), .Y(core__abc_21380_n9911) );
  OR2X2 OR2X2_3746 ( .A(core__abc_21380_n9916), .B(core__abc_21380_n9917), .Y(core__abc_21380_n9918) );
  OR2X2 OR2X2_3747 ( .A(core__abc_21380_n9919), .B(core__abc_21380_n8280), .Y(core__abc_21380_n9920) );
  OR2X2 OR2X2_3748 ( .A(core__abc_21380_n9246_bF_buf2), .B(core__abc_21380_n9920), .Y(core__abc_21380_n9921) );
  OR2X2 OR2X2_3749 ( .A(core__abc_21380_n9914), .B(core__abc_21380_n9921), .Y(core__abc_21380_n9922) );
  OR2X2 OR2X2_375 ( .A(_abc_19068_n1777), .B(_abc_19068_n1776), .Y(_abc_19068_n1778) );
  OR2X2 OR2X2_3750 ( .A(core__abc_21380_n9245_bF_buf1), .B(core_v0_reg_53_), .Y(core__abc_21380_n9923) );
  OR2X2 OR2X2_3751 ( .A(core__abc_21380_n9928), .B(core__abc_21380_n9929), .Y(core__abc_21380_n9930) );
  OR2X2 OR2X2_3752 ( .A(core__abc_21380_n9931), .B(core__abc_21380_n8297), .Y(core__abc_21380_n9932) );
  OR2X2 OR2X2_3753 ( .A(core__abc_21380_n9246_bF_buf1), .B(core__abc_21380_n9932), .Y(core__abc_21380_n9933) );
  OR2X2 OR2X2_3754 ( .A(core__abc_21380_n9926), .B(core__abc_21380_n9933), .Y(core__abc_21380_n9934) );
  OR2X2 OR2X2_3755 ( .A(core__abc_21380_n9245_bF_buf0), .B(core_v0_reg_54_), .Y(core__abc_21380_n9935) );
  OR2X2 OR2X2_3756 ( .A(core__abc_21380_n9940), .B(core__abc_21380_n9941), .Y(core__abc_21380_n9942) );
  OR2X2 OR2X2_3757 ( .A(core__abc_21380_n9943), .B(core__abc_21380_n8312), .Y(core__abc_21380_n9944) );
  OR2X2 OR2X2_3758 ( .A(core__abc_21380_n9246_bF_buf0), .B(core__abc_21380_n9944), .Y(core__abc_21380_n9945) );
  OR2X2 OR2X2_3759 ( .A(core__abc_21380_n9938), .B(core__abc_21380_n9945), .Y(core__abc_21380_n9946) );
  OR2X2 OR2X2_376 ( .A(_abc_19068_n1781), .B(_abc_19068_n1780), .Y(_abc_19068_n1782) );
  OR2X2 OR2X2_3760 ( .A(core__abc_21380_n9245_bF_buf7), .B(core_v0_reg_55_), .Y(core__abc_21380_n9947) );
  OR2X2 OR2X2_3761 ( .A(core__abc_21380_n9952), .B(core__abc_21380_n9953), .Y(core__abc_21380_n9954) );
  OR2X2 OR2X2_3762 ( .A(core__abc_21380_n9955), .B(core__abc_21380_n9957), .Y(core__abc_21380_n9958) );
  OR2X2 OR2X2_3763 ( .A(core__abc_21380_n9246_bF_buf7), .B(core__abc_21380_n9958), .Y(core__abc_21380_n9959) );
  OR2X2 OR2X2_3764 ( .A(core__abc_21380_n9950), .B(core__abc_21380_n9959), .Y(core__abc_21380_n9960) );
  OR2X2 OR2X2_3765 ( .A(core__abc_21380_n9245_bF_buf6), .B(core_v0_reg_56_), .Y(core__abc_21380_n9961) );
  OR2X2 OR2X2_3766 ( .A(core__abc_21380_n9968), .B(core__abc_21380_n9969), .Y(core__abc_21380_n9970) );
  OR2X2 OR2X2_3767 ( .A(core__abc_21380_n9971), .B(core__abc_21380_n9966), .Y(core__abc_21380_n9972) );
  OR2X2 OR2X2_3768 ( .A(core__abc_21380_n9246_bF_buf6), .B(core__abc_21380_n9972), .Y(core__abc_21380_n9973) );
  OR2X2 OR2X2_3769 ( .A(core__abc_21380_n9964), .B(core__abc_21380_n9973), .Y(core__abc_21380_n9974) );
  OR2X2 OR2X2_377 ( .A(_abc_19068_n1785), .B(_abc_19068_n1784), .Y(_abc_19068_n1786) );
  OR2X2 OR2X2_3770 ( .A(core__abc_21380_n9245_bF_buf5), .B(core_v0_reg_57_), .Y(core__abc_21380_n9975) );
  OR2X2 OR2X2_3771 ( .A(core__abc_21380_n9981), .B(core__abc_21380_n9982), .Y(core__abc_21380_n9983) );
  OR2X2 OR2X2_3772 ( .A(core__abc_21380_n9984), .B(core__abc_21380_n9979), .Y(core__abc_21380_n9985) );
  OR2X2 OR2X2_3773 ( .A(core__abc_21380_n9246_bF_buf5), .B(core__abc_21380_n9985), .Y(core__abc_21380_n9986) );
  OR2X2 OR2X2_3774 ( .A(core__abc_21380_n9978), .B(core__abc_21380_n9986), .Y(core__abc_21380_n9987) );
  OR2X2 OR2X2_3775 ( .A(core__abc_21380_n9245_bF_buf4), .B(core_v0_reg_58_), .Y(core__abc_21380_n9988) );
  OR2X2 OR2X2_3776 ( .A(core__abc_21380_n9994), .B(core__abc_21380_n9995), .Y(core__abc_21380_n9996) );
  OR2X2 OR2X2_3777 ( .A(core__abc_21380_n9997), .B(core__abc_21380_n9992), .Y(core__abc_21380_n9998) );
  OR2X2 OR2X2_3778 ( .A(core__abc_21380_n9246_bF_buf4), .B(core__abc_21380_n9998), .Y(core__abc_21380_n9999) );
  OR2X2 OR2X2_3779 ( .A(core__abc_21380_n9991), .B(core__abc_21380_n9999), .Y(core__abc_21380_n10000) );
  OR2X2 OR2X2_378 ( .A(_abc_19068_n1789), .B(_abc_19068_n1788), .Y(_abc_19068_n1790) );
  OR2X2 OR2X2_3780 ( .A(core__abc_21380_n9245_bF_buf3), .B(core_v0_reg_59_), .Y(core__abc_21380_n10001) );
  OR2X2 OR2X2_3781 ( .A(core__abc_21380_n10008), .B(core__abc_21380_n10009), .Y(core__abc_21380_n10010) );
  OR2X2 OR2X2_3782 ( .A(core__abc_21380_n10011), .B(core__abc_21380_n10006), .Y(core__abc_21380_n10012) );
  OR2X2 OR2X2_3783 ( .A(core__abc_21380_n9246_bF_buf3), .B(core__abc_21380_n10012), .Y(core__abc_21380_n10013) );
  OR2X2 OR2X2_3784 ( .A(core__abc_21380_n10004), .B(core__abc_21380_n10013), .Y(core__abc_21380_n10014) );
  OR2X2 OR2X2_3785 ( .A(core__abc_21380_n9245_bF_buf2), .B(core_v0_reg_60_), .Y(core__abc_21380_n10015) );
  OR2X2 OR2X2_3786 ( .A(core__abc_21380_n10020), .B(core__abc_21380_n10021), .Y(core__abc_21380_n10022) );
  OR2X2 OR2X2_3787 ( .A(core__abc_21380_n10023), .B(core__abc_21380_n8408), .Y(core__abc_21380_n10024) );
  OR2X2 OR2X2_3788 ( .A(core__abc_21380_n9246_bF_buf2), .B(core__abc_21380_n10024), .Y(core__abc_21380_n10025) );
  OR2X2 OR2X2_3789 ( .A(core__abc_21380_n10018), .B(core__abc_21380_n10025), .Y(core__abc_21380_n10026) );
  OR2X2 OR2X2_379 ( .A(_abc_19068_n1793), .B(_abc_19068_n1792), .Y(_abc_19068_n1794) );
  OR2X2 OR2X2_3790 ( .A(core__abc_21380_n9245_bF_buf1), .B(core_v0_reg_61_), .Y(core__abc_21380_n10027) );
  OR2X2 OR2X2_3791 ( .A(core__abc_21380_n10032), .B(core__abc_21380_n10033), .Y(core__abc_21380_n10034) );
  OR2X2 OR2X2_3792 ( .A(core__abc_21380_n10035), .B(core__abc_21380_n8425), .Y(core__abc_21380_n10036) );
  OR2X2 OR2X2_3793 ( .A(core__abc_21380_n9246_bF_buf1), .B(core__abc_21380_n10036), .Y(core__abc_21380_n10037) );
  OR2X2 OR2X2_3794 ( .A(core__abc_21380_n10030), .B(core__abc_21380_n10037), .Y(core__abc_21380_n10038) );
  OR2X2 OR2X2_3795 ( .A(core__abc_21380_n9245_bF_buf0), .B(core_v0_reg_62_), .Y(core__abc_21380_n10039) );
  OR2X2 OR2X2_3796 ( .A(core__abc_21380_n10044), .B(core__abc_21380_n10045), .Y(core__abc_21380_n10046) );
  OR2X2 OR2X2_3797 ( .A(core__abc_21380_n10047), .B(core__abc_21380_n8440), .Y(core__abc_21380_n10048) );
  OR2X2 OR2X2_3798 ( .A(core__abc_21380_n9246_bF_buf0), .B(core__abc_21380_n10048), .Y(core__abc_21380_n10049) );
  OR2X2 OR2X2_3799 ( .A(core__abc_21380_n10042), .B(core__abc_21380_n10049), .Y(core__abc_21380_n10050) );
  OR2X2 OR2X2_38 ( .A(_abc_19068_n985_1), .B(_abc_19068_n986), .Y(_abc_19068_n987_1) );
  OR2X2 OR2X2_380 ( .A(_abc_19068_n1797), .B(_abc_19068_n1796), .Y(_abc_19068_n1798) );
  OR2X2 OR2X2_3800 ( .A(core__abc_21380_n9245_bF_buf7), .B(core_v0_reg_63_), .Y(core__abc_21380_n10051) );
  OR2X2 OR2X2_3801 ( .A(core__abc_21380_n10061), .B(core__abc_21380_n1144_1), .Y(core__abc_21380_n10062) );
  OR2X2 OR2X2_3802 ( .A(core__abc_21380_n10063), .B(core__abc_21380_n1241_1), .Y(core__abc_21380_n10064) );
  OR2X2 OR2X2_381 ( .A(_abc_19068_n1801), .B(_abc_19068_n1800), .Y(_abc_19068_n1802) );
  OR2X2 OR2X2_382 ( .A(_abc_19068_n1805), .B(_abc_19068_n1804), .Y(_abc_19068_n1806) );
  OR2X2 OR2X2_383 ( .A(_abc_19068_n1809), .B(_abc_19068_n1808), .Y(_abc_19068_n1810) );
  OR2X2 OR2X2_384 ( .A(_abc_19068_n1813), .B(_abc_19068_n1812), .Y(_abc_19068_n1814) );
  OR2X2 OR2X2_385 ( .A(_abc_19068_n1817), .B(_abc_19068_n1816), .Y(_abc_19068_n1818) );
  OR2X2 OR2X2_386 ( .A(_abc_19068_n1821), .B(_abc_19068_n1820), .Y(_abc_19068_n1822) );
  OR2X2 OR2X2_387 ( .A(_abc_19068_n1825), .B(_abc_19068_n1824), .Y(_abc_19068_n1826) );
  OR2X2 OR2X2_388 ( .A(_abc_19068_n1829), .B(_abc_19068_n1828), .Y(_abc_19068_n1830) );
  OR2X2 OR2X2_389 ( .A(_abc_19068_n1833), .B(_abc_19068_n1832), .Y(_abc_19068_n1834) );
  OR2X2 OR2X2_39 ( .A(_abc_19068_n984_1), .B(_abc_19068_n987_1), .Y(_abc_19068_n988_1) );
  OR2X2 OR2X2_390 ( .A(_abc_19068_n1837), .B(_abc_19068_n1836), .Y(_abc_19068_n1838) );
  OR2X2 OR2X2_391 ( .A(_abc_19068_n1841), .B(_abc_19068_n1840), .Y(_abc_19068_n1842) );
  OR2X2 OR2X2_392 ( .A(_abc_19068_n1845), .B(_abc_19068_n1844), .Y(_abc_19068_n1846) );
  OR2X2 OR2X2_393 ( .A(_abc_19068_n1849), .B(_abc_19068_n1848), .Y(_abc_19068_n1850) );
  OR2X2 OR2X2_394 ( .A(_abc_19068_n1853), .B(_abc_19068_n1852), .Y(_abc_19068_n1854) );
  OR2X2 OR2X2_395 ( .A(_abc_19068_n1857), .B(_abc_19068_n1856), .Y(_abc_19068_n1858) );
  OR2X2 OR2X2_396 ( .A(_abc_19068_n1861), .B(_abc_19068_n1860), .Y(_abc_19068_n1862) );
  OR2X2 OR2X2_397 ( .A(_abc_19068_n1865), .B(_abc_19068_n1864), .Y(_abc_19068_n1866) );
  OR2X2 OR2X2_398 ( .A(_abc_19068_n1869), .B(_abc_19068_n1868), .Y(_abc_19068_n1870) );
  OR2X2 OR2X2_399 ( .A(_abc_19068_n1873), .B(_abc_19068_n1872), .Y(_abc_19068_n1874) );
  OR2X2 OR2X2_4 ( .A(_abc_19068_n903_1), .B(_abc_19068_n897_1_bF_buf4), .Y(_abc_19068_n904_1) );
  OR2X2 OR2X2_40 ( .A(_abc_19068_n988_1), .B(_abc_19068_n981_1), .Y(_abc_19068_n989) );
  OR2X2 OR2X2_400 ( .A(_abc_19068_n1877), .B(_abc_19068_n1876), .Y(_abc_19068_n1878) );
  OR2X2 OR2X2_401 ( .A(_abc_19068_n1881), .B(_abc_19068_n1880), .Y(_abc_19068_n1882) );
  OR2X2 OR2X2_402 ( .A(_abc_19068_n1885), .B(_abc_19068_n1884), .Y(_abc_19068_n1886) );
  OR2X2 OR2X2_403 ( .A(_abc_19068_n1889), .B(_abc_19068_n1888), .Y(_abc_19068_n1890) );
  OR2X2 OR2X2_404 ( .A(_abc_19068_n1893), .B(_abc_19068_n1892), .Y(_abc_19068_n1894) );
  OR2X2 OR2X2_405 ( .A(_abc_19068_n1897), .B(_abc_19068_n1896), .Y(_abc_19068_n1898) );
  OR2X2 OR2X2_406 ( .A(_abc_19068_n1901), .B(_abc_19068_n1900), .Y(_abc_19068_n1902) );
  OR2X2 OR2X2_407 ( .A(_abc_19068_n1905), .B(_abc_19068_n1904), .Y(_abc_19068_n1906) );
  OR2X2 OR2X2_408 ( .A(_abc_19068_n1909), .B(_abc_19068_n1908), .Y(_abc_19068_n1910) );
  OR2X2 OR2X2_409 ( .A(_abc_19068_n1913), .B(_abc_19068_n1912), .Y(_abc_19068_n1914) );
  OR2X2 OR2X2_41 ( .A(_abc_19068_n991_1), .B(_abc_19068_n992), .Y(_abc_19068_n993_1) );
  OR2X2 OR2X2_410 ( .A(_abc_19068_n1917), .B(_abc_19068_n1916), .Y(_abc_19068_n1918) );
  OR2X2 OR2X2_411 ( .A(_abc_19068_n1921), .B(_abc_19068_n1920), .Y(_abc_19068_n1922) );
  OR2X2 OR2X2_412 ( .A(_abc_19068_n1925), .B(_abc_19068_n1924), .Y(_abc_19068_n1926) );
  OR2X2 OR2X2_413 ( .A(_abc_19068_n1929), .B(_abc_19068_n1928), .Y(_abc_19068_n1930) );
  OR2X2 OR2X2_414 ( .A(_abc_19068_n1933), .B(_abc_19068_n1932), .Y(_abc_19068_n1934) );
  OR2X2 OR2X2_415 ( .A(_abc_19068_n1937), .B(_abc_19068_n1936), .Y(_abc_19068_n1938) );
  OR2X2 OR2X2_416 ( .A(_abc_19068_n1941), .B(_abc_19068_n1940), .Y(_abc_19068_n1942) );
  OR2X2 OR2X2_417 ( .A(_abc_19068_n1945), .B(_abc_19068_n1944), .Y(_abc_19068_n1946) );
  OR2X2 OR2X2_418 ( .A(_abc_19068_n1949), .B(_abc_19068_n1948), .Y(_abc_19068_n1950) );
  OR2X2 OR2X2_419 ( .A(_abc_19068_n1953), .B(_abc_19068_n1952), .Y(_abc_19068_n1954) );
  OR2X2 OR2X2_42 ( .A(_abc_19068_n993_1), .B(_abc_19068_n990_1), .Y(_abc_19068_n994_1) );
  OR2X2 OR2X2_420 ( .A(_abc_19068_n1957), .B(_abc_19068_n1956), .Y(_abc_19068_n1958) );
  OR2X2 OR2X2_421 ( .A(_abc_19068_n1961), .B(_abc_19068_n1960), .Y(_abc_19068_n1962) );
  OR2X2 OR2X2_422 ( .A(_abc_19068_n1965), .B(_abc_19068_n1964), .Y(_abc_19068_n1966) );
  OR2X2 OR2X2_423 ( .A(_abc_19068_n1969), .B(_abc_19068_n1968), .Y(_abc_19068_n1970) );
  OR2X2 OR2X2_424 ( .A(_abc_19068_n1973), .B(_abc_19068_n1972), .Y(_abc_19068_n1974) );
  OR2X2 OR2X2_425 ( .A(_abc_19068_n1977), .B(_abc_19068_n1976), .Y(_abc_19068_n1978) );
  OR2X2 OR2X2_426 ( .A(_abc_19068_n1981), .B(_abc_19068_n1980), .Y(_abc_19068_n1982) );
  OR2X2 OR2X2_427 ( .A(_abc_19068_n1985), .B(_abc_19068_n1984), .Y(_abc_19068_n1986) );
  OR2X2 OR2X2_428 ( .A(_abc_19068_n1989), .B(_abc_19068_n1988), .Y(_abc_19068_n1990) );
  OR2X2 OR2X2_429 ( .A(_abc_19068_n1993), .B(_abc_19068_n1992), .Y(_abc_19068_n1994) );
  OR2X2 OR2X2_43 ( .A(_abc_19068_n995), .B(_abc_19068_n996_1), .Y(_abc_19068_n997_1) );
  OR2X2 OR2X2_430 ( .A(_abc_19068_n1997), .B(_abc_19068_n1996), .Y(_abc_19068_n1998) );
  OR2X2 OR2X2_431 ( .A(_abc_19068_n2001), .B(_abc_19068_n2000), .Y(_abc_19068_n2002) );
  OR2X2 OR2X2_432 ( .A(_abc_19068_n2005), .B(_abc_19068_n2004), .Y(_abc_19068_n2006) );
  OR2X2 OR2X2_433 ( .A(_abc_19068_n2009), .B(_abc_19068_n2008), .Y(_abc_19068_n2010) );
  OR2X2 OR2X2_434 ( .A(_abc_19068_n2013), .B(_abc_19068_n2012), .Y(_abc_19068_n2014) );
  OR2X2 OR2X2_435 ( .A(_abc_19068_n2017), .B(_abc_19068_n2016), .Y(_abc_19068_n2018) );
  OR2X2 OR2X2_436 ( .A(_abc_19068_n2021), .B(_abc_19068_n2020), .Y(_abc_19068_n2022) );
  OR2X2 OR2X2_437 ( .A(_abc_19068_n2025), .B(_abc_19068_n2024), .Y(_abc_19068_n2026) );
  OR2X2 OR2X2_438 ( .A(_abc_19068_n2029), .B(_abc_19068_n2028), .Y(_abc_19068_n2030) );
  OR2X2 OR2X2_439 ( .A(_abc_19068_n2033), .B(_abc_19068_n2032), .Y(_abc_19068_n2034) );
  OR2X2 OR2X2_44 ( .A(_abc_19068_n998), .B(_abc_19068_n999_1), .Y(_abc_19068_n1000_1) );
  OR2X2 OR2X2_440 ( .A(_abc_19068_n2037), .B(_abc_19068_n2036), .Y(_abc_19068_n2038) );
  OR2X2 OR2X2_441 ( .A(_abc_19068_n2041), .B(_abc_19068_n2040), .Y(_abc_19068_n2042) );
  OR2X2 OR2X2_442 ( .A(_abc_19068_n2045), .B(_abc_19068_n2044), .Y(_abc_19068_n2046) );
  OR2X2 OR2X2_443 ( .A(_abc_19068_n2049), .B(_abc_19068_n2048), .Y(_abc_19068_n2050) );
  OR2X2 OR2X2_444 ( .A(_abc_19068_n2053), .B(_abc_19068_n2052), .Y(_abc_19068_n2054) );
  OR2X2 OR2X2_445 ( .A(_abc_19068_n2057), .B(_abc_19068_n2056), .Y(_abc_19068_n2058) );
  OR2X2 OR2X2_446 ( .A(_abc_19068_n2061), .B(_abc_19068_n2060), .Y(_abc_19068_n2062) );
  OR2X2 OR2X2_447 ( .A(_abc_19068_n2065), .B(_abc_19068_n2064), .Y(_abc_19068_n2066) );
  OR2X2 OR2X2_448 ( .A(_abc_19068_n2069), .B(_abc_19068_n2068), .Y(_abc_19068_n2070) );
  OR2X2 OR2X2_449 ( .A(_abc_19068_n2073), .B(_abc_19068_n2072), .Y(_abc_19068_n2074) );
  OR2X2 OR2X2_45 ( .A(_abc_19068_n997_1), .B(_abc_19068_n1000_1), .Y(_abc_19068_n1001) );
  OR2X2 OR2X2_450 ( .A(_abc_19068_n2077), .B(_abc_19068_n2076), .Y(_abc_19068_n2078) );
  OR2X2 OR2X2_451 ( .A(_abc_19068_n2081), .B(_abc_19068_n2080), .Y(_abc_19068_n2082) );
  OR2X2 OR2X2_452 ( .A(_abc_19068_n2085), .B(_abc_19068_n2084), .Y(_abc_19068_n2086) );
  OR2X2 OR2X2_453 ( .A(_abc_19068_n2089), .B(_abc_19068_n2088), .Y(_abc_19068_n2090) );
  OR2X2 OR2X2_454 ( .A(_abc_19068_n2093), .B(_abc_19068_n2092), .Y(_abc_19068_n2094) );
  OR2X2 OR2X2_455 ( .A(_abc_19068_n2097), .B(_abc_19068_n2096), .Y(_abc_19068_n2098) );
  OR2X2 OR2X2_456 ( .A(_abc_19068_n2101), .B(_abc_19068_n2100), .Y(_abc_19068_n2102) );
  OR2X2 OR2X2_457 ( .A(_abc_19068_n2105), .B(_abc_19068_n2104), .Y(_abc_19068_n2106) );
  OR2X2 OR2X2_458 ( .A(_abc_19068_n2109), .B(_abc_19068_n2108), .Y(_abc_19068_n2110) );
  OR2X2 OR2X2_459 ( .A(_abc_19068_n2113), .B(_abc_19068_n2112), .Y(_abc_19068_n2114) );
  OR2X2 OR2X2_46 ( .A(_abc_19068_n1001), .B(_abc_19068_n994_1), .Y(_abc_19068_n1002_1) );
  OR2X2 OR2X2_460 ( .A(_abc_19068_n2117), .B(_abc_19068_n2116), .Y(_abc_19068_n2118) );
  OR2X2 OR2X2_461 ( .A(_abc_19068_n2121), .B(_abc_19068_n2120), .Y(_abc_19068_n2122) );
  OR2X2 OR2X2_462 ( .A(_abc_19068_n2125), .B(_abc_19068_n2124), .Y(_abc_19068_n2126) );
  OR2X2 OR2X2_463 ( .A(_abc_19068_n2129), .B(_abc_19068_n2128), .Y(_abc_19068_n2130) );
  OR2X2 OR2X2_464 ( .A(_abc_19068_n2133_bF_buf7), .B(core_mi_32_), .Y(_abc_19068_n2134) );
  OR2X2 OR2X2_465 ( .A(_abc_19068_n2133_bF_buf5), .B(core_mi_33_), .Y(_abc_19068_n2140) );
  OR2X2 OR2X2_466 ( .A(_abc_19068_n2133_bF_buf3), .B(core_mi_34_), .Y(_abc_19068_n2146) );
  OR2X2 OR2X2_467 ( .A(_abc_19068_n2133_bF_buf1), .B(core_mi_35_), .Y(_abc_19068_n2152) );
  OR2X2 OR2X2_468 ( .A(_abc_19068_n2133_bF_buf7), .B(core_mi_36_), .Y(_abc_19068_n2158) );
  OR2X2 OR2X2_469 ( .A(_abc_19068_n2133_bF_buf5), .B(core_mi_37_), .Y(_abc_19068_n2164) );
  OR2X2 OR2X2_47 ( .A(_abc_19068_n989), .B(_abc_19068_n1002_1), .Y(_abc_19068_n1003_1) );
  OR2X2 OR2X2_470 ( .A(_abc_19068_n2133_bF_buf3), .B(core_mi_38_), .Y(_abc_19068_n2170) );
  OR2X2 OR2X2_471 ( .A(_abc_19068_n2133_bF_buf1), .B(core_mi_39_), .Y(_abc_19068_n2176) );
  OR2X2 OR2X2_472 ( .A(_abc_19068_n2133_bF_buf7), .B(core_mi_40_), .Y(_abc_19068_n2182) );
  OR2X2 OR2X2_473 ( .A(_abc_19068_n2133_bF_buf5), .B(core_mi_41_), .Y(_abc_19068_n2188) );
  OR2X2 OR2X2_474 ( .A(_abc_19068_n2133_bF_buf3), .B(core_mi_42_), .Y(_abc_19068_n2194) );
  OR2X2 OR2X2_475 ( .A(_abc_19068_n2133_bF_buf1), .B(core_mi_43_), .Y(_abc_19068_n2200) );
  OR2X2 OR2X2_476 ( .A(_abc_19068_n2133_bF_buf7), .B(core_mi_44_), .Y(_abc_19068_n2206) );
  OR2X2 OR2X2_477 ( .A(_abc_19068_n2133_bF_buf5), .B(core_mi_45_), .Y(_abc_19068_n2212) );
  OR2X2 OR2X2_478 ( .A(_abc_19068_n2133_bF_buf3), .B(core_mi_46_), .Y(_abc_19068_n2218) );
  OR2X2 OR2X2_479 ( .A(_abc_19068_n2133_bF_buf1), .B(core_mi_47_), .Y(_abc_19068_n2224) );
  OR2X2 OR2X2_48 ( .A(_abc_19068_n1005_1), .B(_abc_19068_n1006_1), .Y(_abc_19068_n1007) );
  OR2X2 OR2X2_480 ( .A(_abc_19068_n2133_bF_buf7), .B(core_mi_48_), .Y(_abc_19068_n2230) );
  OR2X2 OR2X2_481 ( .A(_abc_19068_n2133_bF_buf5), .B(core_mi_49_), .Y(_abc_19068_n2236) );
  OR2X2 OR2X2_482 ( .A(_abc_19068_n2133_bF_buf3), .B(core_mi_50_), .Y(_abc_19068_n2242) );
  OR2X2 OR2X2_483 ( .A(_abc_19068_n2133_bF_buf1), .B(core_mi_51_), .Y(_abc_19068_n2248) );
  OR2X2 OR2X2_484 ( .A(_abc_19068_n2133_bF_buf7), .B(core_mi_52_), .Y(_abc_19068_n2254) );
  OR2X2 OR2X2_485 ( .A(_abc_19068_n2133_bF_buf5), .B(core_mi_53_), .Y(_abc_19068_n2260) );
  OR2X2 OR2X2_486 ( .A(_abc_19068_n2133_bF_buf3), .B(core_mi_54_), .Y(_abc_19068_n2266) );
  OR2X2 OR2X2_487 ( .A(_abc_19068_n2133_bF_buf1), .B(core_mi_55_), .Y(_abc_19068_n2272) );
  OR2X2 OR2X2_488 ( .A(_abc_19068_n2133_bF_buf7), .B(core_mi_56_), .Y(_abc_19068_n2278) );
  OR2X2 OR2X2_489 ( .A(_abc_19068_n2133_bF_buf5), .B(core_mi_57_), .Y(_abc_19068_n2284) );
  OR2X2 OR2X2_49 ( .A(_abc_19068_n1008_1), .B(_abc_19068_n1009_1), .Y(_abc_19068_n1010) );
  OR2X2 OR2X2_490 ( .A(_abc_19068_n2133_bF_buf3), .B(core_mi_58_), .Y(_abc_19068_n2290) );
  OR2X2 OR2X2_491 ( .A(_abc_19068_n2133_bF_buf1), .B(core_mi_59_), .Y(_abc_19068_n2296) );
  OR2X2 OR2X2_492 ( .A(_abc_19068_n2133_bF_buf7), .B(core_mi_60_), .Y(_abc_19068_n2302) );
  OR2X2 OR2X2_493 ( .A(_abc_19068_n2133_bF_buf5), .B(core_mi_61_), .Y(_abc_19068_n2308) );
  OR2X2 OR2X2_494 ( .A(_abc_19068_n2133_bF_buf3), .B(core_mi_62_), .Y(_abc_19068_n2314) );
  OR2X2 OR2X2_495 ( .A(_abc_19068_n2133_bF_buf1), .B(core_mi_63_), .Y(_abc_19068_n2320) );
  OR2X2 OR2X2_496 ( .A(_abc_19068_n2326_bF_buf7), .B(core_mi_0_), .Y(_abc_19068_n2327) );
  OR2X2 OR2X2_497 ( .A(_abc_19068_n2326_bF_buf5), .B(core_mi_1_), .Y(_abc_19068_n2332) );
  OR2X2 OR2X2_498 ( .A(_abc_19068_n2326_bF_buf3), .B(core_mi_2_), .Y(_abc_19068_n2337) );
  OR2X2 OR2X2_499 ( .A(_abc_19068_n2326_bF_buf1), .B(core_mi_3_), .Y(_abc_19068_n2342) );
  OR2X2 OR2X2_5 ( .A(_abc_19068_n891_1), .B(_abc_19068_n904_1), .Y(_abc_19068_n905) );
  OR2X2 OR2X2_50 ( .A(_abc_19068_n1007), .B(_abc_19068_n1010), .Y(_abc_19068_n1011_1) );
  OR2X2 OR2X2_500 ( .A(_abc_19068_n2326_bF_buf7), .B(core_mi_4_), .Y(_abc_19068_n2347) );
  OR2X2 OR2X2_501 ( .A(_abc_19068_n2326_bF_buf5), .B(core_mi_5_), .Y(_abc_19068_n2352) );
  OR2X2 OR2X2_502 ( .A(_abc_19068_n2326_bF_buf3), .B(core_mi_6_), .Y(_abc_19068_n2357) );
  OR2X2 OR2X2_503 ( .A(_abc_19068_n2326_bF_buf1), .B(core_mi_7_), .Y(_abc_19068_n2362) );
  OR2X2 OR2X2_504 ( .A(_abc_19068_n2326_bF_buf7), .B(core_mi_8_), .Y(_abc_19068_n2367) );
  OR2X2 OR2X2_505 ( .A(_abc_19068_n2326_bF_buf5), .B(core_mi_9_), .Y(_abc_19068_n2372) );
  OR2X2 OR2X2_506 ( .A(_abc_19068_n2326_bF_buf3), .B(core_mi_10_), .Y(_abc_19068_n2377) );
  OR2X2 OR2X2_507 ( .A(_abc_19068_n2326_bF_buf1), .B(core_mi_11_), .Y(_abc_19068_n2382) );
  OR2X2 OR2X2_508 ( .A(_abc_19068_n2326_bF_buf7), .B(core_mi_12_), .Y(_abc_19068_n2387) );
  OR2X2 OR2X2_509 ( .A(_abc_19068_n2326_bF_buf5), .B(core_mi_13_), .Y(_abc_19068_n2392) );
  OR2X2 OR2X2_51 ( .A(_abc_19068_n1012_1), .B(_abc_19068_n1013), .Y(_abc_19068_n1014_1) );
  OR2X2 OR2X2_510 ( .A(_abc_19068_n2326_bF_buf3), .B(core_mi_14_), .Y(_abc_19068_n2397) );
  OR2X2 OR2X2_511 ( .A(_abc_19068_n2326_bF_buf1), .B(core_mi_15_), .Y(_abc_19068_n2402) );
  OR2X2 OR2X2_512 ( .A(_abc_19068_n2326_bF_buf7), .B(core_mi_16_), .Y(_abc_19068_n2407) );
  OR2X2 OR2X2_513 ( .A(_abc_19068_n2326_bF_buf5), .B(core_mi_17_), .Y(_abc_19068_n2412) );
  OR2X2 OR2X2_514 ( .A(_abc_19068_n2326_bF_buf3), .B(core_mi_18_), .Y(_abc_19068_n2417) );
  OR2X2 OR2X2_515 ( .A(_abc_19068_n2326_bF_buf1), .B(core_mi_19_), .Y(_abc_19068_n2422) );
  OR2X2 OR2X2_516 ( .A(_abc_19068_n2326_bF_buf7), .B(core_mi_20_), .Y(_abc_19068_n2427) );
  OR2X2 OR2X2_517 ( .A(_abc_19068_n2326_bF_buf5), .B(core_mi_21_), .Y(_abc_19068_n2432) );
  OR2X2 OR2X2_518 ( .A(_abc_19068_n2326_bF_buf3), .B(core_mi_22_), .Y(_abc_19068_n2437) );
  OR2X2 OR2X2_519 ( .A(_abc_19068_n2326_bF_buf1), .B(core_mi_23_), .Y(_abc_19068_n2442) );
  OR2X2 OR2X2_52 ( .A(_abc_19068_n1015_1), .B(_abc_19068_n906_1), .Y(_abc_19068_n1016) );
  OR2X2 OR2X2_520 ( .A(_abc_19068_n2326_bF_buf7), .B(core_mi_24_), .Y(_abc_19068_n2447) );
  OR2X2 OR2X2_521 ( .A(_abc_19068_n2326_bF_buf5), .B(core_mi_25_), .Y(_abc_19068_n2452) );
  OR2X2 OR2X2_522 ( .A(_abc_19068_n2326_bF_buf3), .B(core_mi_26_), .Y(_abc_19068_n2457) );
  OR2X2 OR2X2_523 ( .A(_abc_19068_n2326_bF_buf1), .B(core_mi_27_), .Y(_abc_19068_n2462) );
  OR2X2 OR2X2_524 ( .A(_abc_19068_n2326_bF_buf7), .B(core_mi_28_), .Y(_abc_19068_n2467) );
  OR2X2 OR2X2_525 ( .A(_abc_19068_n2326_bF_buf5), .B(core_mi_29_), .Y(_abc_19068_n2472) );
  OR2X2 OR2X2_526 ( .A(_abc_19068_n2326_bF_buf3), .B(core_mi_30_), .Y(_abc_19068_n2477) );
  OR2X2 OR2X2_527 ( .A(_abc_19068_n2326_bF_buf1), .B(core_mi_31_), .Y(_abc_19068_n2482) );
  OR2X2 OR2X2_528 ( .A(_abc_19068_n2487_bF_buf7), .B(core_key_96_), .Y(_abc_19068_n2488) );
  OR2X2 OR2X2_529 ( .A(_abc_19068_n2487_bF_buf5), .B(core_key_97_), .Y(_abc_19068_n2493) );
  OR2X2 OR2X2_53 ( .A(_abc_19068_n1014_1), .B(_abc_19068_n1016), .Y(_abc_19068_n1017_1) );
  OR2X2 OR2X2_530 ( .A(_abc_19068_n2487_bF_buf3), .B(core_key_98_), .Y(_abc_19068_n2498) );
  OR2X2 OR2X2_531 ( .A(_abc_19068_n2487_bF_buf1), .B(core_key_99_), .Y(_abc_19068_n2503) );
  OR2X2 OR2X2_532 ( .A(_abc_19068_n2487_bF_buf7), .B(core_key_100_), .Y(_abc_19068_n2508) );
  OR2X2 OR2X2_533 ( .A(_abc_19068_n2487_bF_buf5), .B(core_key_101_), .Y(_abc_19068_n2513) );
  OR2X2 OR2X2_534 ( .A(_abc_19068_n2487_bF_buf3), .B(core_key_102_), .Y(_abc_19068_n2518) );
  OR2X2 OR2X2_535 ( .A(_abc_19068_n2487_bF_buf1), .B(core_key_103_), .Y(_abc_19068_n2523) );
  OR2X2 OR2X2_536 ( .A(_abc_19068_n2487_bF_buf7), .B(core_key_104_), .Y(_abc_19068_n2528) );
  OR2X2 OR2X2_537 ( .A(_abc_19068_n2487_bF_buf5), .B(core_key_105_), .Y(_abc_19068_n2533) );
  OR2X2 OR2X2_538 ( .A(_abc_19068_n2487_bF_buf3), .B(core_key_106_), .Y(_abc_19068_n2538) );
  OR2X2 OR2X2_539 ( .A(_abc_19068_n2487_bF_buf1), .B(core_key_107_), .Y(_abc_19068_n2543) );
  OR2X2 OR2X2_54 ( .A(_abc_19068_n1011_1), .B(_abc_19068_n1017_1), .Y(_abc_19068_n1018_1) );
  OR2X2 OR2X2_540 ( .A(_abc_19068_n2487_bF_buf7), .B(core_key_108_), .Y(_abc_19068_n2548) );
  OR2X2 OR2X2_541 ( .A(_abc_19068_n2487_bF_buf5), .B(core_key_109_), .Y(_abc_19068_n2553) );
  OR2X2 OR2X2_542 ( .A(_abc_19068_n2487_bF_buf3), .B(core_key_110_), .Y(_abc_19068_n2558) );
  OR2X2 OR2X2_543 ( .A(_abc_19068_n2487_bF_buf1), .B(core_key_111_), .Y(_abc_19068_n2563) );
  OR2X2 OR2X2_544 ( .A(_abc_19068_n2487_bF_buf7), .B(core_key_112_), .Y(_abc_19068_n2568) );
  OR2X2 OR2X2_545 ( .A(_abc_19068_n2487_bF_buf5), .B(core_key_113_), .Y(_abc_19068_n2573) );
  OR2X2 OR2X2_546 ( .A(_abc_19068_n2487_bF_buf3), .B(core_key_114_), .Y(_abc_19068_n2578) );
  OR2X2 OR2X2_547 ( .A(_abc_19068_n2487_bF_buf1), .B(core_key_115_), .Y(_abc_19068_n2583) );
  OR2X2 OR2X2_548 ( .A(_abc_19068_n2487_bF_buf7), .B(core_key_116_), .Y(_abc_19068_n2588) );
  OR2X2 OR2X2_549 ( .A(_abc_19068_n2487_bF_buf5), .B(core_key_117_), .Y(_abc_19068_n2593) );
  OR2X2 OR2X2_55 ( .A(_abc_19068_n1019), .B(_abc_19068_n1020_1), .Y(_abc_19068_n1021_1) );
  OR2X2 OR2X2_550 ( .A(_abc_19068_n2487_bF_buf3), .B(core_key_118_), .Y(_abc_19068_n2598) );
  OR2X2 OR2X2_551 ( .A(_abc_19068_n2487_bF_buf1), .B(core_key_119_), .Y(_abc_19068_n2603) );
  OR2X2 OR2X2_552 ( .A(_abc_19068_n2487_bF_buf7), .B(core_key_120_), .Y(_abc_19068_n2608) );
  OR2X2 OR2X2_553 ( .A(_abc_19068_n2487_bF_buf5), .B(core_key_121_), .Y(_abc_19068_n2613) );
  OR2X2 OR2X2_554 ( .A(_abc_19068_n2487_bF_buf3), .B(core_key_122_), .Y(_abc_19068_n2618) );
  OR2X2 OR2X2_555 ( .A(_abc_19068_n2487_bF_buf1), .B(core_key_123_), .Y(_abc_19068_n2623) );
  OR2X2 OR2X2_556 ( .A(_abc_19068_n2487_bF_buf7), .B(core_key_124_), .Y(_abc_19068_n2628) );
  OR2X2 OR2X2_557 ( .A(_abc_19068_n2487_bF_buf5), .B(core_key_125_), .Y(_abc_19068_n2633) );
  OR2X2 OR2X2_558 ( .A(_abc_19068_n2487_bF_buf3), .B(core_key_126_), .Y(_abc_19068_n2638) );
  OR2X2 OR2X2_559 ( .A(_abc_19068_n2487_bF_buf1), .B(core_key_127_), .Y(_abc_19068_n2643) );
  OR2X2 OR2X2_56 ( .A(_abc_19068_n1022), .B(_abc_19068_n1023_1), .Y(_abc_19068_n1024_1) );
  OR2X2 OR2X2_560 ( .A(_abc_19068_n2648_bF_buf7), .B(core_key_64_), .Y(_abc_19068_n2649) );
  OR2X2 OR2X2_561 ( .A(_abc_19068_n2648_bF_buf5), .B(core_key_65_), .Y(_abc_19068_n2654) );
  OR2X2 OR2X2_562 ( .A(_abc_19068_n2648_bF_buf3), .B(core_key_66_), .Y(_abc_19068_n2659) );
  OR2X2 OR2X2_563 ( .A(_abc_19068_n2648_bF_buf1), .B(core_key_67_), .Y(_abc_19068_n2664) );
  OR2X2 OR2X2_564 ( .A(_abc_19068_n2648_bF_buf7), .B(core_key_68_), .Y(_abc_19068_n2669) );
  OR2X2 OR2X2_565 ( .A(_abc_19068_n2648_bF_buf5), .B(core_key_69_), .Y(_abc_19068_n2674) );
  OR2X2 OR2X2_566 ( .A(_abc_19068_n2648_bF_buf3), .B(core_key_70_), .Y(_abc_19068_n2679) );
  OR2X2 OR2X2_567 ( .A(_abc_19068_n2648_bF_buf1), .B(core_key_71_), .Y(_abc_19068_n2684) );
  OR2X2 OR2X2_568 ( .A(_abc_19068_n2648_bF_buf7), .B(core_key_72_), .Y(_abc_19068_n2689) );
  OR2X2 OR2X2_569 ( .A(_abc_19068_n2648_bF_buf5), .B(core_key_73_), .Y(_abc_19068_n2694) );
  OR2X2 OR2X2_57 ( .A(_abc_19068_n1021_1), .B(_abc_19068_n1024_1), .Y(_abc_19068_n1025) );
  OR2X2 OR2X2_570 ( .A(_abc_19068_n2648_bF_buf3), .B(core_key_74_), .Y(_abc_19068_n2699) );
  OR2X2 OR2X2_571 ( .A(_abc_19068_n2648_bF_buf1), .B(core_key_75_), .Y(_abc_19068_n2704) );
  OR2X2 OR2X2_572 ( .A(_abc_19068_n2648_bF_buf7), .B(core_key_76_), .Y(_abc_19068_n2709) );
  OR2X2 OR2X2_573 ( .A(_abc_19068_n2648_bF_buf5), .B(core_key_77_), .Y(_abc_19068_n2714) );
  OR2X2 OR2X2_574 ( .A(_abc_19068_n2648_bF_buf3), .B(core_key_78_), .Y(_abc_19068_n2719) );
  OR2X2 OR2X2_575 ( .A(_abc_19068_n2648_bF_buf1), .B(core_key_79_), .Y(_abc_19068_n2724) );
  OR2X2 OR2X2_576 ( .A(_abc_19068_n2648_bF_buf7), .B(core_key_80_), .Y(_abc_19068_n2729) );
  OR2X2 OR2X2_577 ( .A(_abc_19068_n2648_bF_buf5), .B(core_key_81_), .Y(_abc_19068_n2734) );
  OR2X2 OR2X2_578 ( .A(_abc_19068_n2648_bF_buf3), .B(core_key_82_), .Y(_abc_19068_n2739) );
  OR2X2 OR2X2_579 ( .A(_abc_19068_n2648_bF_buf1), .B(core_key_83_), .Y(_abc_19068_n2744) );
  OR2X2 OR2X2_58 ( .A(_abc_19068_n1018_1), .B(_abc_19068_n1025), .Y(_abc_19068_n1026_1) );
  OR2X2 OR2X2_580 ( .A(_abc_19068_n2648_bF_buf7), .B(core_key_84_), .Y(_abc_19068_n2749) );
  OR2X2 OR2X2_581 ( .A(_abc_19068_n2648_bF_buf5), .B(core_key_85_), .Y(_abc_19068_n2754) );
  OR2X2 OR2X2_582 ( .A(_abc_19068_n2648_bF_buf3), .B(core_key_86_), .Y(_abc_19068_n2759) );
  OR2X2 OR2X2_583 ( .A(_abc_19068_n2648_bF_buf1), .B(core_key_87_), .Y(_abc_19068_n2764) );
  OR2X2 OR2X2_584 ( .A(_abc_19068_n2648_bF_buf7), .B(core_key_88_), .Y(_abc_19068_n2769) );
  OR2X2 OR2X2_585 ( .A(_abc_19068_n2648_bF_buf5), .B(core_key_89_), .Y(_abc_19068_n2774) );
  OR2X2 OR2X2_586 ( .A(_abc_19068_n2648_bF_buf3), .B(core_key_90_), .Y(_abc_19068_n2779) );
  OR2X2 OR2X2_587 ( .A(_abc_19068_n2648_bF_buf1), .B(core_key_91_), .Y(_abc_19068_n2784) );
  OR2X2 OR2X2_588 ( .A(_abc_19068_n2648_bF_buf7), .B(core_key_92_), .Y(_abc_19068_n2789) );
  OR2X2 OR2X2_589 ( .A(_abc_19068_n2648_bF_buf5), .B(core_key_93_), .Y(_abc_19068_n2794) );
  OR2X2 OR2X2_59 ( .A(_abc_19068_n1028), .B(_abc_19068_n1029_1), .Y(_abc_19068_n1030_1) );
  OR2X2 OR2X2_590 ( .A(_abc_19068_n2648_bF_buf3), .B(core_key_94_), .Y(_abc_19068_n2799) );
  OR2X2 OR2X2_591 ( .A(_abc_19068_n2648_bF_buf1), .B(core_key_95_), .Y(_abc_19068_n2804) );
  OR2X2 OR2X2_592 ( .A(_abc_19068_n2809_bF_buf7), .B(core_key_32_), .Y(_abc_19068_n2810) );
  OR2X2 OR2X2_593 ( .A(_abc_19068_n2809_bF_buf5), .B(core_key_33_), .Y(_abc_19068_n2815) );
  OR2X2 OR2X2_594 ( .A(_abc_19068_n2809_bF_buf3), .B(core_key_34_), .Y(_abc_19068_n2820) );
  OR2X2 OR2X2_595 ( .A(_abc_19068_n2809_bF_buf1), .B(core_key_35_), .Y(_abc_19068_n2825) );
  OR2X2 OR2X2_596 ( .A(_abc_19068_n2809_bF_buf7), .B(core_key_36_), .Y(_abc_19068_n2830) );
  OR2X2 OR2X2_597 ( .A(_abc_19068_n2809_bF_buf5), .B(core_key_37_), .Y(_abc_19068_n2835) );
  OR2X2 OR2X2_598 ( .A(_abc_19068_n2809_bF_buf3), .B(core_key_38_), .Y(_abc_19068_n2840) );
  OR2X2 OR2X2_599 ( .A(_abc_19068_n2809_bF_buf1), .B(core_key_39_), .Y(_abc_19068_n2845) );
  OR2X2 OR2X2_6 ( .A(_abc_19068_n907_1), .B(_abc_19068_n901_1), .Y(_abc_19068_n908) );
  OR2X2 OR2X2_60 ( .A(_abc_19068_n1031), .B(_abc_19068_n1032_1), .Y(_abc_19068_n1033_1) );
  OR2X2 OR2X2_600 ( .A(_abc_19068_n2809_bF_buf7), .B(core_key_40_), .Y(_abc_19068_n2850) );
  OR2X2 OR2X2_601 ( .A(_abc_19068_n2809_bF_buf5), .B(core_key_41_), .Y(_abc_19068_n2855) );
  OR2X2 OR2X2_602 ( .A(_abc_19068_n2809_bF_buf3), .B(core_key_42_), .Y(_abc_19068_n2860) );
  OR2X2 OR2X2_603 ( .A(_abc_19068_n2809_bF_buf1), .B(core_key_43_), .Y(_abc_19068_n2865) );
  OR2X2 OR2X2_604 ( .A(_abc_19068_n2809_bF_buf7), .B(core_key_44_), .Y(_abc_19068_n2870) );
  OR2X2 OR2X2_605 ( .A(_abc_19068_n2809_bF_buf5), .B(core_key_45_), .Y(_abc_19068_n2875) );
  OR2X2 OR2X2_606 ( .A(_abc_19068_n2809_bF_buf3), .B(core_key_46_), .Y(_abc_19068_n2880) );
  OR2X2 OR2X2_607 ( .A(_abc_19068_n2809_bF_buf1), .B(core_key_47_), .Y(_abc_19068_n2885) );
  OR2X2 OR2X2_608 ( .A(_abc_19068_n2809_bF_buf7), .B(core_key_48_), .Y(_abc_19068_n2890) );
  OR2X2 OR2X2_609 ( .A(_abc_19068_n2809_bF_buf5), .B(core_key_49_), .Y(_abc_19068_n2895) );
  OR2X2 OR2X2_61 ( .A(_abc_19068_n1030_1), .B(_abc_19068_n1033_1), .Y(_abc_19068_n1034) );
  OR2X2 OR2X2_610 ( .A(_abc_19068_n2809_bF_buf3), .B(core_key_50_), .Y(_abc_19068_n2900) );
  OR2X2 OR2X2_611 ( .A(_abc_19068_n2809_bF_buf1), .B(core_key_51_), .Y(_abc_19068_n2905) );
  OR2X2 OR2X2_612 ( .A(_abc_19068_n2809_bF_buf7), .B(core_key_52_), .Y(_abc_19068_n2910) );
  OR2X2 OR2X2_613 ( .A(_abc_19068_n2809_bF_buf5), .B(core_key_53_), .Y(_abc_19068_n2915) );
  OR2X2 OR2X2_614 ( .A(_abc_19068_n2809_bF_buf3), .B(core_key_54_), .Y(_abc_19068_n2920) );
  OR2X2 OR2X2_615 ( .A(_abc_19068_n2809_bF_buf1), .B(core_key_55_), .Y(_abc_19068_n2925) );
  OR2X2 OR2X2_616 ( .A(_abc_19068_n2809_bF_buf7), .B(core_key_56_), .Y(_abc_19068_n2930) );
  OR2X2 OR2X2_617 ( .A(_abc_19068_n2809_bF_buf5), .B(core_key_57_), .Y(_abc_19068_n2935) );
  OR2X2 OR2X2_618 ( .A(_abc_19068_n2809_bF_buf3), .B(core_key_58_), .Y(_abc_19068_n2940) );
  OR2X2 OR2X2_619 ( .A(_abc_19068_n2809_bF_buf1), .B(core_key_59_), .Y(_abc_19068_n2945) );
  OR2X2 OR2X2_62 ( .A(_abc_19068_n1035_1), .B(_abc_19068_n1036_1), .Y(_abc_19068_n1037) );
  OR2X2 OR2X2_620 ( .A(_abc_19068_n2809_bF_buf7), .B(core_key_60_), .Y(_abc_19068_n2950) );
  OR2X2 OR2X2_621 ( .A(_abc_19068_n2809_bF_buf5), .B(core_key_61_), .Y(_abc_19068_n2955) );
  OR2X2 OR2X2_622 ( .A(_abc_19068_n2809_bF_buf3), .B(core_key_62_), .Y(_abc_19068_n2960) );
  OR2X2 OR2X2_623 ( .A(_abc_19068_n2809_bF_buf1), .B(core_key_63_), .Y(_abc_19068_n2965) );
  OR2X2 OR2X2_624 ( .A(_abc_19068_n2970_bF_buf7), .B(core_key_0_), .Y(_abc_19068_n2971) );
  OR2X2 OR2X2_625 ( .A(_abc_19068_n2970_bF_buf5), .B(core_key_1_), .Y(_abc_19068_n2976) );
  OR2X2 OR2X2_626 ( .A(_abc_19068_n2970_bF_buf3), .B(core_key_2_), .Y(_abc_19068_n2981) );
  OR2X2 OR2X2_627 ( .A(_abc_19068_n2970_bF_buf1), .B(core_key_3_), .Y(_abc_19068_n2986) );
  OR2X2 OR2X2_628 ( .A(_abc_19068_n2970_bF_buf7), .B(core_key_4_), .Y(_abc_19068_n2991) );
  OR2X2 OR2X2_629 ( .A(_abc_19068_n2970_bF_buf5), .B(core_key_5_), .Y(_abc_19068_n2996) );
  OR2X2 OR2X2_63 ( .A(_abc_19068_n1039_1), .B(_abc_19068_n1038_1), .Y(_abc_19068_n1040) );
  OR2X2 OR2X2_630 ( .A(_abc_19068_n2970_bF_buf3), .B(core_key_6_), .Y(_abc_19068_n3001) );
  OR2X2 OR2X2_631 ( .A(_abc_19068_n2970_bF_buf1), .B(core_key_7_), .Y(_abc_19068_n3006) );
  OR2X2 OR2X2_632 ( .A(_abc_19068_n2970_bF_buf7), .B(core_key_8_), .Y(_abc_19068_n3011) );
  OR2X2 OR2X2_633 ( .A(_abc_19068_n2970_bF_buf5), .B(core_key_9_), .Y(_abc_19068_n3016) );
  OR2X2 OR2X2_634 ( .A(_abc_19068_n2970_bF_buf3), .B(core_key_10_), .Y(_abc_19068_n3021) );
  OR2X2 OR2X2_635 ( .A(_abc_19068_n2970_bF_buf1), .B(core_key_11_), .Y(_abc_19068_n3026) );
  OR2X2 OR2X2_636 ( .A(_abc_19068_n2970_bF_buf7), .B(core_key_12_), .Y(_abc_19068_n3031) );
  OR2X2 OR2X2_637 ( .A(_abc_19068_n2970_bF_buf5), .B(core_key_13_), .Y(_abc_19068_n3036) );
  OR2X2 OR2X2_638 ( .A(_abc_19068_n2970_bF_buf3), .B(core_key_14_), .Y(_abc_19068_n3041) );
  OR2X2 OR2X2_639 ( .A(_abc_19068_n2970_bF_buf1), .B(core_key_15_), .Y(_abc_19068_n3046) );
  OR2X2 OR2X2_64 ( .A(_abc_19068_n1037), .B(_abc_19068_n1040), .Y(_abc_19068_n1041_1) );
  OR2X2 OR2X2_640 ( .A(_abc_19068_n2970_bF_buf7), .B(core_key_16_), .Y(_abc_19068_n3051) );
  OR2X2 OR2X2_641 ( .A(_abc_19068_n2970_bF_buf5), .B(core_key_17_), .Y(_abc_19068_n3056) );
  OR2X2 OR2X2_642 ( .A(_abc_19068_n2970_bF_buf3), .B(core_key_18_), .Y(_abc_19068_n3061) );
  OR2X2 OR2X2_643 ( .A(_abc_19068_n2970_bF_buf1), .B(core_key_19_), .Y(_abc_19068_n3066) );
  OR2X2 OR2X2_644 ( .A(_abc_19068_n2970_bF_buf7), .B(core_key_20_), .Y(_abc_19068_n3071) );
  OR2X2 OR2X2_645 ( .A(_abc_19068_n2970_bF_buf5), .B(core_key_21_), .Y(_abc_19068_n3076) );
  OR2X2 OR2X2_646 ( .A(_abc_19068_n2970_bF_buf3), .B(core_key_22_), .Y(_abc_19068_n3081) );
  OR2X2 OR2X2_647 ( .A(_abc_19068_n2970_bF_buf1), .B(core_key_23_), .Y(_abc_19068_n3086) );
  OR2X2 OR2X2_648 ( .A(_abc_19068_n2970_bF_buf7), .B(core_key_24_), .Y(_abc_19068_n3091) );
  OR2X2 OR2X2_649 ( .A(_abc_19068_n2970_bF_buf5), .B(core_key_25_), .Y(_abc_19068_n3096) );
  OR2X2 OR2X2_65 ( .A(_abc_19068_n1034), .B(_abc_19068_n1041_1), .Y(_abc_19068_n1042_1) );
  OR2X2 OR2X2_650 ( .A(_abc_19068_n2970_bF_buf3), .B(core_key_26_), .Y(_abc_19068_n3101) );
  OR2X2 OR2X2_651 ( .A(_abc_19068_n2970_bF_buf1), .B(core_key_27_), .Y(_abc_19068_n3106) );
  OR2X2 OR2X2_652 ( .A(_abc_19068_n2970_bF_buf7), .B(core_key_28_), .Y(_abc_19068_n3111) );
  OR2X2 OR2X2_653 ( .A(_abc_19068_n2970_bF_buf5), .B(core_key_29_), .Y(_abc_19068_n3116) );
  OR2X2 OR2X2_654 ( .A(_abc_19068_n2970_bF_buf3), .B(core_key_30_), .Y(_abc_19068_n3121) );
  OR2X2 OR2X2_655 ( .A(_abc_19068_n2970_bF_buf1), .B(core_key_31_), .Y(_abc_19068_n3126) );
  OR2X2 OR2X2_656 ( .A(_abc_19068_n3134), .B(_abc_19068_n3132), .Y(_abc_19068_n3135) );
  OR2X2 OR2X2_657 ( .A(_abc_19068_n3139), .B(_abc_19068_n3138), .Y(_abc_19068_n3140) );
  OR2X2 OR2X2_658 ( .A(_abc_19068_n3140), .B(_abc_19068_n3137), .Y(param_reg_1__FF_INPUT) );
  OR2X2 OR2X2_659 ( .A(_abc_19068_n3143), .B(_abc_19068_n3142), .Y(_abc_19068_n3144) );
  OR2X2 OR2X2_66 ( .A(_abc_19068_n1043), .B(_abc_19068_n1044_1), .Y(_abc_19068_n1045_1) );
  OR2X2 OR2X2_660 ( .A(_abc_19068_n3147), .B(_abc_19068_n3146), .Y(_abc_19068_n3148) );
  OR2X2 OR2X2_661 ( .A(_abc_19068_n3151), .B(_abc_19068_n3150), .Y(_abc_19068_n3152) );
  OR2X2 OR2X2_662 ( .A(_abc_19068_n3155), .B(_abc_19068_n3154), .Y(_abc_19068_n3156) );
  OR2X2 OR2X2_663 ( .A(_abc_19068_n3159), .B(_abc_19068_n3138), .Y(_abc_19068_n3160) );
  OR2X2 OR2X2_664 ( .A(_abc_19068_n3160), .B(_abc_19068_n3158), .Y(param_reg_6__FF_INPUT) );
  OR2X2 OR2X2_665 ( .A(_abc_19068_n3163), .B(_abc_19068_n3162), .Y(_abc_19068_n3164) );
  OR2X2 OR2X2_666 ( .A(_abc_19068_n3175), .B(core_long), .Y(_abc_19068_n3178) );
  OR2X2 OR2X2_667 ( .A(core_siphash_ctrl_reg_3_), .B(core_siphash_ctrl_reg_6_), .Y(core__abc_21380_n1140_1) );
  OR2X2 OR2X2_668 ( .A(core__abc_21380_n1140_1), .B(core_siphash_ctrl_reg_4_), .Y(core__abc_21380_n1141_1) );
  OR2X2 OR2X2_669 ( .A(core__abc_21380_n1150_1), .B(core_loop_ctr_reg_1_), .Y(core__abc_21380_n1156_1) );
  OR2X2 OR2X2_67 ( .A(_abc_19068_n1046), .B(_abc_19068_n1047_1), .Y(_abc_19068_n1048_1) );
  OR2X2 OR2X2_670 ( .A(core__abc_21380_n1157_1), .B(core_compression_rounds_1_), .Y(core__abc_21380_n1158_1) );
  OR2X2 OR2X2_671 ( .A(core__abc_21380_n1161_1), .B(core__abc_21380_n1154_1), .Y(core__abc_21380_n1162_1) );
  OR2X2 OR2X2_672 ( .A(core__abc_21380_n1164_1), .B(core__abc_21380_n1163), .Y(core__abc_21380_n1165_1) );
  OR2X2 OR2X2_673 ( .A(core__abc_21380_n1162_1), .B(core__abc_21380_n1165_1), .Y(core__abc_21380_n1166_1) );
  OR2X2 OR2X2_674 ( .A(core__abc_21380_n1152_1), .B(core__abc_21380_n1149_1), .Y(core__abc_21380_n1169_1) );
  OR2X2 OR2X2_675 ( .A(core__abc_21380_n1170_1), .B(core_loop_ctr_reg_2_), .Y(core__abc_21380_n1173_1) );
  OR2X2 OR2X2_676 ( .A(core__abc_21380_n1176_1), .B(core__abc_21380_n1154_1), .Y(core__abc_21380_n1177_1) );
  OR2X2 OR2X2_677 ( .A(core__abc_21380_n1179), .B(core__abc_21380_n1181_1), .Y(core__abc_21380_n1182_1) );
  OR2X2 OR2X2_678 ( .A(core__abc_21380_n1192_1), .B(core__abc_21380_n1193_1), .Y(core__abc_21380_n1194_1) );
  OR2X2 OR2X2_679 ( .A(core__abc_21380_n1157_1), .B(core_final_rounds_1_), .Y(core__abc_21380_n1195) );
  OR2X2 OR2X2_68 ( .A(_abc_19068_n1045_1), .B(_abc_19068_n1048_1), .Y(_abc_19068_n1049) );
  OR2X2 OR2X2_680 ( .A(core__abc_21380_n1188_1), .B(core_loop_ctr_reg_1_), .Y(core__abc_21380_n1196_1) );
  OR2X2 OR2X2_681 ( .A(core__abc_21380_n1199), .B(core__abc_21380_n1200_1), .Y(core__abc_21380_n1201_1) );
  OR2X2 OR2X2_682 ( .A(core__abc_21380_n1201_1), .B(core__abc_21380_n1194_1), .Y(core__abc_21380_n1202_1) );
  OR2X2 OR2X2_683 ( .A(core__abc_21380_n1190_1), .B(core__abc_21380_n1187), .Y(core__abc_21380_n1206_1) );
  OR2X2 OR2X2_684 ( .A(core__abc_21380_n1208_1), .B(core__abc_21380_n1204_1), .Y(core__abc_21380_n1209_1) );
  OR2X2 OR2X2_685 ( .A(core__abc_21380_n1207), .B(core_loop_ctr_reg_2_), .Y(core__abc_21380_n1210_1) );
  OR2X2 OR2X2_686 ( .A(core__abc_21380_n1213_1), .B(core__abc_21380_n1192_1), .Y(core__abc_21380_n1214_1) );
  OR2X2 OR2X2_687 ( .A(core__abc_21380_n1216_1), .B(core__abc_21380_n1217_1), .Y(core__abc_21380_n1218_1) );
  OR2X2 OR2X2_688 ( .A(core__abc_21380_n1221_1), .B(core__abc_21380_n1222_1), .Y(core__abc_21380_n1223) );
  OR2X2 OR2X2_689 ( .A(core__abc_21380_n1223), .B(core__abc_21380_n1185_1), .Y(core__abc_21380_n1224_1) );
  OR2X2 OR2X2_69 ( .A(_abc_19068_n1042_1), .B(_abc_19068_n1049), .Y(_abc_19068_n1050_1) );
  OR2X2 OR2X2_690 ( .A(core__abc_21380_n1224_1), .B(core__abc_21380_n1147), .Y(core__abc_21380_n1225_1) );
  OR2X2 OR2X2_691 ( .A(core__abc_21380_n1233_1), .B(core__abc_21380_n1234_1), .Y(core__abc_21380_n1235) );
  OR2X2 OR2X2_692 ( .A(core__abc_21380_n1235), .B(core__abc_21380_n1231), .Y(core__abc_21380_n1236_1) );
  OR2X2 OR2X2_693 ( .A(core__abc_21380_n1242_1), .B(core_siphash_ctrl_reg_2_), .Y(core__abc_21380_n1243) );
  OR2X2 OR2X2_694 ( .A(core__abc_21380_n1241_1), .B(core__abc_21380_n1243), .Y(core__abc_21380_n1244_1) );
  OR2X2 OR2X2_695 ( .A(core__abc_21380_n1240_1), .B(core__abc_21380_n1244_1), .Y(core__abc_21380_n1245_1) );
  OR2X2 OR2X2_696 ( .A(core__abc_21380_n1245_1), .B(core__abc_21380_n1237_1), .Y(core__abc_21380_n1246_1) );
  OR2X2 OR2X2_697 ( .A(core__abc_21380_n1246_1), .B(core__abc_21380_n1229_1), .Y(core__abc_14829_n1285) );
  OR2X2 OR2X2_698 ( .A(core__abc_21380_n1250_1), .B(core__abc_21380_n1248_1), .Y(core__abc_14829_n1310) );
  OR2X2 OR2X2_699 ( .A(core__abc_21380_n1253_1), .B(core__abc_21380_n1252_1), .Y(core__abc_14829_n1316) );
  OR2X2 OR2X2_7 ( .A(_abc_19068_n909_1), .B(_abc_19068_n906_1), .Y(_abc_19068_n910_1) );
  OR2X2 OR2X2_70 ( .A(_abc_19068_n1052), .B(_abc_19068_n1053_1), .Y(_abc_19068_n1054_1) );
  OR2X2 OR2X2_700 ( .A(core__abc_21380_n1256_1), .B(core__abc_21380_n1257_1), .Y(core__abc_14829_n1330) );
  OR2X2 OR2X2_701 ( .A(core_v0_reg_0_), .B(core_v1_reg_0_), .Y(core__abc_21380_n1259) );
  OR2X2 OR2X2_702 ( .A(core__abc_21380_n1265_1), .B(core__abc_21380_n1266_1), .Y(core__abc_21380_n1267) );
  OR2X2 OR2X2_703 ( .A(core__abc_21380_n1268_1), .B(core__abc_21380_n1262_1), .Y(core__abc_21380_n1269_1) );
  OR2X2 OR2X2_704 ( .A(core__abc_21380_n1270_1), .B(core__abc_21380_n1267), .Y(core__abc_21380_n1271) );
  OR2X2 OR2X2_705 ( .A(core__abc_21380_n1272_1), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n1273_1) );
  OR2X2 OR2X2_706 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_64_), .Y(core__abc_21380_n1274_1) );
  OR2X2 OR2X2_707 ( .A(core_v0_reg_1_), .B(core_v1_reg_1_), .Y(core__abc_21380_n1277_1) );
  OR2X2 OR2X2_708 ( .A(core__abc_21380_n1284_1), .B(core__abc_21380_n1281_1), .Y(core__abc_21380_n1285_1) );
  OR2X2 OR2X2_709 ( .A(core__abc_21380_n1286_1), .B(core__abc_21380_n1280_1), .Y(core__abc_21380_n1287) );
  OR2X2 OR2X2_71 ( .A(_abc_19068_n910_1), .B(_abc_19068_n1054_1), .Y(_abc_19068_n1055) );
  OR2X2 OR2X2_710 ( .A(core__abc_21380_n1290), .B(core__abc_21380_n1278_1), .Y(core__abc_21380_n1291) );
  OR2X2 OR2X2_711 ( .A(core__abc_21380_n1291), .B(core__abc_21380_n1285_1), .Y(core__abc_21380_n1292) );
  OR2X2 OR2X2_712 ( .A(core__abc_21380_n1293), .B(core__abc_21380_n1134_1_bF_buf5), .Y(core__abc_21380_n1294) );
  OR2X2 OR2X2_713 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_65_), .Y(core__abc_21380_n1295) );
  OR2X2 OR2X2_714 ( .A(core__abc_21380_n1300), .B(core__abc_21380_n1301), .Y(core__abc_21380_n1302) );
  OR2X2 OR2X2_715 ( .A(core__abc_21380_n1307), .B(core__abc_21380_n1304), .Y(core__abc_21380_n1308) );
  OR2X2 OR2X2_716 ( .A(core__abc_21380_n1303), .B(core__abc_21380_n1309), .Y(core__abc_21380_n1310) );
  OR2X2 OR2X2_717 ( .A(core__abc_21380_n1302), .B(core__abc_21380_n1308), .Y(core__abc_21380_n1311) );
  OR2X2 OR2X2_718 ( .A(core__abc_21380_n1312), .B(core__abc_21380_n1134_1_bF_buf4), .Y(core__abc_21380_n1313) );
  OR2X2 OR2X2_719 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_66_), .Y(core__abc_21380_n1314) );
  OR2X2 OR2X2_72 ( .A(_abc_19068_n1057_1), .B(_abc_19068_n1058), .Y(_abc_19068_n1059_1) );
  OR2X2 OR2X2_720 ( .A(core__abc_21380_n1320), .B(core__abc_21380_n1317), .Y(core__abc_21380_n1321) );
  OR2X2 OR2X2_721 ( .A(core__abc_21380_n1326), .B(core__abc_21380_n1323), .Y(core__abc_21380_n1327) );
  OR2X2 OR2X2_722 ( .A(core__abc_21380_n1328), .B(core__abc_21380_n1330), .Y(core__abc_21380_n1331) );
  OR2X2 OR2X2_723 ( .A(core__abc_21380_n1331), .B(core__abc_21380_n1134_1_bF_buf3), .Y(core__abc_21380_n1332) );
  OR2X2 OR2X2_724 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_67_), .Y(core__abc_21380_n1333) );
  OR2X2 OR2X2_725 ( .A(core_v0_reg_4_), .B(core_v1_reg_4_), .Y(core__abc_21380_n1336) );
  OR2X2 OR2X2_726 ( .A(core__abc_21380_n1343), .B(core__abc_21380_n1340), .Y(core__abc_21380_n1344) );
  OR2X2 OR2X2_727 ( .A(core__abc_21380_n1345), .B(core__abc_21380_n1339), .Y(core__abc_21380_n1346) );
  OR2X2 OR2X2_728 ( .A(core__abc_21380_n1347), .B(core__abc_21380_n1344), .Y(core__abc_21380_n1348) );
  OR2X2 OR2X2_729 ( .A(core__abc_21380_n1349), .B(core__abc_21380_n1134_1_bF_buf2), .Y(core__abc_21380_n1350) );
  OR2X2 OR2X2_73 ( .A(_abc_19068_n1059_1), .B(_abc_19068_n1056_1), .Y(_abc_19068_n1060_1) );
  OR2X2 OR2X2_730 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_68_), .Y(core__abc_21380_n1351) );
  OR2X2 OR2X2_731 ( .A(core__abc_21380_n1357), .B(core__abc_21380_n1354), .Y(core__abc_21380_n1358) );
  OR2X2 OR2X2_732 ( .A(core__abc_21380_n1363), .B(core__abc_21380_n1360), .Y(core__abc_21380_n1364) );
  OR2X2 OR2X2_733 ( .A(core__abc_21380_n1367), .B(core__abc_21380_n1365), .Y(core__abc_21380_n1368) );
  OR2X2 OR2X2_734 ( .A(core__abc_21380_n1368), .B(core__abc_21380_n1134_1_bF_buf1), .Y(core__abc_21380_n1369) );
  OR2X2 OR2X2_735 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_69_), .Y(core__abc_21380_n1370) );
  OR2X2 OR2X2_736 ( .A(core__abc_21380_n1375), .B(core__abc_21380_n1376), .Y(core__abc_21380_n1377) );
  OR2X2 OR2X2_737 ( .A(core__abc_21380_n1382), .B(core__abc_21380_n1379), .Y(core__abc_21380_n1383) );
  OR2X2 OR2X2_738 ( .A(core__abc_21380_n1384), .B(core__abc_21380_n1378), .Y(core__abc_21380_n1385) );
  OR2X2 OR2X2_739 ( .A(core__abc_21380_n1377), .B(core__abc_21380_n1383), .Y(core__abc_21380_n1386) );
  OR2X2 OR2X2_74 ( .A(_abc_19068_n1055), .B(_abc_19068_n1060_1), .Y(_abc_19068_n1061) );
  OR2X2 OR2X2_740 ( .A(core__abc_21380_n1387), .B(core__abc_21380_n1134_1_bF_buf0), .Y(core__abc_21380_n1388) );
  OR2X2 OR2X2_741 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_70_), .Y(core__abc_21380_n1389) );
  OR2X2 OR2X2_742 ( .A(core__abc_21380_n1394), .B(core__abc_21380_n1395), .Y(core__abc_21380_n1396) );
  OR2X2 OR2X2_743 ( .A(core__abc_21380_n1401), .B(core__abc_21380_n1398), .Y(core__abc_21380_n1402) );
  OR2X2 OR2X2_744 ( .A(core__abc_21380_n1403), .B(core__abc_21380_n1397), .Y(core__abc_21380_n1404) );
  OR2X2 OR2X2_745 ( .A(core__abc_21380_n1396), .B(core__abc_21380_n1402), .Y(core__abc_21380_n1405) );
  OR2X2 OR2X2_746 ( .A(core__abc_21380_n1406), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n1407) );
  OR2X2 OR2X2_747 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_71_), .Y(core__abc_21380_n1408) );
  OR2X2 OR2X2_748 ( .A(core_v0_reg_8_), .B(core_v1_reg_8_), .Y(core__abc_21380_n1413) );
  OR2X2 OR2X2_749 ( .A(core_v2_reg_8_), .B(core_v3_reg_8_), .Y(core__abc_21380_n1417) );
  OR2X2 OR2X2_75 ( .A(_abc_19068_n1062_1), .B(_abc_19068_n1063_1), .Y(_abc_19068_n1064) );
  OR2X2 OR2X2_750 ( .A(core__abc_21380_n1420), .B(core__abc_21380_n1422), .Y(core__abc_21380_n1423) );
  OR2X2 OR2X2_751 ( .A(core__abc_21380_n1423), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n1424) );
  OR2X2 OR2X2_752 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_72_), .Y(core__abc_21380_n1425) );
  OR2X2 OR2X2_753 ( .A(core_v2_reg_9_), .B(core_v3_reg_9_), .Y(core__abc_21380_n1437) );
  OR2X2 OR2X2_754 ( .A(core__abc_21380_n1442), .B(core__abc_21380_n1440), .Y(core__abc_21380_n1443) );
  OR2X2 OR2X2_755 ( .A(core__abc_21380_n1443), .B(core__abc_21380_n1134_1_bF_buf5), .Y(core__abc_21380_n1444) );
  OR2X2 OR2X2_756 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_73_), .Y(core__abc_21380_n1445) );
  OR2X2 OR2X2_757 ( .A(core_v0_reg_10_), .B(core_v1_reg_10_), .Y(core__abc_21380_n1448) );
  OR2X2 OR2X2_758 ( .A(core_v3_reg_10_), .B(core_v2_reg_10_), .Y(core__abc_21380_n1454) );
  OR2X2 OR2X2_759 ( .A(core__abc_21380_n1451), .B(core__abc_21380_n1455), .Y(core__abc_21380_n1456) );
  OR2X2 OR2X2_76 ( .A(_abc_19068_n1065_1), .B(_abc_19068_n1066_1), .Y(_abc_19068_n1067) );
  OR2X2 OR2X2_760 ( .A(core__abc_21380_n1458), .B(core__abc_21380_n1457), .Y(core__abc_21380_n1459) );
  OR2X2 OR2X2_761 ( .A(core__abc_21380_n1460), .B(core__abc_21380_n1134_1_bF_buf4), .Y(core__abc_21380_n1461) );
  OR2X2 OR2X2_762 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_74_), .Y(core__abc_21380_n1462) );
  OR2X2 OR2X2_763 ( .A(core_v0_reg_11_), .B(core_v1_reg_11_), .Y(core__abc_21380_n1465) );
  OR2X2 OR2X2_764 ( .A(core_v3_reg_11_), .B(core_v2_reg_11_), .Y(core__abc_21380_n1471) );
  OR2X2 OR2X2_765 ( .A(core__abc_21380_n1468), .B(core__abc_21380_n1472), .Y(core__abc_21380_n1473) );
  OR2X2 OR2X2_766 ( .A(core__abc_21380_n1475), .B(core__abc_21380_n1474), .Y(core__abc_21380_n1476) );
  OR2X2 OR2X2_767 ( .A(core__abc_21380_n1477), .B(core__abc_21380_n1134_1_bF_buf3), .Y(core__abc_21380_n1478) );
  OR2X2 OR2X2_768 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_75_), .Y(core__abc_21380_n1479) );
  OR2X2 OR2X2_769 ( .A(core__abc_21380_n1485), .B(core__abc_21380_n1482), .Y(core__abc_21380_n1486) );
  OR2X2 OR2X2_77 ( .A(_abc_19068_n1068_1), .B(_abc_19068_n1069_1), .Y(_abc_19068_n1070) );
  OR2X2 OR2X2_770 ( .A(core_v2_reg_12_), .B(core_v3_reg_12_), .Y(core__abc_21380_n1490) );
  OR2X2 OR2X2_771 ( .A(core__abc_21380_n1493), .B(core__abc_21380_n1494), .Y(core__abc_21380_n1495) );
  OR2X2 OR2X2_772 ( .A(core__abc_21380_n1495), .B(core__abc_21380_n1134_1_bF_buf2), .Y(core__abc_21380_n1496) );
  OR2X2 OR2X2_773 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_76_), .Y(core__abc_21380_n1497) );
  OR2X2 OR2X2_774 ( .A(core__abc_21380_n1502), .B(core__abc_21380_n1503), .Y(core__abc_21380_n1504) );
  OR2X2 OR2X2_775 ( .A(core_v3_reg_13_), .B(core_v2_reg_13_), .Y(core__abc_21380_n1508) );
  OR2X2 OR2X2_776 ( .A(core__abc_21380_n1505), .B(core__abc_21380_n1509), .Y(core__abc_21380_n1510) );
  OR2X2 OR2X2_777 ( .A(core__abc_21380_n1511), .B(core__abc_21380_n1504), .Y(core__abc_21380_n1512) );
  OR2X2 OR2X2_778 ( .A(core__abc_21380_n1513), .B(core__abc_21380_n1134_1_bF_buf1), .Y(core__abc_21380_n1514) );
  OR2X2 OR2X2_779 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_77_), .Y(core__abc_21380_n1515) );
  OR2X2 OR2X2_78 ( .A(_abc_19068_n1067), .B(_abc_19068_n1070), .Y(_abc_19068_n1071_1) );
  OR2X2 OR2X2_780 ( .A(core__abc_21380_n1520), .B(core__abc_21380_n1521), .Y(core__abc_21380_n1522) );
  OR2X2 OR2X2_781 ( .A(core_v3_reg_14_), .B(core_v2_reg_14_), .Y(core__abc_21380_n1526) );
  OR2X2 OR2X2_782 ( .A(core__abc_21380_n1523), .B(core__abc_21380_n1527), .Y(core__abc_21380_n1528) );
  OR2X2 OR2X2_783 ( .A(core__abc_21380_n1529), .B(core__abc_21380_n1522), .Y(core__abc_21380_n1530) );
  OR2X2 OR2X2_784 ( .A(core__abc_21380_n1531), .B(core__abc_21380_n1134_1_bF_buf0), .Y(core__abc_21380_n1532) );
  OR2X2 OR2X2_785 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_78_), .Y(core__abc_21380_n1533) );
  OR2X2 OR2X2_786 ( .A(core_v3_reg_15_), .B(core_v2_reg_15_), .Y(core__abc_21380_n1545) );
  OR2X2 OR2X2_787 ( .A(core__abc_21380_n1542), .B(core__abc_21380_n1546), .Y(core__abc_21380_n1547) );
  OR2X2 OR2X2_788 ( .A(core__abc_21380_n1548), .B(core__abc_21380_n1549), .Y(core__abc_21380_n1550) );
  OR2X2 OR2X2_789 ( .A(core__abc_21380_n1551), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n1552) );
  OR2X2 OR2X2_79 ( .A(_abc_19068_n1071_1), .B(_abc_19068_n1064), .Y(_abc_19068_n1072_1) );
  OR2X2 OR2X2_790 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_79_), .Y(core__abc_21380_n1553) );
  OR2X2 OR2X2_791 ( .A(core__abc_21380_n1559), .B(core__abc_21380_n1556), .Y(core__abc_21380_n1560) );
  OR2X2 OR2X2_792 ( .A(core_v2_reg_16_), .B(core_v3_reg_16_), .Y(core__abc_21380_n1564) );
  OR2X2 OR2X2_793 ( .A(core__abc_21380_n1567), .B(core__abc_21380_n1568), .Y(core__abc_21380_n1569) );
  OR2X2 OR2X2_794 ( .A(core__abc_21380_n1569), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n1570) );
  OR2X2 OR2X2_795 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_80_), .Y(core__abc_21380_n1571) );
  OR2X2 OR2X2_796 ( .A(core_v2_reg_17_), .B(core_v3_reg_17_), .Y(core__abc_21380_n1583) );
  OR2X2 OR2X2_797 ( .A(core__abc_21380_n1588), .B(core__abc_21380_n1586), .Y(core__abc_21380_n1589) );
  OR2X2 OR2X2_798 ( .A(core__abc_21380_n1589), .B(core__abc_21380_n1134_1_bF_buf5), .Y(core__abc_21380_n1590) );
  OR2X2 OR2X2_799 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_81_), .Y(core__abc_21380_n1591) );
  OR2X2 OR2X2_8 ( .A(_abc_19068_n888_1), .B(_abc_19068_n893), .Y(_abc_19068_n913_1) );
  OR2X2 OR2X2_80 ( .A(_abc_19068_n1061), .B(_abc_19068_n1072_1), .Y(_abc_19068_n1073) );
  OR2X2 OR2X2_800 ( .A(core_v0_reg_18_), .B(core_v1_reg_18_), .Y(core__abc_21380_n1594) );
  OR2X2 OR2X2_801 ( .A(core_v3_reg_18_), .B(core_v2_reg_18_), .Y(core__abc_21380_n1600) );
  OR2X2 OR2X2_802 ( .A(core__abc_21380_n1597), .B(core__abc_21380_n1601), .Y(core__abc_21380_n1602) );
  OR2X2 OR2X2_803 ( .A(core__abc_21380_n1604), .B(core__abc_21380_n1603), .Y(core__abc_21380_n1605) );
  OR2X2 OR2X2_804 ( .A(core__abc_21380_n1606), .B(core__abc_21380_n1134_1_bF_buf4), .Y(core__abc_21380_n1607) );
  OR2X2 OR2X2_805 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_82_), .Y(core__abc_21380_n1608) );
  OR2X2 OR2X2_806 ( .A(core_v0_reg_19_), .B(core_v1_reg_19_), .Y(core__abc_21380_n1613) );
  OR2X2 OR2X2_807 ( .A(core_v2_reg_19_), .B(core_v3_reg_19_), .Y(core__abc_21380_n1617) );
  OR2X2 OR2X2_808 ( .A(core__abc_21380_n1620), .B(core__abc_21380_n1622), .Y(core__abc_21380_n1623) );
  OR2X2 OR2X2_809 ( .A(core__abc_21380_n1623), .B(core__abc_21380_n1134_1_bF_buf3), .Y(core__abc_21380_n1624) );
  OR2X2 OR2X2_81 ( .A(_abc_19068_n1075_1), .B(_abc_19068_n1076), .Y(_abc_19068_n1077_1) );
  OR2X2 OR2X2_810 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_83_), .Y(core__abc_21380_n1625) );
  OR2X2 OR2X2_811 ( .A(core__abc_21380_n1630), .B(core__abc_21380_n1631), .Y(core__abc_21380_n1632) );
  OR2X2 OR2X2_812 ( .A(core_v3_reg_20_), .B(core_v2_reg_20_), .Y(core__abc_21380_n1636) );
  OR2X2 OR2X2_813 ( .A(core__abc_21380_n1633), .B(core__abc_21380_n1637), .Y(core__abc_21380_n1638) );
  OR2X2 OR2X2_814 ( .A(core__abc_21380_n1639), .B(core__abc_21380_n1632), .Y(core__abc_21380_n1640) );
  OR2X2 OR2X2_815 ( .A(core__abc_21380_n1641), .B(core__abc_21380_n1134_1_bF_buf2), .Y(core__abc_21380_n1642) );
  OR2X2 OR2X2_816 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_84_), .Y(core__abc_21380_n1643) );
  OR2X2 OR2X2_817 ( .A(core__abc_21380_n1648), .B(core__abc_21380_n1649_1), .Y(core__abc_21380_n1650) );
  OR2X2 OR2X2_818 ( .A(core_v3_reg_21_), .B(core_v2_reg_21_), .Y(core__abc_21380_n1654) );
  OR2X2 OR2X2_819 ( .A(core__abc_21380_n1651), .B(core__abc_21380_n1655_1), .Y(core__abc_21380_n1656) );
  OR2X2 OR2X2_82 ( .A(_abc_19068_n1078_1), .B(_abc_19068_n1079), .Y(_abc_19068_n1080_1) );
  OR2X2 OR2X2_820 ( .A(core__abc_21380_n1657), .B(core__abc_21380_n1650), .Y(core__abc_21380_n1658) );
  OR2X2 OR2X2_821 ( .A(core__abc_21380_n1659), .B(core__abc_21380_n1134_1_bF_buf1), .Y(core__abc_21380_n1660) );
  OR2X2 OR2X2_822 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_85_), .Y(core__abc_21380_n1661) );
  OR2X2 OR2X2_823 ( .A(core__abc_21380_n1666), .B(core__abc_21380_n1667), .Y(core__abc_21380_n1668) );
  OR2X2 OR2X2_824 ( .A(core_v3_reg_22_), .B(core_v2_reg_22_), .Y(core__abc_21380_n1672) );
  OR2X2 OR2X2_825 ( .A(core__abc_21380_n1669), .B(core__abc_21380_n1673), .Y(core__abc_21380_n1674) );
  OR2X2 OR2X2_826 ( .A(core__abc_21380_n1675), .B(core__abc_21380_n1668), .Y(core__abc_21380_n1676) );
  OR2X2 OR2X2_827 ( .A(core__abc_21380_n1677), .B(core__abc_21380_n1134_1_bF_buf0), .Y(core__abc_21380_n1678) );
  OR2X2 OR2X2_828 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_86_), .Y(core__abc_21380_n1679) );
  OR2X2 OR2X2_829 ( .A(core_v3_reg_23_), .B(core_v2_reg_23_), .Y(core__abc_21380_n1691) );
  OR2X2 OR2X2_83 ( .A(_abc_19068_n1077_1), .B(_abc_19068_n1080_1), .Y(_abc_19068_n1081_1) );
  OR2X2 OR2X2_830 ( .A(core__abc_21380_n1688), .B(core__abc_21380_n1692), .Y(core__abc_21380_n1693) );
  OR2X2 OR2X2_831 ( .A(core__abc_21380_n1694), .B(core__abc_21380_n1695), .Y(core__abc_21380_n1696) );
  OR2X2 OR2X2_832 ( .A(core__abc_21380_n1697), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n1698) );
  OR2X2 OR2X2_833 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_87_), .Y(core__abc_21380_n1699) );
  OR2X2 OR2X2_834 ( .A(core__abc_21380_n1704), .B(core__abc_21380_n1705), .Y(core__abc_21380_n1706) );
  OR2X2 OR2X2_835 ( .A(core_v3_reg_24_), .B(core_v2_reg_24_), .Y(core__abc_21380_n1710) );
  OR2X2 OR2X2_836 ( .A(core__abc_21380_n1707), .B(core__abc_21380_n1711), .Y(core__abc_21380_n1712) );
  OR2X2 OR2X2_837 ( .A(core__abc_21380_n1713), .B(core__abc_21380_n1706), .Y(core__abc_21380_n1714) );
  OR2X2 OR2X2_838 ( .A(core__abc_21380_n1715), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n1716) );
  OR2X2 OR2X2_839 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_88_), .Y(core__abc_21380_n1717) );
  OR2X2 OR2X2_84 ( .A(_abc_19068_n1082), .B(_abc_19068_n1083_1), .Y(_abc_19068_n1084_1) );
  OR2X2 OR2X2_840 ( .A(core_v3_reg_25_), .B(core_v2_reg_25_), .Y(core__abc_21380_n1729) );
  OR2X2 OR2X2_841 ( .A(core__abc_21380_n1726), .B(core__abc_21380_n1730), .Y(core__abc_21380_n1731) );
  OR2X2 OR2X2_842 ( .A(core__abc_21380_n1732), .B(core__abc_21380_n1733), .Y(core__abc_21380_n1734) );
  OR2X2 OR2X2_843 ( .A(core__abc_21380_n1735), .B(core__abc_21380_n1134_1_bF_buf5), .Y(core__abc_21380_n1736) );
  OR2X2 OR2X2_844 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_89_), .Y(core__abc_21380_n1737) );
  OR2X2 OR2X2_845 ( .A(core_v0_reg_26_), .B(core_v1_reg_26_), .Y(core__abc_21380_n1740) );
  OR2X2 OR2X2_846 ( .A(core_v3_reg_26_), .B(core_v2_reg_26_), .Y(core__abc_21380_n1746) );
  OR2X2 OR2X2_847 ( .A(core__abc_21380_n1743), .B(core__abc_21380_n1747), .Y(core__abc_21380_n1748) );
  OR2X2 OR2X2_848 ( .A(core__abc_21380_n1749), .B(core__abc_21380_n1750), .Y(core__abc_21380_n1751) );
  OR2X2 OR2X2_849 ( .A(core__abc_21380_n1752), .B(core__abc_21380_n1134_1_bF_buf4), .Y(core__abc_21380_n1753) );
  OR2X2 OR2X2_85 ( .A(_abc_19068_n1085), .B(_abc_19068_n906_1), .Y(_abc_19068_n1086_1) );
  OR2X2 OR2X2_850 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_90_), .Y(core__abc_21380_n1754_1) );
  OR2X2 OR2X2_851 ( .A(core_v3_reg_27_), .B(core_v2_reg_27_), .Y(core__abc_21380_n1766) );
  OR2X2 OR2X2_852 ( .A(core__abc_21380_n1763), .B(core__abc_21380_n1767), .Y(core__abc_21380_n1768) );
  OR2X2 OR2X2_853 ( .A(core__abc_21380_n1769), .B(core__abc_21380_n1770), .Y(core__abc_21380_n1771) );
  OR2X2 OR2X2_854 ( .A(core__abc_21380_n1772), .B(core__abc_21380_n1134_1_bF_buf3), .Y(core__abc_21380_n1773) );
  OR2X2 OR2X2_855 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_91_), .Y(core__abc_21380_n1774) );
  OR2X2 OR2X2_856 ( .A(core__abc_21380_n1779), .B(core__abc_21380_n1780), .Y(core__abc_21380_n1781) );
  OR2X2 OR2X2_857 ( .A(core_v3_reg_28_), .B(core_v2_reg_28_), .Y(core__abc_21380_n1785) );
  OR2X2 OR2X2_858 ( .A(core__abc_21380_n1782_1), .B(core__abc_21380_n1786_1), .Y(core__abc_21380_n1787) );
  OR2X2 OR2X2_859 ( .A(core__abc_21380_n1788), .B(core__abc_21380_n1781), .Y(core__abc_21380_n1789) );
  OR2X2 OR2X2_86 ( .A(_abc_19068_n1084_1), .B(_abc_19068_n1086_1), .Y(_abc_19068_n1087_1) );
  OR2X2 OR2X2_860 ( .A(core__abc_21380_n1790), .B(core__abc_21380_n1134_1_bF_buf2), .Y(core__abc_21380_n1791) );
  OR2X2 OR2X2_861 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_92_), .Y(core__abc_21380_n1792) );
  OR2X2 OR2X2_862 ( .A(core_v3_reg_29_), .B(core_v2_reg_29_), .Y(core__abc_21380_n1804) );
  OR2X2 OR2X2_863 ( .A(core__abc_21380_n1801), .B(core__abc_21380_n1805), .Y(core__abc_21380_n1806) );
  OR2X2 OR2X2_864 ( .A(core__abc_21380_n1807), .B(core__abc_21380_n1808), .Y(core__abc_21380_n1809) );
  OR2X2 OR2X2_865 ( .A(core__abc_21380_n1810), .B(core__abc_21380_n1134_1_bF_buf1), .Y(core__abc_21380_n1811) );
  OR2X2 OR2X2_866 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_93_), .Y(core__abc_21380_n1812_1) );
  OR2X2 OR2X2_867 ( .A(core__abc_21380_n1817), .B(core__abc_21380_n1818), .Y(core__abc_21380_n1819) );
  OR2X2 OR2X2_868 ( .A(core_v3_reg_30_), .B(core_v2_reg_30_), .Y(core__abc_21380_n1823) );
  OR2X2 OR2X2_869 ( .A(core__abc_21380_n1820), .B(core__abc_21380_n1824), .Y(core__abc_21380_n1825) );
  OR2X2 OR2X2_87 ( .A(_abc_19068_n1081_1), .B(_abc_19068_n1087_1), .Y(_abc_19068_n1088) );
  OR2X2 OR2X2_870 ( .A(core__abc_21380_n1826), .B(core__abc_21380_n1819), .Y(core__abc_21380_n1827) );
  OR2X2 OR2X2_871 ( .A(core__abc_21380_n1828), .B(core__abc_21380_n1134_1_bF_buf0), .Y(core__abc_21380_n1829) );
  OR2X2 OR2X2_872 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_94_), .Y(core__abc_21380_n1830) );
  OR2X2 OR2X2_873 ( .A(core_v3_reg_31_), .B(core_v2_reg_31_), .Y(core__abc_21380_n1842) );
  OR2X2 OR2X2_874 ( .A(core__abc_21380_n1839), .B(core__abc_21380_n1843), .Y(core__abc_21380_n1844) );
  OR2X2 OR2X2_875 ( .A(core__abc_21380_n1845), .B(core__abc_21380_n1846_1), .Y(core__abc_21380_n1847) );
  OR2X2 OR2X2_876 ( .A(core__abc_21380_n1848), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n1849) );
  OR2X2 OR2X2_877 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_95_), .Y(core__abc_21380_n1850) );
  OR2X2 OR2X2_878 ( .A(core__abc_21380_n1855), .B(core__abc_21380_n1856), .Y(core__abc_21380_n1857) );
  OR2X2 OR2X2_879 ( .A(core_v3_reg_32_), .B(core_v2_reg_32_), .Y(core__abc_21380_n1861) );
  OR2X2 OR2X2_88 ( .A(_abc_19068_n1089_1), .B(_abc_19068_n1090_1), .Y(_abc_19068_n1091) );
  OR2X2 OR2X2_880 ( .A(core__abc_21380_n1858), .B(core__abc_21380_n1862), .Y(core__abc_21380_n1863) );
  OR2X2 OR2X2_881 ( .A(core__abc_21380_n1864), .B(core__abc_21380_n1857), .Y(core__abc_21380_n1865) );
  OR2X2 OR2X2_882 ( .A(core__abc_21380_n1866), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n1867) );
  OR2X2 OR2X2_883 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_96_), .Y(core__abc_21380_n1868) );
  OR2X2 OR2X2_884 ( .A(core__abc_21380_n1873), .B(core__abc_21380_n1874), .Y(core__abc_21380_n1875) );
  OR2X2 OR2X2_885 ( .A(core_v3_reg_33_), .B(core_v2_reg_33_), .Y(core__abc_21380_n1879) );
  OR2X2 OR2X2_886 ( .A(core__abc_21380_n1876), .B(core__abc_21380_n1880), .Y(core__abc_21380_n1881) );
  OR2X2 OR2X2_887 ( .A(core__abc_21380_n1882), .B(core__abc_21380_n1875), .Y(core__abc_21380_n1883) );
  OR2X2 OR2X2_888 ( .A(core__abc_21380_n1884), .B(core__abc_21380_n1134_1_bF_buf5), .Y(core__abc_21380_n1885) );
  OR2X2 OR2X2_889 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_97_), .Y(core__abc_21380_n1886) );
  OR2X2 OR2X2_89 ( .A(_abc_19068_n1092_1), .B(_abc_19068_n1093_1), .Y(_abc_19068_n1094) );
  OR2X2 OR2X2_890 ( .A(core__abc_21380_n1891), .B(core__abc_21380_n1892), .Y(core__abc_21380_n1893) );
  OR2X2 OR2X2_891 ( .A(core_v3_reg_34_), .B(core_v2_reg_34_), .Y(core__abc_21380_n1897) );
  OR2X2 OR2X2_892 ( .A(core__abc_21380_n1894_1), .B(core__abc_21380_n1898), .Y(core__abc_21380_n1899) );
  OR2X2 OR2X2_893 ( .A(core__abc_21380_n1900), .B(core__abc_21380_n1893), .Y(core__abc_21380_n1901) );
  OR2X2 OR2X2_894 ( .A(core__abc_21380_n1902), .B(core__abc_21380_n1134_1_bF_buf4), .Y(core__abc_21380_n1903) );
  OR2X2 OR2X2_895 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_98_), .Y(core__abc_21380_n1904) );
  OR2X2 OR2X2_896 ( .A(core_v3_reg_35_), .B(core_v2_reg_35_), .Y(core__abc_21380_n1916) );
  OR2X2 OR2X2_897 ( .A(core__abc_21380_n1913), .B(core__abc_21380_n1917), .Y(core__abc_21380_n1918) );
  OR2X2 OR2X2_898 ( .A(core__abc_21380_n1919), .B(core__abc_21380_n1920), .Y(core__abc_21380_n1921) );
  OR2X2 OR2X2_899 ( .A(core__abc_21380_n1922), .B(core__abc_21380_n1134_1_bF_buf3), .Y(core__abc_21380_n1923) );
  OR2X2 OR2X2_9 ( .A(_abc_19068_n915_1_bF_buf4), .B(_abc_19068_n916_1_bF_buf4), .Y(_abc_19068_n917) );
  OR2X2 OR2X2_90 ( .A(_abc_19068_n1091), .B(_abc_19068_n1094), .Y(_abc_19068_n1095_1) );
  OR2X2 OR2X2_900 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_99_), .Y(core__abc_21380_n1924) );
  OR2X2 OR2X2_901 ( .A(core__abc_21380_n1930), .B(core__abc_21380_n1927), .Y(core__abc_21380_n1931) );
  OR2X2 OR2X2_902 ( .A(core_v3_reg_36_), .B(core_v2_reg_36_), .Y(core__abc_21380_n1934_1) );
  OR2X2 OR2X2_903 ( .A(core__abc_21380_n1939), .B(core__abc_21380_n1936), .Y(core__abc_21380_n1940) );
  OR2X2 OR2X2_904 ( .A(core__abc_21380_n1940), .B(core__abc_21380_n1134_1_bF_buf2), .Y(core__abc_21380_n1941) );
  OR2X2 OR2X2_905 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_100_), .Y(core__abc_21380_n1942) );
  OR2X2 OR2X2_906 ( .A(core_v3_reg_37_), .B(core_v2_reg_37_), .Y(core__abc_21380_n1954) );
  OR2X2 OR2X2_907 ( .A(core__abc_21380_n1959), .B(core__abc_21380_n1957), .Y(core__abc_21380_n1960) );
  OR2X2 OR2X2_908 ( .A(core__abc_21380_n1960), .B(core__abc_21380_n1134_1_bF_buf1), .Y(core__abc_21380_n1961_1) );
  OR2X2 OR2X2_909 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_101_), .Y(core__abc_21380_n1962) );
  OR2X2 OR2X2_91 ( .A(_abc_19068_n1088), .B(_abc_19068_n1095_1), .Y(_abc_19068_n1096_1) );
  OR2X2 OR2X2_910 ( .A(core__abc_21380_n1967), .B(core__abc_21380_n1968), .Y(core__abc_21380_n1969) );
  OR2X2 OR2X2_911 ( .A(core_v3_reg_38_), .B(core_v2_reg_38_), .Y(core__abc_21380_n1973) );
  OR2X2 OR2X2_912 ( .A(core__abc_21380_n1970), .B(core__abc_21380_n1974), .Y(core__abc_21380_n1975) );
  OR2X2 OR2X2_913 ( .A(core__abc_21380_n1976), .B(core__abc_21380_n1969), .Y(core__abc_21380_n1977) );
  OR2X2 OR2X2_914 ( .A(core__abc_21380_n1978), .B(core__abc_21380_n1134_1_bF_buf0), .Y(core__abc_21380_n1979) );
  OR2X2 OR2X2_915 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_102_), .Y(core__abc_21380_n1980) );
  OR2X2 OR2X2_916 ( .A(core_v3_reg_39_), .B(core_v2_reg_39_), .Y(core__abc_21380_n1992) );
  OR2X2 OR2X2_917 ( .A(core__abc_21380_n1989), .B(core__abc_21380_n1993), .Y(core__abc_21380_n1994) );
  OR2X2 OR2X2_918 ( .A(core__abc_21380_n1995_1), .B(core__abc_21380_n1996), .Y(core__abc_21380_n1997) );
  OR2X2 OR2X2_919 ( .A(core__abc_21380_n1998), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n1999) );
  OR2X2 OR2X2_92 ( .A(_abc_19068_n1098_1), .B(_abc_19068_n1099_1), .Y(_abc_19068_n1100) );
  OR2X2 OR2X2_920 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_103_), .Y(core__abc_21380_n2000) );
  OR2X2 OR2X2_921 ( .A(core__abc_21380_n2006), .B(core__abc_21380_n2003), .Y(core__abc_21380_n2007) );
  OR2X2 OR2X2_922 ( .A(core_v3_reg_40_), .B(core_v2_reg_40_), .Y(core__abc_21380_n2011) );
  OR2X2 OR2X2_923 ( .A(core__abc_21380_n2014), .B(core__abc_21380_n2015), .Y(core__abc_21380_n2016) );
  OR2X2 OR2X2_924 ( .A(core__abc_21380_n2016), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n2017) );
  OR2X2 OR2X2_925 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_104_), .Y(core__abc_21380_n2018) );
  OR2X2 OR2X2_926 ( .A(core__abc_21380_n2024), .B(core__abc_21380_n2021), .Y(core__abc_21380_n2025) );
  OR2X2 OR2X2_927 ( .A(core_v3_reg_41_), .B(core_v2_reg_41_), .Y(core__abc_21380_n2028) );
  OR2X2 OR2X2_928 ( .A(core__abc_21380_n2033), .B(core__abc_21380_n2030), .Y(core__abc_21380_n2034) );
  OR2X2 OR2X2_929 ( .A(core__abc_21380_n2034), .B(core__abc_21380_n1134_1_bF_buf5), .Y(core__abc_21380_n2035_1) );
  OR2X2 OR2X2_93 ( .A(_abc_19068_n1101_1), .B(_abc_19068_n1102_1), .Y(_abc_19068_n1103) );
  OR2X2 OR2X2_930 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_105_), .Y(core__abc_21380_n2036) );
  OR2X2 OR2X2_931 ( .A(core__abc_21380_n2041), .B(core__abc_21380_n2042), .Y(core__abc_21380_n2043) );
  OR2X2 OR2X2_932 ( .A(core_v3_reg_42_), .B(core_v2_reg_42_), .Y(core__abc_21380_n2047) );
  OR2X2 OR2X2_933 ( .A(core__abc_21380_n2044), .B(core__abc_21380_n2048), .Y(core__abc_21380_n2049) );
  OR2X2 OR2X2_934 ( .A(core__abc_21380_n2050), .B(core__abc_21380_n2043), .Y(core__abc_21380_n2051) );
  OR2X2 OR2X2_935 ( .A(core__abc_21380_n2052), .B(core__abc_21380_n1134_1_bF_buf4), .Y(core__abc_21380_n2053) );
  OR2X2 OR2X2_936 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_106_), .Y(core__abc_21380_n2054) );
  OR2X2 OR2X2_937 ( .A(core_v3_reg_43_), .B(core_v2_reg_43_), .Y(core__abc_21380_n2064) );
  OR2X2 OR2X2_938 ( .A(core__abc_21380_n2063), .B(core__abc_21380_n2067_1), .Y(core__abc_21380_n2068) );
  OR2X2 OR2X2_939 ( .A(core__abc_21380_n2069), .B(core__abc_21380_n2070), .Y(core__abc_21380_n2071) );
  OR2X2 OR2X2_94 ( .A(_abc_19068_n1100), .B(_abc_19068_n1103), .Y(_abc_19068_n1104_1) );
  OR2X2 OR2X2_940 ( .A(core__abc_21380_n2072), .B(core__abc_21380_n1134_1_bF_buf3), .Y(core__abc_21380_n2073_1) );
  OR2X2 OR2X2_941 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_107_), .Y(core__abc_21380_n2074) );
  OR2X2 OR2X2_942 ( .A(core__abc_21380_n2080), .B(core__abc_21380_n2077), .Y(core__abc_21380_n2081) );
  OR2X2 OR2X2_943 ( .A(core_v2_reg_44_), .B(core_v3_reg_44_), .Y(core__abc_21380_n2082) );
  OR2X2 OR2X2_944 ( .A(core__abc_21380_n2089), .B(core__abc_21380_n2086), .Y(core__abc_21380_n2090) );
  OR2X2 OR2X2_945 ( .A(core__abc_21380_n2090), .B(core__abc_21380_n1134_1_bF_buf2), .Y(core__abc_21380_n2091) );
  OR2X2 OR2X2_946 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_108_), .Y(core__abc_21380_n2092) );
  OR2X2 OR2X2_947 ( .A(core_v3_reg_45_), .B(core_v2_reg_45_), .Y(core__abc_21380_n2102) );
  OR2X2 OR2X2_948 ( .A(core__abc_21380_n2101), .B(core__abc_21380_n2105), .Y(core__abc_21380_n2106) );
  OR2X2 OR2X2_949 ( .A(core__abc_21380_n2107), .B(core__abc_21380_n2108), .Y(core__abc_21380_n2109) );
  OR2X2 OR2X2_95 ( .A(_abc_19068_n1106), .B(_abc_19068_n1107_1), .Y(_abc_19068_n1108_1) );
  OR2X2 OR2X2_950 ( .A(core__abc_21380_n2110), .B(core__abc_21380_n1134_1_bF_buf1), .Y(core__abc_21380_n2111) );
  OR2X2 OR2X2_951 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_109_), .Y(core__abc_21380_n2112) );
  OR2X2 OR2X2_952 ( .A(core__abc_21380_n2118), .B(core__abc_21380_n2115), .Y(core__abc_21380_n2119) );
  OR2X2 OR2X2_953 ( .A(core_v2_reg_46_), .B(core_v3_reg_46_), .Y(core__abc_21380_n2120) );
  OR2X2 OR2X2_954 ( .A(core__abc_21380_n2127), .B(core__abc_21380_n2124), .Y(core__abc_21380_n2128) );
  OR2X2 OR2X2_955 ( .A(core__abc_21380_n2128), .B(core__abc_21380_n1134_1_bF_buf0), .Y(core__abc_21380_n2129) );
  OR2X2 OR2X2_956 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_110_), .Y(core__abc_21380_n2130) );
  OR2X2 OR2X2_957 ( .A(core_v2_reg_47_), .B(core_v3_reg_47_), .Y(core__abc_21380_n2141) );
  OR2X2 OR2X2_958 ( .A(core__abc_21380_n2145), .B(core__abc_21380_n2147), .Y(core__abc_21380_n2148) );
  OR2X2 OR2X2_959 ( .A(core__abc_21380_n2148), .B(core__abc_21380_n1134_1_bF_buf7), .Y(core__abc_21380_n2149) );
  OR2X2 OR2X2_96 ( .A(_abc_19068_n1108_1), .B(_abc_19068_n1105_1), .Y(_abc_19068_n1109) );
  OR2X2 OR2X2_960 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_111_), .Y(core__abc_21380_n2150) );
  OR2X2 OR2X2_961 ( .A(core__abc_21380_n2155), .B(core__abc_21380_n2156), .Y(core__abc_21380_n2157) );
  OR2X2 OR2X2_962 ( .A(core_v2_reg_48_), .B(core_v3_reg_48_), .Y(core__abc_21380_n2159) );
  OR2X2 OR2X2_963 ( .A(core__abc_21380_n2158), .B(core__abc_21380_n2162), .Y(core__abc_21380_n2163) );
  OR2X2 OR2X2_964 ( .A(core__abc_21380_n2164), .B(core__abc_21380_n2157), .Y(core__abc_21380_n2165) );
  OR2X2 OR2X2_965 ( .A(core__abc_21380_n2166), .B(core__abc_21380_n1134_1_bF_buf6), .Y(core__abc_21380_n2167) );
  OR2X2 OR2X2_966 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_112_), .Y(core__abc_21380_n2168) );
  OR2X2 OR2X2_967 ( .A(core__abc_21380_n2174), .B(core__abc_21380_n2171), .Y(core__abc_21380_n2175) );
  OR2X2 OR2X2_968 ( .A(core_v2_reg_49_), .B(core_v3_reg_49_), .Y(core__abc_21380_n2176) );
  OR2X2 OR2X2_969 ( .A(core__abc_21380_n2183), .B(core__abc_21380_n2180), .Y(core__abc_21380_n2184) );
  OR2X2 OR2X2_97 ( .A(_abc_19068_n1110_1), .B(_abc_19068_n1111_1), .Y(_abc_19068_n1112) );
  OR2X2 OR2X2_970 ( .A(core__abc_21380_n2184), .B(core__abc_21380_n1134_1_bF_buf5), .Y(core__abc_21380_n2185_1) );
  OR2X2 OR2X2_971 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_113_), .Y(core__abc_21380_n2186) );
  OR2X2 OR2X2_972 ( .A(core__abc_21380_n2192), .B(core__abc_21380_n2189), .Y(core__abc_21380_n2193) );
  OR2X2 OR2X2_973 ( .A(core_v2_reg_50_), .B(core_v3_reg_50_), .Y(core__abc_21380_n2194) );
  OR2X2 OR2X2_974 ( .A(core__abc_21380_n2201), .B(core__abc_21380_n2198), .Y(core__abc_21380_n2202) );
  OR2X2 OR2X2_975 ( .A(core__abc_21380_n2202), .B(core__abc_21380_n1134_1_bF_buf4), .Y(core__abc_21380_n2203) );
  OR2X2 OR2X2_976 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_114_), .Y(core__abc_21380_n2204) );
  OR2X2 OR2X2_977 ( .A(core_v3_reg_51_), .B(core_v2_reg_51_), .Y(core__abc_21380_n2215) );
  OR2X2 OR2X2_978 ( .A(core__abc_21380_n2219_1), .B(core__abc_21380_n2221), .Y(core__abc_21380_n2222) );
  OR2X2 OR2X2_979 ( .A(core__abc_21380_n2222), .B(core__abc_21380_n1134_1_bF_buf3), .Y(core__abc_21380_n2223) );
  OR2X2 OR2X2_98 ( .A(_abc_19068_n1113_1), .B(_abc_19068_n1114_1), .Y(_abc_19068_n1115) );
  OR2X2 OR2X2_980 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_115_), .Y(core__abc_21380_n2224) );
  OR2X2 OR2X2_981 ( .A(core_v0_reg_52_), .B(core_v1_reg_52_), .Y(core__abc_21380_n2227) );
  OR2X2 OR2X2_982 ( .A(core_v3_reg_52_), .B(core_v2_reg_52_), .Y(core__abc_21380_n2231) );
  OR2X2 OR2X2_983 ( .A(core__abc_21380_n2230), .B(core__abc_21380_n2234), .Y(core__abc_21380_n2235) );
  OR2X2 OR2X2_984 ( .A(core__abc_21380_n2236), .B(core__abc_21380_n2237), .Y(core__abc_21380_n2238) );
  OR2X2 OR2X2_985 ( .A(core__abc_21380_n2239), .B(core__abc_21380_n1134_1_bF_buf2), .Y(core__abc_21380_n2240) );
  OR2X2 OR2X2_986 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_116_), .Y(core__abc_21380_n2241) );
  OR2X2 OR2X2_987 ( .A(core_v3_reg_53_), .B(core_v2_reg_53_), .Y(core__abc_21380_n2252) );
  OR2X2 OR2X2_988 ( .A(core__abc_21380_n2256), .B(core__abc_21380_n2258), .Y(core__abc_21380_n2259) );
  OR2X2 OR2X2_989 ( .A(core__abc_21380_n2259), .B(core__abc_21380_n1134_1_bF_buf1), .Y(core__abc_21380_n2260) );
  OR2X2 OR2X2_99 ( .A(_abc_19068_n1112), .B(_abc_19068_n1115), .Y(_abc_19068_n1116_1) );
  OR2X2 OR2X2_990 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_117_), .Y(core__abc_21380_n2261) );
  OR2X2 OR2X2_991 ( .A(core__abc_21380_n2266), .B(core__abc_21380_n2267), .Y(core__abc_21380_n2268) );
  OR2X2 OR2X2_992 ( .A(core_v3_reg_54_), .B(core_v2_reg_54_), .Y(core__abc_21380_n2270) );
  OR2X2 OR2X2_993 ( .A(core__abc_21380_n2269), .B(core__abc_21380_n2273), .Y(core__abc_21380_n2274) );
  OR2X2 OR2X2_994 ( .A(core__abc_21380_n2275), .B(core__abc_21380_n2268), .Y(core__abc_21380_n2276) );
  OR2X2 OR2X2_995 ( .A(core__abc_21380_n2277), .B(core__abc_21380_n1134_1_bF_buf0), .Y(core__abc_21380_n2278) );
  OR2X2 OR2X2_996 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_118_), .Y(core__abc_21380_n2279) );
  OR2X2 OR2X2_997 ( .A(core_v3_reg_55_), .B(core_v2_reg_55_), .Y(core__abc_21380_n2289) );
  OR2X2 OR2X2_998 ( .A(core__abc_21380_n2288), .B(core__abc_21380_n2292), .Y(core__abc_21380_n2293) );
  OR2X2 OR2X2_999 ( .A(core__abc_21380_n2294_1), .B(core__abc_21380_n2295), .Y(core__abc_21380_n2296) );
endmodule
