module b14_reset(clock, RESET_G, nRESET_G, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_, ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_, ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_, ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_, DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_, DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_, DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_, DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_, DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_, DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_, DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_, DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG);
  output ADDR_REG_0_;
  output ADDR_REG_10_;
  output ADDR_REG_11_;
  output ADDR_REG_12_;
  output ADDR_REG_13_;
  output ADDR_REG_14_;
  output ADDR_REG_15_;
  output ADDR_REG_16_;
  output ADDR_REG_17_;
  output ADDR_REG_18_;
  output ADDR_REG_19_;
  output ADDR_REG_1_;
  output ADDR_REG_2_;
  output ADDR_REG_3_;
  output ADDR_REG_4_;
  output ADDR_REG_5_;
  output ADDR_REG_6_;
  output ADDR_REG_7_;
  output ADDR_REG_8_;
  output ADDR_REG_9_;
  wire B_REG;
  input DATAI_0_;
  input DATAI_10_;
  input DATAI_11_;
  input DATAI_12_;
  input DATAI_13_;
  input DATAI_14_;
  input DATAI_15_;
  input DATAI_16_;
  input DATAI_17_;
  input DATAI_18_;
  input DATAI_19_;
  input DATAI_1_;
  input DATAI_20_;
  input DATAI_21_;
  input DATAI_22_;
  input DATAI_23_;
  input DATAI_24_;
  input DATAI_25_;
  input DATAI_26_;
  input DATAI_27_;
  input DATAI_28_;
  input DATAI_29_;
  input DATAI_2_;
  input DATAI_30_;
  input DATAI_31_;
  input DATAI_3_;
  input DATAI_4_;
  input DATAI_5_;
  input DATAI_6_;
  input DATAI_7_;
  input DATAI_8_;
  input DATAI_9_;
  output DATAO_REG_0_;
  output DATAO_REG_10_;
  output DATAO_REG_11_;
  output DATAO_REG_12_;
  output DATAO_REG_13_;
  output DATAO_REG_14_;
  output DATAO_REG_15_;
  output DATAO_REG_16_;
  output DATAO_REG_17_;
  output DATAO_REG_18_;
  output DATAO_REG_19_;
  output DATAO_REG_1_;
  output DATAO_REG_20_;
  output DATAO_REG_21_;
  output DATAO_REG_22_;
  output DATAO_REG_23_;
  output DATAO_REG_24_;
  output DATAO_REG_25_;
  output DATAO_REG_26_;
  output DATAO_REG_27_;
  output DATAO_REG_28_;
  output DATAO_REG_29_;
  output DATAO_REG_2_;
  output DATAO_REG_30_;
  output DATAO_REG_31_;
  output DATAO_REG_3_;
  output DATAO_REG_4_;
  output DATAO_REG_5_;
  output DATAO_REG_6_;
  output DATAO_REG_7_;
  output DATAO_REG_8_;
  output DATAO_REG_9_;
  wire D_REG_0_;
  wire D_REG_10_;
  wire D_REG_11_;
  wire D_REG_12_;
  wire D_REG_13_;
  wire D_REG_14_;
  wire D_REG_15_;
  wire D_REG_16_;
  wire D_REG_17_;
  wire D_REG_18_;
  wire D_REG_19_;
  wire D_REG_1_;
  wire D_REG_20_;
  wire D_REG_21_;
  wire D_REG_22_;
  wire D_REG_23_;
  wire D_REG_24_;
  wire D_REG_25_;
  wire D_REG_26_;
  wire D_REG_27_;
  wire D_REG_28_;
  wire D_REG_29_;
  wire D_REG_2_;
  wire D_REG_30_;
  wire D_REG_31_;
  wire D_REG_3_;
  wire D_REG_4_;
  wire D_REG_5_;
  wire D_REG_6_;
  wire D_REG_7_;
  wire D_REG_8_;
  wire D_REG_9_;
  wire IR_REG_0_;
  wire IR_REG_10_;
  wire IR_REG_11_;
  wire IR_REG_12_;
  wire IR_REG_13_;
  wire IR_REG_14_;
  wire IR_REG_15_;
  wire IR_REG_16_;
  wire IR_REG_17_;
  wire IR_REG_18_;
  wire IR_REG_19_;
  wire IR_REG_1_;
  wire IR_REG_20_;
  wire IR_REG_21_;
  wire IR_REG_22_;
  wire IR_REG_23_;
  wire IR_REG_24_;
  wire IR_REG_25_;
  wire IR_REG_26_;
  wire IR_REG_27_;
  wire IR_REG_28_;
  wire IR_REG_29_;
  wire IR_REG_2_;
  wire IR_REG_30_;
  wire IR_REG_31_;
  wire IR_REG_31__bF_buf0;
  wire IR_REG_31__bF_buf1;
  wire IR_REG_31__bF_buf2;
  wire IR_REG_31__bF_buf3;
  wire IR_REG_31__bF_buf4;
  wire IR_REG_3_;
  wire IR_REG_4_;
  wire IR_REG_5_;
  wire IR_REG_6_;
  wire IR_REG_7_;
  wire IR_REG_8_;
  wire IR_REG_9_;
  output RD_REG;
  wire REG0_REG_0_;
  wire REG0_REG_10_;
  wire REG0_REG_11_;
  wire REG0_REG_12_;
  wire REG0_REG_13_;
  wire REG0_REG_14_;
  wire REG0_REG_15_;
  wire REG0_REG_16_;
  wire REG0_REG_17_;
  wire REG0_REG_18_;
  wire REG0_REG_19_;
  wire REG0_REG_1_;
  wire REG0_REG_20_;
  wire REG0_REG_21_;
  wire REG0_REG_22_;
  wire REG0_REG_23_;
  wire REG0_REG_24_;
  wire REG0_REG_25_;
  wire REG0_REG_26_;
  wire REG0_REG_27_;
  wire REG0_REG_28_;
  wire REG0_REG_29_;
  wire REG0_REG_2_;
  wire REG0_REG_30_;
  wire REG0_REG_31_;
  wire REG0_REG_3_;
  wire REG0_REG_4_;
  wire REG0_REG_5_;
  wire REG0_REG_6_;
  wire REG0_REG_7_;
  wire REG0_REG_8_;
  wire REG0_REG_9_;
  wire REG1_REG_0_;
  wire REG1_REG_10_;
  wire REG1_REG_11_;
  wire REG1_REG_12_;
  wire REG1_REG_13_;
  wire REG1_REG_14_;
  wire REG1_REG_15_;
  wire REG1_REG_16_;
  wire REG1_REG_17_;
  wire REG1_REG_18_;
  wire REG1_REG_19_;
  wire REG1_REG_1_;
  wire REG1_REG_20_;
  wire REG1_REG_21_;
  wire REG1_REG_22_;
  wire REG1_REG_23_;
  wire REG1_REG_24_;
  wire REG1_REG_25_;
  wire REG1_REG_26_;
  wire REG1_REG_27_;
  wire REG1_REG_28_;
  wire REG1_REG_29_;
  wire REG1_REG_2_;
  wire REG1_REG_30_;
  wire REG1_REG_31_;
  wire REG1_REG_3_;
  wire REG1_REG_4_;
  wire REG1_REG_5_;
  wire REG1_REG_6_;
  wire REG1_REG_7_;
  wire REG1_REG_8_;
  wire REG1_REG_9_;
  wire REG2_REG_0_;
  wire REG2_REG_10_;
  wire REG2_REG_11_;
  wire REG2_REG_12_;
  wire REG2_REG_13_;
  wire REG2_REG_14_;
  wire REG2_REG_15_;
  wire REG2_REG_16_;
  wire REG2_REG_17_;
  wire REG2_REG_18_;
  wire REG2_REG_19_;
  wire REG2_REG_1_;
  wire REG2_REG_20_;
  wire REG2_REG_21_;
  wire REG2_REG_22_;
  wire REG2_REG_23_;
  wire REG2_REG_24_;
  wire REG2_REG_25_;
  wire REG2_REG_26_;
  wire REG2_REG_27_;
  wire REG2_REG_28_;
  wire REG2_REG_29_;
  wire REG2_REG_2_;
  wire REG2_REG_30_;
  wire REG2_REG_31_;
  wire REG2_REG_3_;
  wire REG2_REG_4_;
  wire REG2_REG_5_;
  wire REG2_REG_6_;
  wire REG2_REG_7_;
  wire REG2_REG_8_;
  wire REG2_REG_9_;
  wire REG3_REG_0_;
  wire REG3_REG_10_;
  wire REG3_REG_11_;
  wire REG3_REG_12_;
  wire REG3_REG_13_;
  wire REG3_REG_14_;
  wire REG3_REG_15_;
  wire REG3_REG_16_;
  wire REG3_REG_17_;
  wire REG3_REG_18_;
  wire REG3_REG_19_;
  wire REG3_REG_1_;
  wire REG3_REG_20_;
  wire REG3_REG_21_;
  wire REG3_REG_22_;
  wire REG3_REG_23_;
  wire REG3_REG_24_;
  wire REG3_REG_25_;
  wire REG3_REG_26_;
  wire REG3_REG_27_;
  wire REG3_REG_28_;
  wire REG3_REG_2_;
  wire REG3_REG_3_;
  wire REG3_REG_4_;
  wire REG3_REG_5_;
  wire REG3_REG_6_;
  wire REG3_REG_7_;
  wire REG3_REG_8_;
  wire REG3_REG_9_;
  input RESET_G;
  wire STATE_REG;
  output WR_REG;
  wire _abc_40344_n1000;
  wire _abc_40344_n1001;
  wire _abc_40344_n1002;
  wire _abc_40344_n1003;
  wire _abc_40344_n1004;
  wire _abc_40344_n1005;
  wire _abc_40344_n1005_bF_buf0;
  wire _abc_40344_n1005_bF_buf1;
  wire _abc_40344_n1005_bF_buf2;
  wire _abc_40344_n1005_bF_buf3;
  wire _abc_40344_n1005_bF_buf4;
  wire _abc_40344_n1006;
  wire _abc_40344_n1007;
  wire _abc_40344_n1008;
  wire _abc_40344_n1009;
  wire _abc_40344_n1010;
  wire _abc_40344_n1011;
  wire _abc_40344_n1012;
  wire _abc_40344_n1013;
  wire _abc_40344_n1014;
  wire _abc_40344_n1015;
  wire _abc_40344_n1016;
  wire _abc_40344_n1017;
  wire _abc_40344_n1018;
  wire _abc_40344_n1019;
  wire _abc_40344_n1020;
  wire _abc_40344_n1021;
  wire _abc_40344_n1022;
  wire _abc_40344_n1023_1;
  wire _abc_40344_n1023_1_bF_buf0;
  wire _abc_40344_n1023_1_bF_buf1;
  wire _abc_40344_n1023_1_bF_buf2;
  wire _abc_40344_n1023_1_bF_buf3;
  wire _abc_40344_n1023_1_bF_buf4;
  wire _abc_40344_n1024;
  wire _abc_40344_n1025;
  wire _abc_40344_n1026;
  wire _abc_40344_n1027_1;
  wire _abc_40344_n1028;
  wire _abc_40344_n1029_1;
  wire _abc_40344_n1030_1;
  wire _abc_40344_n1031;
  wire _abc_40344_n1031_bF_buf0;
  wire _abc_40344_n1031_bF_buf1;
  wire _abc_40344_n1031_bF_buf2;
  wire _abc_40344_n1031_bF_buf3;
  wire _abc_40344_n1032;
  wire _abc_40344_n1032_bF_buf0;
  wire _abc_40344_n1032_bF_buf1;
  wire _abc_40344_n1032_bF_buf2;
  wire _abc_40344_n1032_bF_buf3;
  wire _abc_40344_n1032_bF_buf4;
  wire _abc_40344_n1033;
  wire _abc_40344_n1033_bF_buf0;
  wire _abc_40344_n1033_bF_buf1;
  wire _abc_40344_n1033_bF_buf2;
  wire _abc_40344_n1033_bF_buf3;
  wire _abc_40344_n1033_bF_buf4;
  wire _abc_40344_n1034_1;
  wire _abc_40344_n1035;
  wire _abc_40344_n1036;
  wire _abc_40344_n1037;
  wire _abc_40344_n1039;
  wire _abc_40344_n1040;
  wire _abc_40344_n1041;
  wire _abc_40344_n1042;
  wire _abc_40344_n1043;
  wire _abc_40344_n1044;
  wire _abc_40344_n1045_1;
  wire _abc_40344_n1046;
  wire _abc_40344_n1047;
  wire _abc_40344_n1048;
  wire _abc_40344_n1049_1;
  wire _abc_40344_n1050;
  wire _abc_40344_n1051_1;
  wire _abc_40344_n1052_1;
  wire _abc_40344_n1053;
  wire _abc_40344_n1054;
  wire _abc_40344_n1055;
  wire _abc_40344_n1056;
  wire _abc_40344_n1057;
  wire _abc_40344_n1058;
  wire _abc_40344_n1059;
  wire _abc_40344_n1060;
  wire _abc_40344_n1061;
  wire _abc_40344_n1062;
  wire _abc_40344_n1063;
  wire _abc_40344_n1064;
  wire _abc_40344_n1065;
  wire _abc_40344_n1066_1;
  wire _abc_40344_n1067;
  wire _abc_40344_n1068;
  wire _abc_40344_n1069;
  wire _abc_40344_n1070;
  wire _abc_40344_n1071;
  wire _abc_40344_n1072;
  wire _abc_40344_n1073;
  wire _abc_40344_n1074;
  wire _abc_40344_n1075;
  wire _abc_40344_n1076;
  wire _abc_40344_n1077;
  wire _abc_40344_n1078_1;
  wire _abc_40344_n1079;
  wire _abc_40344_n1080;
  wire _abc_40344_n1081;
  wire _abc_40344_n1082;
  wire _abc_40344_n1083;
  wire _abc_40344_n1084;
  wire _abc_40344_n1085;
  wire _abc_40344_n1086;
  wire _abc_40344_n1087;
  wire _abc_40344_n1088;
  wire _abc_40344_n1089;
  wire _abc_40344_n1090_1;
  wire _abc_40344_n1091;
  wire _abc_40344_n1092;
  wire _abc_40344_n1093;
  wire _abc_40344_n1094;
  wire _abc_40344_n1095;
  wire _abc_40344_n1096;
  wire _abc_40344_n1097;
  wire _abc_40344_n1098;
  wire _abc_40344_n1099;
  wire _abc_40344_n1100;
  wire _abc_40344_n1101;
  wire _abc_40344_n1102;
  wire _abc_40344_n1103_1;
  wire _abc_40344_n1104;
  wire _abc_40344_n1105;
  wire _abc_40344_n1106;
  wire _abc_40344_n1107;
  wire _abc_40344_n1108;
  wire _abc_40344_n1109;
  wire _abc_40344_n1110;
  wire _abc_40344_n1111;
  wire _abc_40344_n1112;
  wire _abc_40344_n1113;
  wire _abc_40344_n1114;
  wire _abc_40344_n1115;
  wire _abc_40344_n1116;
  wire _abc_40344_n1117;
  wire _abc_40344_n1118_1;
  wire _abc_40344_n1119;
  wire _abc_40344_n1120;
  wire _abc_40344_n1121;
  wire _abc_40344_n1122;
  wire _abc_40344_n1123;
  wire _abc_40344_n1124;
  wire _abc_40344_n1125;
  wire _abc_40344_n1126;
  wire _abc_40344_n1127;
  wire _abc_40344_n1128;
  wire _abc_40344_n1129;
  wire _abc_40344_n1130;
  wire _abc_40344_n1131;
  wire _abc_40344_n1132_1;
  wire _abc_40344_n1133;
  wire _abc_40344_n1134;
  wire _abc_40344_n1135_1;
  wire _abc_40344_n1136;
  wire _abc_40344_n1137;
  wire _abc_40344_n1138;
  wire _abc_40344_n1139;
  wire _abc_40344_n1140;
  wire _abc_40344_n1141;
  wire _abc_40344_n1142;
  wire _abc_40344_n1143;
  wire _abc_40344_n1144;
  wire _abc_40344_n1145;
  wire _abc_40344_n1146;
  wire _abc_40344_n1147;
  wire _abc_40344_n1148;
  wire _abc_40344_n1149;
  wire _abc_40344_n1150;
  wire _abc_40344_n1151;
  wire _abc_40344_n1152_1;
  wire _abc_40344_n1153;
  wire _abc_40344_n1154_1;
  wire _abc_40344_n1155_1;
  wire _abc_40344_n1156;
  wire _abc_40344_n1157;
  wire _abc_40344_n1158;
  wire _abc_40344_n1159;
  wire _abc_40344_n1160;
  wire _abc_40344_n1161;
  wire _abc_40344_n1162;
  wire _abc_40344_n1163;
  wire _abc_40344_n1164;
  wire _abc_40344_n1165;
  wire _abc_40344_n1166_1;
  wire _abc_40344_n1167;
  wire _abc_40344_n1168;
  wire _abc_40344_n1169;
  wire _abc_40344_n1170;
  wire _abc_40344_n1171;
  wire _abc_40344_n1172;
  wire _abc_40344_n1173;
  wire _abc_40344_n1174;
  wire _abc_40344_n1175;
  wire _abc_40344_n1176;
  wire _abc_40344_n1177;
  wire _abc_40344_n1178;
  wire _abc_40344_n1179;
  wire _abc_40344_n1180_1;
  wire _abc_40344_n1181;
  wire _abc_40344_n1182;
  wire _abc_40344_n1183;
  wire _abc_40344_n1184;
  wire _abc_40344_n1185;
  wire _abc_40344_n1186;
  wire _abc_40344_n1187;
  wire _abc_40344_n1188;
  wire _abc_40344_n1189;
  wire _abc_40344_n1190;
  wire _abc_40344_n1191;
  wire _abc_40344_n1192;
  wire _abc_40344_n1193_1;
  wire _abc_40344_n1194;
  wire _abc_40344_n1195;
  wire _abc_40344_n1196;
  wire _abc_40344_n1197;
  wire _abc_40344_n1198;
  wire _abc_40344_n1199;
  wire _abc_40344_n1200;
  wire _abc_40344_n1201;
  wire _abc_40344_n1202;
  wire _abc_40344_n1203;
  wire _abc_40344_n1204;
  wire _abc_40344_n1205;
  wire _abc_40344_n1206;
  wire _abc_40344_n1207;
  wire _abc_40344_n1208;
  wire _abc_40344_n1209_1;
  wire _abc_40344_n1210;
  wire _abc_40344_n1211;
  wire _abc_40344_n1212;
  wire _abc_40344_n1213;
  wire _abc_40344_n1214;
  wire _abc_40344_n1215;
  wire _abc_40344_n1216;
  wire _abc_40344_n1217;
  wire _abc_40344_n1218;
  wire _abc_40344_n1219;
  wire _abc_40344_n1220;
  wire _abc_40344_n1221;
  wire _abc_40344_n1222;
  wire _abc_40344_n1223;
  wire _abc_40344_n1224;
  wire _abc_40344_n1225_1;
  wire _abc_40344_n1226;
  wire _abc_40344_n1227;
  wire _abc_40344_n1228;
  wire _abc_40344_n1229;
  wire _abc_40344_n1230;
  wire _abc_40344_n1231;
  wire _abc_40344_n1232;
  wire _abc_40344_n1233;
  wire _abc_40344_n1234;
  wire _abc_40344_n1235;
  wire _abc_40344_n1236;
  wire _abc_40344_n1237;
  wire _abc_40344_n1238;
  wire _abc_40344_n1239;
  wire _abc_40344_n1240_1;
  wire _abc_40344_n1241;
  wire _abc_40344_n1242;
  wire _abc_40344_n1243;
  wire _abc_40344_n1244;
  wire _abc_40344_n1245;
  wire _abc_40344_n1246;
  wire _abc_40344_n1247;
  wire _abc_40344_n1248;
  wire _abc_40344_n1249;
  wire _abc_40344_n1250;
  wire _abc_40344_n1251;
  wire _abc_40344_n1252;
  wire _abc_40344_n1253;
  wire _abc_40344_n1254_1;
  wire _abc_40344_n1255;
  wire _abc_40344_n1256;
  wire _abc_40344_n1257;
  wire _abc_40344_n1258;
  wire _abc_40344_n1259;
  wire _abc_40344_n1260;
  wire _abc_40344_n1261;
  wire _abc_40344_n1262;
  wire _abc_40344_n1263;
  wire _abc_40344_n1264;
  wire _abc_40344_n1265_1;
  wire _abc_40344_n1266;
  wire _abc_40344_n1267;
  wire _abc_40344_n1268;
  wire _abc_40344_n1269;
  wire _abc_40344_n1270;
  wire _abc_40344_n1271;
  wire _abc_40344_n1272;
  wire _abc_40344_n1273;
  wire _abc_40344_n1274;
  wire _abc_40344_n1275;
  wire _abc_40344_n1276;
  wire _abc_40344_n1277;
  wire _abc_40344_n1278;
  wire _abc_40344_n1279;
  wire _abc_40344_n1280;
  wire _abc_40344_n1281;
  wire _abc_40344_n1282_1;
  wire _abc_40344_n1283;
  wire _abc_40344_n1284;
  wire _abc_40344_n1285;
  wire _abc_40344_n1286;
  wire _abc_40344_n1287;
  wire _abc_40344_n1288;
  wire _abc_40344_n1289;
  wire _abc_40344_n1290;
  wire _abc_40344_n1291;
  wire _abc_40344_n1292;
  wire _abc_40344_n1293_1;
  wire _abc_40344_n1294;
  wire _abc_40344_n1295;
  wire _abc_40344_n1296;
  wire _abc_40344_n1297;
  wire _abc_40344_n1298;
  wire _abc_40344_n1299;
  wire _abc_40344_n1300;
  wire _abc_40344_n1301;
  wire _abc_40344_n1302;
  wire _abc_40344_n1303;
  wire _abc_40344_n1304_1;
  wire _abc_40344_n1305;
  wire _abc_40344_n1306;
  wire _abc_40344_n1307;
  wire _abc_40344_n1308;
  wire _abc_40344_n1309;
  wire _abc_40344_n1310;
  wire _abc_40344_n1311;
  wire _abc_40344_n1312;
  wire _abc_40344_n1313;
  wire _abc_40344_n1314;
  wire _abc_40344_n1315;
  wire _abc_40344_n1316;
  wire _abc_40344_n1317_1;
  wire _abc_40344_n1318;
  wire _abc_40344_n1319;
  wire _abc_40344_n1320;
  wire _abc_40344_n1321;
  wire _abc_40344_n1322;
  wire _abc_40344_n1323;
  wire _abc_40344_n1324;
  wire _abc_40344_n1325;
  wire _abc_40344_n1326;
  wire _abc_40344_n1327;
  wire _abc_40344_n1328;
  wire _abc_40344_n1329;
  wire _abc_40344_n1330;
  wire _abc_40344_n1331_1;
  wire _abc_40344_n1332;
  wire _abc_40344_n1333;
  wire _abc_40344_n1334;
  wire _abc_40344_n1335;
  wire _abc_40344_n1336;
  wire _abc_40344_n1337;
  wire _abc_40344_n1338;
  wire _abc_40344_n1339;
  wire _abc_40344_n1340;
  wire _abc_40344_n1341;
  wire _abc_40344_n1342;
  wire _abc_40344_n1343_1;
  wire _abc_40344_n1344;
  wire _abc_40344_n1345;
  wire _abc_40344_n1346;
  wire _abc_40344_n1347;
  wire _abc_40344_n1348;
  wire _abc_40344_n1349;
  wire _abc_40344_n1350;
  wire _abc_40344_n1351;
  wire _abc_40344_n1352;
  wire _abc_40344_n1353;
  wire _abc_40344_n1354;
  wire _abc_40344_n1355;
  wire _abc_40344_n1356;
  wire _abc_40344_n1357;
  wire _abc_40344_n1358;
  wire _abc_40344_n1359_1;
  wire _abc_40344_n1360;
  wire _abc_40344_n1361;
  wire _abc_40344_n1362;
  wire _abc_40344_n1363;
  wire _abc_40344_n1364;
  wire _abc_40344_n1365;
  wire _abc_40344_n1366;
  wire _abc_40344_n1367;
  wire _abc_40344_n1368;
  wire _abc_40344_n1369;
  wire _abc_40344_n1370;
  wire _abc_40344_n1371_1;
  wire _abc_40344_n1372;
  wire _abc_40344_n1373;
  wire _abc_40344_n1374;
  wire _abc_40344_n1375;
  wire _abc_40344_n1376;
  wire _abc_40344_n1377;
  wire _abc_40344_n1378;
  wire _abc_40344_n1379;
  wire _abc_40344_n1380;
  wire _abc_40344_n1381;
  wire _abc_40344_n1382;
  wire _abc_40344_n1383_1;
  wire _abc_40344_n1384;
  wire _abc_40344_n1385;
  wire _abc_40344_n1386;
  wire _abc_40344_n1387;
  wire _abc_40344_n1388;
  wire _abc_40344_n1389;
  wire _abc_40344_n1390;
  wire _abc_40344_n1391;
  wire _abc_40344_n1392;
  wire _abc_40344_n1393;
  wire _abc_40344_n1394;
  wire _abc_40344_n1395;
  wire _abc_40344_n1396_1;
  wire _abc_40344_n1397;
  wire _abc_40344_n1398;
  wire _abc_40344_n1399;
  wire _abc_40344_n1400;
  wire _abc_40344_n1401;
  wire _abc_40344_n1402;
  wire _abc_40344_n1403;
  wire _abc_40344_n1404;
  wire _abc_40344_n1405;
  wire _abc_40344_n1406;
  wire _abc_40344_n1407;
  wire _abc_40344_n1408;
  wire _abc_40344_n1409_1;
  wire _abc_40344_n1410;
  wire _abc_40344_n1411;
  wire _abc_40344_n1412;
  wire _abc_40344_n1413;
  wire _abc_40344_n1414;
  wire _abc_40344_n1415;
  wire _abc_40344_n1416;
  wire _abc_40344_n1417;
  wire _abc_40344_n1418;
  wire _abc_40344_n1419;
  wire _abc_40344_n1420;
  wire _abc_40344_n1421_1;
  wire _abc_40344_n1422;
  wire _abc_40344_n1423;
  wire _abc_40344_n1424;
  wire _abc_40344_n1425;
  wire _abc_40344_n1426;
  wire _abc_40344_n1427;
  wire _abc_40344_n1428;
  wire _abc_40344_n1429;
  wire _abc_40344_n1430;
  wire _abc_40344_n1431;
  wire _abc_40344_n1432;
  wire _abc_40344_n1433;
  wire _abc_40344_n1434;
  wire _abc_40344_n1435;
  wire _abc_40344_n1436;
  wire _abc_40344_n1437;
  wire _abc_40344_n1438;
  wire _abc_40344_n1439_1;
  wire _abc_40344_n1440;
  wire _abc_40344_n1441;
  wire _abc_40344_n1442;
  wire _abc_40344_n1443;
  wire _abc_40344_n1444;
  wire _abc_40344_n1445;
  wire _abc_40344_n1446;
  wire _abc_40344_n1447;
  wire _abc_40344_n1448;
  wire _abc_40344_n1449;
  wire _abc_40344_n1450;
  wire _abc_40344_n1451_1;
  wire _abc_40344_n1452;
  wire _abc_40344_n1453;
  wire _abc_40344_n1454;
  wire _abc_40344_n1455;
  wire _abc_40344_n1456;
  wire _abc_40344_n1457;
  wire _abc_40344_n1458;
  wire _abc_40344_n1459;
  wire _abc_40344_n1460;
  wire _abc_40344_n1461;
  wire _abc_40344_n1462;
  wire _abc_40344_n1463;
  wire _abc_40344_n1464;
  wire _abc_40344_n1465;
  wire _abc_40344_n1466;
  wire _abc_40344_n1467;
  wire _abc_40344_n1468;
  wire _abc_40344_n1469;
  wire _abc_40344_n1470;
  wire _abc_40344_n1471;
  wire _abc_40344_n1472;
  wire _abc_40344_n1473;
  wire _abc_40344_n1474;
  wire _abc_40344_n1475;
  wire _abc_40344_n1476;
  wire _abc_40344_n1477;
  wire _abc_40344_n1478;
  wire _abc_40344_n1479;
  wire _abc_40344_n1480;
  wire _abc_40344_n1481;
  wire _abc_40344_n1482;
  wire _abc_40344_n1483;
  wire _abc_40344_n1484;
  wire _abc_40344_n1485;
  wire _abc_40344_n1486;
  wire _abc_40344_n1487;
  wire _abc_40344_n1488;
  wire _abc_40344_n1489;
  wire _abc_40344_n1490;
  wire _abc_40344_n1491;
  wire _abc_40344_n1492;
  wire _abc_40344_n1493;
  wire _abc_40344_n1494;
  wire _abc_40344_n1495;
  wire _abc_40344_n1496;
  wire _abc_40344_n1497;
  wire _abc_40344_n1498;
  wire _abc_40344_n1499;
  wire _abc_40344_n1500;
  wire _abc_40344_n1501;
  wire _abc_40344_n1502;
  wire _abc_40344_n1503_1;
  wire _abc_40344_n1504;
  wire _abc_40344_n1505_1;
  wire _abc_40344_n1506;
  wire _abc_40344_n1507_1;
  wire _abc_40344_n1508_1;
  wire _abc_40344_n1509;
  wire _abc_40344_n1510;
  wire _abc_40344_n1511_1;
  wire _abc_40344_n1512;
  wire _abc_40344_n1513;
  wire _abc_40344_n1514_1;
  wire _abc_40344_n1515;
  wire _abc_40344_n1516_1;
  wire _abc_40344_n1517_1;
  wire _abc_40344_n1518;
  wire _abc_40344_n1519;
  wire _abc_40344_n1520_1;
  wire _abc_40344_n1521;
  wire _abc_40344_n1522;
  wire _abc_40344_n1523;
  wire _abc_40344_n1524;
  wire _abc_40344_n1525;
  wire _abc_40344_n1526;
  wire _abc_40344_n1527;
  wire _abc_40344_n1528;
  wire _abc_40344_n1529;
  wire _abc_40344_n1530;
  wire _abc_40344_n1531;
  wire _abc_40344_n1532;
  wire _abc_40344_n1533;
  wire _abc_40344_n1534;
  wire _abc_40344_n1535;
  wire _abc_40344_n1536;
  wire _abc_40344_n1537;
  wire _abc_40344_n1537_bF_buf0;
  wire _abc_40344_n1537_bF_buf1;
  wire _abc_40344_n1537_bF_buf2;
  wire _abc_40344_n1537_bF_buf3;
  wire _abc_40344_n1538;
  wire _abc_40344_n1539;
  wire _abc_40344_n1540;
  wire _abc_40344_n1541;
  wire _abc_40344_n1542;
  wire _abc_40344_n1543;
  wire _abc_40344_n1544;
  wire _abc_40344_n1545;
  wire _abc_40344_n1546;
  wire _abc_40344_n1547;
  wire _abc_40344_n1548;
  wire _abc_40344_n1549;
  wire _abc_40344_n1550;
  wire _abc_40344_n1550_bF_buf0;
  wire _abc_40344_n1550_bF_buf1;
  wire _abc_40344_n1550_bF_buf2;
  wire _abc_40344_n1550_bF_buf3;
  wire _abc_40344_n1551;
  wire _abc_40344_n1552;
  wire _abc_40344_n1553;
  wire _abc_40344_n1554;
  wire _abc_40344_n1555;
  wire _abc_40344_n1555_bF_buf0;
  wire _abc_40344_n1555_bF_buf1;
  wire _abc_40344_n1555_bF_buf2;
  wire _abc_40344_n1555_bF_buf3;
  wire _abc_40344_n1556;
  wire _abc_40344_n1557;
  wire _abc_40344_n1559;
  wire _abc_40344_n1560;
  wire _abc_40344_n1561;
  wire _abc_40344_n1562;
  wire _abc_40344_n1563;
  wire _abc_40344_n1564;
  wire _abc_40344_n1565;
  wire _abc_40344_n1566;
  wire _abc_40344_n1567;
  wire _abc_40344_n1568;
  wire _abc_40344_n1569;
  wire _abc_40344_n1571;
  wire _abc_40344_n1572;
  wire _abc_40344_n1573;
  wire _abc_40344_n1574;
  wire _abc_40344_n1575;
  wire _abc_40344_n1576;
  wire _abc_40344_n1577;
  wire _abc_40344_n1578;
  wire _abc_40344_n1579;
  wire _abc_40344_n1580;
  wire _abc_40344_n1581;
  wire _abc_40344_n1582;
  wire _abc_40344_n1583;
  wire _abc_40344_n1584;
  wire _abc_40344_n1586;
  wire _abc_40344_n1587;
  wire _abc_40344_n1588;
  wire _abc_40344_n1589;
  wire _abc_40344_n1590;
  wire _abc_40344_n1591;
  wire _abc_40344_n1592;
  wire _abc_40344_n1593;
  wire _abc_40344_n1594;
  wire _abc_40344_n1595;
  wire _abc_40344_n1596;
  wire _abc_40344_n1597;
  wire _abc_40344_n1599;
  wire _abc_40344_n1600;
  wire _abc_40344_n1601;
  wire _abc_40344_n1602;
  wire _abc_40344_n1603;
  wire _abc_40344_n1604;
  wire _abc_40344_n1605;
  wire _abc_40344_n1606;
  wire _abc_40344_n1607;
  wire _abc_40344_n1608;
  wire _abc_40344_n1609;
  wire _abc_40344_n1610;
  wire _abc_40344_n1611;
  wire _abc_40344_n1612;
  wire _abc_40344_n1613;
  wire _abc_40344_n1614;
  wire _abc_40344_n1616;
  wire _abc_40344_n1617;
  wire _abc_40344_n1618;
  wire _abc_40344_n1619;
  wire _abc_40344_n1620;
  wire _abc_40344_n1621;
  wire _abc_40344_n1622;
  wire _abc_40344_n1623;
  wire _abc_40344_n1624;
  wire _abc_40344_n1625;
  wire _abc_40344_n1626;
  wire _abc_40344_n1628;
  wire _abc_40344_n1629;
  wire _abc_40344_n1630;
  wire _abc_40344_n1631;
  wire _abc_40344_n1632;
  wire _abc_40344_n1633;
  wire _abc_40344_n1634;
  wire _abc_40344_n1635;
  wire _abc_40344_n1636;
  wire _abc_40344_n1637;
  wire _abc_40344_n1638;
  wire _abc_40344_n1639;
  wire _abc_40344_n1640;
  wire _abc_40344_n1641;
  wire _abc_40344_n1642;
  wire _abc_40344_n1643;
  wire _abc_40344_n1644;
  wire _abc_40344_n1645;
  wire _abc_40344_n1646;
  wire _abc_40344_n1647;
  wire _abc_40344_n1648;
  wire _abc_40344_n1649;
  wire _abc_40344_n1650;
  wire _abc_40344_n1651;
  wire _abc_40344_n1652;
  wire _abc_40344_n1653;
  wire _abc_40344_n1655;
  wire _abc_40344_n1656;
  wire _abc_40344_n1657;
  wire _abc_40344_n1658;
  wire _abc_40344_n1659;
  wire _abc_40344_n1660;
  wire _abc_40344_n1661;
  wire _abc_40344_n1662;
  wire _abc_40344_n1663;
  wire _abc_40344_n1664;
  wire _abc_40344_n1665;
  wire _abc_40344_n1666;
  wire _abc_40344_n1667;
  wire _abc_40344_n1668;
  wire _abc_40344_n1669;
  wire _abc_40344_n1671;
  wire _abc_40344_n1672;
  wire _abc_40344_n1673;
  wire _abc_40344_n1674;
  wire _abc_40344_n1675;
  wire _abc_40344_n1676;
  wire _abc_40344_n1677;
  wire _abc_40344_n1678;
  wire _abc_40344_n1679;
  wire _abc_40344_n1680;
  wire _abc_40344_n1681;
  wire _abc_40344_n1682;
  wire _abc_40344_n1684;
  wire _abc_40344_n1685;
  wire _abc_40344_n1686;
  wire _abc_40344_n1687;
  wire _abc_40344_n1688;
  wire _abc_40344_n1689;
  wire _abc_40344_n1690;
  wire _abc_40344_n1691;
  wire _abc_40344_n1692;
  wire _abc_40344_n1693;
  wire _abc_40344_n1694;
  wire _abc_40344_n1695;
  wire _abc_40344_n1696;
  wire _abc_40344_n1697;
  wire _abc_40344_n1698;
  wire _abc_40344_n1699;
  wire _abc_40344_n1701;
  wire _abc_40344_n1702;
  wire _abc_40344_n1703;
  wire _abc_40344_n1704;
  wire _abc_40344_n1705;
  wire _abc_40344_n1706;
  wire _abc_40344_n1707;
  wire _abc_40344_n1708;
  wire _abc_40344_n1709;
  wire _abc_40344_n1710;
  wire _abc_40344_n1711;
  wire _abc_40344_n1712;
  wire _abc_40344_n1713;
  wire _abc_40344_n1715;
  wire _abc_40344_n1716;
  wire _abc_40344_n1717;
  wire _abc_40344_n1718;
  wire _abc_40344_n1719;
  wire _abc_40344_n1720;
  wire _abc_40344_n1721;
  wire _abc_40344_n1722;
  wire _abc_40344_n1723;
  wire _abc_40344_n1724;
  wire _abc_40344_n1725;
  wire _abc_40344_n1726;
  wire _abc_40344_n1727;
  wire _abc_40344_n1728;
  wire _abc_40344_n1729;
  wire _abc_40344_n1730;
  wire _abc_40344_n1732;
  wire _abc_40344_n1733;
  wire _abc_40344_n1734;
  wire _abc_40344_n1735;
  wire _abc_40344_n1736;
  wire _abc_40344_n1737;
  wire _abc_40344_n1738;
  wire _abc_40344_n1739;
  wire _abc_40344_n1740;
  wire _abc_40344_n1742;
  wire _abc_40344_n1743;
  wire _abc_40344_n1744;
  wire _abc_40344_n1745;
  wire _abc_40344_n1746;
  wire _abc_40344_n1747;
  wire _abc_40344_n1748;
  wire _abc_40344_n1750;
  wire _abc_40344_n1751;
  wire _abc_40344_n1752;
  wire _abc_40344_n1753;
  wire _abc_40344_n1754;
  wire _abc_40344_n1755;
  wire _abc_40344_n1756;
  wire _abc_40344_n1757;
  wire _abc_40344_n1758;
  wire _abc_40344_n1759;
  wire _abc_40344_n1760;
  wire _abc_40344_n1761;
  wire _abc_40344_n1763;
  wire _abc_40344_n1764;
  wire _abc_40344_n1765;
  wire _abc_40344_n1766;
  wire _abc_40344_n1767;
  wire _abc_40344_n1768;
  wire _abc_40344_n1769;
  wire _abc_40344_n1770;
  wire _abc_40344_n1771;
  wire _abc_40344_n1773;
  wire _abc_40344_n1774;
  wire _abc_40344_n1775;
  wire _abc_40344_n1776;
  wire _abc_40344_n1777;
  wire _abc_40344_n1778;
  wire _abc_40344_n1779;
  wire _abc_40344_n1780;
  wire _abc_40344_n1782;
  wire _abc_40344_n1783;
  wire _abc_40344_n1784;
  wire _abc_40344_n1785;
  wire _abc_40344_n1786;
  wire _abc_40344_n1787;
  wire _abc_40344_n1788;
  wire _abc_40344_n1789;
  wire _abc_40344_n1790;
  wire _abc_40344_n1791;
  wire _abc_40344_n1792;
  wire _abc_40344_n1794;
  wire _abc_40344_n1795;
  wire _abc_40344_n1796;
  wire _abc_40344_n1797;
  wire _abc_40344_n1798;
  wire _abc_40344_n1799;
  wire _abc_40344_n1800;
  wire _abc_40344_n1801;
  wire _abc_40344_n1802;
  wire _abc_40344_n1803;
  wire _abc_40344_n1804;
  wire _abc_40344_n1805;
  wire _abc_40344_n1807;
  wire _abc_40344_n1808;
  wire _abc_40344_n1809;
  wire _abc_40344_n1810;
  wire _abc_40344_n1811;
  wire _abc_40344_n1812;
  wire _abc_40344_n1813;
  wire _abc_40344_n1814;
  wire _abc_40344_n1815;
  wire _abc_40344_n1816;
  wire _abc_40344_n1818;
  wire _abc_40344_n1819;
  wire _abc_40344_n1820;
  wire _abc_40344_n1821;
  wire _abc_40344_n1822;
  wire _abc_40344_n1823;
  wire _abc_40344_n1824;
  wire _abc_40344_n1825;
  wire _abc_40344_n1826;
  wire _abc_40344_n1827;
  wire _abc_40344_n1828;
  wire _abc_40344_n1829;
  wire _abc_40344_n1831;
  wire _abc_40344_n1832;
  wire _abc_40344_n1833;
  wire _abc_40344_n1834;
  wire _abc_40344_n1835;
  wire _abc_40344_n1836;
  wire _abc_40344_n1837;
  wire _abc_40344_n1838;
  wire _abc_40344_n1840;
  wire _abc_40344_n1841;
  wire _abc_40344_n1842;
  wire _abc_40344_n1843;
  wire _abc_40344_n1844;
  wire _abc_40344_n1845;
  wire _abc_40344_n1846;
  wire _abc_40344_n1847;
  wire _abc_40344_n1848;
  wire _abc_40344_n1849;
  wire _abc_40344_n1851;
  wire _abc_40344_n1852;
  wire _abc_40344_n1853;
  wire _abc_40344_n1854;
  wire _abc_40344_n1855;
  wire _abc_40344_n1856;
  wire _abc_40344_n1857;
  wire _abc_40344_n1858;
  wire _abc_40344_n1860;
  wire _abc_40344_n1861;
  wire _abc_40344_n1862;
  wire _abc_40344_n1863;
  wire _abc_40344_n1864;
  wire _abc_40344_n1865;
  wire _abc_40344_n1866;
  wire _abc_40344_n1867;
  wire _abc_40344_n1869;
  wire _abc_40344_n1870;
  wire _abc_40344_n1871;
  wire _abc_40344_n1872;
  wire _abc_40344_n1873;
  wire _abc_40344_n1874;
  wire _abc_40344_n1875;
  wire _abc_40344_n1876;
  wire _abc_40344_n1878;
  wire _abc_40344_n1879;
  wire _abc_40344_n1880;
  wire _abc_40344_n1881;
  wire _abc_40344_n1882;
  wire _abc_40344_n1883;
  wire _abc_40344_n1884;
  wire _abc_40344_n1885;
  wire _abc_40344_n1886;
  wire _abc_40344_n1887;
  wire _abc_40344_n1888;
  wire _abc_40344_n1889;
  wire _abc_40344_n1890;
  wire _abc_40344_n1891;
  wire _abc_40344_n1892;
  wire _abc_40344_n1894;
  wire _abc_40344_n1895;
  wire _abc_40344_n1896;
  wire _abc_40344_n1897;
  wire _abc_40344_n1898;
  wire _abc_40344_n1899;
  wire _abc_40344_n1900;
  wire _abc_40344_n1901;
  wire _abc_40344_n1902;
  wire _abc_40344_n1904;
  wire _abc_40344_n1905;
  wire _abc_40344_n1906;
  wire _abc_40344_n1907;
  wire _abc_40344_n1908;
  wire _abc_40344_n1909;
  wire _abc_40344_n1910;
  wire _abc_40344_n1911;
  wire _abc_40344_n1912;
  wire _abc_40344_n1913;
  wire _abc_40344_n1914;
  wire _abc_40344_n1915;
  wire _abc_40344_n1916;
  wire _abc_40344_n1917;
  wire _abc_40344_n1918;
  wire _abc_40344_n1919;
  wire _abc_40344_n1920;
  wire _abc_40344_n1921;
  wire _abc_40344_n1922;
  wire _abc_40344_n1923;
  wire _abc_40344_n1924;
  wire _abc_40344_n1925;
  wire _abc_40344_n1926;
  wire _abc_40344_n1927;
  wire _abc_40344_n1928;
  wire _abc_40344_n1929;
  wire _abc_40344_n1930;
  wire _abc_40344_n1931;
  wire _abc_40344_n1932;
  wire _abc_40344_n1933;
  wire _abc_40344_n1934;
  wire _abc_40344_n1935;
  wire _abc_40344_n1936;
  wire _abc_40344_n1937;
  wire _abc_40344_n1938;
  wire _abc_40344_n1939;
  wire _abc_40344_n1940;
  wire _abc_40344_n1941;
  wire _abc_40344_n1942;
  wire _abc_40344_n1943;
  wire _abc_40344_n1944;
  wire _abc_40344_n1945;
  wire _abc_40344_n1946;
  wire _abc_40344_n1947;
  wire _abc_40344_n1948;
  wire _abc_40344_n1949;
  wire _abc_40344_n1950;
  wire _abc_40344_n1951;
  wire _abc_40344_n1952;
  wire _abc_40344_n1953;
  wire _abc_40344_n1954;
  wire _abc_40344_n1955;
  wire _abc_40344_n1956;
  wire _abc_40344_n1957;
  wire _abc_40344_n1958;
  wire _abc_40344_n1959;
  wire _abc_40344_n1960;
  wire _abc_40344_n1961;
  wire _abc_40344_n1962;
  wire _abc_40344_n1963;
  wire _abc_40344_n1964;
  wire _abc_40344_n1965;
  wire _abc_40344_n1966;
  wire _abc_40344_n1967;
  wire _abc_40344_n1968;
  wire _abc_40344_n1969;
  wire _abc_40344_n1970;
  wire _abc_40344_n1971;
  wire _abc_40344_n1972;
  wire _abc_40344_n1973;
  wire _abc_40344_n1974;
  wire _abc_40344_n1975;
  wire _abc_40344_n1976;
  wire _abc_40344_n1977;
  wire _abc_40344_n1978;
  wire _abc_40344_n1979;
  wire _abc_40344_n1980;
  wire _abc_40344_n1981;
  wire _abc_40344_n1982;
  wire _abc_40344_n1983;
  wire _abc_40344_n1984;
  wire _abc_40344_n1985;
  wire _abc_40344_n1986;
  wire _abc_40344_n1987;
  wire _abc_40344_n1988;
  wire _abc_40344_n1989;
  wire _abc_40344_n1990;
  wire _abc_40344_n1991;
  wire _abc_40344_n1992;
  wire _abc_40344_n1993;
  wire _abc_40344_n1994;
  wire _abc_40344_n1995;
  wire _abc_40344_n1996;
  wire _abc_40344_n1997;
  wire _abc_40344_n1998;
  wire _abc_40344_n1999;
  wire _abc_40344_n2000;
  wire _abc_40344_n2001;
  wire _abc_40344_n2002;
  wire _abc_40344_n2003;
  wire _abc_40344_n2004;
  wire _abc_40344_n2005;
  wire _abc_40344_n2006;
  wire _abc_40344_n2007;
  wire _abc_40344_n2008;
  wire _abc_40344_n2009;
  wire _abc_40344_n2010;
  wire _abc_40344_n2011;
  wire _abc_40344_n2012;
  wire _abc_40344_n2013;
  wire _abc_40344_n2014;
  wire _abc_40344_n2015;
  wire _abc_40344_n2016;
  wire _abc_40344_n2017;
  wire _abc_40344_n2018;
  wire _abc_40344_n2019;
  wire _abc_40344_n2020;
  wire _abc_40344_n2021;
  wire _abc_40344_n2022;
  wire _abc_40344_n2023;
  wire _abc_40344_n2024;
  wire _abc_40344_n2025;
  wire _abc_40344_n2026;
  wire _abc_40344_n2027;
  wire _abc_40344_n2028;
  wire _abc_40344_n2029;
  wire _abc_40344_n2030;
  wire _abc_40344_n2031;
  wire _abc_40344_n2032;
  wire _abc_40344_n2033;
  wire _abc_40344_n2034;
  wire _abc_40344_n2035;
  wire _abc_40344_n2036;
  wire _abc_40344_n2037;
  wire _abc_40344_n2038;
  wire _abc_40344_n2039;
  wire _abc_40344_n2040;
  wire _abc_40344_n2041;
  wire _abc_40344_n2042;
  wire _abc_40344_n2043;
  wire _abc_40344_n2044;
  wire _abc_40344_n2045;
  wire _abc_40344_n2046;
  wire _abc_40344_n2047;
  wire _abc_40344_n2048;
  wire _abc_40344_n2049;
  wire _abc_40344_n2050;
  wire _abc_40344_n2051;
  wire _abc_40344_n2052;
  wire _abc_40344_n2053;
  wire _abc_40344_n2054;
  wire _abc_40344_n2055;
  wire _abc_40344_n2056;
  wire _abc_40344_n2057;
  wire _abc_40344_n2058;
  wire _abc_40344_n2059;
  wire _abc_40344_n2060;
  wire _abc_40344_n2061;
  wire _abc_40344_n2062;
  wire _abc_40344_n2063;
  wire _abc_40344_n2064;
  wire _abc_40344_n2065;
  wire _abc_40344_n2066;
  wire _abc_40344_n2067;
  wire _abc_40344_n2068;
  wire _abc_40344_n2069;
  wire _abc_40344_n2070;
  wire _abc_40344_n2071;
  wire _abc_40344_n2072;
  wire _abc_40344_n2073;
  wire _abc_40344_n2074;
  wire _abc_40344_n2075;
  wire _abc_40344_n2076;
  wire _abc_40344_n2077;
  wire _abc_40344_n2078;
  wire _abc_40344_n2079;
  wire _abc_40344_n2080;
  wire _abc_40344_n2081;
  wire _abc_40344_n2082;
  wire _abc_40344_n2083;
  wire _abc_40344_n2084;
  wire _abc_40344_n2085;
  wire _abc_40344_n2086;
  wire _abc_40344_n2087;
  wire _abc_40344_n2088;
  wire _abc_40344_n2089;
  wire _abc_40344_n2090;
  wire _abc_40344_n2091;
  wire _abc_40344_n2092;
  wire _abc_40344_n2093;
  wire _abc_40344_n2094;
  wire _abc_40344_n2095;
  wire _abc_40344_n2096;
  wire _abc_40344_n2097;
  wire _abc_40344_n2098;
  wire _abc_40344_n2099;
  wire _abc_40344_n2100;
  wire _abc_40344_n2101;
  wire _abc_40344_n2102;
  wire _abc_40344_n2103;
  wire _abc_40344_n2104;
  wire _abc_40344_n2105;
  wire _abc_40344_n2106;
  wire _abc_40344_n2107;
  wire _abc_40344_n2108;
  wire _abc_40344_n2109;
  wire _abc_40344_n2110;
  wire _abc_40344_n2111;
  wire _abc_40344_n2112;
  wire _abc_40344_n2113;
  wire _abc_40344_n2114;
  wire _abc_40344_n2115;
  wire _abc_40344_n2116;
  wire _abc_40344_n2117;
  wire _abc_40344_n2118;
  wire _abc_40344_n2119;
  wire _abc_40344_n2120;
  wire _abc_40344_n2121;
  wire _abc_40344_n2122;
  wire _abc_40344_n2123;
  wire _abc_40344_n2124;
  wire _abc_40344_n2125;
  wire _abc_40344_n2126;
  wire _abc_40344_n2127;
  wire _abc_40344_n2128;
  wire _abc_40344_n2129;
  wire _abc_40344_n2130;
  wire _abc_40344_n2131;
  wire _abc_40344_n2132;
  wire _abc_40344_n2133;
  wire _abc_40344_n2134;
  wire _abc_40344_n2135;
  wire _abc_40344_n2136;
  wire _abc_40344_n2137;
  wire _abc_40344_n2138;
  wire _abc_40344_n2139;
  wire _abc_40344_n2140;
  wire _abc_40344_n2141;
  wire _abc_40344_n2142;
  wire _abc_40344_n2143;
  wire _abc_40344_n2144;
  wire _abc_40344_n2145;
  wire _abc_40344_n2146;
  wire _abc_40344_n2147;
  wire _abc_40344_n2148;
  wire _abc_40344_n2149;
  wire _abc_40344_n2150;
  wire _abc_40344_n2151;
  wire _abc_40344_n2152;
  wire _abc_40344_n2153;
  wire _abc_40344_n2154;
  wire _abc_40344_n2155;
  wire _abc_40344_n2156;
  wire _abc_40344_n2157;
  wire _abc_40344_n2158;
  wire _abc_40344_n2159;
  wire _abc_40344_n2160;
  wire _abc_40344_n2161;
  wire _abc_40344_n2161_bF_buf0;
  wire _abc_40344_n2161_bF_buf1;
  wire _abc_40344_n2161_bF_buf2;
  wire _abc_40344_n2161_bF_buf3;
  wire _abc_40344_n2162;
  wire _abc_40344_n2162_bF_buf0;
  wire _abc_40344_n2162_bF_buf1;
  wire _abc_40344_n2162_bF_buf2;
  wire _abc_40344_n2162_bF_buf3;
  wire _abc_40344_n2163;
  wire _abc_40344_n2164;
  wire _abc_40344_n2165;
  wire _abc_40344_n2165_bF_buf0;
  wire _abc_40344_n2165_bF_buf1;
  wire _abc_40344_n2165_bF_buf2;
  wire _abc_40344_n2165_bF_buf3;
  wire _abc_40344_n2165_bF_buf4;
  wire _abc_40344_n2165_bF_buf5;
  wire _abc_40344_n2165_bF_buf6;
  wire _abc_40344_n2166;
  wire _abc_40344_n2167;
  wire _abc_40344_n2168;
  wire _abc_40344_n2169;
  wire _abc_40344_n2170;
  wire _abc_40344_n2171;
  wire _abc_40344_n2172;
  wire _abc_40344_n2173;
  wire _abc_40344_n2173_bF_buf0;
  wire _abc_40344_n2173_bF_buf1;
  wire _abc_40344_n2173_bF_buf2;
  wire _abc_40344_n2173_bF_buf3;
  wire _abc_40344_n2173_bF_buf4;
  wire _abc_40344_n2174;
  wire _abc_40344_n2175;
  wire _abc_40344_n2176;
  wire _abc_40344_n2177;
  wire _abc_40344_n2178;
  wire _abc_40344_n2179;
  wire _abc_40344_n2179_bF_buf0;
  wire _abc_40344_n2179_bF_buf1;
  wire _abc_40344_n2179_bF_buf2;
  wire _abc_40344_n2179_bF_buf3;
  wire _abc_40344_n2179_bF_buf4;
  wire _abc_40344_n2180;
  wire _abc_40344_n2181;
  wire _abc_40344_n2182;
  wire _abc_40344_n2183;
  wire _abc_40344_n2184;
  wire _abc_40344_n2185;
  wire _abc_40344_n2186;
  wire _abc_40344_n2187;
  wire _abc_40344_n2188;
  wire _abc_40344_n2189;
  wire _abc_40344_n2190;
  wire _abc_40344_n2191;
  wire _abc_40344_n2192;
  wire _abc_40344_n2193;
  wire _abc_40344_n2194;
  wire _abc_40344_n2195;
  wire _abc_40344_n2196;
  wire _abc_40344_n2197;
  wire _abc_40344_n2198;
  wire _abc_40344_n2199;
  wire _abc_40344_n2200;
  wire _abc_40344_n2201;
  wire _abc_40344_n2202;
  wire _abc_40344_n2203;
  wire _abc_40344_n2204;
  wire _abc_40344_n2205;
  wire _abc_40344_n2206;
  wire _abc_40344_n2207;
  wire _abc_40344_n2208;
  wire _abc_40344_n2209;
  wire _abc_40344_n2210;
  wire _abc_40344_n2211;
  wire _abc_40344_n2212;
  wire _abc_40344_n2213;
  wire _abc_40344_n2214;
  wire _abc_40344_n2215;
  wire _abc_40344_n2216;
  wire _abc_40344_n2217;
  wire _abc_40344_n2218;
  wire _abc_40344_n2219;
  wire _abc_40344_n2220;
  wire _abc_40344_n2221;
  wire _abc_40344_n2222;
  wire _abc_40344_n2223;
  wire _abc_40344_n2224;
  wire _abc_40344_n2225;
  wire _abc_40344_n2226;
  wire _abc_40344_n2227;
  wire _abc_40344_n2228;
  wire _abc_40344_n2229;
  wire _abc_40344_n2230;
  wire _abc_40344_n2231;
  wire _abc_40344_n2232;
  wire _abc_40344_n2233;
  wire _abc_40344_n2234;
  wire _abc_40344_n2235;
  wire _abc_40344_n2236;
  wire _abc_40344_n2237;
  wire _abc_40344_n2238;
  wire _abc_40344_n2239;
  wire _abc_40344_n2240;
  wire _abc_40344_n2241;
  wire _abc_40344_n2242;
  wire _abc_40344_n2243;
  wire _abc_40344_n2244;
  wire _abc_40344_n2245;
  wire _abc_40344_n2246;
  wire _abc_40344_n2247;
  wire _abc_40344_n2248;
  wire _abc_40344_n2249;
  wire _abc_40344_n2250;
  wire _abc_40344_n2251;
  wire _abc_40344_n2252;
  wire _abc_40344_n2253_1;
  wire _abc_40344_n2254;
  wire _abc_40344_n2255;
  wire _abc_40344_n2256;
  wire _abc_40344_n2257;
  wire _abc_40344_n2258;
  wire _abc_40344_n2259;
  wire _abc_40344_n2260;
  wire _abc_40344_n2261;
  wire _abc_40344_n2262;
  wire _abc_40344_n2263;
  wire _abc_40344_n2264;
  wire _abc_40344_n2265;
  wire _abc_40344_n2266;
  wire _abc_40344_n2267;
  wire _abc_40344_n2268;
  wire _abc_40344_n2269;
  wire _abc_40344_n2270;
  wire _abc_40344_n2271;
  wire _abc_40344_n2272;
  wire _abc_40344_n2273;
  wire _abc_40344_n2274;
  wire _abc_40344_n2275;
  wire _abc_40344_n2276;
  wire _abc_40344_n2277_1;
  wire _abc_40344_n2278;
  wire _abc_40344_n2279;
  wire _abc_40344_n2280;
  wire _abc_40344_n2281;
  wire _abc_40344_n2282;
  wire _abc_40344_n2283;
  wire _abc_40344_n2284;
  wire _abc_40344_n2285;
  wire _abc_40344_n2286;
  wire _abc_40344_n2287;
  wire _abc_40344_n2288_1;
  wire _abc_40344_n2289;
  wire _abc_40344_n2290;
  wire _abc_40344_n2291;
  wire _abc_40344_n2292;
  wire _abc_40344_n2293;
  wire _abc_40344_n2294;
  wire _abc_40344_n2295;
  wire _abc_40344_n2296;
  wire _abc_40344_n2297;
  wire _abc_40344_n2298;
  wire _abc_40344_n2299;
  wire _abc_40344_n2300;
  wire _abc_40344_n2301;
  wire _abc_40344_n2302;
  wire _abc_40344_n2303;
  wire _abc_40344_n2304;
  wire _abc_40344_n2305;
  wire _abc_40344_n2306;
  wire _abc_40344_n2307;
  wire _abc_40344_n2308_1;
  wire _abc_40344_n2309;
  wire _abc_40344_n2310;
  wire _abc_40344_n2311;
  wire _abc_40344_n2312;
  wire _abc_40344_n2313;
  wire _abc_40344_n2314_1;
  wire _abc_40344_n2315;
  wire _abc_40344_n2316;
  wire _abc_40344_n2317;
  wire _abc_40344_n2318;
  wire _abc_40344_n2319;
  wire _abc_40344_n2320;
  wire _abc_40344_n2321;
  wire _abc_40344_n2322;
  wire _abc_40344_n2323;
  wire _abc_40344_n2324;
  wire _abc_40344_n2325;
  wire _abc_40344_n2326;
  wire _abc_40344_n2327;
  wire _abc_40344_n2328;
  wire _abc_40344_n2329;
  wire _abc_40344_n2330;
  wire _abc_40344_n2331_1;
  wire _abc_40344_n2332;
  wire _abc_40344_n2333;
  wire _abc_40344_n2334;
  wire _abc_40344_n2335;
  wire _abc_40344_n2336;
  wire _abc_40344_n2337;
  wire _abc_40344_n2338;
  wire _abc_40344_n2339;
  wire _abc_40344_n2340_1;
  wire _abc_40344_n2341;
  wire _abc_40344_n2342;
  wire _abc_40344_n2343;
  wire _abc_40344_n2344;
  wire _abc_40344_n2345;
  wire _abc_40344_n2346;
  wire _abc_40344_n2347;
  wire _abc_40344_n2348;
  wire _abc_40344_n2349;
  wire _abc_40344_n2350;
  wire _abc_40344_n2351;
  wire _abc_40344_n2352;
  wire _abc_40344_n2353;
  wire _abc_40344_n2354;
  wire _abc_40344_n2355;
  wire _abc_40344_n2356;
  wire _abc_40344_n2357;
  wire _abc_40344_n2358;
  wire _abc_40344_n2359;
  wire _abc_40344_n2360;
  wire _abc_40344_n2361;
  wire _abc_40344_n2362_1;
  wire _abc_40344_n2363;
  wire _abc_40344_n2364;
  wire _abc_40344_n2365;
  wire _abc_40344_n2366;
  wire _abc_40344_n2367;
  wire _abc_40344_n2368;
  wire _abc_40344_n2369_1;
  wire _abc_40344_n2370;
  wire _abc_40344_n2371;
  wire _abc_40344_n2372;
  wire _abc_40344_n2373;
  wire _abc_40344_n2374;
  wire _abc_40344_n2375;
  wire _abc_40344_n2376;
  wire _abc_40344_n2377;
  wire _abc_40344_n2378;
  wire _abc_40344_n2379;
  wire _abc_40344_n2380_1;
  wire _abc_40344_n2381;
  wire _abc_40344_n2382;
  wire _abc_40344_n2383;
  wire _abc_40344_n2384;
  wire _abc_40344_n2385;
  wire _abc_40344_n2386;
  wire _abc_40344_n2387;
  wire _abc_40344_n2388;
  wire _abc_40344_n2389_1;
  wire _abc_40344_n2390;
  wire _abc_40344_n2391;
  wire _abc_40344_n2392;
  wire _abc_40344_n2393;
  wire _abc_40344_n2394;
  wire _abc_40344_n2395;
  wire _abc_40344_n2396;
  wire _abc_40344_n2397;
  wire _abc_40344_n2398;
  wire _abc_40344_n2399;
  wire _abc_40344_n2400;
  wire _abc_40344_n2401;
  wire _abc_40344_n2402;
  wire _abc_40344_n2403;
  wire _abc_40344_n2404;
  wire _abc_40344_n2405;
  wire _abc_40344_n2406;
  wire _abc_40344_n2407;
  wire _abc_40344_n2408_1;
  wire _abc_40344_n2409;
  wire _abc_40344_n2410;
  wire _abc_40344_n2411;
  wire _abc_40344_n2412;
  wire _abc_40344_n2413;
  wire _abc_40344_n2414;
  wire _abc_40344_n2415;
  wire _abc_40344_n2416_1;
  wire _abc_40344_n2417;
  wire _abc_40344_n2418;
  wire _abc_40344_n2419;
  wire _abc_40344_n2420;
  wire _abc_40344_n2421;
  wire _abc_40344_n2422;
  wire _abc_40344_n2423;
  wire _abc_40344_n2424;
  wire _abc_40344_n2425;
  wire _abc_40344_n2426;
  wire _abc_40344_n2427;
  wire _abc_40344_n2428_1;
  wire _abc_40344_n2429;
  wire _abc_40344_n2430;
  wire _abc_40344_n2431;
  wire _abc_40344_n2432;
  wire _abc_40344_n2433;
  wire _abc_40344_n2434;
  wire _abc_40344_n2435_1;
  wire _abc_40344_n2436;
  wire _abc_40344_n2437;
  wire _abc_40344_n2438;
  wire _abc_40344_n2439;
  wire _abc_40344_n2440;
  wire _abc_40344_n2441;
  wire _abc_40344_n2442;
  wire _abc_40344_n2443;
  wire _abc_40344_n2444;
  wire _abc_40344_n2445;
  wire _abc_40344_n2446;
  wire _abc_40344_n2447;
  wire _abc_40344_n2448;
  wire _abc_40344_n2449;
  wire _abc_40344_n2450;
  wire _abc_40344_n2451_1;
  wire _abc_40344_n2452;
  wire _abc_40344_n2453;
  wire _abc_40344_n2454;
  wire _abc_40344_n2455;
  wire _abc_40344_n2456;
  wire _abc_40344_n2457;
  wire _abc_40344_n2458_1;
  wire _abc_40344_n2459;
  wire _abc_40344_n2460;
  wire _abc_40344_n2461;
  wire _abc_40344_n2462;
  wire _abc_40344_n2463;
  wire _abc_40344_n2464;
  wire _abc_40344_n2465;
  wire _abc_40344_n2466;
  wire _abc_40344_n2467;
  wire _abc_40344_n2468;
  wire _abc_40344_n2469;
  wire _abc_40344_n2470;
  wire _abc_40344_n2471;
  wire _abc_40344_n2472;
  wire _abc_40344_n2473;
  wire _abc_40344_n2474;
  wire _abc_40344_n2475;
  wire _abc_40344_n2476;
  wire _abc_40344_n2477;
  wire _abc_40344_n2478_1;
  wire _abc_40344_n2479;
  wire _abc_40344_n2480;
  wire _abc_40344_n2481;
  wire _abc_40344_n2482;
  wire _abc_40344_n2483;
  wire _abc_40344_n2484_1;
  wire _abc_40344_n2485;
  wire _abc_40344_n2486;
  wire _abc_40344_n2487;
  wire _abc_40344_n2488;
  wire _abc_40344_n2489;
  wire _abc_40344_n2490;
  wire _abc_40344_n2491;
  wire _abc_40344_n2492;
  wire _abc_40344_n2493;
  wire _abc_40344_n2494;
  wire _abc_40344_n2495;
  wire _abc_40344_n2496_1;
  wire _abc_40344_n2497;
  wire _abc_40344_n2498;
  wire _abc_40344_n2499;
  wire _abc_40344_n2500;
  wire _abc_40344_n2501;
  wire _abc_40344_n2502_1;
  wire _abc_40344_n2503;
  wire _abc_40344_n2504;
  wire _abc_40344_n2505;
  wire _abc_40344_n2506;
  wire _abc_40344_n2507;
  wire _abc_40344_n2508;
  wire _abc_40344_n2509;
  wire _abc_40344_n2510;
  wire _abc_40344_n2511;
  wire _abc_40344_n2512;
  wire _abc_40344_n2513;
  wire _abc_40344_n2514;
  wire _abc_40344_n2515;
  wire _abc_40344_n2516;
  wire _abc_40344_n2517;
  wire _abc_40344_n2518;
  wire _abc_40344_n2519;
  wire _abc_40344_n2520;
  wire _abc_40344_n2521;
  wire _abc_40344_n2522;
  wire _abc_40344_n2523_1;
  wire _abc_40344_n2524;
  wire _abc_40344_n2525;
  wire _abc_40344_n2526;
  wire _abc_40344_n2527;
  wire _abc_40344_n2528;
  wire _abc_40344_n2529_1;
  wire _abc_40344_n2530;
  wire _abc_40344_n2531;
  wire _abc_40344_n2532;
  wire _abc_40344_n2533;
  wire _abc_40344_n2534;
  wire _abc_40344_n2535;
  wire _abc_40344_n2536;
  wire _abc_40344_n2537;
  wire _abc_40344_n2538;
  wire _abc_40344_n2539;
  wire _abc_40344_n2540;
  wire _abc_40344_n2541;
  wire _abc_40344_n2542;
  wire _abc_40344_n2543_1;
  wire _abc_40344_n2544;
  wire _abc_40344_n2545;
  wire _abc_40344_n2546;
  wire _abc_40344_n2547;
  wire _abc_40344_n2548;
  wire _abc_40344_n2549_1;
  wire _abc_40344_n2550;
  wire _abc_40344_n2551;
  wire _abc_40344_n2552;
  wire _abc_40344_n2553;
  wire _abc_40344_n2554;
  wire _abc_40344_n2555;
  wire _abc_40344_n2556;
  wire _abc_40344_n2557;
  wire _abc_40344_n2558;
  wire _abc_40344_n2559;
  wire _abc_40344_n2560;
  wire _abc_40344_n2561;
  wire _abc_40344_n2562;
  wire _abc_40344_n2563;
  wire _abc_40344_n2564;
  wire _abc_40344_n2565;
  wire _abc_40344_n2566;
  wire _abc_40344_n2567_1;
  wire _abc_40344_n2568;
  wire _abc_40344_n2569;
  wire _abc_40344_n2570;
  wire _abc_40344_n2571;
  wire _abc_40344_n2572;
  wire _abc_40344_n2573_1;
  wire _abc_40344_n2574;
  wire _abc_40344_n2575;
  wire _abc_40344_n2576;
  wire _abc_40344_n2577;
  wire _abc_40344_n2578;
  wire _abc_40344_n2579;
  wire _abc_40344_n2580;
  wire _abc_40344_n2581;
  wire _abc_40344_n2582;
  wire _abc_40344_n2583;
  wire _abc_40344_n2584;
  wire _abc_40344_n2585;
  wire _abc_40344_n2586;
  wire _abc_40344_n2587;
  wire _abc_40344_n2588;
  wire _abc_40344_n2589;
  wire _abc_40344_n2590;
  wire _abc_40344_n2591;
  wire _abc_40344_n2592;
  wire _abc_40344_n2593_1;
  wire _abc_40344_n2594;
  wire _abc_40344_n2595;
  wire _abc_40344_n2596;
  wire _abc_40344_n2597;
  wire _abc_40344_n2598;
  wire _abc_40344_n2599_1;
  wire _abc_40344_n2600;
  wire _abc_40344_n2601;
  wire _abc_40344_n2602;
  wire _abc_40344_n2603;
  wire _abc_40344_n2604;
  wire _abc_40344_n2605;
  wire _abc_40344_n2606;
  wire _abc_40344_n2607;
  wire _abc_40344_n2608;
  wire _abc_40344_n2609;
  wire _abc_40344_n2610;
  wire _abc_40344_n2611;
  wire _abc_40344_n2612;
  wire _abc_40344_n2613;
  wire _abc_40344_n2614;
  wire _abc_40344_n2615;
  wire _abc_40344_n2616;
  wire _abc_40344_n2617;
  wire _abc_40344_n2618;
  wire _abc_40344_n2619_1;
  wire _abc_40344_n2620;
  wire _abc_40344_n2621;
  wire _abc_40344_n2622;
  wire _abc_40344_n2623;
  wire _abc_40344_n2624;
  wire _abc_40344_n2625_1;
  wire _abc_40344_n2626;
  wire _abc_40344_n2627;
  wire _abc_40344_n2628;
  wire _abc_40344_n2629;
  wire _abc_40344_n2630;
  wire _abc_40344_n2631;
  wire _abc_40344_n2632;
  wire _abc_40344_n2633;
  wire _abc_40344_n2634;
  wire _abc_40344_n2635;
  wire _abc_40344_n2636;
  wire _abc_40344_n2637;
  wire _abc_40344_n2638;
  wire _abc_40344_n2639;
  wire _abc_40344_n2640;
  wire _abc_40344_n2641;
  wire _abc_40344_n2642;
  wire _abc_40344_n2643;
  wire _abc_40344_n2644_1;
  wire _abc_40344_n2645;
  wire _abc_40344_n2646;
  wire _abc_40344_n2647;
  wire _abc_40344_n2648;
  wire _abc_40344_n2649;
  wire _abc_40344_n2650_1;
  wire _abc_40344_n2651;
  wire _abc_40344_n2652;
  wire _abc_40344_n2653;
  wire _abc_40344_n2654;
  wire _abc_40344_n2655;
  wire _abc_40344_n2656;
  wire _abc_40344_n2657;
  wire _abc_40344_n2658;
  wire _abc_40344_n2659;
  wire _abc_40344_n2660;
  wire _abc_40344_n2661;
  wire _abc_40344_n2662;
  wire _abc_40344_n2663;
  wire _abc_40344_n2664;
  wire _abc_40344_n2665;
  wire _abc_40344_n2666_1;
  wire _abc_40344_n2667;
  wire _abc_40344_n2668;
  wire _abc_40344_n2669;
  wire _abc_40344_n2670;
  wire _abc_40344_n2671;
  wire _abc_40344_n2673;
  wire _abc_40344_n2674;
  wire _abc_40344_n2675;
  wire _abc_40344_n2676;
  wire _abc_40344_n2677;
  wire _abc_40344_n2678;
  wire _abc_40344_n2679;
  wire _abc_40344_n2680;
  wire _abc_40344_n2681;
  wire _abc_40344_n2682;
  wire _abc_40344_n2683;
  wire _abc_40344_n2684;
  wire _abc_40344_n2685;
  wire _abc_40344_n2687;
  wire _abc_40344_n2688;
  wire _abc_40344_n2689;
  wire _abc_40344_n2690;
  wire _abc_40344_n2691;
  wire _abc_40344_n2692_1;
  wire _abc_40344_n2693;
  wire _abc_40344_n2694;
  wire _abc_40344_n2695;
  wire _abc_40344_n2696;
  wire _abc_40344_n2697;
  wire _abc_40344_n2698_1;
  wire _abc_40344_n2699;
  wire _abc_40344_n2700;
  wire _abc_40344_n2701;
  wire _abc_40344_n2702;
  wire _abc_40344_n2703;
  wire _abc_40344_n2704;
  wire _abc_40344_n2705;
  wire _abc_40344_n2706;
  wire _abc_40344_n2708;
  wire _abc_40344_n2709;
  wire _abc_40344_n2710;
  wire _abc_40344_n2711;
  wire _abc_40344_n2712;
  wire _abc_40344_n2713;
  wire _abc_40344_n2714;
  wire _abc_40344_n2715;
  wire _abc_40344_n2716;
  wire _abc_40344_n2717;
  wire _abc_40344_n2718;
  wire _abc_40344_n2719;
  wire _abc_40344_n2720;
  wire _abc_40344_n2721;
  wire _abc_40344_n2722_1;
  wire _abc_40344_n2723;
  wire _abc_40344_n2724;
  wire _abc_40344_n2725;
  wire _abc_40344_n2727;
  wire _abc_40344_n2728;
  wire _abc_40344_n2729;
  wire _abc_40344_n2730_1;
  wire _abc_40344_n2731;
  wire _abc_40344_n2732;
  wire _abc_40344_n2733;
  wire _abc_40344_n2734;
  wire _abc_40344_n2735;
  wire _abc_40344_n2736;
  wire _abc_40344_n2737;
  wire _abc_40344_n2738;
  wire _abc_40344_n2739;
  wire _abc_40344_n2740;
  wire _abc_40344_n2741;
  wire _abc_40344_n2742;
  wire _abc_40344_n2743;
  wire _abc_40344_n2744;
  wire _abc_40344_n2746;
  wire _abc_40344_n2747;
  wire _abc_40344_n2748;
  wire _abc_40344_n2749;
  wire _abc_40344_n2750;
  wire _abc_40344_n2751;
  wire _abc_40344_n2752;
  wire _abc_40344_n2753;
  wire _abc_40344_n2754;
  wire _abc_40344_n2755;
  wire _abc_40344_n2756;
  wire _abc_40344_n2757;
  wire _abc_40344_n2758;
  wire _abc_40344_n2760_1;
  wire _abc_40344_n2761;
  wire _abc_40344_n2762;
  wire _abc_40344_n2763;
  wire _abc_40344_n2764;
  wire _abc_40344_n2765;
  wire _abc_40344_n2766;
  wire _abc_40344_n2767;
  wire _abc_40344_n2768_1;
  wire _abc_40344_n2769;
  wire _abc_40344_n2770;
  wire _abc_40344_n2771;
  wire _abc_40344_n2772;
  wire _abc_40344_n2774;
  wire _abc_40344_n2775;
  wire _abc_40344_n2776;
  wire _abc_40344_n2777;
  wire _abc_40344_n2778;
  wire _abc_40344_n2779;
  wire _abc_40344_n2780;
  wire _abc_40344_n2781;
  wire _abc_40344_n2782;
  wire _abc_40344_n2783;
  wire _abc_40344_n2784;
  wire _abc_40344_n2785;
  wire _abc_40344_n2786;
  wire _abc_40344_n2787;
  wire _abc_40344_n2788;
  wire _abc_40344_n2789;
  wire _abc_40344_n2790;
  wire _abc_40344_n2791;
  wire _abc_40344_n2792;
  wire _abc_40344_n2793;
  wire _abc_40344_n2795;
  wire _abc_40344_n2796;
  wire _abc_40344_n2797;
  wire _abc_40344_n2798;
  wire _abc_40344_n2799;
  wire _abc_40344_n2800;
  wire _abc_40344_n2801;
  wire _abc_40344_n2802;
  wire _abc_40344_n2803;
  wire _abc_40344_n2804;
  wire _abc_40344_n2805;
  wire _abc_40344_n2806;
  wire _abc_40344_n2807;
  wire _abc_40344_n2808;
  wire _abc_40344_n2809;
  wire _abc_40344_n2810;
  wire _abc_40344_n2812;
  wire _abc_40344_n2813;
  wire _abc_40344_n2814;
  wire _abc_40344_n2815;
  wire _abc_40344_n2816_1;
  wire _abc_40344_n2817;
  wire _abc_40344_n2818;
  wire _abc_40344_n2819;
  wire _abc_40344_n2820;
  wire _abc_40344_n2821;
  wire _abc_40344_n2822;
  wire _abc_40344_n2823_1;
  wire _abc_40344_n2824;
  wire _abc_40344_n2825;
  wire _abc_40344_n2826;
  wire _abc_40344_n2828;
  wire _abc_40344_n2829;
  wire _abc_40344_n2830;
  wire _abc_40344_n2831;
  wire _abc_40344_n2832;
  wire _abc_40344_n2833;
  wire _abc_40344_n2834;
  wire _abc_40344_n2835;
  wire _abc_40344_n2836;
  wire _abc_40344_n2837;
  wire _abc_40344_n2838;
  wire _abc_40344_n2839;
  wire _abc_40344_n2840;
  wire _abc_40344_n2841;
  wire _abc_40344_n2843;
  wire _abc_40344_n2844;
  wire _abc_40344_n2845;
  wire _abc_40344_n2846;
  wire _abc_40344_n2847;
  wire _abc_40344_n2848;
  wire _abc_40344_n2849;
  wire _abc_40344_n2850;
  wire _abc_40344_n2851;
  wire _abc_40344_n2852;
  wire _abc_40344_n2853;
  wire _abc_40344_n2854;
  wire _abc_40344_n2855;
  wire _abc_40344_n2856;
  wire _abc_40344_n2857;
  wire _abc_40344_n2858;
  wire _abc_40344_n2859;
  wire _abc_40344_n2860;
  wire _abc_40344_n2861;
  wire _abc_40344_n2863;
  wire _abc_40344_n2864;
  wire _abc_40344_n2865;
  wire _abc_40344_n2866;
  wire _abc_40344_n2867;
  wire _abc_40344_n2868;
  wire _abc_40344_n2869;
  wire _abc_40344_n2870;
  wire _abc_40344_n2871;
  wire _abc_40344_n2872;
  wire _abc_40344_n2873;
  wire _abc_40344_n2874;
  wire _abc_40344_n2875;
  wire _abc_40344_n2876;
  wire _abc_40344_n2877;
  wire _abc_40344_n2878;
  wire _abc_40344_n2879;
  wire _abc_40344_n2880;
  wire _abc_40344_n2882;
  wire _abc_40344_n2883;
  wire _abc_40344_n2884;
  wire _abc_40344_n2885;
  wire _abc_40344_n2886;
  wire _abc_40344_n2887;
  wire _abc_40344_n2888;
  wire _abc_40344_n2889;
  wire _abc_40344_n2890;
  wire _abc_40344_n2891;
  wire _abc_40344_n2892;
  wire _abc_40344_n2893;
  wire _abc_40344_n2894;
  wire _abc_40344_n2895;
  wire _abc_40344_n2896;
  wire _abc_40344_n2897;
  wire _abc_40344_n2898;
  wire _abc_40344_n2899;
  wire _abc_40344_n2900;
  wire _abc_40344_n2901;
  wire _abc_40344_n2902;
  wire _abc_40344_n2904;
  wire _abc_40344_n2905;
  wire _abc_40344_n2906;
  wire _abc_40344_n2907;
  wire _abc_40344_n2908;
  wire _abc_40344_n2909;
  wire _abc_40344_n2910;
  wire _abc_40344_n2911;
  wire _abc_40344_n2912;
  wire _abc_40344_n2913;
  wire _abc_40344_n2914;
  wire _abc_40344_n2915;
  wire _abc_40344_n2916;
  wire _abc_40344_n2917;
  wire _abc_40344_n2918;
  wire _abc_40344_n2919;
  wire _abc_40344_n2920;
  wire _abc_40344_n2921;
  wire _abc_40344_n2922;
  wire _abc_40344_n2923;
  wire _abc_40344_n2925;
  wire _abc_40344_n2926;
  wire _abc_40344_n2927;
  wire _abc_40344_n2928;
  wire _abc_40344_n2929;
  wire _abc_40344_n2930;
  wire _abc_40344_n2931;
  wire _abc_40344_n2932;
  wire _abc_40344_n2933;
  wire _abc_40344_n2934;
  wire _abc_40344_n2935;
  wire _abc_40344_n2936;
  wire _abc_40344_n2937;
  wire _abc_40344_n2938;
  wire _abc_40344_n2939;
  wire _abc_40344_n2940;
  wire _abc_40344_n2941;
  wire _abc_40344_n2942;
  wire _abc_40344_n2943;
  wire _abc_40344_n2944;
  wire _abc_40344_n2945;
  wire _abc_40344_n2946;
  wire _abc_40344_n2947;
  wire _abc_40344_n2949;
  wire _abc_40344_n2950;
  wire _abc_40344_n2951;
  wire _abc_40344_n2952;
  wire _abc_40344_n2953;
  wire _abc_40344_n2954;
  wire _abc_40344_n2955;
  wire _abc_40344_n2956;
  wire _abc_40344_n2957;
  wire _abc_40344_n2958;
  wire _abc_40344_n2959;
  wire _abc_40344_n2960;
  wire _abc_40344_n2961;
  wire _abc_40344_n2962;
  wire _abc_40344_n2963;
  wire _abc_40344_n2964;
  wire _abc_40344_n2965;
  wire _abc_40344_n2966;
  wire _abc_40344_n2967;
  wire _abc_40344_n2968;
  wire _abc_40344_n2970;
  wire _abc_40344_n2971;
  wire _abc_40344_n2972;
  wire _abc_40344_n2973;
  wire _abc_40344_n2974;
  wire _abc_40344_n2975;
  wire _abc_40344_n2976;
  wire _abc_40344_n2977;
  wire _abc_40344_n2978;
  wire _abc_40344_n2979;
  wire _abc_40344_n2980;
  wire _abc_40344_n2981;
  wire _abc_40344_n2982;
  wire _abc_40344_n2983;
  wire _abc_40344_n2984;
  wire _abc_40344_n2985;
  wire _abc_40344_n2986;
  wire _abc_40344_n2987;
  wire _abc_40344_n2988;
  wire _abc_40344_n2989;
  wire _abc_40344_n2991;
  wire _abc_40344_n2992;
  wire _abc_40344_n2993;
  wire _abc_40344_n2994;
  wire _abc_40344_n2995;
  wire _abc_40344_n2996;
  wire _abc_40344_n2997;
  wire _abc_40344_n2998;
  wire _abc_40344_n2999;
  wire _abc_40344_n3000;
  wire _abc_40344_n3001;
  wire _abc_40344_n3002;
  wire _abc_40344_n3003;
  wire _abc_40344_n3004;
  wire _abc_40344_n3005;
  wire _abc_40344_n3006;
  wire _abc_40344_n3007;
  wire _abc_40344_n3008;
  wire _abc_40344_n3009;
  wire _abc_40344_n3010;
  wire _abc_40344_n3011;
  wire _abc_40344_n3012;
  wire _abc_40344_n3014;
  wire _abc_40344_n3015;
  wire _abc_40344_n3016;
  wire _abc_40344_n3017;
  wire _abc_40344_n3018;
  wire _abc_40344_n3019;
  wire _abc_40344_n3020;
  wire _abc_40344_n3021;
  wire _abc_40344_n3022;
  wire _abc_40344_n3023;
  wire _abc_40344_n3024;
  wire _abc_40344_n3025;
  wire _abc_40344_n3026;
  wire _abc_40344_n3027;
  wire _abc_40344_n3028;
  wire _abc_40344_n3029;
  wire _abc_40344_n3030;
  wire _abc_40344_n3031;
  wire _abc_40344_n3032;
  wire _abc_40344_n3034;
  wire _abc_40344_n3035;
  wire _abc_40344_n3036;
  wire _abc_40344_n3037;
  wire _abc_40344_n3038;
  wire _abc_40344_n3039;
  wire _abc_40344_n3040;
  wire _abc_40344_n3041_1;
  wire _abc_40344_n3042;
  wire _abc_40344_n3043;
  wire _abc_40344_n3044;
  wire _abc_40344_n3045;
  wire _abc_40344_n3046;
  wire _abc_40344_n3047;
  wire _abc_40344_n3048;
  wire _abc_40344_n3049;
  wire _abc_40344_n3050;
  wire _abc_40344_n3051;
  wire _abc_40344_n3052;
  wire _abc_40344_n3053;
  wire _abc_40344_n3054;
  wire _abc_40344_n3055;
  wire _abc_40344_n3056;
  wire _abc_40344_n3057;
  wire _abc_40344_n3058;
  wire _abc_40344_n3059;
  wire _abc_40344_n3061;
  wire _abc_40344_n3062;
  wire _abc_40344_n3063;
  wire _abc_40344_n3064;
  wire _abc_40344_n3065;
  wire _abc_40344_n3066;
  wire _abc_40344_n3066_bF_buf0;
  wire _abc_40344_n3066_bF_buf1;
  wire _abc_40344_n3066_bF_buf2;
  wire _abc_40344_n3066_bF_buf3;
  wire _abc_40344_n3066_bF_buf4;
  wire _abc_40344_n3066_bF_buf5;
  wire _abc_40344_n3067;
  wire _abc_40344_n3067_bF_buf0;
  wire _abc_40344_n3067_bF_buf1;
  wire _abc_40344_n3067_bF_buf2;
  wire _abc_40344_n3067_bF_buf3;
  wire _abc_40344_n3067_bF_buf4;
  wire _abc_40344_n3067_bF_buf5;
  wire _abc_40344_n3068;
  wire _abc_40344_n3069;
  wire _abc_40344_n3070;
  wire _abc_40344_n3071;
  wire _abc_40344_n3072;
  wire _abc_40344_n3073;
  wire _abc_40344_n3074;
  wire _abc_40344_n3075;
  wire _abc_40344_n3076;
  wire _abc_40344_n3077;
  wire _abc_40344_n3078;
  wire _abc_40344_n3079;
  wire _abc_40344_n3080;
  wire _abc_40344_n3081_1;
  wire _abc_40344_n3082;
  wire _abc_40344_n3083;
  wire _abc_40344_n3084;
  wire _abc_40344_n3085;
  wire _abc_40344_n3086;
  wire _abc_40344_n3087;
  wire _abc_40344_n3088;
  wire _abc_40344_n3089;
  wire _abc_40344_n3090;
  wire _abc_40344_n3091;
  wire _abc_40344_n3092;
  wire _abc_40344_n3093;
  wire _abc_40344_n3094;
  wire _abc_40344_n3095;
  wire _abc_40344_n3096;
  wire _abc_40344_n3097;
  wire _abc_40344_n3098;
  wire _abc_40344_n3099;
  wire _abc_40344_n3100;
  wire _abc_40344_n3101;
  wire _abc_40344_n3102;
  wire _abc_40344_n3103;
  wire _abc_40344_n3103_bF_buf0;
  wire _abc_40344_n3103_bF_buf1;
  wire _abc_40344_n3103_bF_buf2;
  wire _abc_40344_n3103_bF_buf3;
  wire _abc_40344_n3104;
  wire _abc_40344_n3105;
  wire _abc_40344_n3106;
  wire _abc_40344_n3107;
  wire _abc_40344_n3108;
  wire _abc_40344_n3109;
  wire _abc_40344_n3109_bF_buf0;
  wire _abc_40344_n3109_bF_buf1;
  wire _abc_40344_n3109_bF_buf2;
  wire _abc_40344_n3109_bF_buf3;
  wire _abc_40344_n3110;
  wire _abc_40344_n3111;
  wire _abc_40344_n3112;
  wire _abc_40344_n3114;
  wire _abc_40344_n3115;
  wire _abc_40344_n3116;
  wire _abc_40344_n3117;
  wire _abc_40344_n3118;
  wire _abc_40344_n3120;
  wire _abc_40344_n3121;
  wire _abc_40344_n3122;
  wire _abc_40344_n3123;
  wire _abc_40344_n3124;
  wire _abc_40344_n3125_1;
  wire _abc_40344_n3126;
  wire _abc_40344_n3127;
  wire _abc_40344_n3128;
  wire _abc_40344_n3129;
  wire _abc_40344_n3130;
  wire _abc_40344_n3131;
  wire _abc_40344_n3132;
  wire _abc_40344_n3133;
  wire _abc_40344_n3134;
  wire _abc_40344_n3135;
  wire _abc_40344_n3136;
  wire _abc_40344_n3137;
  wire _abc_40344_n3138;
  wire _abc_40344_n3139;
  wire _abc_40344_n3140;
  wire _abc_40344_n3141;
  wire _abc_40344_n3142;
  wire _abc_40344_n3143;
  wire _abc_40344_n3144;
  wire _abc_40344_n3145;
  wire _abc_40344_n3146;
  wire _abc_40344_n3147_1;
  wire _abc_40344_n3148;
  wire _abc_40344_n3149;
  wire _abc_40344_n3150;
  wire _abc_40344_n3151;
  wire _abc_40344_n3152;
  wire _abc_40344_n3153;
  wire _abc_40344_n3154;
  wire _abc_40344_n3155;
  wire _abc_40344_n3156;
  wire _abc_40344_n3157;
  wire _abc_40344_n3158;
  wire _abc_40344_n3159;
  wire _abc_40344_n3160;
  wire _abc_40344_n3161;
  wire _abc_40344_n3162;
  wire _abc_40344_n3163;
  wire _abc_40344_n3164;
  wire _abc_40344_n3165;
  wire _abc_40344_n3166;
  wire _abc_40344_n3167;
  wire _abc_40344_n3168;
  wire _abc_40344_n3169;
  wire _abc_40344_n3170;
  wire _abc_40344_n3171;
  wire _abc_40344_n3172_1;
  wire _abc_40344_n3173;
  wire _abc_40344_n3174;
  wire _abc_40344_n3175;
  wire _abc_40344_n3176;
  wire _abc_40344_n3177;
  wire _abc_40344_n3178;
  wire _abc_40344_n3179;
  wire _abc_40344_n3180;
  wire _abc_40344_n3181;
  wire _abc_40344_n3182;
  wire _abc_40344_n3183;
  wire _abc_40344_n3184;
  wire _abc_40344_n3185;
  wire _abc_40344_n3186;
  wire _abc_40344_n3187;
  wire _abc_40344_n3188;
  wire _abc_40344_n3189;
  wire _abc_40344_n3190;
  wire _abc_40344_n3191;
  wire _abc_40344_n3192;
  wire _abc_40344_n3193;
  wire _abc_40344_n3194;
  wire _abc_40344_n3195;
  wire _abc_40344_n3196;
  wire _abc_40344_n3197;
  wire _abc_40344_n3198;
  wire _abc_40344_n3199;
  wire _abc_40344_n3200;
  wire _abc_40344_n3201;
  wire _abc_40344_n3202;
  wire _abc_40344_n3203;
  wire _abc_40344_n3204;
  wire _abc_40344_n3205;
  wire _abc_40344_n3206;
  wire _abc_40344_n3207;
  wire _abc_40344_n3208;
  wire _abc_40344_n3209;
  wire _abc_40344_n3210;
  wire _abc_40344_n3211;
  wire _abc_40344_n3212;
  wire _abc_40344_n3213;
  wire _abc_40344_n3214;
  wire _abc_40344_n3215;
  wire _abc_40344_n3216;
  wire _abc_40344_n3217;
  wire _abc_40344_n3218;
  wire _abc_40344_n3219;
  wire _abc_40344_n3220;
  wire _abc_40344_n3220_bF_buf0;
  wire _abc_40344_n3220_bF_buf1;
  wire _abc_40344_n3220_bF_buf2;
  wire _abc_40344_n3220_bF_buf3;
  wire _abc_40344_n3220_bF_buf4;
  wire _abc_40344_n3221_1;
  wire _abc_40344_n3222;
  wire _abc_40344_n3223;
  wire _abc_40344_n3223_bF_buf0;
  wire _abc_40344_n3223_bF_buf1;
  wire _abc_40344_n3223_bF_buf2;
  wire _abc_40344_n3223_bF_buf3;
  wire _abc_40344_n3224;
  wire _abc_40344_n3225;
  wire _abc_40344_n3226;
  wire _abc_40344_n3227;
  wire _abc_40344_n3228;
  wire _abc_40344_n3228_bF_buf0;
  wire _abc_40344_n3228_bF_buf1;
  wire _abc_40344_n3228_bF_buf2;
  wire _abc_40344_n3228_bF_buf3;
  wire _abc_40344_n3229;
  wire _abc_40344_n3230;
  wire _abc_40344_n3231;
  wire _abc_40344_n3232;
  wire _abc_40344_n3233;
  wire _abc_40344_n3234;
  wire _abc_40344_n3235;
  wire _abc_40344_n3236;
  wire _abc_40344_n3237;
  wire _abc_40344_n3238;
  wire _abc_40344_n3239;
  wire _abc_40344_n3240;
  wire _abc_40344_n3241;
  wire _abc_40344_n3242;
  wire _abc_40344_n3244;
  wire _abc_40344_n3245;
  wire _abc_40344_n3246;
  wire _abc_40344_n3247;
  wire _abc_40344_n3248;
  wire _abc_40344_n3249;
  wire _abc_40344_n3250;
  wire _abc_40344_n3251;
  wire _abc_40344_n3252;
  wire _abc_40344_n3253;
  wire _abc_40344_n3254;
  wire _abc_40344_n3255;
  wire _abc_40344_n3256;
  wire _abc_40344_n3257;
  wire _abc_40344_n3258;
  wire _abc_40344_n3259;
  wire _abc_40344_n3261;
  wire _abc_40344_n3262;
  wire _abc_40344_n3263;
  wire _abc_40344_n3264;
  wire _abc_40344_n3265;
  wire _abc_40344_n3266;
  wire _abc_40344_n3267;
  wire _abc_40344_n3268;
  wire _abc_40344_n3269_1;
  wire _abc_40344_n3270;
  wire _abc_40344_n3271;
  wire _abc_40344_n3272;
  wire _abc_40344_n3273;
  wire _abc_40344_n3274;
  wire _abc_40344_n3275;
  wire _abc_40344_n3276;
  wire _abc_40344_n3277;
  wire _abc_40344_n3278;
  wire _abc_40344_n3279;
  wire _abc_40344_n3280;
  wire _abc_40344_n3281;
  wire _abc_40344_n3283;
  wire _abc_40344_n3284;
  wire _abc_40344_n3285;
  wire _abc_40344_n3286;
  wire _abc_40344_n3287;
  wire _abc_40344_n3288;
  wire _abc_40344_n3289;
  wire _abc_40344_n3290;
  wire _abc_40344_n3291;
  wire _abc_40344_n3292;
  wire _abc_40344_n3293;
  wire _abc_40344_n3294;
  wire _abc_40344_n3296;
  wire _abc_40344_n3297;
  wire _abc_40344_n3298;
  wire _abc_40344_n3299;
  wire _abc_40344_n3300;
  wire _abc_40344_n3301;
  wire _abc_40344_n3302;
  wire _abc_40344_n3303;
  wire _abc_40344_n3304;
  wire _abc_40344_n3305;
  wire _abc_40344_n3306;
  wire _abc_40344_n3307;
  wire _abc_40344_n3308;
  wire _abc_40344_n3309;
  wire _abc_40344_n3310;
  wire _abc_40344_n3311;
  wire _abc_40344_n3312;
  wire _abc_40344_n3313;
  wire _abc_40344_n3314_1;
  wire _abc_40344_n3315;
  wire _abc_40344_n3316;
  wire _abc_40344_n3317;
  wire _abc_40344_n3318;
  wire _abc_40344_n3319;
  wire _abc_40344_n3320;
  wire _abc_40344_n3321;
  wire _abc_40344_n3322;
  wire _abc_40344_n3323;
  wire _abc_40344_n3324;
  wire _abc_40344_n3325;
  wire _abc_40344_n3326;
  wire _abc_40344_n3327;
  wire _abc_40344_n3328;
  wire _abc_40344_n3329;
  wire _abc_40344_n3330;
  wire _abc_40344_n3331;
  wire _abc_40344_n3332;
  wire _abc_40344_n3333;
  wire _abc_40344_n3334;
  wire _abc_40344_n3335_1;
  wire _abc_40344_n3336;
  wire _abc_40344_n3337;
  wire _abc_40344_n3338;
  wire _abc_40344_n3339;
  wire _abc_40344_n3340;
  wire _abc_40344_n3341;
  wire _abc_40344_n3342;
  wire _abc_40344_n3343;
  wire _abc_40344_n3344;
  wire _abc_40344_n3345;
  wire _abc_40344_n3346;
  wire _abc_40344_n3347;
  wire _abc_40344_n3348;
  wire _abc_40344_n3349;
  wire _abc_40344_n3351;
  wire _abc_40344_n3352;
  wire _abc_40344_n3353;
  wire _abc_40344_n3354;
  wire _abc_40344_n3355;
  wire _abc_40344_n3356;
  wire _abc_40344_n3357;
  wire _abc_40344_n3358;
  wire _abc_40344_n3359_1;
  wire _abc_40344_n3360;
  wire _abc_40344_n3361;
  wire _abc_40344_n3362;
  wire _abc_40344_n3363;
  wire _abc_40344_n3364;
  wire _abc_40344_n3365;
  wire _abc_40344_n3366;
  wire _abc_40344_n3367;
  wire _abc_40344_n3368;
  wire _abc_40344_n3369;
  wire _abc_40344_n3370;
  wire _abc_40344_n3371;
  wire _abc_40344_n3372;
  wire _abc_40344_n3373;
  wire _abc_40344_n3374;
  wire _abc_40344_n3375;
  wire _abc_40344_n3376;
  wire _abc_40344_n3377;
  wire _abc_40344_n3379;
  wire _abc_40344_n3380;
  wire _abc_40344_n3381;
  wire _abc_40344_n3382;
  wire _abc_40344_n3383;
  wire _abc_40344_n3384;
  wire _abc_40344_n3385;
  wire _abc_40344_n3386;
  wire _abc_40344_n3387;
  wire _abc_40344_n3388_1;
  wire _abc_40344_n3389;
  wire _abc_40344_n3390;
  wire _abc_40344_n3391;
  wire _abc_40344_n3392;
  wire _abc_40344_n3393;
  wire _abc_40344_n3394;
  wire _abc_40344_n3396;
  wire _abc_40344_n3397;
  wire _abc_40344_n3398;
  wire _abc_40344_n3399;
  wire _abc_40344_n3400;
  wire _abc_40344_n3401;
  wire _abc_40344_n3402;
  wire _abc_40344_n3403;
  wire _abc_40344_n3404;
  wire _abc_40344_n3405;
  wire _abc_40344_n3406;
  wire _abc_40344_n3407;
  wire _abc_40344_n3408;
  wire _abc_40344_n3409;
  wire _abc_40344_n3410;
  wire _abc_40344_n3411_1;
  wire _abc_40344_n3412;
  wire _abc_40344_n3413;
  wire _abc_40344_n3414;
  wire _abc_40344_n3415;
  wire _abc_40344_n3416;
  wire _abc_40344_n3417;
  wire _abc_40344_n3418;
  wire _abc_40344_n3419;
  wire _abc_40344_n3420;
  wire _abc_40344_n3421;
  wire _abc_40344_n3423;
  wire _abc_40344_n3424;
  wire _abc_40344_n3425;
  wire _abc_40344_n3426;
  wire _abc_40344_n3427;
  wire _abc_40344_n3428;
  wire _abc_40344_n3429;
  wire _abc_40344_n3430;
  wire _abc_40344_n3431_1;
  wire _abc_40344_n3432;
  wire _abc_40344_n3433;
  wire _abc_40344_n3434;
  wire _abc_40344_n3435;
  wire _abc_40344_n3436;
  wire _abc_40344_n3437;
  wire _abc_40344_n3438;
  wire _abc_40344_n3439;
  wire _abc_40344_n3440;
  wire _abc_40344_n3441;
  wire _abc_40344_n3442;
  wire _abc_40344_n3443;
  wire _abc_40344_n3445;
  wire _abc_40344_n3446;
  wire _abc_40344_n3447;
  wire _abc_40344_n3448;
  wire _abc_40344_n3449;
  wire _abc_40344_n3450;
  wire _abc_40344_n3451;
  wire _abc_40344_n3452;
  wire _abc_40344_n3453;
  wire _abc_40344_n3454;
  wire _abc_40344_n3455;
  wire _abc_40344_n3456;
  wire _abc_40344_n3457_1;
  wire _abc_40344_n3459;
  wire _abc_40344_n3460;
  wire _abc_40344_n3461;
  wire _abc_40344_n3462;
  wire _abc_40344_n3463;
  wire _abc_40344_n3464;
  wire _abc_40344_n3465;
  wire _abc_40344_n3466;
  wire _abc_40344_n3467;
  wire _abc_40344_n3468;
  wire _abc_40344_n3469;
  wire _abc_40344_n3470;
  wire _abc_40344_n3471;
  wire _abc_40344_n3472;
  wire _abc_40344_n3473;
  wire _abc_40344_n3474;
  wire _abc_40344_n3475;
  wire _abc_40344_n3476;
  wire _abc_40344_n3478_1;
  wire _abc_40344_n3479;
  wire _abc_40344_n3480;
  wire _abc_40344_n3481;
  wire _abc_40344_n3482;
  wire _abc_40344_n3483;
  wire _abc_40344_n3484;
  wire _abc_40344_n3485;
  wire _abc_40344_n3486;
  wire _abc_40344_n3487;
  wire _abc_40344_n3488;
  wire _abc_40344_n3489;
  wire _abc_40344_n3490;
  wire _abc_40344_n3491;
  wire _abc_40344_n3492;
  wire _abc_40344_n3493;
  wire _abc_40344_n3494;
  wire _abc_40344_n3495;
  wire _abc_40344_n3496;
  wire _abc_40344_n3497;
  wire _abc_40344_n3498;
  wire _abc_40344_n3500;
  wire _abc_40344_n3501;
  wire _abc_40344_n3502;
  wire _abc_40344_n3503;
  wire _abc_40344_n3504;
  wire _abc_40344_n3505;
  wire _abc_40344_n3506_1;
  wire _abc_40344_n3507;
  wire _abc_40344_n3508;
  wire _abc_40344_n3509;
  wire _abc_40344_n3510;
  wire _abc_40344_n3511;
  wire _abc_40344_n3512;
  wire _abc_40344_n3513;
  wire _abc_40344_n3514;
  wire _abc_40344_n3515;
  wire _abc_40344_n3516;
  wire _abc_40344_n3518;
  wire _abc_40344_n3519;
  wire _abc_40344_n3520;
  wire _abc_40344_n3521;
  wire _abc_40344_n3522;
  wire _abc_40344_n3523;
  wire _abc_40344_n3524;
  wire _abc_40344_n3525;
  wire _abc_40344_n3526;
  wire _abc_40344_n3527;
  wire _abc_40344_n3528;
  wire _abc_40344_n3529;
  wire _abc_40344_n3530;
  wire _abc_40344_n3531;
  wire _abc_40344_n3532;
  wire _abc_40344_n3533;
  wire _abc_40344_n3534;
  wire _abc_40344_n3535_1;
  wire _abc_40344_n3536;
  wire _abc_40344_n3537;
  wire _abc_40344_n3539;
  wire _abc_40344_n3540;
  wire _abc_40344_n3541;
  wire _abc_40344_n3542;
  wire _abc_40344_n3543;
  wire _abc_40344_n3544;
  wire _abc_40344_n3545;
  wire _abc_40344_n3546;
  wire _abc_40344_n3547;
  wire _abc_40344_n3548;
  wire _abc_40344_n3549;
  wire _abc_40344_n3550;
  wire _abc_40344_n3551;
  wire _abc_40344_n3552;
  wire _abc_40344_n3553;
  wire _abc_40344_n3554;
  wire _abc_40344_n3555_1;
  wire _abc_40344_n3557;
  wire _abc_40344_n3558;
  wire _abc_40344_n3559;
  wire _abc_40344_n3560;
  wire _abc_40344_n3561;
  wire _abc_40344_n3562;
  wire _abc_40344_n3563;
  wire _abc_40344_n3564;
  wire _abc_40344_n3565;
  wire _abc_40344_n3566;
  wire _abc_40344_n3567;
  wire _abc_40344_n3568;
  wire _abc_40344_n3569;
  wire _abc_40344_n3570;
  wire _abc_40344_n3571;
  wire _abc_40344_n3572;
  wire _abc_40344_n3574;
  wire _abc_40344_n3575;
  wire _abc_40344_n3576;
  wire _abc_40344_n3577;
  wire _abc_40344_n3578;
  wire _abc_40344_n3579;
  wire _abc_40344_n3580;
  wire _abc_40344_n3581_1;
  wire _abc_40344_n3582;
  wire _abc_40344_n3583;
  wire _abc_40344_n3584;
  wire _abc_40344_n3585;
  wire _abc_40344_n3586;
  wire _abc_40344_n3587;
  wire _abc_40344_n3588;
  wire _abc_40344_n3589;
  wire _abc_40344_n3590;
  wire _abc_40344_n3591;
  wire _abc_40344_n3593;
  wire _abc_40344_n3594;
  wire _abc_40344_n3595;
  wire _abc_40344_n3596;
  wire _abc_40344_n3597;
  wire _abc_40344_n3598;
  wire _abc_40344_n3599;
  wire _abc_40344_n3600;
  wire _abc_40344_n3601;
  wire _abc_40344_n3602;
  wire _abc_40344_n3603;
  wire _abc_40344_n3604_1;
  wire _abc_40344_n3605;
  wire _abc_40344_n3606;
  wire _abc_40344_n3607;
  wire _abc_40344_n3608;
  wire _abc_40344_n3610;
  wire _abc_40344_n3611;
  wire _abc_40344_n3612;
  wire _abc_40344_n3613;
  wire _abc_40344_n3614;
  wire _abc_40344_n3615;
  wire _abc_40344_n3616;
  wire _abc_40344_n3617;
  wire _abc_40344_n3618;
  wire _abc_40344_n3619;
  wire _abc_40344_n3620;
  wire _abc_40344_n3621;
  wire _abc_40344_n3622;
  wire _abc_40344_n3623;
  wire _abc_40344_n3624;
  wire _abc_40344_n3625;
  wire _abc_40344_n3626;
  wire _abc_40344_n3627;
  wire _abc_40344_n3628;
  wire _abc_40344_n3629;
  wire _abc_40344_n3630;
  wire _abc_40344_n3631;
  wire _abc_40344_n3632_1;
  wire _abc_40344_n3633;
  wire _abc_40344_n3635;
  wire _abc_40344_n3636;
  wire _abc_40344_n3637;
  wire _abc_40344_n3638;
  wire _abc_40344_n3639;
  wire _abc_40344_n3640;
  wire _abc_40344_n3641;
  wire _abc_40344_n3642;
  wire _abc_40344_n3643;
  wire _abc_40344_n3644;
  wire _abc_40344_n3645;
  wire _abc_40344_n3646;
  wire _abc_40344_n3647;
  wire _abc_40344_n3648;
  wire _abc_40344_n3649;
  wire _abc_40344_n3651;
  wire _abc_40344_n3652;
  wire _abc_40344_n3653;
  wire _abc_40344_n3654;
  wire _abc_40344_n3655;
  wire _abc_40344_n3656;
  wire _abc_40344_n3657;
  wire _abc_40344_n3658;
  wire _abc_40344_n3659;
  wire _abc_40344_n3660;
  wire _abc_40344_n3661;
  wire _abc_40344_n3662_1;
  wire _abc_40344_n3663;
  wire _abc_40344_n3664;
  wire _abc_40344_n3665;
  wire _abc_40344_n3666;
  wire _abc_40344_n3667;
  wire _abc_40344_n3668;
  wire _abc_40344_n3670;
  wire _abc_40344_n3671;
  wire _abc_40344_n3672;
  wire _abc_40344_n3673;
  wire _abc_40344_n3674;
  wire _abc_40344_n3675;
  wire _abc_40344_n3676;
  wire _abc_40344_n3677;
  wire _abc_40344_n3678;
  wire _abc_40344_n3679;
  wire _abc_40344_n3680;
  wire _abc_40344_n3681;
  wire _abc_40344_n3682_1;
  wire _abc_40344_n3683;
  wire _abc_40344_n3684;
  wire _abc_40344_n3686;
  wire _abc_40344_n3687;
  wire _abc_40344_n3688;
  wire _abc_40344_n3689;
  wire _abc_40344_n3690;
  wire _abc_40344_n3691;
  wire _abc_40344_n3692;
  wire _abc_40344_n3693;
  wire _abc_40344_n3694;
  wire _abc_40344_n3695;
  wire _abc_40344_n3696;
  wire _abc_40344_n3697;
  wire _abc_40344_n3698;
  wire _abc_40344_n3699;
  wire _abc_40344_n3700;
  wire _abc_40344_n3701;
  wire _abc_40344_n3703;
  wire _abc_40344_n3704;
  wire _abc_40344_n3705;
  wire _abc_40344_n3706_1;
  wire _abc_40344_n3707;
  wire _abc_40344_n3708;
  wire _abc_40344_n3709;
  wire _abc_40344_n3710;
  wire _abc_40344_n3711;
  wire _abc_40344_n3712;
  wire _abc_40344_n3713;
  wire _abc_40344_n3714;
  wire _abc_40344_n3715;
  wire _abc_40344_n3716;
  wire _abc_40344_n3717;
  wire _abc_40344_n3718;
  wire _abc_40344_n3719;
  wire _abc_40344_n3720;
  wire _abc_40344_n3721;
  wire _abc_40344_n3722;
  wire _abc_40344_n3724;
  wire _abc_40344_n3725;
  wire _abc_40344_n3725_bF_buf0;
  wire _abc_40344_n3725_bF_buf1;
  wire _abc_40344_n3725_bF_buf2;
  wire _abc_40344_n3725_bF_buf3;
  wire _abc_40344_n3726;
  wire _abc_40344_n3727_1;
  wire _abc_40344_n3728;
  wire _abc_40344_n3729;
  wire _abc_40344_n3730;
  wire _abc_40344_n3731;
  wire _abc_40344_n3732;
  wire _abc_40344_n3733;
  wire _abc_40344_n3734;
  wire _abc_40344_n3735;
  wire _abc_40344_n3736;
  wire _abc_40344_n3737;
  wire _abc_40344_n3739;
  wire _abc_40344_n3740;
  wire _abc_40344_n3741;
  wire _abc_40344_n3742;
  wire _abc_40344_n3743;
  wire _abc_40344_n3744;
  wire _abc_40344_n3745;
  wire _abc_40344_n3746;
  wire _abc_40344_n3747;
  wire _abc_40344_n3748;
  wire _abc_40344_n3749_1;
  wire _abc_40344_n3750;
  wire _abc_40344_n3751;
  wire _abc_40344_n3752;
  wire _abc_40344_n3753;
  wire _abc_40344_n3754;
  wire _abc_40344_n3756;
  wire _abc_40344_n3757;
  wire _abc_40344_n3758;
  wire _abc_40344_n3759;
  wire _abc_40344_n3760;
  wire _abc_40344_n3761;
  wire _abc_40344_n3762;
  wire _abc_40344_n3763;
  wire _abc_40344_n3764;
  wire _abc_40344_n3765;
  wire _abc_40344_n3766_1;
  wire _abc_40344_n3767;
  wire _abc_40344_n3768;
  wire _abc_40344_n3770_1;
  wire _abc_40344_n3771_1;
  wire _abc_40344_n3772_1;
  wire _abc_40344_n3773_1;
  wire _abc_40344_n3774_1;
  wire _abc_40344_n3775_1;
  wire _abc_40344_n3776_1;
  wire _abc_40344_n3777_1;
  wire _abc_40344_n3778_1;
  wire _abc_40344_n3779_1;
  wire _abc_40344_n3780_1;
  wire _abc_40344_n3781_1;
  wire _abc_40344_n3782_1;
  wire _abc_40344_n3784_1;
  wire _abc_40344_n3785_1;
  wire _abc_40344_n3786_1;
  wire _abc_40344_n3787_1;
  wire _abc_40344_n3788_1;
  wire _abc_40344_n3789_1;
  wire _abc_40344_n3790_1;
  wire _abc_40344_n3791_1;
  wire _abc_40344_n3792_1;
  wire _abc_40344_n3794_1;
  wire _abc_40344_n3795_1;
  wire _abc_40344_n3795_1_bF_buf0;
  wire _abc_40344_n3795_1_bF_buf1;
  wire _abc_40344_n3795_1_bF_buf2;
  wire _abc_40344_n3795_1_bF_buf3;
  wire _abc_40344_n3795_1_bF_buf4;
  wire _abc_40344_n3796_1;
  wire _abc_40344_n3798_1;
  wire _abc_40344_n3800;
  wire _abc_40344_n3802;
  wire _abc_40344_n3804;
  wire _abc_40344_n3806;
  wire _abc_40344_n3808;
  wire _abc_40344_n3810_1;
  wire _abc_40344_n3812;
  wire _abc_40344_n3814;
  wire _abc_40344_n3816;
  wire _abc_40344_n3818;
  wire _abc_40344_n3820;
  wire _abc_40344_n3822;
  wire _abc_40344_n3824_1;
  wire _abc_40344_n3826;
  wire _abc_40344_n3828;
  wire _abc_40344_n3830_1;
  wire _abc_40344_n3832;
  wire _abc_40344_n3834;
  wire _abc_40344_n3836_1;
  wire _abc_40344_n3838;
  wire _abc_40344_n3840;
  wire _abc_40344_n3842_1;
  wire _abc_40344_n3844;
  wire _abc_40344_n3846_1;
  wire _abc_40344_n3848;
  wire _abc_40344_n3850;
  wire _abc_40344_n3852_1;
  wire _abc_40344_n3854;
  wire _abc_40344_n3856;
  wire _abc_40344_n3857;
  wire _abc_40344_n3857_bF_buf0;
  wire _abc_40344_n3857_bF_buf1;
  wire _abc_40344_n3857_bF_buf2;
  wire _abc_40344_n3857_bF_buf3;
  wire _abc_40344_n3857_bF_buf4;
  wire _abc_40344_n3858_1;
  wire _abc_40344_n3860;
  wire _abc_40344_n3861_1;
  wire _abc_40344_n3861_1_bF_buf0;
  wire _abc_40344_n3861_1_bF_buf1;
  wire _abc_40344_n3861_1_bF_buf2;
  wire _abc_40344_n3861_1_bF_buf3;
  wire _abc_40344_n3862;
  wire _abc_40344_n3863;
  wire _abc_40344_n3864_1;
  wire _abc_40344_n3866;
  wire _abc_40344_n3867;
  wire _abc_40344_n3868_1;
  wire _abc_40344_n3869;
  wire _abc_40344_n3871_1;
  wire _abc_40344_n3872;
  wire _abc_40344_n3874_1;
  wire _abc_40344_n3875;
  wire _abc_40344_n3876;
  wire _abc_40344_n3877_1;
  wire _abc_40344_n3879;
  wire _abc_40344_n3880_1;
  wire _abc_40344_n3881;
  wire _abc_40344_n3882;
  wire _abc_40344_n3884;
  wire _abc_40344_n3885;
  wire _abc_40344_n3886_1;
  wire _abc_40344_n3887;
  wire _abc_40344_n3889;
  wire _abc_40344_n3890_1;
  wire _abc_40344_n3891;
  wire _abc_40344_n3892;
  wire _abc_40344_n3893_1;
  wire _abc_40344_n3895;
  wire _abc_40344_n3897_1;
  wire _abc_40344_n3898;
  wire _abc_40344_n3899;
  wire _abc_40344_n3900_1;
  wire _abc_40344_n3902;
  wire _abc_40344_n3903;
  wire _abc_40344_n3904;
  wire _abc_40344_n3906;
  wire _abc_40344_n3907;
  wire _abc_40344_n3908_1;
  wire _abc_40344_n3909;
  wire _abc_40344_n3910;
  wire _abc_40344_n3912;
  wire _abc_40344_n3913;
  wire _abc_40344_n3914;
  wire _abc_40344_n3916;
  wire _abc_40344_n3917;
  wire _abc_40344_n3918;
  wire _abc_40344_n3919;
  wire _abc_40344_n3921;
  wire _abc_40344_n3922;
  wire _abc_40344_n3923;
  wire _abc_40344_n3924;
  wire _abc_40344_n3926;
  wire _abc_40344_n3927;
  wire _abc_40344_n3928;
  wire _abc_40344_n3929;
  wire _abc_40344_n3931;
  wire _abc_40344_n3932;
  wire _abc_40344_n3933;
  wire _abc_40344_n3935;
  wire _abc_40344_n3936;
  wire _abc_40344_n3937;
  wire _abc_40344_n3938;
  wire _abc_40344_n3940;
  wire _abc_40344_n3941;
  wire _abc_40344_n3942;
  wire _abc_40344_n3943;
  wire _abc_40344_n3945;
  wire _abc_40344_n3946;
  wire _abc_40344_n3947;
  wire _abc_40344_n3949;
  wire _abc_40344_n3950;
  wire _abc_40344_n3951_1;
  wire _abc_40344_n3952;
  wire _abc_40344_n3954;
  wire _abc_40344_n3955;
  wire _abc_40344_n3956_1;
  wire _abc_40344_n3958_1;
  wire _abc_40344_n3959;
  wire _abc_40344_n3960;
  wire _abc_40344_n3961;
  wire _abc_40344_n3963;
  wire _abc_40344_n3964;
  wire _abc_40344_n3965;
  wire _abc_40344_n3967;
  wire _abc_40344_n3968;
  wire _abc_40344_n3969;
  wire _abc_40344_n3971;
  wire _abc_40344_n3972_1;
  wire _abc_40344_n3973;
  wire _abc_40344_n3975;
  wire _abc_40344_n3976;
  wire _abc_40344_n3977;
  wire _abc_40344_n3979_1;
  wire _abc_40344_n3980;
  wire _abc_40344_n3981;
  wire _abc_40344_n3983;
  wire _abc_40344_n3984;
  wire _abc_40344_n3985_1;
  wire _abc_40344_n3987;
  wire _abc_40344_n3988;
  wire _abc_40344_n3989;
  wire _abc_40344_n3991;
  wire _abc_40344_n3992_1;
  wire _abc_40344_n3993;
  wire _abc_40344_n3995;
  wire _abc_40344_n3997;
  wire _abc_40344_n3998;
  wire _abc_40344_n3999_1;
  wire _abc_40344_n4000;
  wire _abc_40344_n4001;
  wire _abc_40344_n4002;
  wire _abc_40344_n4003;
  wire _abc_40344_n4004;
  wire _abc_40344_n4005;
  wire _abc_40344_n4006_1;
  wire _abc_40344_n4007;
  wire _abc_40344_n4008;
  wire _abc_40344_n4009;
  wire _abc_40344_n4010;
  wire _abc_40344_n4011;
  wire _abc_40344_n4012;
  wire _abc_40344_n4013_1;
  wire _abc_40344_n4014;
  wire _abc_40344_n4015;
  wire _abc_40344_n4016;
  wire _abc_40344_n4017;
  wire _abc_40344_n4018;
  wire _abc_40344_n4019;
  wire _abc_40344_n4020_1;
  wire _abc_40344_n4021;
  wire _abc_40344_n4022;
  wire _abc_40344_n4023;
  wire _abc_40344_n4024;
  wire _abc_40344_n4025;
  wire _abc_40344_n4026_1;
  wire _abc_40344_n4027;
  wire _abc_40344_n4028;
  wire _abc_40344_n4029;
  wire _abc_40344_n4031;
  wire _abc_40344_n4032;
  wire _abc_40344_n4033_1;
  wire _abc_40344_n4035;
  wire _abc_40344_n4036;
  wire _abc_40344_n4038;
  wire _abc_40344_n4039;
  wire _abc_40344_n4040_1;
  wire _abc_40344_n4041;
  wire _abc_40344_n4042;
  wire _abc_40344_n4042_bF_buf0;
  wire _abc_40344_n4042_bF_buf1;
  wire _abc_40344_n4042_bF_buf2;
  wire _abc_40344_n4042_bF_buf3;
  wire _abc_40344_n4042_bF_buf4;
  wire _abc_40344_n4042_bF_buf5;
  wire _abc_40344_n4043;
  wire _abc_40344_n4044;
  wire _abc_40344_n4045;
  wire _abc_40344_n4046_1;
  wire _abc_40344_n4048;
  wire _abc_40344_n4049;
  wire _abc_40344_n4049_bF_buf0;
  wire _abc_40344_n4049_bF_buf1;
  wire _abc_40344_n4049_bF_buf2;
  wire _abc_40344_n4049_bF_buf3;
  wire _abc_40344_n4050;
  wire _abc_40344_n4051;
  wire _abc_40344_n4052_1;
  wire _abc_40344_n4053;
  wire _abc_40344_n4055;
  wire _abc_40344_n4056;
  wire _abc_40344_n4057;
  wire _abc_40344_n4058_1;
  wire _abc_40344_n4059;
  wire _abc_40344_n4061;
  wire _abc_40344_n4062;
  wire _abc_40344_n4063;
  wire _abc_40344_n4064_1;
  wire _abc_40344_n4066;
  wire _abc_40344_n4067;
  wire _abc_40344_n4068;
  wire _abc_40344_n4070_1;
  wire _abc_40344_n4071;
  wire _abc_40344_n4072;
  wire _abc_40344_n4074;
  wire _abc_40344_n4075;
  wire _abc_40344_n4076;
  wire _abc_40344_n4077_1;
  wire _abc_40344_n4078;
  wire _abc_40344_n4080;
  wire _abc_40344_n4081;
  wire _abc_40344_n4082;
  wire _abc_40344_n4083_1;
  wire _abc_40344_n4084;
  wire _abc_40344_n4086;
  wire _abc_40344_n4087;
  wire _abc_40344_n4088;
  wire _abc_40344_n4089_1;
  wire _abc_40344_n4090;
  wire _abc_40344_n4092;
  wire _abc_40344_n4093;
  wire _abc_40344_n4094;
  wire _abc_40344_n4095_1;
  wire _abc_40344_n4096;
  wire _abc_40344_n4098;
  wire _abc_40344_n4099;
  wire _abc_40344_n4100;
  wire _abc_40344_n4101_1;
  wire _abc_40344_n4102;
  wire _abc_40344_n4104;
  wire _abc_40344_n4105;
  wire _abc_40344_n4106;
  wire _abc_40344_n4107_1;
  wire _abc_40344_n4108;
  wire _abc_40344_n4110;
  wire _abc_40344_n4111;
  wire _abc_40344_n4112;
  wire _abc_40344_n4113_1;
  wire _abc_40344_n4114;
  wire _abc_40344_n4116;
  wire _abc_40344_n4117;
  wire _abc_40344_n4118;
  wire _abc_40344_n4119_1;
  wire _abc_40344_n4120;
  wire _abc_40344_n4121;
  wire _abc_40344_n4123;
  wire _abc_40344_n4124;
  wire _abc_40344_n4125_1;
  wire _abc_40344_n4126;
  wire _abc_40344_n4127;
  wire _abc_40344_n4128;
  wire _abc_40344_n4130;
  wire _abc_40344_n4131_1;
  wire _abc_40344_n4132;
  wire _abc_40344_n4133;
  wire _abc_40344_n4134;
  wire _abc_40344_n4135;
  wire _abc_40344_n4137_1;
  wire _abc_40344_n4138;
  wire _abc_40344_n4139;
  wire _abc_40344_n4140;
  wire _abc_40344_n4141;
  wire _abc_40344_n4142;
  wire _abc_40344_n4144;
  wire _abc_40344_n4145;
  wire _abc_40344_n4146;
  wire _abc_40344_n4147;
  wire _abc_40344_n4148;
  wire _abc_40344_n4149_1;
  wire _abc_40344_n4151;
  wire _abc_40344_n4152;
  wire _abc_40344_n4153;
  wire _abc_40344_n4154;
  wire _abc_40344_n4156;
  wire _abc_40344_n4157;
  wire _abc_40344_n4158_1;
  wire _abc_40344_n4159;
  wire _abc_40344_n4160;
  wire _abc_40344_n4161;
  wire _abc_40344_n4162;
  wire _abc_40344_n4164;
  wire _abc_40344_n4165;
  wire _abc_40344_n4166;
  wire _abc_40344_n4167_1;
  wire _abc_40344_n4168;
  wire _abc_40344_n4170;
  wire _abc_40344_n4171_1;
  wire _abc_40344_n4172;
  wire _abc_40344_n4173_1;
  wire _abc_40344_n4174;
  wire _abc_40344_n4176;
  wire _abc_40344_n4177_1;
  wire _abc_40344_n4178;
  wire _abc_40344_n4179_1;
  wire _abc_40344_n4180;
  wire _abc_40344_n4182;
  wire _abc_40344_n4183_1;
  wire _abc_40344_n4184;
  wire _abc_40344_n4185_1;
  wire _abc_40344_n4186;
  wire _abc_40344_n4187_1;
  wire _abc_40344_n4189_1;
  wire _abc_40344_n4190;
  wire _abc_40344_n4191_1;
  wire _abc_40344_n4192;
  wire _abc_40344_n4193_1;
  wire _abc_40344_n4195_1;
  wire _abc_40344_n4196;
  wire _abc_40344_n4197_1;
  wire _abc_40344_n4198;
  wire _abc_40344_n4199_1;
  wire _abc_40344_n4201_1;
  wire _abc_40344_n4202;
  wire _abc_40344_n4203_1;
  wire _abc_40344_n4204;
  wire _abc_40344_n4205_1;
  wire _abc_40344_n4207_1;
  wire _abc_40344_n4208;
  wire _abc_40344_n4209_1;
  wire _abc_40344_n4210;
  wire _abc_40344_n4211_1;
  wire _abc_40344_n4213_1;
  wire _abc_40344_n4214;
  wire _abc_40344_n4215_1;
  wire _abc_40344_n4216;
  wire _abc_40344_n4217_1;
  wire _abc_40344_n4219_1;
  wire _abc_40344_n4220;
  wire _abc_40344_n4221_1;
  wire _abc_40344_n4222;
  wire _abc_40344_n4223_1;
  wire _abc_40344_n4224;
  wire _abc_40344_n4225_1;
  wire _abc_40344_n4227_1;
  wire _abc_40344_n4228;
  wire _abc_40344_n4229_1;
  wire _abc_40344_n4230;
  wire _abc_40344_n4232;
  wire _abc_40344_n4233_1;
  wire _abc_40344_n4234;
  wire _abc_40344_n4235;
  wire _abc_40344_n4237;
  wire _abc_40344_n4237_bF_buf0;
  wire _abc_40344_n4237_bF_buf1;
  wire _abc_40344_n4237_bF_buf2;
  wire _abc_40344_n4237_bF_buf3;
  wire _abc_40344_n4237_bF_buf4;
  wire _abc_40344_n4237_bF_buf5;
  wire _abc_40344_n4237_bF_buf6;
  wire _abc_40344_n4238_1;
  wire _abc_40344_n4239_1;
  wire _abc_40344_n4241_1;
  wire _abc_40344_n4242_1;
  wire _abc_40344_n4244_1;
  wire _abc_40344_n4246;
  wire _abc_40344_n4247_1;
  wire _abc_40344_n4249;
  wire _abc_40344_n4250_1;
  wire _abc_40344_n4252;
  wire _abc_40344_n4254_1;
  wire _abc_40344_n4255;
  wire _abc_40344_n4257_1;
  wire _abc_40344_n4258;
  wire _abc_40344_n4260_1;
  wire _abc_40344_n4261;
  wire _abc_40344_n4263_1;
  wire _abc_40344_n4264;
  wire _abc_40344_n4266_1;
  wire _abc_40344_n4268_1;
  wire _abc_40344_n4269_1;
  wire _abc_40344_n4271_1;
  wire _abc_40344_n4272_1;
  wire _abc_40344_n4274_1;
  wire _abc_40344_n4275_1;
  wire _abc_40344_n4277_1;
  wire _abc_40344_n4278_1;
  wire _abc_40344_n4280_1;
  wire _abc_40344_n4281_1;
  wire _abc_40344_n4283_1;
  wire _abc_40344_n4284_1;
  wire _abc_40344_n4286_1;
  wire _abc_40344_n4288;
  wire _abc_40344_n4289_1;
  wire _abc_40344_n4291;
  wire _abc_40344_n4292_1;
  wire _abc_40344_n4294;
  wire _abc_40344_n4295_1;
  wire _abc_40344_n4297;
  wire _abc_40344_n4298_1;
  wire _abc_40344_n4300;
  wire _abc_40344_n4302_1;
  wire _abc_40344_n4303;
  wire _abc_40344_n4305_1;
  wire _abc_40344_n4306;
  wire _abc_40344_n4308_1;
  wire _abc_40344_n4309;
  wire _abc_40344_n4311_1;
  wire _abc_40344_n4312;
  wire _abc_40344_n4314_1;
  wire _abc_40344_n4315;
  wire _abc_40344_n4317_1;
  wire _abc_40344_n4318;
  wire _abc_40344_n4320_1;
  wire _abc_40344_n4321;
  wire _abc_40344_n4323_1;
  wire _abc_40344_n4324;
  wire _abc_40344_n4326_1;
  wire _abc_40344_n4327;
  wire _abc_40344_n4329_1;
  wire _abc_40344_n4329_1_bF_buf0;
  wire _abc_40344_n4329_1_bF_buf1;
  wire _abc_40344_n4329_1_bF_buf2;
  wire _abc_40344_n4329_1_bF_buf3;
  wire _abc_40344_n4329_1_bF_buf4;
  wire _abc_40344_n4330;
  wire _abc_40344_n4332;
  wire _abc_40344_n4334;
  wire _abc_40344_n4336;
  wire _abc_40344_n4338;
  wire _abc_40344_n4340;
  wire _abc_40344_n4342;
  wire _abc_40344_n4344;
  wire _abc_40344_n4346;
  wire _abc_40344_n4348;
  wire _abc_40344_n4350;
  wire _abc_40344_n4352;
  wire _abc_40344_n4354;
  wire _abc_40344_n4356;
  wire _abc_40344_n4358;
  wire _abc_40344_n4360;
  wire _abc_40344_n4362;
  wire _abc_40344_n4364;
  wire _abc_40344_n4366;
  wire _abc_40344_n4368;
  wire _abc_40344_n4370;
  wire _abc_40344_n4372;
  wire _abc_40344_n4374;
  wire _abc_40344_n4376;
  wire _abc_40344_n4378;
  wire _abc_40344_n4380;
  wire _abc_40344_n4382;
  wire _abc_40344_n4384;
  wire _abc_40344_n4386;
  wire _abc_40344_n4388;
  wire _abc_40344_n4390;
  wire _abc_40344_n4392;
  wire _abc_40344_n523;
  wire _abc_40344_n524;
  wire _abc_40344_n525;
  wire _abc_40344_n526;
  wire _abc_40344_n527;
  wire _abc_40344_n528;
  wire _abc_40344_n529;
  wire _abc_40344_n530;
  wire _abc_40344_n531;
  wire _abc_40344_n532;
  wire _abc_40344_n533;
  wire _abc_40344_n534;
  wire _abc_40344_n535;
  wire _abc_40344_n536;
  wire _abc_40344_n537_1;
  wire _abc_40344_n538_1;
  wire _abc_40344_n539;
  wire _abc_40344_n540;
  wire _abc_40344_n541_1;
  wire _abc_40344_n542_1;
  wire _abc_40344_n543;
  wire _abc_40344_n544;
  wire _abc_40344_n545_1;
  wire _abc_40344_n546_1;
  wire _abc_40344_n547;
  wire _abc_40344_n548;
  wire _abc_40344_n549_1;
  wire _abc_40344_n550_1;
  wire _abc_40344_n551;
  wire _abc_40344_n552;
  wire _abc_40344_n553_1;
  wire _abc_40344_n554_1;
  wire _abc_40344_n555;
  wire _abc_40344_n556;
  wire _abc_40344_n557_1;
  wire _abc_40344_n558;
  wire _abc_40344_n559_1;
  wire _abc_40344_n559_1_bF_buf0;
  wire _abc_40344_n559_1_bF_buf1;
  wire _abc_40344_n559_1_bF_buf2;
  wire _abc_40344_n559_1_bF_buf3;
  wire _abc_40344_n559_1_bF_buf4;
  wire _abc_40344_n559_1_bF_buf5;
  wire _abc_40344_n560;
  wire _abc_40344_n561_1;
  wire _abc_40344_n562;
  wire _abc_40344_n563_1;
  wire _abc_40344_n564;
  wire _abc_40344_n565_1;
  wire _abc_40344_n566;
  wire _abc_40344_n567_1;
  wire _abc_40344_n568;
  wire _abc_40344_n569_1;
  wire _abc_40344_n570;
  wire _abc_40344_n571_1;
  wire _abc_40344_n572;
  wire _abc_40344_n573_1;
  wire _abc_40344_n574;
  wire _abc_40344_n575_1;
  wire _abc_40344_n576;
  wire _abc_40344_n577_1;
  wire _abc_40344_n578_1;
  wire _abc_40344_n579;
  wire _abc_40344_n580;
  wire _abc_40344_n581;
  wire _abc_40344_n582;
  wire _abc_40344_n583;
  wire _abc_40344_n584_1;
  wire _abc_40344_n585;
  wire _abc_40344_n585_bF_buf0;
  wire _abc_40344_n585_bF_buf1;
  wire _abc_40344_n585_bF_buf2;
  wire _abc_40344_n585_bF_buf3;
  wire _abc_40344_n586;
  wire _abc_40344_n586_bF_buf0;
  wire _abc_40344_n586_bF_buf1;
  wire _abc_40344_n586_bF_buf2;
  wire _abc_40344_n586_bF_buf3;
  wire _abc_40344_n586_bF_buf4;
  wire _abc_40344_n587;
  wire _abc_40344_n588;
  wire _abc_40344_n589;
  wire _abc_40344_n589_bF_buf0;
  wire _abc_40344_n589_bF_buf1;
  wire _abc_40344_n589_bF_buf2;
  wire _abc_40344_n589_bF_buf3;
  wire _abc_40344_n589_bF_buf4;
  wire _abc_40344_n592;
  wire _abc_40344_n593_1;
  wire _abc_40344_n594;
  wire _abc_40344_n595_1;
  wire _abc_40344_n596_1;
  wire _abc_40344_n597;
  wire _abc_40344_n598;
  wire _abc_40344_n599;
  wire _abc_40344_n600_1;
  wire _abc_40344_n601;
  wire _abc_40344_n602;
  wire _abc_40344_n602_bF_buf0;
  wire _abc_40344_n602_bF_buf1;
  wire _abc_40344_n602_bF_buf2;
  wire _abc_40344_n602_bF_buf3;
  wire _abc_40344_n603;
  wire _abc_40344_n603_bF_buf0;
  wire _abc_40344_n603_bF_buf1;
  wire _abc_40344_n603_bF_buf2;
  wire _abc_40344_n603_bF_buf3;
  wire _abc_40344_n603_bF_buf4;
  wire _abc_40344_n604;
  wire _abc_40344_n605;
  wire _abc_40344_n606;
  wire _abc_40344_n607;
  wire _abc_40344_n608_1;
  wire _abc_40344_n609;
  wire _abc_40344_n610_1;
  wire _abc_40344_n610_1_bF_buf0;
  wire _abc_40344_n610_1_bF_buf1;
  wire _abc_40344_n610_1_bF_buf2;
  wire _abc_40344_n610_1_bF_buf3;
  wire _abc_40344_n611_1;
  wire _abc_40344_n611_1_bF_buf0;
  wire _abc_40344_n611_1_bF_buf1;
  wire _abc_40344_n611_1_bF_buf2;
  wire _abc_40344_n611_1_bF_buf3;
  wire _abc_40344_n612;
  wire _abc_40344_n613;
  wire _abc_40344_n614;
  wire _abc_40344_n615;
  wire _abc_40344_n616;
  wire _abc_40344_n617_1;
  wire _abc_40344_n618;
  wire _abc_40344_n619;
  wire _abc_40344_n620;
  wire _abc_40344_n621;
  wire _abc_40344_n622;
  wire _abc_40344_n623;
  wire _abc_40344_n624;
  wire _abc_40344_n625;
  wire _abc_40344_n626;
  wire _abc_40344_n627;
  wire _abc_40344_n628;
  wire _abc_40344_n629;
  wire _abc_40344_n630_1;
  wire _abc_40344_n630_1_bF_buf0;
  wire _abc_40344_n630_1_bF_buf1;
  wire _abc_40344_n630_1_bF_buf2;
  wire _abc_40344_n630_1_bF_buf3;
  wire _abc_40344_n630_1_bF_buf4;
  wire _abc_40344_n630_1_bF_buf5;
  wire _abc_40344_n630_1_bF_buf6;
  wire _abc_40344_n630_1_bF_buf7;
  wire _abc_40344_n630_1_bF_buf8;
  wire _abc_40344_n630_1_bF_buf9;
  wire _abc_40344_n631;
  wire _abc_40344_n633_1;
  wire _abc_40344_n634;
  wire _abc_40344_n635;
  wire _abc_40344_n636;
  wire _abc_40344_n637;
  wire _abc_40344_n638;
  wire _abc_40344_n639_1;
  wire _abc_40344_n640;
  wire _abc_40344_n641;
  wire _abc_40344_n642;
  wire _abc_40344_n643;
  wire _abc_40344_n644;
  wire _abc_40344_n645;
  wire _abc_40344_n646;
  wire _abc_40344_n647;
  wire _abc_40344_n648;
  wire _abc_40344_n649_1;
  wire _abc_40344_n650;
  wire _abc_40344_n650_bF_buf0;
  wire _abc_40344_n650_bF_buf1;
  wire _abc_40344_n650_bF_buf2;
  wire _abc_40344_n650_bF_buf3;
  wire _abc_40344_n651_1;
  wire _abc_40344_n652_1;
  wire _abc_40344_n653;
  wire _abc_40344_n654;
  wire _abc_40344_n655;
  wire _abc_40344_n656;
  wire _abc_40344_n657;
  wire _abc_40344_n658_1;
  wire _abc_40344_n659;
  wire _abc_40344_n660;
  wire _abc_40344_n661;
  wire _abc_40344_n662;
  wire _abc_40344_n663;
  wire _abc_40344_n664;
  wire _abc_40344_n665;
  wire _abc_40344_n666_1;
  wire _abc_40344_n667;
  wire _abc_40344_n668_1;
  wire _abc_40344_n669;
  wire _abc_40344_n670;
  wire _abc_40344_n671_1;
  wire _abc_40344_n672;
  wire _abc_40344_n673;
  wire _abc_40344_n673_bF_buf0;
  wire _abc_40344_n673_bF_buf1;
  wire _abc_40344_n673_bF_buf2;
  wire _abc_40344_n673_bF_buf3;
  wire _abc_40344_n674_1;
  wire _abc_40344_n675;
  wire _abc_40344_n676;
  wire _abc_40344_n677;
  wire _abc_40344_n678;
  wire _abc_40344_n679;
  wire _abc_40344_n680;
  wire _abc_40344_n681;
  wire _abc_40344_n682;
  wire _abc_40344_n683_1;
  wire _abc_40344_n684;
  wire _abc_40344_n685_1;
  wire _abc_40344_n686;
  wire _abc_40344_n687;
  wire _abc_40344_n688_1;
  wire _abc_40344_n689;
  wire _abc_40344_n690;
  wire _abc_40344_n691;
  wire _abc_40344_n692;
  wire _abc_40344_n693;
  wire _abc_40344_n694_1;
  wire _abc_40344_n695;
  wire _abc_40344_n695_bF_buf0;
  wire _abc_40344_n695_bF_buf1;
  wire _abc_40344_n695_bF_buf2;
  wire _abc_40344_n695_bF_buf3;
  wire _abc_40344_n696;
  wire _abc_40344_n697;
  wire _abc_40344_n698;
  wire _abc_40344_n699;
  wire _abc_40344_n700;
  wire _abc_40344_n700_bF_buf0;
  wire _abc_40344_n700_bF_buf1;
  wire _abc_40344_n700_bF_buf2;
  wire _abc_40344_n700_bF_buf3;
  wire _abc_40344_n700_bF_buf4;
  wire _abc_40344_n700_bF_buf5;
  wire _abc_40344_n701;
  wire _abc_40344_n702;
  wire _abc_40344_n703;
  wire _abc_40344_n704;
  wire _abc_40344_n705_1;
  wire _abc_40344_n705_1_bF_buf0;
  wire _abc_40344_n705_1_bF_buf1;
  wire _abc_40344_n705_1_bF_buf2;
  wire _abc_40344_n705_1_bF_buf3;
  wire _abc_40344_n705_1_bF_buf4;
  wire _abc_40344_n705_1_bF_buf5;
  wire _abc_40344_n705_1_bF_buf6;
  wire _abc_40344_n706;
  wire _abc_40344_n707_1;
  wire _abc_40344_n708;
  wire _abc_40344_n709;
  wire _abc_40344_n710_1;
  wire _abc_40344_n711;
  wire _abc_40344_n712;
  wire _abc_40344_n713_1;
  wire _abc_40344_n714;
  wire _abc_40344_n715;
  wire _abc_40344_n716;
  wire _abc_40344_n717;
  wire _abc_40344_n718;
  wire _abc_40344_n719;
  wire _abc_40344_n719_bF_buf0;
  wire _abc_40344_n719_bF_buf1;
  wire _abc_40344_n719_bF_buf2;
  wire _abc_40344_n719_bF_buf3;
  wire _abc_40344_n720;
  wire _abc_40344_n720_bF_buf0;
  wire _abc_40344_n720_bF_buf1;
  wire _abc_40344_n720_bF_buf2;
  wire _abc_40344_n720_bF_buf3;
  wire _abc_40344_n721;
  wire _abc_40344_n722;
  wire _abc_40344_n723;
  wire _abc_40344_n724;
  wire _abc_40344_n725;
  wire _abc_40344_n726;
  wire _abc_40344_n727_1;
  wire _abc_40344_n728;
  wire _abc_40344_n729_1;
  wire _abc_40344_n730;
  wire _abc_40344_n731;
  wire _abc_40344_n732_1;
  wire _abc_40344_n733;
  wire _abc_40344_n734;
  wire _abc_40344_n735;
  wire _abc_40344_n736;
  wire _abc_40344_n737;
  wire _abc_40344_n738_1;
  wire _abc_40344_n739;
  wire _abc_40344_n740;
  wire _abc_40344_n741;
  wire _abc_40344_n742;
  wire _abc_40344_n743;
  wire _abc_40344_n744;
  wire _abc_40344_n745;
  wire _abc_40344_n745_bF_buf0;
  wire _abc_40344_n745_bF_buf1;
  wire _abc_40344_n745_bF_buf2;
  wire _abc_40344_n745_bF_buf3;
  wire _abc_40344_n745_bF_buf4;
  wire _abc_40344_n746;
  wire _abc_40344_n747;
  wire _abc_40344_n748;
  wire _abc_40344_n749_1;
  wire _abc_40344_n750;
  wire _abc_40344_n751_1;
  wire _abc_40344_n752;
  wire _abc_40344_n753;
  wire _abc_40344_n754_1;
  wire _abc_40344_n755;
  wire _abc_40344_n756;
  wire _abc_40344_n757;
  wire _abc_40344_n758;
  wire _abc_40344_n759;
  wire _abc_40344_n760;
  wire _abc_40344_n761_1;
  wire _abc_40344_n761_1_bF_buf0;
  wire _abc_40344_n761_1_bF_buf1;
  wire _abc_40344_n761_1_bF_buf2;
  wire _abc_40344_n761_1_bF_buf3;
  wire _abc_40344_n761_1_bF_buf4;
  wire _abc_40344_n762;
  wire _abc_40344_n763;
  wire _abc_40344_n764;
  wire _abc_40344_n765;
  wire _abc_40344_n766;
  wire _abc_40344_n767;
  wire _abc_40344_n768;
  wire _abc_40344_n769;
  wire _abc_40344_n770;
  wire _abc_40344_n771;
  wire _abc_40344_n772;
  wire _abc_40344_n773;
  wire _abc_40344_n774;
  wire _abc_40344_n775_1;
  wire _abc_40344_n776;
  wire _abc_40344_n777_1;
  wire _abc_40344_n778;
  wire _abc_40344_n779;
  wire _abc_40344_n780_1;
  wire _abc_40344_n781;
  wire _abc_40344_n782;
  wire _abc_40344_n783;
  wire _abc_40344_n784;
  wire _abc_40344_n785;
  wire _abc_40344_n786;
  wire _abc_40344_n787_1;
  wire _abc_40344_n788;
  wire _abc_40344_n789;
  wire _abc_40344_n790;
  wire _abc_40344_n791;
  wire _abc_40344_n792;
  wire _abc_40344_n793;
  wire _abc_40344_n794;
  wire _abc_40344_n795;
  wire _abc_40344_n796;
  wire _abc_40344_n797;
  wire _abc_40344_n798;
  wire _abc_40344_n799;
  wire _abc_40344_n800_1;
  wire _abc_40344_n801_1;
  wire _abc_40344_n802;
  wire _abc_40344_n802_bF_buf0;
  wire _abc_40344_n802_bF_buf1;
  wire _abc_40344_n802_bF_buf2;
  wire _abc_40344_n802_bF_buf3;
  wire _abc_40344_n803;
  wire _abc_40344_n804;
  wire _abc_40344_n805;
  wire _abc_40344_n806;
  wire _abc_40344_n807_1;
  wire _abc_40344_n808;
  wire _abc_40344_n809;
  wire _abc_40344_n810;
  wire _abc_40344_n811;
  wire _abc_40344_n812;
  wire _abc_40344_n813;
  wire _abc_40344_n814;
  wire _abc_40344_n815;
  wire _abc_40344_n816;
  wire _abc_40344_n817;
  wire _abc_40344_n818_1;
  wire _abc_40344_n819;
  wire _abc_40344_n820;
  wire _abc_40344_n821;
  wire _abc_40344_n822;
  wire _abc_40344_n823;
  wire _abc_40344_n824_1;
  wire _abc_40344_n825;
  wire _abc_40344_n826_1;
  wire _abc_40344_n827;
  wire _abc_40344_n828;
  wire _abc_40344_n829_1;
  wire _abc_40344_n830;
  wire _abc_40344_n831;
  wire _abc_40344_n832;
  wire _abc_40344_n833;
  wire _abc_40344_n834;
  wire _abc_40344_n835_1;
  wire _abc_40344_n836;
  wire _abc_40344_n837;
  wire _abc_40344_n838;
  wire _abc_40344_n839;
  wire _abc_40344_n840;
  wire _abc_40344_n841;
  wire _abc_40344_n842;
  wire _abc_40344_n843;
  wire _abc_40344_n844;
  wire _abc_40344_n845;
  wire _abc_40344_n846;
  wire _abc_40344_n847;
  wire _abc_40344_n848;
  wire _abc_40344_n849_1;
  wire _abc_40344_n850_1;
  wire _abc_40344_n851;
  wire _abc_40344_n852;
  wire _abc_40344_n853;
  wire _abc_40344_n854_1;
  wire _abc_40344_n855;
  wire _abc_40344_n856;
  wire _abc_40344_n857;
  wire _abc_40344_n858;
  wire _abc_40344_n859;
  wire _abc_40344_n860;
  wire _abc_40344_n861;
  wire _abc_40344_n862;
  wire _abc_40344_n863;
  wire _abc_40344_n864;
  wire _abc_40344_n865;
  wire _abc_40344_n866_1;
  wire _abc_40344_n867;
  wire _abc_40344_n868;
  wire _abc_40344_n869;
  wire _abc_40344_n870;
  wire _abc_40344_n871;
  wire _abc_40344_n872;
  wire _abc_40344_n873;
  wire _abc_40344_n874;
  wire _abc_40344_n875;
  wire _abc_40344_n876;
  wire _abc_40344_n877_1;
  wire _abc_40344_n878;
  wire _abc_40344_n879;
  wire _abc_40344_n880;
  wire _abc_40344_n881;
  wire _abc_40344_n882;
  wire _abc_40344_n883;
  wire _abc_40344_n884;
  wire _abc_40344_n885;
  wire _abc_40344_n886;
  wire _abc_40344_n887;
  wire _abc_40344_n888;
  wire _abc_40344_n889;
  wire _abc_40344_n890;
  wire _abc_40344_n891;
  wire _abc_40344_n892;
  wire _abc_40344_n893;
  wire _abc_40344_n894;
  wire _abc_40344_n895;
  wire _abc_40344_n896;
  wire _abc_40344_n897;
  wire _abc_40344_n898;
  wire _abc_40344_n899;
  wire _abc_40344_n900;
  wire _abc_40344_n901;
  wire _abc_40344_n902_1;
  wire _abc_40344_n903_1;
  wire _abc_40344_n904;
  wire _abc_40344_n905;
  wire _abc_40344_n906_1;
  wire _abc_40344_n907;
  wire _abc_40344_n908;
  wire _abc_40344_n909;
  wire _abc_40344_n910;
  wire _abc_40344_n911;
  wire _abc_40344_n912;
  wire _abc_40344_n913;
  wire _abc_40344_n914;
  wire _abc_40344_n915_1;
  wire _abc_40344_n916;
  wire _abc_40344_n917;
  wire _abc_40344_n918;
  wire _abc_40344_n919;
  wire _abc_40344_n920;
  wire _abc_40344_n921;
  wire _abc_40344_n921_bF_buf0;
  wire _abc_40344_n921_bF_buf1;
  wire _abc_40344_n921_bF_buf2;
  wire _abc_40344_n921_bF_buf3;
  wire _abc_40344_n922_1;
  wire _abc_40344_n923_1;
  wire _abc_40344_n924;
  wire _abc_40344_n925;
  wire _abc_40344_n926;
  wire _abc_40344_n927_1;
  wire _abc_40344_n928;
  wire _abc_40344_n929;
  wire _abc_40344_n930;
  wire _abc_40344_n931;
  wire _abc_40344_n932;
  wire _abc_40344_n933;
  wire _abc_40344_n934;
  wire _abc_40344_n935_1;
  wire _abc_40344_n936;
  wire _abc_40344_n937;
  wire _abc_40344_n938;
  wire _abc_40344_n939;
  wire _abc_40344_n940;
  wire _abc_40344_n941;
  wire _abc_40344_n942;
  wire _abc_40344_n943_1;
  wire _abc_40344_n944;
  wire _abc_40344_n945_1;
  wire _abc_40344_n946;
  wire _abc_40344_n947;
  wire _abc_40344_n948_1;
  wire _abc_40344_n949;
  wire _abc_40344_n950;
  wire _abc_40344_n951;
  wire _abc_40344_n952;
  wire _abc_40344_n953;
  wire _abc_40344_n954;
  wire _abc_40344_n955_1;
  wire _abc_40344_n956;
  wire _abc_40344_n957;
  wire _abc_40344_n958;
  wire _abc_40344_n959;
  wire _abc_40344_n960;
  wire _abc_40344_n961;
  wire _abc_40344_n962;
  wire _abc_40344_n963;
  wire _abc_40344_n964;
  wire _abc_40344_n965;
  wire _abc_40344_n966;
  wire _abc_40344_n967;
  wire _abc_40344_n968;
  wire _abc_40344_n969;
  wire _abc_40344_n970_1;
  wire _abc_40344_n971;
  wire _abc_40344_n972_1;
  wire _abc_40344_n973;
  wire _abc_40344_n974;
  wire _abc_40344_n975_1;
  wire _abc_40344_n976;
  wire _abc_40344_n977;
  wire _abc_40344_n978;
  wire _abc_40344_n979;
  wire _abc_40344_n980;
  wire _abc_40344_n981_1;
  wire _abc_40344_n982;
  wire _abc_40344_n983;
  wire _abc_40344_n984;
  wire _abc_40344_n985;
  wire _abc_40344_n986;
  wire _abc_40344_n987;
  wire _abc_40344_n988;
  wire _abc_40344_n989;
  wire _abc_40344_n990;
  wire _abc_40344_n991;
  wire _abc_40344_n992;
  wire _abc_40344_n993;
  wire _abc_40344_n993_bF_buf0;
  wire _abc_40344_n993_bF_buf1;
  wire _abc_40344_n993_bF_buf2;
  wire _abc_40344_n993_bF_buf3;
  wire _abc_40344_n994;
  wire _abc_40344_n995;
  wire _abc_40344_n996;
  wire _abc_40344_n997;
  wire _abc_40344_n998;
  wire _abc_40344_n999;
  input clock;
  wire clock_bF_buf0;
  wire clock_bF_buf1;
  wire clock_bF_buf10;
  wire clock_bF_buf10_bF_buf0;
  wire clock_bF_buf10_bF_buf1;
  wire clock_bF_buf10_bF_buf2;
  wire clock_bF_buf10_bF_buf3;
  wire clock_bF_buf11;
  wire clock_bF_buf11_bF_buf0;
  wire clock_bF_buf11_bF_buf1;
  wire clock_bF_buf11_bF_buf2;
  wire clock_bF_buf11_bF_buf3;
  wire clock_bF_buf12;
  wire clock_bF_buf12_bF_buf0;
  wire clock_bF_buf12_bF_buf1;
  wire clock_bF_buf12_bF_buf2;
  wire clock_bF_buf12_bF_buf3;
  wire clock_bF_buf13;
  wire clock_bF_buf13_bF_buf0;
  wire clock_bF_buf13_bF_buf1;
  wire clock_bF_buf13_bF_buf2;
  wire clock_bF_buf13_bF_buf3;
  wire clock_bF_buf14;
  wire clock_bF_buf14_bF_buf0;
  wire clock_bF_buf14_bF_buf1;
  wire clock_bF_buf14_bF_buf2;
  wire clock_bF_buf14_bF_buf3;
  wire clock_bF_buf2;
  wire clock_bF_buf3;
  wire clock_bF_buf4;
  wire clock_bF_buf5;
  wire clock_bF_buf6;
  wire clock_bF_buf7;
  wire clock_bF_buf8;
  wire clock_bF_buf9;
  wire n1002;
  wire n1006;
  wire n1010;
  wire n1014;
  wire n1018;
  wire n1022;
  wire n1026;
  wire n1030;
  wire n1034;
  wire n1038;
  wire n1042;
  wire n1046;
  wire n1050;
  wire n1054;
  wire n1058;
  wire n1062;
  wire n1066;
  wire n1070;
  wire n1074;
  wire n1078;
  wire n1082;
  wire n1086;
  wire n1090;
  wire n1094;
  wire n1098;
  wire n1102;
  wire n1106;
  wire n1110;
  wire n1114;
  wire n1118;
  wire n1122;
  wire n1126;
  wire n1130;
  wire n1134;
  wire n1138;
  wire n1142;
  wire n1146;
  wire n1150;
  wire n1154;
  wire n1158;
  wire n1162;
  wire n1166;
  wire n1170;
  wire n1174;
  wire n1178;
  wire n1182;
  wire n1186;
  wire n1191;
  wire n1196;
  wire n1201;
  wire n1206;
  wire n1211;
  wire n1216;
  wire n1221;
  wire n1226;
  wire n1231;
  wire n1236;
  wire n1241;
  wire n1246;
  wire n1251;
  wire n1256;
  wire n1261;
  wire n1266;
  wire n1271;
  wire n1276;
  wire n1281;
  wire n1286;
  wire n1291;
  wire n1296;
  wire n1301;
  wire n1306;
  wire n1311;
  wire n1316;
  wire n1321;
  wire n1326;
  wire n1331;
  wire n1336;
  wire n1336_bF_buf0;
  wire n1336_bF_buf1;
  wire n1336_bF_buf2;
  wire n1336_bF_buf3;
  wire n1336_bF_buf4;
  wire n1341;
  wire n1345;
  wire n178;
  wire n183;
  wire n188;
  wire n193;
  wire n198;
  wire n203;
  wire n208;
  wire n213;
  wire n218;
  wire n223;
  wire n228;
  wire n233;
  wire n238;
  wire n243;
  wire n248;
  wire n253;
  wire n258;
  wire n263;
  wire n268;
  wire n273;
  wire n278;
  wire n283;
  wire n288;
  wire n293;
  wire n298;
  wire n303;
  wire n308;
  wire n313;
  wire n318;
  wire n323;
  wire n328;
  wire n333;
  wire n338;
  wire n343;
  wire n348;
  wire n353;
  wire n358;
  wire n363;
  wire n368;
  wire n373;
  wire n378;
  wire n383;
  wire n388;
  wire n393;
  wire n398;
  wire n403;
  wire n408;
  wire n413;
  wire n418;
  wire n423;
  wire n428;
  wire n433;
  wire n438;
  wire n443;
  wire n448;
  wire n453;
  wire n458;
  wire n463;
  wire n468;
  wire n473;
  wire n478;
  wire n483;
  wire n488;
  wire n493;
  wire n498;
  wire n503;
  wire n508;
  wire n513;
  wire n518;
  wire n523;
  wire n528;
  wire n533;
  wire n538;
  wire n543;
  wire n548;
  wire n553;
  wire n558;
  wire n563;
  wire n568;
  wire n573;
  wire n578;
  wire n583;
  wire n588;
  wire n593;
  wire n598;
  wire n603;
  wire n608;
  wire n613;
  wire n618;
  wire n623;
  wire n628;
  wire n633;
  wire n638;
  wire n643;
  wire n648;
  wire n653;
  wire n658;
  wire n663;
  wire n668;
  wire n673;
  wire n678;
  wire n683;
  wire n688;
  wire n693;
  wire n698;
  wire n703;
  wire n708;
  wire n713;
  wire n718;
  wire n723;
  wire n728;
  wire n733;
  wire n738;
  wire n743;
  wire n748;
  wire n753;
  wire n758;
  wire n763;
  wire n768;
  wire n773;
  wire n778;
  wire n783;
  wire n788;
  wire n793;
  wire n798;
  wire n803;
  wire n808;
  wire n813;
  wire n818;
  wire n823;
  wire n828;
  wire n833;
  wire n838;
  wire n843;
  wire n848;
  wire n853;
  wire n858;
  wire n863;
  wire n868;
  wire n873;
  wire n878;
  wire n883;
  wire n888;
  wire n893;
  wire n898;
  wire n903;
  wire n908;
  wire n913;
  wire n918;
  wire n923;
  wire n928;
  wire n933;
  wire n938;
  wire n943;
  wire n948;
  wire n953;
  wire n958;
  wire n963;
  wire n968;
  wire n973;
  wire n978;
  wire n982;
  wire n986;
  wire n990;
  wire n994;
  wire n998;
  input nRESET_G;
  wire nRESET_G_bF_buf0;
  wire nRESET_G_bF_buf1;
  wire nRESET_G_bF_buf2;
  wire nRESET_G_bF_buf3;
  wire nRESET_G_bF_buf4;
  wire nRESET_G_bF_buf5;
  wire nRESET_G_bF_buf6;
  wire nRESET_G_bF_buf7;
  wire nRESET_G_bF_buf8;
  AND2X2 AND2X2_1 ( .A(_abc_40344_n558), .B(_abc_40344_n560), .Y(_abc_40344_n561_1) );
  AND2X2 AND2X2_10 ( .A(_abc_40344_n1159), .B(_abc_40344_n1157), .Y(_abc_40344_n1160) );
  AND2X2 AND2X2_100 ( .A(_abc_40344_n4077_1), .B(nRESET_G), .Y(_abc_40344_n4078) );
  AND2X2 AND2X2_101 ( .A(_abc_40344_n4083_1), .B(nRESET_G), .Y(_abc_40344_n4084) );
  AND2X2 AND2X2_102 ( .A(_abc_40344_n4089_1), .B(nRESET_G), .Y(_abc_40344_n4090) );
  AND2X2 AND2X2_103 ( .A(_abc_40344_n4095_1), .B(nRESET_G), .Y(_abc_40344_n4096) );
  AND2X2 AND2X2_104 ( .A(_abc_40344_n4107_1), .B(nRESET_G), .Y(_abc_40344_n4108) );
  AND2X2 AND2X2_105 ( .A(_abc_40344_n4113_1), .B(nRESET_G), .Y(_abc_40344_n4114) );
  AND2X2 AND2X2_106 ( .A(_abc_40344_n3564), .B(_abc_40344_n4048), .Y(_abc_40344_n4116) );
  AND2X2 AND2X2_107 ( .A(_abc_40344_n4120), .B(nRESET_G), .Y(_abc_40344_n4121) );
  AND2X2 AND2X2_108 ( .A(_abc_40344_n3385), .B(_abc_40344_n4178), .Y(_abc_40344_n4179_1) );
  AND2X2 AND2X2_109 ( .A(_abc_40344_n3296), .B(_abc_40344_n4048), .Y(_abc_40344_n4189_1) );
  AND2X2 AND2X2_11 ( .A(_abc_40344_n1192), .B(_abc_40344_n1145), .Y(_abc_40344_n1193_1) );
  AND2X2 AND2X2_110 ( .A(_abc_40344_n4241_1), .B(nRESET_G), .Y(_abc_40344_n4242_1) );
  AND2X2 AND2X2_111 ( .A(_abc_40344_n4246), .B(nRESET_G), .Y(_abc_40344_n4247_1) );
  AND2X2 AND2X2_112 ( .A(_abc_40344_n4249), .B(nRESET_G), .Y(_abc_40344_n4250_1) );
  AND2X2 AND2X2_113 ( .A(_abc_40344_n4254_1), .B(nRESET_G), .Y(_abc_40344_n4255) );
  AND2X2 AND2X2_114 ( .A(_abc_40344_n4257_1), .B(nRESET_G), .Y(_abc_40344_n4258) );
  AND2X2 AND2X2_115 ( .A(_abc_40344_n4260_1), .B(nRESET_G), .Y(_abc_40344_n4261) );
  AND2X2 AND2X2_116 ( .A(_abc_40344_n4263_1), .B(nRESET_G), .Y(_abc_40344_n4264) );
  AND2X2 AND2X2_117 ( .A(_abc_40344_n4268_1), .B(nRESET_G), .Y(_abc_40344_n4269_1) );
  AND2X2 AND2X2_118 ( .A(_abc_40344_n4271_1), .B(nRESET_G), .Y(_abc_40344_n4272_1) );
  AND2X2 AND2X2_119 ( .A(_abc_40344_n4274_1), .B(nRESET_G), .Y(_abc_40344_n4275_1) );
  AND2X2 AND2X2_12 ( .A(_abc_40344_n1156), .B(_abc_40344_n1226), .Y(_abc_40344_n1227) );
  AND2X2 AND2X2_120 ( .A(_abc_40344_n4277_1), .B(nRESET_G), .Y(_abc_40344_n4278_1) );
  AND2X2 AND2X2_121 ( .A(_abc_40344_n4280_1), .B(nRESET_G), .Y(_abc_40344_n4281_1) );
  AND2X2 AND2X2_122 ( .A(_abc_40344_n4283_1), .B(nRESET_G), .Y(_abc_40344_n4284_1) );
  AND2X2 AND2X2_123 ( .A(_abc_40344_n4288), .B(nRESET_G), .Y(_abc_40344_n4289_1) );
  AND2X2 AND2X2_124 ( .A(_abc_40344_n4291), .B(nRESET_G), .Y(_abc_40344_n4292_1) );
  AND2X2 AND2X2_125 ( .A(_abc_40344_n4323_1), .B(nRESET_G), .Y(_abc_40344_n4324) );
  AND2X2 AND2X2_13 ( .A(_abc_40344_n1300), .B(_abc_40344_n1055), .Y(_abc_40344_n1301) );
  AND2X2 AND2X2_14 ( .A(_abc_40344_n1314), .B(_abc_40344_n1313), .Y(_abc_40344_n1315) );
  AND2X2 AND2X2_15 ( .A(_abc_40344_n1342), .B(_abc_40344_n1343_1), .Y(_abc_40344_n1344) );
  AND2X2 AND2X2_16 ( .A(_abc_40344_n1357), .B(_abc_40344_n1355), .Y(_abc_40344_n1358) );
  AND2X2 AND2X2_17 ( .A(_abc_40344_n1060), .B(_abc_40344_n1406), .Y(_abc_40344_n1407) );
  AND2X2 AND2X2_18 ( .A(_abc_40344_n1103_1), .B(_abc_40344_n1435), .Y(_abc_40344_n1436) );
  AND2X2 AND2X2_19 ( .A(_abc_40344_n1453), .B(_abc_40344_n1454), .Y(_abc_40344_n1455) );
  AND2X2 AND2X2_2 ( .A(_abc_40344_n674_1), .B(_abc_40344_n675), .Y(_abc_40344_n781) );
  AND2X2 AND2X2_20 ( .A(_abc_40344_n1480), .B(_abc_40344_n1478), .Y(_abc_40344_n1481) );
  AND2X2 AND2X2_21 ( .A(_abc_40344_n1067), .B(_abc_40344_n1538), .Y(_abc_40344_n1539) );
  AND2X2 AND2X2_22 ( .A(_abc_40344_n1541), .B(_abc_40344_n685_1), .Y(_abc_40344_n1542) );
  AND2X2 AND2X2_23 ( .A(_abc_40344_n1098), .B(_abc_40344_n1096), .Y(_abc_40344_n1573) );
  AND2X2 AND2X2_24 ( .A(_abc_40344_n1572), .B(_abc_40344_n1573), .Y(_abc_40344_n1574) );
  AND2X2 AND2X2_25 ( .A(_abc_40344_n1583), .B(_abc_40344_n1579), .Y(_abc_40344_n1584) );
  AND2X2 AND2X2_26 ( .A(_abc_40344_n894), .B(_abc_40344_n874), .Y(_abc_40344_n1600) );
  AND2X2 AND2X2_27 ( .A(_abc_40344_n1613), .B(_abc_40344_n1606), .Y(_abc_40344_n1614) );
  AND2X2 AND2X2_28 ( .A(_abc_40344_n1452), .B(_abc_40344_n1618), .Y(_abc_40344_n1619) );
  AND2X2 AND2X2_29 ( .A(_abc_40344_n1617), .B(_abc_40344_n1619), .Y(_abc_40344_n1620) );
  AND2X2 AND2X2_3 ( .A(_abc_40344_n851), .B(_abc_40344_n852), .Y(_abc_40344_n853) );
  AND2X2 AND2X2_30 ( .A(_abc_40344_n1634), .B(_abc_40344_n1079), .Y(_abc_40344_n1638) );
  AND2X2 AND2X2_31 ( .A(_abc_40344_n874), .B(_abc_40344_n876), .Y(_abc_40344_n1672) );
  AND2X2 AND2X2_32 ( .A(_abc_40344_n1672), .B(_abc_40344_n1671), .Y(_abc_40344_n1673) );
  AND2X2 AND2X2_33 ( .A(_abc_40344_n1338), .B(_abc_40344_n1336), .Y(_abc_40344_n1702) );
  AND2X2 AND2X2_34 ( .A(_abc_40344_n1706), .B(_abc_40344_n1701), .Y(_abc_40344_n1707) );
  AND2X2 AND2X2_35 ( .A(_abc_40344_n1725), .B(_abc_40344_n1729), .Y(_abc_40344_n1730) );
  AND2X2 AND2X2_36 ( .A(_abc_40344_n1525), .B(_abc_40344_n1733), .Y(_abc_40344_n1734) );
  AND2X2 AND2X2_37 ( .A(_abc_40344_n1389), .B(_abc_40344_n1386), .Y(_abc_40344_n1782) );
  AND2X2 AND2X2_38 ( .A(_abc_40344_n1685), .B(_abc_40344_n1808), .Y(_abc_40344_n1809) );
  AND2X2 AND2X2_39 ( .A(_abc_40344_n1706), .B(_abc_40344_n1314), .Y(_abc_40344_n1827) );
  AND2X2 AND2X2_4 ( .A(_abc_40344_n880), .B(_abc_40344_n888), .Y(_abc_40344_n889) );
  AND2X2 AND2X2_40 ( .A(_abc_40344_n1908), .B(_abc_40344_n1907), .Y(_abc_40344_n1909) );
  AND2X2 AND2X2_41 ( .A(_abc_40344_n695), .B(REG2_REG_31_), .Y(_abc_40344_n1910) );
  AND2X2 AND2X2_42 ( .A(_abc_40344_n695), .B(REG2_REG_30_), .Y(_abc_40344_n1918) );
  AND2X2 AND2X2_43 ( .A(_abc_40344_n1960), .B(_abc_40344_n1964), .Y(_abc_40344_n1965) );
  AND2X2 AND2X2_44 ( .A(_abc_40344_n1945), .B(_abc_40344_n1942), .Y(_abc_40344_n2031) );
  AND2X2 AND2X2_45 ( .A(_abc_40344_n2145), .B(_abc_40344_n2147), .Y(_abc_40344_n2148) );
  AND2X2 AND2X2_46 ( .A(_abc_40344_n585), .B(_abc_40344_n2161), .Y(_abc_40344_n2165) );
  AND2X2 AND2X2_47 ( .A(_abc_40344_n2166), .B(_abc_40344_n2164), .Y(_abc_40344_n2198) );
  AND2X2 AND2X2_48 ( .A(_abc_40344_n2218), .B(_abc_40344_n2217), .Y(_abc_40344_n2219) );
  AND2X2 AND2X2_49 ( .A(_abc_40344_n2212), .B(_abc_40344_n2213), .Y(_abc_40344_n2227) );
  AND2X2 AND2X2_5 ( .A(_abc_40344_n909), .B(_abc_40344_n911), .Y(_abc_40344_n912) );
  AND2X2 AND2X2_50 ( .A(_abc_40344_n2251), .B(_abc_40344_n2252), .Y(_abc_40344_n2271) );
  AND2X2 AND2X2_51 ( .A(_abc_40344_n2280), .B(_abc_40344_n2284), .Y(_abc_40344_n2285) );
  AND2X2 AND2X2_52 ( .A(_abc_40344_n2280), .B(_abc_40344_n2288_1), .Y(_abc_40344_n2289) );
  AND2X2 AND2X2_53 ( .A(_abc_40344_n2332), .B(_abc_40344_n2333), .Y(_abc_40344_n2334) );
  AND2X2 AND2X2_54 ( .A(_abc_40344_n2185), .B(_abc_40344_n2256), .Y(_abc_40344_n2423) );
  AND2X2 AND2X2_55 ( .A(_abc_40344_n2188), .B(_abc_40344_n2257), .Y(_abc_40344_n2424) );
  AND2X2 AND2X2_56 ( .A(_abc_40344_n2170), .B(_abc_40344_n2171), .Y(_abc_40344_n2426) );
  AND2X2 AND2X2_57 ( .A(_abc_40344_n2271), .B(_abc_40344_n2269), .Y(_abc_40344_n2446) );
  AND2X2 AND2X2_58 ( .A(_abc_40344_n2489), .B(_abc_40344_n2495), .Y(_abc_40344_n2496_1) );
  AND2X2 AND2X2_59 ( .A(_abc_40344_n2574), .B(_abc_40344_n2511), .Y(_abc_40344_n2578) );
  AND2X2 AND2X2_6 ( .A(_abc_40344_n960), .B(_abc_40344_n961), .Y(_abc_40344_n962) );
  AND2X2 AND2X2_60 ( .A(_abc_40344_n2578), .B(_abc_40344_n2583), .Y(_abc_40344_n2584) );
  AND2X2 AND2X2_61 ( .A(_abc_40344_n2584), .B(_abc_40344_n2585), .Y(_abc_40344_n2586) );
  AND2X2 AND2X2_62 ( .A(_abc_40344_n2698_1), .B(_abc_40344_n853), .Y(_abc_40344_n2700) );
  AND2X2 AND2X2_63 ( .A(_abc_40344_n1800), .B(_abc_40344_n2708), .Y(_abc_40344_n2709) );
  AND2X2 AND2X2_64 ( .A(_abc_40344_n2767), .B(_abc_40344_n2752), .Y(_abc_40344_n2768_1) );
  AND2X2 AND2X2_65 ( .A(_abc_40344_n2925), .B(_abc_40344_n2906), .Y(_abc_40344_n2926) );
  AND2X2 AND2X2_66 ( .A(_abc_40344_n2941), .B(_abc_40344_n2939), .Y(_abc_40344_n2942) );
  AND2X2 AND2X2_67 ( .A(_abc_40344_n2953), .B(_abc_40344_n1197), .Y(_abc_40344_n2954) );
  AND2X2 AND2X2_68 ( .A(_abc_40344_n3143), .B(_abc_40344_n3138), .Y(_abc_40344_n3144) );
  AND2X2 AND2X2_69 ( .A(_abc_40344_n3145), .B(_abc_40344_n3146), .Y(_abc_40344_n3147_1) );
  AND2X2 AND2X2_7 ( .A(_abc_40344_n969), .B(_abc_40344_n970_1), .Y(_abc_40344_n971) );
  AND2X2 AND2X2_70 ( .A(_abc_40344_n3148), .B(_abc_40344_n3139), .Y(_abc_40344_n3149) );
  AND2X2 AND2X2_71 ( .A(_abc_40344_n3208), .B(_abc_40344_n3199), .Y(_abc_40344_n3209) );
  AND2X2 AND2X2_72 ( .A(_abc_40344_n3238), .B(_abc_40344_n3097), .Y(_abc_40344_n3239) );
  AND2X2 AND2X2_73 ( .A(_abc_40344_n3273), .B(_abc_40344_n3237), .Y(_abc_40344_n3274) );
  AND2X2 AND2X2_74 ( .A(_abc_40344_n2030), .B(_abc_40344_n3329), .Y(_abc_40344_n3330) );
  AND2X2 AND2X2_75 ( .A(_abc_40344_n3328), .B(_abc_40344_n3335_1), .Y(_abc_40344_n3336) );
  AND2X2 AND2X2_76 ( .A(_abc_40344_n3336), .B(_abc_40344_n2521), .Y(_abc_40344_n3337) );
  AND2X2 AND2X2_77 ( .A(_abc_40344_n3387), .B(_abc_40344_n3091), .Y(_abc_40344_n3388_1) );
  AND2X2 AND2X2_78 ( .A(_abc_40344_n3440), .B(_abc_40344_n3438), .Y(_abc_40344_n3441) );
  AND2X2 AND2X2_79 ( .A(_abc_40344_n3467), .B(_abc_40344_n3423), .Y(_abc_40344_n3468) );
  AND2X2 AND2X2_8 ( .A(_abc_40344_n1014), .B(_abc_40344_n1013), .Y(_abc_40344_n1015) );
  AND2X2 AND2X2_80 ( .A(_abc_40344_n3480), .B(_abc_40344_n3223), .Y(_abc_40344_n3481) );
  AND2X2 AND2X2_81 ( .A(_abc_40344_n3319), .B(_abc_40344_n3306), .Y(_abc_40344_n3482) );
  AND2X2 AND2X2_82 ( .A(_abc_40344_n3529), .B(_abc_40344_n3525), .Y(_abc_40344_n3530) );
  AND2X2 AND2X2_83 ( .A(_abc_40344_n3546), .B(_abc_40344_n3082), .Y(_abc_40344_n3547) );
  AND2X2 AND2X2_84 ( .A(_abc_40344_n3552), .B(_abc_40344_n3550), .Y(_abc_40344_n3553) );
  AND2X2 AND2X2_85 ( .A(_abc_40344_n3320), .B(_abc_40344_n2545), .Y(_abc_40344_n3559) );
  AND2X2 AND2X2_86 ( .A(_abc_40344_n3526), .B(_abc_40344_n3604_1), .Y(_abc_40344_n3605) );
  AND2X2 AND2X2_87 ( .A(_abc_40344_n3574), .B(_abc_40344_n3624), .Y(_abc_40344_n3625) );
  AND2X2 AND2X2_88 ( .A(_abc_40344_n3078), .B(_abc_40344_n3635), .Y(_abc_40344_n3636) );
  AND2X2 AND2X2_89 ( .A(_abc_40344_n3646), .B(_abc_40344_n3644), .Y(_abc_40344_n3647) );
  AND2X2 AND2X2_9 ( .A(_abc_40344_n1125), .B(_abc_40344_n1126), .Y(_abc_40344_n1127) );
  AND2X2 AND2X2_90 ( .A(_abc_40344_n3623), .B(_abc_40344_n3664), .Y(_abc_40344_n3665) );
  AND2X2 AND2X2_91 ( .A(_abc_40344_n3076), .B(_abc_40344_n3670), .Y(_abc_40344_n3671) );
  AND2X2 AND2X2_92 ( .A(_abc_40344_n3691), .B(_abc_40344_n2482), .Y(_abc_40344_n3709) );
  AND2X2 AND2X2_93 ( .A(_abc_40344_n3074), .B(_abc_40344_n3717), .Y(_abc_40344_n3718) );
  AND2X2 AND2X2_94 ( .A(_abc_40344_n3756), .B(_abc_40344_n2546), .Y(_abc_40344_n3757) );
  AND2X2 AND2X2_95 ( .A(_abc_40344_n2558), .B(_abc_40344_n2555), .Y(_abc_40344_n4013_1) );
  AND2X2 AND2X2_96 ( .A(_abc_40344_n3777_1), .B(_abc_40344_n3775_1), .Y(_abc_40344_n4050) );
  AND2X2 AND2X2_97 ( .A(_abc_40344_n4052_1), .B(nRESET_G), .Y(_abc_40344_n4053) );
  AND2X2 AND2X2_98 ( .A(_abc_40344_n3749_1), .B(_abc_40344_n3739), .Y(_abc_40344_n4061) );
  AND2X2 AND2X2_99 ( .A(_abc_40344_n4063), .B(nRESET_G), .Y(_abc_40344_n4064_1) );
  AOI21X1 AOI21X1_1 ( .A(_abc_40344_n621), .B(_abc_40344_n546_1), .C(_abc_40344_n613), .Y(_abc_40344_n638) );
  AOI21X1 AOI21X1_10 ( .A(_abc_40344_n682), .B(_abc_40344_n676), .C(_abc_40344_n559_1), .Y(_abc_40344_n753) );
  AOI21X1 AOI21X1_100 ( .A(_abc_40344_n1894), .B(_abc_40344_n1895), .C(_abc_40344_n1590), .Y(_abc_40344_n1896) );
  AOI21X1 AOI21X1_101 ( .A(_abc_40344_n1032), .B(_abc_40344_n1201), .C(_abc_40344_n1899), .Y(_abc_40344_n1900) );
  AOI21X1 AOI21X1_102 ( .A(_abc_40344_n1005), .B(_abc_40344_n1898), .C(_abc_40344_n1901), .Y(_abc_40344_n1902) );
  AOI21X1 AOI21X1_103 ( .A(_abc_40344_n1040), .B(_abc_40344_n1073), .C(_abc_40344_n1928), .Y(_abc_40344_n1929) );
  AOI21X1 AOI21X1_104 ( .A(_abc_40344_n1961), .B(_abc_40344_n1234), .C(_abc_40344_n1963), .Y(_abc_40344_n1964) );
  AOI21X1 AOI21X1_105 ( .A(_abc_40344_n1477), .B(_abc_40344_n1488), .C(_abc_40344_n2002), .Y(_abc_40344_n2003) );
  AOI21X1 AOI21X1_106 ( .A(_abc_40344_n2027), .B(_abc_40344_n1548), .C(_abc_40344_n1649), .Y(_abc_40344_n2028) );
  AOI21X1 AOI21X1_107 ( .A(_abc_40344_n1110), .B(_abc_40344_n1100), .C(_abc_40344_n2029), .Y(_abc_40344_n2030) );
  AOI21X1 AOI21X1_108 ( .A(_abc_40344_n2030), .B(_abc_40344_n2031), .C(_abc_40344_n2028), .Y(_abc_40344_n2032) );
  AOI21X1 AOI21X1_109 ( .A(_abc_40344_n2075), .B(_abc_40344_n2079), .C(_abc_40344_n2011), .Y(_abc_40344_n2080) );
  AOI21X1 AOI21X1_11 ( .A(_abc_40344_n765), .B(_abc_40344_n766), .C(_abc_40344_n743), .Y(_abc_40344_n767) );
  AOI21X1 AOI21X1_110 ( .A(_abc_40344_n1645), .B(_abc_40344_n1926), .C(_abc_40344_n2103), .Y(_abc_40344_n2104) );
  AOI21X1 AOI21X1_111 ( .A(_abc_40344_n1550), .B(_abc_40344_n2104), .C(_abc_40344_n2101), .Y(_abc_40344_n2105) );
  AOI21X1 AOI21X1_112 ( .A(_abc_40344_n2113), .B(_abc_40344_n2034), .C(_abc_40344_n2109), .Y(_abc_40344_n2114) );
  AOI21X1 AOI21X1_113 ( .A(_abc_40344_n2060), .B(_abc_40344_n1998), .C(_abc_40344_n2144), .Y(_abc_40344_n2145) );
  AOI21X1 AOI21X1_114 ( .A(_abc_40344_n2176), .B(_abc_40344_n2175), .C(_abc_40344_n2161), .Y(_abc_40344_n2199) );
  AOI21X1 AOI21X1_115 ( .A(_abc_40344_n2169), .B(_abc_40344_n775_1), .C(_abc_40344_n2179), .Y(_abc_40344_n2208) );
  AOI21X1 AOI21X1_116 ( .A(_abc_40344_n825), .B(_abc_40344_n2162), .C(_abc_40344_n2214), .Y(_abc_40344_n2215) );
  AOI21X1 AOI21X1_117 ( .A(_abc_40344_n2162), .B(_abc_40344_n908), .C(_abc_40344_n2234), .Y(_abc_40344_n2235) );
  AOI21X1 AOI21X1_118 ( .A(_abc_40344_n1327), .B(_abc_40344_n2162), .C(_abc_40344_n2240), .Y(_abc_40344_n2241) );
  AOI21X1 AOI21X1_119 ( .A(_abc_40344_n1350), .B(_abc_40344_n2162), .C(_abc_40344_n2245), .Y(_abc_40344_n2246) );
  AOI21X1 AOI21X1_12 ( .A(_abc_40344_n817), .B(_abc_40344_n845), .C(_abc_40344_n846), .Y(_abc_40344_n847) );
  AOI21X1 AOI21X1_120 ( .A(_abc_40344_n2162), .B(_abc_40344_n1665), .C(_abc_40344_n2250), .Y(_abc_40344_n2251) );
  AOI21X1 AOI21X1_121 ( .A(_abc_40344_n2237), .B(_abc_40344_n2262), .C(_abc_40344_n2254), .Y(_abc_40344_n2263) );
  AOI21X1 AOI21X1_122 ( .A(_abc_40344_n2264), .B(_abc_40344_n1326), .C(_abc_40344_n2161), .Y(_abc_40344_n2265) );
  AOI21X1 AOI21X1_123 ( .A(_abc_40344_n2267), .B(_abc_40344_n1968), .C(_abc_40344_n2179), .Y(_abc_40344_n2268) );
  AOI21X1 AOI21X1_124 ( .A(_abc_40344_n1251), .B(_abc_40344_n2162), .C(_abc_40344_n2274), .Y(_abc_40344_n2275) );
  AOI21X1 AOI21X1_125 ( .A(_abc_40344_n1308), .B(_abc_40344_n2162), .C(_abc_40344_n2278), .Y(_abc_40344_n2279) );
  AOI21X1 AOI21X1_126 ( .A(_abc_40344_n1273), .B(_abc_40344_n2162), .C(_abc_40344_n2282), .Y(_abc_40344_n2283) );
  AOI21X1 AOI21X1_127 ( .A(_abc_40344_n2232), .B(_abc_40344_n2263), .C(_abc_40344_n2286), .Y(_abc_40344_n2287) );
  AOI21X1 AOI21X1_128 ( .A(_abc_40344_n2308_1), .B(_abc_40344_n2315), .C(_abc_40344_n2321), .Y(_abc_40344_n2322) );
  AOI21X1 AOI21X1_129 ( .A(_abc_40344_n2037), .B(_abc_40344_n2165), .C(_abc_40344_n2336), .Y(_abc_40344_n2337) );
  AOI21X1 AOI21X1_13 ( .A(_abc_40344_n889), .B(_abc_40344_n720), .C(_abc_40344_n892), .Y(_abc_40344_n893) );
  AOI21X1 AOI21X1_130 ( .A(_abc_40344_n2335), .B(_abc_40344_n2340_1), .C(_abc_40344_n2346), .Y(_abc_40344_n2347) );
  AOI21X1 AOI21X1_131 ( .A(_abc_40344_n2363), .B(_abc_40344_n2369_1), .C(_abc_40344_n2374), .Y(_abc_40344_n2375) );
  AOI21X1 AOI21X1_132 ( .A(_abc_40344_n2388), .B(_abc_40344_n2393), .C(_abc_40344_n2399), .Y(_abc_40344_n2400) );
  AOI21X1 AOI21X1_133 ( .A(_abc_40344_n2162), .B(_abc_40344_n714), .C(_abc_40344_n2420), .Y(_abc_40344_n2421) );
  AOI21X1 AOI21X1_134 ( .A(_abc_40344_n776), .B(_abc_40344_n2165), .C(_abc_40344_n2207), .Y(_abc_40344_n2427) );
  AOI21X1 AOI21X1_135 ( .A(_abc_40344_n856), .B(_abc_40344_n2162), .C(_abc_40344_n2432), .Y(_abc_40344_n2433) );
  AOI21X1 AOI21X1_136 ( .A(_abc_40344_n2438), .B(_abc_40344_n2430), .C(_abc_40344_n2429), .Y(_abc_40344_n2439) );
  AOI21X1 AOI21X1_137 ( .A(_abc_40344_n2446), .B(_abc_40344_n2270), .C(_abc_40344_n2447), .Y(_abc_40344_n2448) );
  AOI21X1 AOI21X1_138 ( .A(_abc_40344_n2449), .B(_abc_40344_n2450), .C(_abc_40344_n2306), .Y(_abc_40344_n2451_1) );
  AOI21X1 AOI21X1_139 ( .A(_abc_40344_n2453), .B(_abc_40344_n2454), .C(_abc_40344_n2455), .Y(_abc_40344_n2456) );
  AOI21X1 AOI21X1_14 ( .A(_abc_40344_n929), .B(_abc_40344_n931), .C(_abc_40344_n916), .Y(_abc_40344_n932) );
  AOI21X1 AOI21X1_140 ( .A(_abc_40344_n2458_1), .B(_abc_40344_n2354), .C(_abc_40344_n2361), .Y(_abc_40344_n2459) );
  AOI21X1 AOI21X1_141 ( .A(_abc_40344_n2461), .B(_abc_40344_n2380_1), .C(_abc_40344_n2386), .Y(_abc_40344_n2462) );
  AOI21X1 AOI21X1_142 ( .A(_abc_40344_n2465), .B(_abc_40344_n2406), .C(_abc_40344_n2410), .Y(_abc_40344_n2466) );
  AOI21X1 AOI21X1_143 ( .A(_abc_40344_n2568), .B(_abc_40344_n2401), .C(_abc_40344_n2101), .Y(_abc_40344_n2569) );
  AOI21X1 AOI21X1_144 ( .A(_abc_40344_n2580), .B(_abc_40344_n2565), .C(_abc_40344_n2576), .Y(_abc_40344_n2581) );
  AOI21X1 AOI21X1_145 ( .A(_abc_40344_n2515), .B(_abc_40344_n2594), .C(_abc_40344_n1935), .Y(_abc_40344_n2595) );
  AOI21X1 AOI21X1_146 ( .A(_abc_40344_n2593_1), .B(_abc_40344_n2589), .C(_abc_40344_n2597), .Y(_abc_40344_n2598) );
  AOI21X1 AOI21X1_147 ( .A(_abc_40344_n2618), .B(_abc_40344_n2620), .C(_abc_40344_n2609), .Y(_abc_40344_n2621) );
  AOI21X1 AOI21X1_148 ( .A(_abc_40344_n2640), .B(_abc_40344_n2581), .C(_abc_40344_n2641), .Y(_abc_40344_n2642) );
  AOI21X1 AOI21X1_149 ( .A(_abc_40344_n2646), .B(_abc_40344_n2635), .C(_abc_40344_n2587), .Y(_abc_40344_n2647) );
  AOI21X1 AOI21X1_15 ( .A(_abc_40344_n901), .B(_abc_40344_n727_1), .C(_abc_40344_n936), .Y(_abc_40344_n937) );
  AOI21X1 AOI21X1_150 ( .A(_abc_40344_n2650_1), .B(_abc_40344_n2653), .C(_abc_40344_n2654), .Y(_abc_40344_n2655) );
  AOI21X1 AOI21X1_151 ( .A(_abc_40344_n2563), .B(_abc_40344_n2415), .C(_abc_40344_n2662), .Y(_abc_40344_n2663) );
  AOI21X1 AOI21X1_152 ( .A(_abc_40344_n585), .B(_abc_40344_n625), .C(_abc_40344_n523), .Y(_abc_40344_n2669) );
  AOI21X1 AOI21X1_153 ( .A(_abc_40344_n2670), .B(B_REG), .C(_abc_40344_n630_1), .Y(_abc_40344_n2671) );
  AOI21X1 AOI21X1_154 ( .A(_abc_40344_n2675), .B(ADDR_REG_0_), .C(_abc_40344_n1802), .Y(_abc_40344_n2676) );
  AOI21X1 AOI21X1_155 ( .A(_abc_40344_n538_1), .B(_abc_40344_n885), .C(_abc_40344_n2678), .Y(_abc_40344_n2679) );
  AOI21X1 AOI21X1_156 ( .A(_abc_40344_n2675), .B(ADDR_REG_1_), .C(_abc_40344_n1679), .Y(_abc_40344_n2687) );
  AOI21X1 AOI21X1_157 ( .A(_abc_40344_n2666_1), .B(_abc_40344_n2693), .C(_abc_40344_n2702), .Y(_abc_40344_n2703) );
  AOI21X1 AOI21X1_158 ( .A(_abc_40344_n2675), .B(ADDR_REG_2_), .C(_abc_40344_n1855), .Y(_abc_40344_n2711) );
  AOI21X1 AOI21X1_159 ( .A(_abc_40344_n2675), .B(ADDR_REG_3_), .C(_abc_40344_n1610), .Y(_abc_40344_n2727) );
  AOI21X1 AOI21X1_16 ( .A(_abc_40344_n945_1), .B(_abc_40344_n565_1), .C(_abc_40344_n561_1), .Y(_abc_40344_n946) );
  AOI21X1 AOI21X1_160 ( .A(_abc_40344_n2738), .B(_abc_40344_n2736), .C(_abc_40344_n1607), .Y(_abc_40344_n2741) );
  AOI21X1 AOI21X1_161 ( .A(_abc_40344_n2666_1), .B(_abc_40344_n2733), .C(_abc_40344_n2743), .Y(_abc_40344_n2744) );
  AOI21X1 AOI21X1_162 ( .A(_abc_40344_n2675), .B(ADDR_REG_4_), .C(_abc_40344_n1776), .Y(_abc_40344_n2746) );
  AOI21X1 AOI21X1_163 ( .A(_abc_40344_n2747), .B(_abc_40344_n2749), .C(_abc_40344_n2750), .Y(_abc_40344_n2751) );
  AOI21X1 AOI21X1_164 ( .A(_abc_40344_n2675), .B(ADDR_REG_5_), .C(_abc_40344_n1745), .Y(_abc_40344_n2760_1) );
  AOI21X1 AOI21X1_165 ( .A(_abc_40344_n748), .B(_abc_40344_n2763), .C(_abc_40344_n2764), .Y(_abc_40344_n2765) );
  AOI21X1 AOI21X1_166 ( .A(_abc_40344_n2768_1), .B(_abc_40344_n2766), .C(_abc_40344_n2667), .Y(_abc_40344_n2769) );
  AOI21X1 AOI21X1_167 ( .A(_abc_40344_n2675), .B(ADDR_REG_7_), .C(_abc_40344_n1034_1), .Y(_abc_40344_n2795) );
  AOI21X1 AOI21X1_168 ( .A(_abc_40344_n2803), .B(_abc_40344_n2805), .C(_abc_40344_n2804), .Y(_abc_40344_n2806) );
  AOI21X1 AOI21X1_169 ( .A(_abc_40344_n610_1), .B(_abc_40344_n2801), .C(_abc_40344_n2809), .Y(_abc_40344_n2810) );
  AOI21X1 AOI21X1_17 ( .A(_abc_40344_n1019), .B(_abc_40344_n1020), .C(_abc_40344_n1024), .Y(_abc_40344_n1025) );
  AOI21X1 AOI21X1_170 ( .A(_abc_40344_n2812), .B(_abc_40344_n2798), .C(_abc_40344_n1007), .Y(_abc_40344_n2813) );
  AOI21X1 AOI21X1_171 ( .A(_abc_40344_n1372), .B(_abc_40344_n2816_1), .C(_abc_40344_n2819), .Y(_abc_40344_n2820) );
  AOI21X1 AOI21X1_172 ( .A(_abc_40344_n2675), .B(ADDR_REG_8_), .C(_abc_40344_n1666), .Y(_abc_40344_n2821) );
  AOI21X1 AOI21X1_173 ( .A(_abc_40344_n2804), .B(_abc_40344_n2805), .C(_abc_40344_n2802), .Y(_abc_40344_n2823_1) );
  AOI21X1 AOI21X1_174 ( .A(_abc_40344_n2829), .B(_abc_40344_n2831), .C(_abc_40344_n2832), .Y(_abc_40344_n2833) );
  AOI21X1 AOI21X1_175 ( .A(_abc_40344_n602), .B(_abc_40344_n1348), .C(_abc_40344_n2833), .Y(_abc_40344_n2834) );
  AOI21X1 AOI21X1_176 ( .A(_abc_40344_n1372), .B(_abc_40344_n2814), .C(_abc_40344_n2813), .Y(_abc_40344_n2838) );
  AOI21X1 AOI21X1_177 ( .A(_abc_40344_n2840), .B(_abc_40344_n2705), .C(_abc_40344_n1789), .Y(_abc_40344_n2841) );
  AOI21X1 AOI21X1_178 ( .A(_abc_40344_n2675), .B(ADDR_REG_10_), .C(_abc_40344_n1594), .Y(_abc_40344_n2843) );
  AOI21X1 AOI21X1_179 ( .A(_abc_40344_n610_1), .B(_abc_40344_n2852), .C(_abc_40344_n2860), .Y(_abc_40344_n2861) );
  AOI21X1 AOI21X1_18 ( .A(_abc_40344_n1032), .B(_abc_40344_n908), .C(_abc_40344_n1034_1), .Y(_abc_40344_n1035) );
  AOI21X1 AOI21X1_180 ( .A(_abc_40344_n2675), .B(ADDR_REG_11_), .C(_abc_40344_n1842), .Y(_abc_40344_n2877) );
  AOI21X1 AOI21X1_181 ( .A(_abc_40344_n2876), .B(_abc_40344_n2871), .C(_abc_40344_n2879), .Y(_abc_40344_n2880) );
  AOI21X1 AOI21X1_182 ( .A(_abc_40344_n2675), .B(ADDR_REG_12_), .C(_abc_40344_n1710), .Y(_abc_40344_n2899) );
  AOI21X1 AOI21X1_183 ( .A(_abc_40344_n2896), .B(_abc_40344_n2871), .C(_abc_40344_n2901), .Y(_abc_40344_n2902) );
  AOI21X1 AOI21X1_184 ( .A(_abc_40344_n2677), .B(_abc_40344_n2918), .C(_abc_40344_n1820), .Y(_abc_40344_n2921) );
  AOI21X1 AOI21X1_185 ( .A(_abc_40344_n2917), .B(_abc_40344_n2871), .C(_abc_40344_n2922), .Y(_abc_40344_n2923) );
  AOI21X1 AOI21X1_186 ( .A(_abc_40344_n2927), .B(_abc_40344_n2929), .C(_abc_40344_n1222), .Y(_abc_40344_n2930) );
  AOI21X1 AOI21X1_187 ( .A(_abc_40344_n1232), .B(_abc_40344_n2926), .C(_abc_40344_n2931), .Y(_abc_40344_n2932) );
  AOI21X1 AOI21X1_188 ( .A(_abc_40344_n2938), .B(_abc_40344_n2942), .C(_abc_40344_n2943), .Y(_abc_40344_n2944) );
  AOI21X1 AOI21X1_189 ( .A(_abc_40344_n2675), .B(ADDR_REG_14_), .C(_abc_40344_n1566), .Y(_abc_40344_n2945) );
  AOI21X1 AOI21X1_19 ( .A(_abc_40344_n912), .B(_abc_40344_n1001), .C(_abc_40344_n1036), .Y(_abc_40344_n1037) );
  AOI21X1 AOI21X1_190 ( .A(_abc_40344_n2949), .B(_abc_40344_n2929), .C(_abc_40344_n1206), .Y(_abc_40344_n2950) );
  AOI21X1 AOI21X1_191 ( .A(_abc_40344_n2967), .B(_abc_40344_n2705), .C(_abc_40344_n2958), .Y(_abc_40344_n2968) );
  AOI21X1 AOI21X1_192 ( .A(_abc_40344_n2983), .B(_abc_40344_n2981), .C(_abc_40344_n2870), .Y(_abc_40344_n2984) );
  AOI21X1 AOI21X1_193 ( .A(_abc_40344_n2675), .B(ADDR_REG_16_), .C(_abc_40344_n1737), .Y(_abc_40344_n2987) );
  AOI21X1 AOI21X1_194 ( .A(_abc_40344_n2998), .B(_abc_40344_n2995), .C(_abc_40344_n2817), .Y(_abc_40344_n2999) );
  AOI21X1 AOI21X1_195 ( .A(_abc_40344_n3005), .B(_abc_40344_n3004), .C(_abc_40344_n2870), .Y(_abc_40344_n3006) );
  AOI21X1 AOI21X1_196 ( .A(_abc_40344_n3008), .B(_abc_40344_n2991), .C(_abc_40344_n3011), .Y(_abc_40344_n3012) );
  AOI21X1 AOI21X1_197 ( .A(_abc_40344_n2675), .B(ADDR_REG_18_), .C(_abc_40344_n1864), .Y(_abc_40344_n3014) );
  AOI21X1 AOI21X1_198 ( .A(_abc_40344_n3024), .B(_abc_40344_n2871), .C(_abc_40344_n3015), .Y(_abc_40344_n3025) );
  AOI21X1 AOI21X1_199 ( .A(_abc_40344_n3029), .B(_abc_40344_n2993), .C(_abc_40344_n3028), .Y(_abc_40344_n3030) );
  AOI21X1 AOI21X1_2 ( .A(_abc_40344_n646), .B(_abc_40344_n625), .C(_abc_40344_n641), .Y(_abc_40344_n647) );
  AOI21X1 AOI21X1_20 ( .A(REG0_REG_27_), .B(_abc_40344_n673), .C(_abc_40344_n1071), .Y(_abc_40344_n1072) );
  AOI21X1 AOI21X1_200 ( .A(_abc_40344_n2675), .B(ADDR_REG_19_), .C(_abc_40344_n1623), .Y(_abc_40344_n3036) );
  AOI21X1 AOI21X1_201 ( .A(_abc_40344_n1411), .B(_abc_40344_n648), .C(_abc_40344_n3042), .Y(_abc_40344_n3043) );
  AOI21X1 AOI21X1_202 ( .A(_abc_40344_n3044), .B(_abc_40344_n3041_1), .C(_abc_40344_n3018), .Y(_abc_40344_n3045) );
  AOI21X1 AOI21X1_203 ( .A(_abc_40344_n3046), .B(_abc_40344_n2871), .C(_abc_40344_n3037), .Y(_abc_40344_n3047) );
  AOI21X1 AOI21X1_204 ( .A(_abc_40344_n3050), .B(_abc_40344_n2992), .C(_abc_40344_n3027), .Y(_abc_40344_n3051) );
  AOI21X1 AOI21X1_205 ( .A(_abc_40344_n3029), .B(_abc_40344_n2993), .C(_abc_40344_n3026), .Y(_abc_40344_n3052) );
  AOI21X1 AOI21X1_206 ( .A(_abc_40344_n3101), .B(_abc_40344_n3100), .C(_abc_40344_n3069), .Y(_abc_40344_n3102) );
  AOI21X1 AOI21X1_207 ( .A(REG2_REG_31_), .B(_abc_40344_n3067), .C(_abc_40344_n3107), .Y(_abc_40344_n3108) );
  AOI21X1 AOI21X1_208 ( .A(_abc_40344_n3115), .B(_abc_40344_n3114), .C(_abc_40344_n3069), .Y(_abc_40344_n3116) );
  AOI21X1 AOI21X1_209 ( .A(REG2_REG_30_), .B(_abc_40344_n3067), .C(_abc_40344_n3107), .Y(_abc_40344_n3117) );
  AOI21X1 AOI21X1_21 ( .A(_abc_40344_n1086), .B(_abc_40344_n685_1), .C(_abc_40344_n1089), .Y(_abc_40344_n1090_1) );
  AOI21X1 AOI21X1_210 ( .A(_abc_40344_n1251), .B(_abc_40344_n1260), .C(_abc_40344_n2501), .Y(_abc_40344_n3165) );
  AOI21X1 AOI21X1_211 ( .A(_abc_40344_n3159), .B(_abc_40344_n3175), .C(_abc_40344_n3170), .Y(_abc_40344_n3176) );
  AOI21X1 AOI21X1_212 ( .A(_abc_40344_n1418), .B(_abc_40344_n1414), .C(_abc_40344_n3179), .Y(_abc_40344_n3180) );
  AOI21X1 AOI21X1_213 ( .A(_abc_40344_n3182), .B(_abc_40344_n3183), .C(_abc_40344_n3179), .Y(_abc_40344_n3184) );
  AOI21X1 AOI21X1_214 ( .A(_abc_40344_n1434), .B(_abc_40344_n1441), .C(_abc_40344_n3184), .Y(_abc_40344_n3185) );
  AOI21X1 AOI21X1_215 ( .A(_abc_40344_n3189), .B(_abc_40344_n2541), .C(_abc_40344_n2540), .Y(_abc_40344_n3190) );
  AOI21X1 AOI21X1_216 ( .A(_abc_40344_n1495), .B(_abc_40344_n1507_1), .C(_abc_40344_n3206), .Y(_abc_40344_n3207) );
  AOI21X1 AOI21X1_217 ( .A(_abc_40344_n3226), .B(_abc_40344_n3120), .C(_abc_40344_n3228), .Y(_abc_40344_n3229) );
  AOI21X1 AOI21X1_218 ( .A(_abc_40344_n3067), .B(REG2_REG_28_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3234) );
  AOI21X1 AOI21X1_219 ( .A(_abc_40344_n1645), .B(_abc_40344_n3233), .C(_abc_40344_n3235), .Y(_abc_40344_n3236) );
  AOI21X1 AOI21X1_22 ( .A(_abc_40344_n1247), .B(IR_REG_13_), .C(_abc_40344_n574), .Y(_abc_40344_n1248) );
  AOI21X1 AOI21X1_220 ( .A(_abc_40344_n3231), .B(_abc_40344_n3066), .C(_abc_40344_n3241), .Y(_abc_40344_n3242) );
  AOI21X1 AOI21X1_221 ( .A(_abc_40344_n3225), .B(_abc_40344_n3248), .C(_abc_40344_n3228), .Y(_abc_40344_n3249) );
  AOI21X1 AOI21X1_222 ( .A(_abc_40344_n3067), .B(REG2_REG_27_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3254) );
  AOI21X1 AOI21X1_223 ( .A(_abc_40344_n3252), .B(_abc_40344_n3068), .C(_abc_40344_n3256), .Y(_abc_40344_n3257) );
  AOI21X1 AOI21X1_224 ( .A(_abc_40344_n3251), .B(_abc_40344_n3066), .C(_abc_40344_n3258), .Y(_abc_40344_n3259) );
  AOI21X1 AOI21X1_225 ( .A(_abc_40344_n3067), .B(REG2_REG_26_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3276) );
  AOI21X1 AOI21X1_226 ( .A(_abc_40344_n3274), .B(_abc_40344_n3068), .C(_abc_40344_n3278), .Y(_abc_40344_n3279) );
  AOI21X1 AOI21X1_227 ( .A(_abc_40344_n3270), .B(_abc_40344_n3066), .C(_abc_40344_n3280), .Y(_abc_40344_n3281) );
  AOI21X1 AOI21X1_228 ( .A(_abc_40344_n2647), .B(_abc_40344_n2514), .C(_abc_40344_n3228), .Y(_abc_40344_n3285) );
  AOI21X1 AOI21X1_229 ( .A(_abc_40344_n3067), .B(REG2_REG_25_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3288) );
  AOI21X1 AOI21X1_23 ( .A(_abc_40344_n705_1), .B(_abc_40344_n1249), .C(_abc_40344_n1250), .Y(_abc_40344_n1251) );
  AOI21X1 AOI21X1_230 ( .A(_abc_40344_n1507_1), .B(_abc_40344_n3233), .C(_abc_40344_n3289), .Y(_abc_40344_n3290) );
  AOI21X1 AOI21X1_231 ( .A(_abc_40344_n3066), .B(_abc_40344_n3287), .C(_abc_40344_n3293), .Y(_abc_40344_n3294) );
  AOI21X1 AOI21X1_232 ( .A(_abc_40344_n3307), .B(_abc_40344_n2490), .C(_abc_40344_n2628), .Y(_abc_40344_n3308) );
  AOI21X1 AOI21X1_233 ( .A(_abc_40344_n3310), .B(_abc_40344_n3311), .C(_abc_40344_n3312), .Y(_abc_40344_n3313) );
  AOI21X1 AOI21X1_234 ( .A(_abc_40344_n3320), .B(_abc_40344_n1938), .C(_abc_40344_n2068), .Y(_abc_40344_n3321) );
  AOI21X1 AOI21X1_235 ( .A(_abc_40344_n3067), .B(REG2_REG_24_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3345) );
  AOI21X1 AOI21X1_236 ( .A(_abc_40344_n3344), .B(_abc_40344_n3066), .C(_abc_40344_n3346), .Y(_abc_40344_n3347) );
  AOI21X1 AOI21X1_237 ( .A(_abc_40344_n3218), .B(_abc_40344_n3296), .C(_abc_40344_n3348), .Y(_abc_40344_n3349) );
  AOI21X1 AOI21X1_238 ( .A(_abc_40344_n3067), .B(REG2_REG_23_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3373) );
  AOI21X1 AOI21X1_239 ( .A(_abc_40344_n1030_1), .B(_abc_40344_n1086), .C(_abc_40344_n3374), .Y(_abc_40344_n3375) );
  AOI21X1 AOI21X1_24 ( .A(_abc_40344_n705_1), .B(_abc_40344_n1271), .C(_abc_40344_n1272), .Y(_abc_40344_n1273) );
  AOI21X1 AOI21X1_240 ( .A(_abc_40344_n3372), .B(_abc_40344_n3068), .C(_abc_40344_n3376), .Y(_abc_40344_n3377) );
  AOI21X1 AOI21X1_241 ( .A(_abc_40344_n3383), .B(_abc_40344_n3382), .C(_abc_40344_n3228), .Y(_abc_40344_n3384) );
  AOI21X1 AOI21X1_242 ( .A(_abc_40344_n3067), .B(REG2_REG_22_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3390) );
  AOI21X1 AOI21X1_243 ( .A(_abc_40344_n3388_1), .B(_abc_40344_n3068), .C(_abc_40344_n3393), .Y(_abc_40344_n3394) );
  AOI21X1 AOI21X1_244 ( .A(_abc_40344_n3398), .B(_abc_40344_n3399), .C(_abc_40344_n3400), .Y(_abc_40344_n3401) );
  AOI21X1 AOI21X1_245 ( .A(_abc_40344_n3067), .B(REG2_REG_21_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3417) );
  AOI21X1 AOI21X1_246 ( .A(_abc_40344_n3415), .B(_abc_40344_n3066), .C(_abc_40344_n3420), .Y(_abc_40344_n3421) );
  AOI21X1 AOI21X1_247 ( .A(_abc_40344_n3355), .B(_abc_40344_n2064), .C(_abc_40344_n2471), .Y(_abc_40344_n3426) );
  AOI21X1 AOI21X1_248 ( .A(_abc_40344_n3426), .B(_abc_40344_n2527), .C(_abc_40344_n3228), .Y(_abc_40344_n3427) );
  AOI21X1 AOI21X1_249 ( .A(_abc_40344_n3067), .B(REG2_REG_20_), .C(_abc_40344_n3439), .Y(_abc_40344_n3440) );
  AOI21X1 AOI21X1_25 ( .A(_abc_40344_n1051_1), .B(REG3_REG_10_), .C(REG3_REG_11_), .Y(_abc_40344_n1277) );
  AOI21X1 AOI21X1_250 ( .A(_abc_40344_n3436), .B(_abc_40344_n3066), .C(_abc_40344_n3442), .Y(_abc_40344_n3443) );
  AOI21X1 AOI21X1_251 ( .A(_abc_40344_n3067), .B(REG2_REG_19_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3448) );
  AOI21X1 AOI21X1_252 ( .A(_abc_40344_n3445), .B(_abc_40344_n3218), .C(_abc_40344_n3451), .Y(_abc_40344_n3452) );
  AOI21X1 AOI21X1_253 ( .A(_abc_40344_n2473), .B(_abc_40344_n3326), .C(_abc_40344_n3453), .Y(_abc_40344_n3454) );
  AOI21X1 AOI21X1_254 ( .A(_abc_40344_n3066), .B(_abc_40344_n3464), .C(_abc_40344_n3475), .Y(_abc_40344_n3476) );
  AOI21X1 AOI21X1_255 ( .A(_abc_40344_n3484), .B(_abc_40344_n3478_1), .C(_abc_40344_n3228), .Y(_abc_40344_n3485) );
  AOI21X1 AOI21X1_256 ( .A(_abc_40344_n3066), .B(_abc_40344_n3493), .C(_abc_40344_n3494), .Y(_abc_40344_n3495) );
  AOI21X1 AOI21X1_257 ( .A(_abc_40344_n3218), .B(_abc_40344_n3480), .C(_abc_40344_n3497), .Y(_abc_40344_n3498) );
  AOI21X1 AOI21X1_258 ( .A(_abc_40344_n3502), .B(_abc_40344_n2537), .C(_abc_40344_n1963), .Y(_abc_40344_n3503) );
  AOI21X1 AOI21X1_259 ( .A(_abc_40344_n3110), .B(_abc_40344_n1153), .C(_abc_40344_n3513), .Y(_abc_40344_n3514) );
  AOI21X1 AOI21X1_26 ( .A(_abc_40344_n705_1), .B(_abc_40344_n1293_1), .C(_abc_40344_n1307), .Y(_abc_40344_n1308) );
  AOI21X1 AOI21X1_260 ( .A(_abc_40344_n3510), .B(_abc_40344_n3068), .C(_abc_40344_n3515), .Y(_abc_40344_n3516) );
  AOI21X1 AOI21X1_261 ( .A(_abc_40344_n3067), .B(REG2_REG_15_), .C(_abc_40344_n3532), .Y(_abc_40344_n3533) );
  AOI21X1 AOI21X1_262 ( .A(_abc_40344_n1168), .B(_abc_40344_n3233), .C(_abc_40344_n3534), .Y(_abc_40344_n3535_1) );
  AOI21X1 AOI21X1_263 ( .A(_abc_40344_n3218), .B(_abc_40344_n3520), .C(_abc_40344_n3536), .Y(_abc_40344_n3537) );
  AOI21X1 AOI21X1_264 ( .A(_abc_40344_n3110), .B(_abc_40344_n1224), .C(_abc_40344_n3551), .Y(_abc_40344_n3552) );
  AOI21X1 AOI21X1_265 ( .A(_abc_40344_n3218), .B(_abc_40344_n3541), .C(_abc_40344_n3554), .Y(_abc_40344_n3555_1) );
  AOI21X1 AOI21X1_266 ( .A(_abc_40344_n3110), .B(_abc_40344_n1251), .C(_abc_40344_n3569), .Y(_abc_40344_n3570) );
  AOI21X1 AOI21X1_267 ( .A(_abc_40344_n3566), .B(_abc_40344_n3066), .C(_abc_40344_n3571), .Y(_abc_40344_n3572) );
  AOI21X1 AOI21X1_268 ( .A(_abc_40344_n3304), .B(_abc_40344_n3306), .C(_abc_40344_n3319), .Y(_abc_40344_n3577) );
  AOI21X1 AOI21X1_269 ( .A(_abc_40344_n3067), .B(REG2_REG_12_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3587) );
  AOI21X1 AOI21X1_27 ( .A(_abc_40344_n1385), .B(_abc_40344_n1380), .C(_abc_40344_n1383_1), .Y(_abc_40344_n1386) );
  AOI21X1 AOI21X1_270 ( .A(_abc_40344_n3583), .B(_abc_40344_n3066), .C(_abc_40344_n3590), .Y(_abc_40344_n3591) );
  AOI21X1 AOI21X1_271 ( .A(_abc_40344_n3067), .B(REG2_REG_11_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3601) );
  AOI21X1 AOI21X1_272 ( .A(_abc_40344_n3600), .B(_abc_40344_n3066), .C(_abc_40344_n3607), .Y(_abc_40344_n3608) );
  AOI21X1 AOI21X1_273 ( .A(_abc_40344_n3619), .B(_abc_40344_n3218), .C(_abc_40344_n3632_1), .Y(_abc_40344_n3633) );
  AOI21X1 AOI21X1_274 ( .A(_abc_40344_n3233), .B(_abc_40344_n1335), .C(_abc_40344_n3645), .Y(_abc_40344_n3646) );
  AOI21X1 AOI21X1_275 ( .A(_abc_40344_n3642), .B(_abc_40344_n3066), .C(_abc_40344_n3648), .Y(_abc_40344_n3649) );
  AOI21X1 AOI21X1_276 ( .A(_abc_40344_n3067), .B(REG2_REG_8_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3659) );
  AOI21X1 AOI21X1_277 ( .A(_abc_40344_n3067), .B(REG2_REG_7_), .C(_abc_40344_n3679), .Y(_abc_40344_n3680) );
  AOI21X1 AOI21X1_278 ( .A(_abc_40344_n908), .B(_abc_40344_n3110), .C(_abc_40344_n3681), .Y(_abc_40344_n3682_1) );
  AOI21X1 AOI21X1_279 ( .A(_abc_40344_n3677), .B(_abc_40344_n3066), .C(_abc_40344_n3683), .Y(_abc_40344_n3684) );
  AOI21X1 AOI21X1_28 ( .A(_abc_40344_n1336), .B(_abc_40344_n1338), .C(_abc_40344_n1319), .Y(_abc_40344_n1392) );
  AOI21X1 AOI21X1_280 ( .A(_abc_40344_n3067), .B(REG2_REG_6_), .C(_abc_40344_n3696), .Y(_abc_40344_n3697) );
  AOI21X1 AOI21X1_281 ( .A(_abc_40344_n714), .B(_abc_40344_n3110), .C(_abc_40344_n3698), .Y(_abc_40344_n3699) );
  AOI21X1 AOI21X1_282 ( .A(_abc_40344_n3694), .B(_abc_40344_n3066), .C(_abc_40344_n3700), .Y(_abc_40344_n3701) );
  AOI21X1 AOI21X1_283 ( .A(_abc_40344_n3705), .B(_abc_40344_n3139), .C(_abc_40344_n3152), .Y(_abc_40344_n3706_1) );
  AOI21X1 AOI21X1_284 ( .A(_abc_40344_n3068), .B(_abc_40344_n3718), .C(_abc_40344_n3721), .Y(_abc_40344_n3722) );
  AOI21X1 AOI21X1_285 ( .A(_abc_40344_n3072), .B(_abc_40344_n777_1), .C(_abc_40344_n3726), .Y(_abc_40344_n3727_1) );
  AOI21X1 AOI21X1_286 ( .A(_abc_40344_n777_1), .B(_abc_40344_n995), .C(_abc_40344_n3732), .Y(_abc_40344_n3733) );
  AOI21X1 AOI21X1_287 ( .A(_abc_40344_n2018), .B(_abc_40344_n2490), .C(_abc_40344_n3307), .Y(_abc_40344_n3740) );
  AOI21X1 AOI21X1_288 ( .A(_abc_40344_n3071), .B(_abc_40344_n1609), .C(_abc_40344_n3726), .Y(_abc_40344_n3748) );
  AOI21X1 AOI21X1_289 ( .A(_abc_40344_n3067), .B(REG2_REG_2_), .C(_abc_40344_n3767), .Y(_abc_40344_n3768) );
  AOI21X1 AOI21X1_29 ( .A(_abc_40344_n1395), .B(_abc_40344_n1216), .C(_abc_40344_n1191), .Y(_abc_40344_n1396_1) );
  AOI21X1 AOI21X1_290 ( .A(_abc_40344_n2631), .B(_abc_40344_n2488), .C(_abc_40344_n3771_1), .Y(_abc_40344_n3772_1) );
  AOI21X1 AOI21X1_291 ( .A(_abc_40344_n887), .B(_abc_40344_n3220), .C(_abc_40344_n3772_1), .Y(_abc_40344_n3773_1) );
  AOI21X1 AOI21X1_292 ( .A(_abc_40344_n869), .B(_abc_40344_n1797), .C(_abc_40344_n3726), .Y(_abc_40344_n3776_1) );
  AOI21X1 AOI21X1_293 ( .A(_abc_40344_n3067), .B(REG2_REG_1_), .C(_abc_40344_n3781_1), .Y(_abc_40344_n3782_1) );
  AOI21X1 AOI21X1_294 ( .A(_abc_40344_n3066), .B(_abc_40344_n3790_1), .C(_abc_40344_n630_1), .Y(_abc_40344_n3791_1) );
  AOI21X1 AOI21X1_295 ( .A(n1336), .B(DATAI_31_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3858_1) );
  AOI21X1 AOI21X1_296 ( .A(n1336), .B(DATAI_30_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3862) );
  AOI21X1 AOI21X1_297 ( .A(n1336), .B(DATAI_29_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3867) );
  AOI21X1 AOI21X1_298 ( .A(_abc_40344_n3860), .B(IR_REG_27_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3875) );
  AOI21X1 AOI21X1_299 ( .A(n1336), .B(DATAI_26_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3880_1) );
  AOI21X1 AOI21X1_3 ( .A(_abc_40344_n596_1), .B(_abc_40344_n574), .C(_abc_40344_n670), .Y(_abc_40344_n671_1) );
  AOI21X1 AOI21X1_30 ( .A(_abc_40344_n1399), .B(_abc_40344_n1400), .C(_abc_40344_n1397), .Y(_abc_40344_n1401) );
  AOI21X1 AOI21X1_300 ( .A(n1336), .B(DATAI_25_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3885) );
  AOI21X1 AOI21X1_301 ( .A(n1336), .B(DATAI_24_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3891) );
  AOI21X1 AOI21X1_302 ( .A(n1336), .B(DATAI_23_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3895) );
  AOI21X1 AOI21X1_303 ( .A(n1336), .B(DATAI_22_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3898) );
  AOI21X1 AOI21X1_304 ( .A(n1336), .B(DATAI_21_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3902) );
  AOI21X1 AOI21X1_305 ( .A(n1336), .B(DATAI_20_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3908_1) );
  AOI21X1 AOI21X1_306 ( .A(n1336), .B(DATAI_18_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3917) );
  AOI21X1 AOI21X1_307 ( .A(n1336), .B(DATAI_17_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3922) );
  AOI21X1 AOI21X1_308 ( .A(n1336), .B(DATAI_16_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3927) );
  AOI21X1 AOI21X1_309 ( .A(_abc_40344_n3860), .B(IR_REG_15_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3931) );
  AOI21X1 AOI21X1_31 ( .A(_abc_40344_n1436), .B(_abc_40344_n685_1), .C(_abc_40344_n1439_1), .Y(_abc_40344_n1440) );
  AOI21X1 AOI21X1_310 ( .A(n1336), .B(DATAI_14_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3936) );
  AOI21X1 AOI21X1_311 ( .A(n1336), .B(DATAI_13_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3941) );
  AOI21X1 AOI21X1_312 ( .A(n1336), .B(DATAI_11_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3950) );
  AOI21X1 AOI21X1_313 ( .A(n1336), .B(DATAI_10_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3954) );
  AOI21X1 AOI21X1_314 ( .A(n1336), .B(DATAI_9_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3959) );
  AOI21X1 AOI21X1_315 ( .A(n1336), .B(DATAI_8_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3963) );
  AOI21X1 AOI21X1_316 ( .A(_abc_40344_n3860), .B(IR_REG_7_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3967) );
  AOI21X1 AOI21X1_317 ( .A(_abc_40344_n3860), .B(IR_REG_6_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3971) );
  AOI21X1 AOI21X1_318 ( .A(_abc_40344_n3860), .B(IR_REG_5_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3975) );
  AOI21X1 AOI21X1_319 ( .A(_abc_40344_n3860), .B(IR_REG_4_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3979_1) );
  AOI21X1 AOI21X1_32 ( .A(_abc_40344_n1402), .B(_abc_40344_n1141), .C(_abc_40344_n1448), .Y(_abc_40344_n1449) );
  AOI21X1 AOI21X1_320 ( .A(_abc_40344_n3860), .B(IR_REG_3_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3983) );
  AOI21X1 AOI21X1_321 ( .A(n1336), .B(DATAI_2_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3987) );
  AOI21X1 AOI21X1_322 ( .A(n1336), .B(DATAI_1_), .C(_abc_40344_n630_1), .Y(_abc_40344_n3991) );
  AOI21X1 AOI21X1_323 ( .A(IR_REG_0_), .B(STATE_REG), .C(_abc_40344_n630_1), .Y(_abc_40344_n3995) );
  AOI21X1 AOI21X1_324 ( .A(_abc_40344_n2637), .B(_abc_40344_n1932), .C(_abc_40344_n2648), .Y(_abc_40344_n4012) );
  AOI21X1 AOI21X1_325 ( .A(_abc_40344_n4014), .B(_abc_40344_n4018), .C(_abc_40344_n3228), .Y(_abc_40344_n4019) );
  AOI21X1 AOI21X1_326 ( .A(_abc_40344_n3067), .B(REG2_REG_29_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4025) );
  AOI21X1 AOI21X1_327 ( .A(_abc_40344_n2394), .B(_abc_40344_n3110), .C(_abc_40344_n4026_1), .Y(_abc_40344_n4027) );
  AOI21X1 AOI21X1_328 ( .A(_abc_40344_n3068), .B(_abc_40344_n4023), .C(_abc_40344_n4028), .Y(_abc_40344_n4029) );
  AOI21X1 AOI21X1_329 ( .A(_abc_40344_n3794_1), .B(_abc_40344_n4032), .C(_abc_40344_n630_1), .Y(_abc_40344_n4033_1) );
  AOI21X1 AOI21X1_33 ( .A(REG0_REG_24_), .B(_abc_40344_n673), .C(_abc_40344_n1469), .Y(_abc_40344_n1470) );
  AOI21X1 AOI21X1_330 ( .A(_abc_40344_n3794_1), .B(_abc_40344_n944), .C(_abc_40344_n630_1), .Y(_abc_40344_n4036) );
  AOI21X1 AOI21X1_331 ( .A(_abc_40344_n2529_1), .B(_abc_40344_n4044), .C(_abc_40344_n3788_1), .Y(_abc_40344_n4045) );
  AOI21X1 AOI21X1_332 ( .A(_abc_40344_n4043), .B(REG0_REG_0_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4046_1) );
  AOI21X1 AOI21X1_333 ( .A(_abc_40344_n4058_1), .B(_abc_40344_n4042), .C(_abc_40344_n630_1), .Y(_abc_40344_n4059) );
  AOI21X1 AOI21X1_334 ( .A(_abc_40344_n4071), .B(_abc_40344_n4042), .C(_abc_40344_n630_1), .Y(_abc_40344_n4072) );
  AOI21X1 AOI21X1_335 ( .A(_abc_40344_n3671), .B(_abc_40344_n3725), .C(_abc_40344_n4080), .Y(_abc_40344_n4081) );
  AOI21X1 AOI21X1_336 ( .A(_abc_40344_n3665), .B(_abc_40344_n3725), .C(_abc_40344_n4086), .Y(_abc_40344_n4087) );
  AOI21X1 AOI21X1_337 ( .A(_abc_40344_n3636), .B(_abc_40344_n3725), .C(_abc_40344_n4092), .Y(_abc_40344_n4093) );
  AOI21X1 AOI21X1_338 ( .A(_abc_40344_n3619), .B(_abc_40344_n4048), .C(_abc_40344_n4099), .Y(_abc_40344_n4100) );
  AOI21X1 AOI21X1_339 ( .A(_abc_40344_n4101_1), .B(_abc_40344_n4042), .C(_abc_40344_n630_1), .Y(_abc_40344_n4102) );
  AOI21X1 AOI21X1_34 ( .A(_abc_40344_n1496), .B(_abc_40344_n1497), .C(_abc_40344_n921), .Y(_abc_40344_n1498) );
  AOI21X1 AOI21X1_340 ( .A(_abc_40344_n3605), .B(_abc_40344_n3725), .C(_abc_40344_n4104), .Y(_abc_40344_n4105) );
  AOI21X1 AOI21X1_341 ( .A(_abc_40344_n1260), .B(_abc_40344_n3103), .C(_abc_40344_n4110), .Y(_abc_40344_n4111) );
  AOI21X1 AOI21X1_342 ( .A(_abc_40344_n995), .B(_abc_40344_n1224), .C(_abc_40344_n4124), .Y(_abc_40344_n4125_1) );
  AOI21X1 AOI21X1_343 ( .A(_abc_40344_n3490), .B(_abc_40344_n3725), .C(_abc_40344_n4146), .Y(_abc_40344_n4147) );
  AOI21X1 AOI21X1_344 ( .A(_abc_40344_n4148), .B(_abc_40344_n4042), .C(_abc_40344_n630_1), .Y(_abc_40344_n4149_1) );
  AOI21X1 AOI21X1_345 ( .A(_abc_40344_n3468), .B(_abc_40344_n3725), .C(_abc_40344_n3470), .Y(_abc_40344_n4151) );
  AOI21X1 AOI21X1_346 ( .A(_abc_40344_n4157), .B(_abc_40344_n3725), .C(_abc_40344_n4158_1), .Y(_abc_40344_n4159) );
  AOI21X1 AOI21X1_347 ( .A(_abc_40344_n4164), .B(_abc_40344_n3725), .C(_abc_40344_n3437), .Y(_abc_40344_n4165) );
  AOI21X1 AOI21X1_348 ( .A(_abc_40344_n4043), .B(REG0_REG_20_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4168) );
  AOI21X1 AOI21X1_349 ( .A(_abc_40344_n3396), .B(_abc_40344_n3725), .C(_abc_40344_n4170), .Y(_abc_40344_n4171_1) );
  AOI21X1 AOI21X1_35 ( .A(_abc_40344_n1532), .B(_abc_40344_n1098), .C(_abc_40344_n1514_1), .Y(_abc_40344_n1533) );
  AOI21X1 AOI21X1_350 ( .A(_abc_40344_n4043), .B(REG0_REG_21_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4174) );
  AOI21X1 AOI21X1_351 ( .A(_abc_40344_n3388_1), .B(_abc_40344_n3725), .C(_abc_40344_n4177_1), .Y(_abc_40344_n4178) );
  AOI21X1 AOI21X1_352 ( .A(_abc_40344_n4043), .B(REG0_REG_22_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4180) );
  AOI21X1 AOI21X1_353 ( .A(_abc_40344_n4043), .B(REG0_REG_23_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4187_1) );
  AOI21X1 AOI21X1_354 ( .A(_abc_40344_n4043), .B(REG0_REG_24_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4193_1) );
  AOI21X1 AOI21X1_355 ( .A(_abc_40344_n3291), .B(_abc_40344_n3725), .C(_abc_40344_n4195_1), .Y(_abc_40344_n4196) );
  AOI21X1 AOI21X1_356 ( .A(_abc_40344_n4043), .B(REG0_REG_25_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4199_1) );
  AOI21X1 AOI21X1_357 ( .A(_abc_40344_n3274), .B(_abc_40344_n3725), .C(_abc_40344_n4201_1), .Y(_abc_40344_n4202) );
  AOI21X1 AOI21X1_358 ( .A(_abc_40344_n4043), .B(REG0_REG_26_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4205_1) );
  AOI21X1 AOI21X1_359 ( .A(_abc_40344_n3252), .B(_abc_40344_n3725), .C(_abc_40344_n4207_1), .Y(_abc_40344_n4208) );
  AOI21X1 AOI21X1_36 ( .A(_abc_40344_n1032), .B(_abc_40344_n1076), .C(_abc_40344_n1552), .Y(_abc_40344_n1553) );
  AOI21X1 AOI21X1_360 ( .A(_abc_40344_n4043), .B(REG0_REG_27_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4211_1) );
  AOI21X1 AOI21X1_361 ( .A(_abc_40344_n3239), .B(_abc_40344_n3725), .C(_abc_40344_n4213_1), .Y(_abc_40344_n4214) );
  AOI21X1 AOI21X1_362 ( .A(_abc_40344_n4043), .B(REG0_REG_28_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4217_1) );
  AOI21X1 AOI21X1_363 ( .A(_abc_40344_n4021), .B(_abc_40344_n4022), .C(_abc_40344_n3726), .Y(_abc_40344_n4221_1) );
  AOI21X1 AOI21X1_364 ( .A(_abc_40344_n4043), .B(REG0_REG_29_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4225_1) );
  AOI21X1 AOI21X1_365 ( .A(_abc_40344_n3115), .B(_abc_40344_n3114), .C(_abc_40344_n3726), .Y(_abc_40344_n4227_1) );
  AOI21X1 AOI21X1_366 ( .A(_abc_40344_n4043), .B(REG0_REG_30_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4230) );
  AOI21X1 AOI21X1_367 ( .A(_abc_40344_n3101), .B(_abc_40344_n3100), .C(_abc_40344_n3726), .Y(_abc_40344_n4232) );
  AOI21X1 AOI21X1_368 ( .A(_abc_40344_n4238_1), .B(REG1_REG_0_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4239_1) );
  AOI21X1 AOI21X1_369 ( .A(_abc_40344_n4058_1), .B(_abc_40344_n4237), .C(_abc_40344_n630_1), .Y(_abc_40344_n4244_1) );
  AOI21X1 AOI21X1_37 ( .A(_abc_40344_n1551), .B(_abc_40344_n1005), .C(_abc_40344_n1556), .Y(_abc_40344_n1557) );
  AOI21X1 AOI21X1_370 ( .A(_abc_40344_n4071), .B(_abc_40344_n4237), .C(_abc_40344_n630_1), .Y(_abc_40344_n4252) );
  AOI21X1 AOI21X1_371 ( .A(_abc_40344_n4101_1), .B(_abc_40344_n4237), .C(_abc_40344_n630_1), .Y(_abc_40344_n4266_1) );
  AOI21X1 AOI21X1_372 ( .A(_abc_40344_n4148), .B(_abc_40344_n4237), .C(_abc_40344_n630_1), .Y(_abc_40344_n4286_1) );
  AOI21X1 AOI21X1_373 ( .A(_abc_40344_n4238_1), .B(REG1_REG_20_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4295_1) );
  AOI21X1 AOI21X1_374 ( .A(_abc_40344_n4238_1), .B(REG1_REG_21_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4298_1) );
  AOI21X1 AOI21X1_375 ( .A(_abc_40344_n4238_1), .B(REG1_REG_22_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4300) );
  AOI21X1 AOI21X1_376 ( .A(_abc_40344_n4238_1), .B(REG1_REG_23_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4303) );
  AOI21X1 AOI21X1_377 ( .A(_abc_40344_n4238_1), .B(REG1_REG_24_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4306) );
  AOI21X1 AOI21X1_378 ( .A(_abc_40344_n4238_1), .B(REG1_REG_25_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4309) );
  AOI21X1 AOI21X1_379 ( .A(_abc_40344_n4238_1), .B(REG1_REG_26_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4312) );
  AOI21X1 AOI21X1_38 ( .A(_abc_40344_n1032), .B(_abc_40344_n1224), .C(_abc_40344_n1566), .Y(_abc_40344_n1567) );
  AOI21X1 AOI21X1_380 ( .A(_abc_40344_n4238_1), .B(REG1_REG_27_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4315) );
  AOI21X1 AOI21X1_381 ( .A(_abc_40344_n4238_1), .B(REG1_REG_28_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4318) );
  AOI21X1 AOI21X1_382 ( .A(_abc_40344_n4238_1), .B(REG1_REG_29_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4321) );
  AOI21X1 AOI21X1_383 ( .A(_abc_40344_n589), .B(DATAO_REG_0_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4330) );
  AOI21X1 AOI21X1_384 ( .A(_abc_40344_n589), .B(DATAO_REG_1_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4332) );
  AOI21X1 AOI21X1_385 ( .A(_abc_40344_n589), .B(DATAO_REG_2_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4334) );
  AOI21X1 AOI21X1_386 ( .A(_abc_40344_n589), .B(DATAO_REG_3_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4336) );
  AOI21X1 AOI21X1_387 ( .A(_abc_40344_n589), .B(DATAO_REG_4_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4338) );
  AOI21X1 AOI21X1_388 ( .A(_abc_40344_n589), .B(DATAO_REG_5_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4340) );
  AOI21X1 AOI21X1_389 ( .A(_abc_40344_n589), .B(DATAO_REG_6_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4342) );
  AOI21X1 AOI21X1_39 ( .A(_abc_40344_n1005), .B(_abc_40344_n1565), .C(_abc_40344_n1568), .Y(_abc_40344_n1569) );
  AOI21X1 AOI21X1_390 ( .A(_abc_40344_n589), .B(DATAO_REG_7_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4344) );
  AOI21X1 AOI21X1_391 ( .A(_abc_40344_n589), .B(DATAO_REG_8_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4346) );
  AOI21X1 AOI21X1_392 ( .A(_abc_40344_n589), .B(DATAO_REG_9_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4348) );
  AOI21X1 AOI21X1_393 ( .A(_abc_40344_n589), .B(DATAO_REG_10_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4350) );
  AOI21X1 AOI21X1_394 ( .A(_abc_40344_n589), .B(DATAO_REG_11_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4352) );
  AOI21X1 AOI21X1_395 ( .A(_abc_40344_n589), .B(DATAO_REG_12_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4354) );
  AOI21X1 AOI21X1_396 ( .A(_abc_40344_n589), .B(DATAO_REG_13_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4356) );
  AOI21X1 AOI21X1_397 ( .A(_abc_40344_n589), .B(DATAO_REG_14_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4358) );
  AOI21X1 AOI21X1_398 ( .A(_abc_40344_n589), .B(DATAO_REG_15_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4360) );
  AOI21X1 AOI21X1_399 ( .A(_abc_40344_n589), .B(DATAO_REG_16_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4362) );
  AOI21X1 AOI21X1_4 ( .A(_abc_40344_n689), .B(REG3_REG_5_), .C(REG3_REG_6_), .Y(_abc_40344_n692) );
  AOI21X1 AOI21X1_40 ( .A(n1336), .B(REG3_REG_23_), .C(_abc_40344_n630_1), .Y(_abc_40344_n1581) );
  AOI21X1 AOI21X1_400 ( .A(_abc_40344_n589), .B(DATAO_REG_17_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4364) );
  AOI21X1 AOI21X1_401 ( .A(_abc_40344_n589), .B(DATAO_REG_18_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4366) );
  AOI21X1 AOI21X1_402 ( .A(_abc_40344_n589), .B(DATAO_REG_19_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4368) );
  AOI21X1 AOI21X1_403 ( .A(_abc_40344_n589), .B(DATAO_REG_20_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4370) );
  AOI21X1 AOI21X1_404 ( .A(_abc_40344_n589), .B(DATAO_REG_21_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4372) );
  AOI21X1 AOI21X1_405 ( .A(_abc_40344_n589), .B(DATAO_REG_22_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4374) );
  AOI21X1 AOI21X1_406 ( .A(_abc_40344_n589), .B(DATAO_REG_23_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4376) );
  AOI21X1 AOI21X1_407 ( .A(_abc_40344_n589), .B(DATAO_REG_24_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4378) );
  AOI21X1 AOI21X1_408 ( .A(_abc_40344_n589), .B(DATAO_REG_25_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4380) );
  AOI21X1 AOI21X1_409 ( .A(_abc_40344_n589), .B(DATAO_REG_26_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4382) );
  AOI21X1 AOI21X1_41 ( .A(_abc_40344_n1086), .B(_abc_40344_n1554), .C(_abc_40344_n1582), .Y(_abc_40344_n1583) );
  AOI21X1 AOI21X1_410 ( .A(_abc_40344_n589), .B(DATAO_REG_27_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4384) );
  AOI21X1 AOI21X1_411 ( .A(_abc_40344_n589), .B(DATAO_REG_28_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4386) );
  AOI21X1 AOI21X1_412 ( .A(_abc_40344_n589), .B(DATAO_REG_29_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4388) );
  AOI21X1 AOI21X1_413 ( .A(_abc_40344_n589), .B(DATAO_REG_30_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4390) );
  AOI21X1 AOI21X1_414 ( .A(_abc_40344_n589), .B(DATAO_REG_31_), .C(_abc_40344_n630_1), .Y(_abc_40344_n4392) );
  AOI21X1 AOI21X1_42 ( .A(_abc_40344_n1586), .B(_abc_40344_n1589), .C(_abc_40344_n1590), .Y(_abc_40344_n1591) );
  AOI21X1 AOI21X1_43 ( .A(_abc_40344_n1032), .B(_abc_40344_n1327), .C(_abc_40344_n1594), .Y(_abc_40344_n1595) );
  AOI21X1 AOI21X1_44 ( .A(_abc_40344_n1005), .B(_abc_40344_n1593), .C(_abc_40344_n1596), .Y(_abc_40344_n1597) );
  AOI21X1 AOI21X1_45 ( .A(_abc_40344_n688_1), .B(_abc_40344_n1554), .C(_abc_40344_n1612), .Y(_abc_40344_n1613) );
  AOI21X1 AOI21X1_46 ( .A(_abc_40344_n1032), .B(_abc_40344_n1404), .C(_abc_40344_n1623), .Y(_abc_40344_n1624) );
  AOI21X1 AOI21X1_47 ( .A(_abc_40344_n1005), .B(_abc_40344_n1622), .C(_abc_40344_n1625), .Y(_abc_40344_n1626) );
  AOI21X1 AOI21X1_48 ( .A(REG0_REG_29_), .B(_abc_40344_n673), .C(_abc_40344_n1643), .Y(_abc_40344_n1644) );
  AOI21X1 AOI21X1_49 ( .A(_abc_40344_n1032), .B(_abc_40344_n1649), .C(_abc_40344_n1650), .Y(_abc_40344_n1651) );
  AOI21X1 AOI21X1_5 ( .A(_abc_40344_n637), .B(_abc_40344_n633_1), .C(_abc_40344_n699), .Y(_abc_40344_n700) );
  AOI21X1 AOI21X1_50 ( .A(_abc_40344_n1647), .B(_abc_40344_n1005), .C(_abc_40344_n1652), .Y(_abc_40344_n1653) );
  AOI21X1 AOI21X1_51 ( .A(_abc_40344_n1032), .B(_abc_40344_n1665), .C(_abc_40344_n1666), .Y(_abc_40344_n1667) );
  AOI21X1 AOI21X1_52 ( .A(_abc_40344_n1005), .B(_abc_40344_n1662), .C(_abc_40344_n1668), .Y(_abc_40344_n1669) );
  AOI21X1 AOI21X1_53 ( .A(_abc_40344_n1032), .B(_abc_40344_n856), .C(_abc_40344_n1679), .Y(_abc_40344_n1680) );
  AOI21X1 AOI21X1_54 ( .A(_abc_40344_n1005), .B(_abc_40344_n1677), .C(_abc_40344_n1681), .Y(_abc_40344_n1682) );
  AOI21X1 AOI21X1_55 ( .A(_abc_40344_n1445), .B(_abc_40344_n1453), .C(_abc_40344_n1687), .Y(_abc_40344_n1688) );
  AOI21X1 AOI21X1_56 ( .A(_abc_40344_n1020), .B(_abc_40344_n1111), .C(_abc_40344_n1694), .Y(_abc_40344_n1695) );
  AOI21X1 AOI21X1_57 ( .A(_abc_40344_n1032), .B(_abc_40344_n1434), .C(_abc_40344_n1696), .Y(_abc_40344_n1697) );
  AOI21X1 AOI21X1_58 ( .A(_abc_40344_n1001), .B(_abc_40344_n1436), .C(_abc_40344_n1698), .Y(_abc_40344_n1699) );
  AOI21X1 AOI21X1_59 ( .A(_abc_40344_n1032), .B(_abc_40344_n1308), .C(_abc_40344_n1710), .Y(_abc_40344_n1711) );
  AOI21X1 AOI21X1_6 ( .A(_abc_40344_n556), .B(_abc_40344_n597), .C(_abc_40344_n600_1), .Y(_abc_40344_n703) );
  AOI21X1 AOI21X1_60 ( .A(_abc_40344_n1005), .B(_abc_40344_n1709), .C(_abc_40344_n1712), .Y(_abc_40344_n1713) );
  AOI21X1 AOI21X1_61 ( .A(_abc_40344_n1532), .B(_abc_40344_n1098), .C(_abc_40344_n1476), .Y(_abc_40344_n1720) );
  AOI21X1 AOI21X1_62 ( .A(n1336), .B(REG3_REG_25_), .C(_abc_40344_n630_1), .Y(_abc_40344_n1727) );
  AOI21X1 AOI21X1_63 ( .A(_abc_40344_n1726), .B(_abc_40344_n1554), .C(_abc_40344_n1728), .Y(_abc_40344_n1729) );
  AOI21X1 AOI21X1_64 ( .A(_abc_40344_n1032), .B(_abc_40344_n1153), .C(_abc_40344_n1737), .Y(_abc_40344_n1738) );
  AOI21X1 AOI21X1_65 ( .A(_abc_40344_n1005), .B(_abc_40344_n1736), .C(_abc_40344_n1739), .Y(_abc_40344_n1740) );
  AOI21X1 AOI21X1_66 ( .A(_abc_40344_n1032), .B(_abc_40344_n734), .C(_abc_40344_n1745), .Y(_abc_40344_n1746) );
  AOI21X1 AOI21X1_67 ( .A(_abc_40344_n1005), .B(_abc_40344_n1744), .C(_abc_40344_n1747), .Y(_abc_40344_n1748) );
  AOI21X1 AOI21X1_68 ( .A(_abc_40344_n1395), .B(_abc_40344_n1216), .C(_abc_40344_n1732), .Y(_abc_40344_n1753) );
  AOI21X1 AOI21X1_69 ( .A(_abc_40344_n1032), .B(_abc_40344_n1178), .C(_abc_40344_n1758), .Y(_abc_40344_n1759) );
  AOI21X1 AOI21X1_7 ( .A(_abc_40344_n646), .B(_abc_40344_n625), .C(_abc_40344_n618), .Y(_abc_40344_n718) );
  AOI21X1 AOI21X1_70 ( .A(_abc_40344_n1005), .B(_abc_40344_n1756), .C(_abc_40344_n1760), .Y(_abc_40344_n1761) );
  AOI21X1 AOI21X1_71 ( .A(_abc_40344_n1460), .B(_abc_40344_n1096), .C(_abc_40344_n1763), .Y(_abc_40344_n1764) );
  AOI21X1 AOI21X1_72 ( .A(_abc_40344_n1032), .B(_abc_40344_n1463), .C(_abc_40344_n1768), .Y(_abc_40344_n1769) );
  AOI21X1 AOI21X1_73 ( .A(_abc_40344_n1767), .B(_abc_40344_n1005), .C(_abc_40344_n1770), .Y(_abc_40344_n1771) );
  AOI21X1 AOI21X1_74 ( .A(_abc_40344_n1032), .B(_abc_40344_n777_1), .C(_abc_40344_n1776), .Y(_abc_40344_n1777) );
  AOI21X1 AOI21X1_75 ( .A(_abc_40344_n779), .B(_abc_40344_n1554), .C(_abc_40344_n1779), .Y(_abc_40344_n1780) );
  AOI21X1 AOI21X1_76 ( .A(_abc_40344_n1032), .B(_abc_40344_n1350), .C(_abc_40344_n1789), .Y(_abc_40344_n1790) );
  AOI21X1 AOI21X1_77 ( .A(_abc_40344_n1005), .B(_abc_40344_n1788), .C(_abc_40344_n1791), .Y(_abc_40344_n1792) );
  AOI21X1 AOI21X1_78 ( .A(_abc_40344_n1020), .B(_abc_40344_n1801), .C(_abc_40344_n1802), .Y(_abc_40344_n1803) );
  AOI21X1 AOI21X1_79 ( .A(_abc_40344_n993), .B(_abc_40344_n1800), .C(_abc_40344_n1804), .Y(_abc_40344_n1805) );
  AOI21X1 AOI21X1_8 ( .A(_abc_40344_n725), .B(_abc_40344_n724), .C(_abc_40344_n715), .Y(_abc_40344_n726) );
  AOI21X1 AOI21X1_80 ( .A(_abc_40344_n1032), .B(_abc_40344_n1812), .C(_abc_40344_n1813), .Y(_abc_40344_n1814) );
  AOI21X1 AOI21X1_81 ( .A(_abc_40344_n1005), .B(_abc_40344_n1811), .C(_abc_40344_n1815), .Y(_abc_40344_n1816) );
  AOI21X1 AOI21X1_82 ( .A(_abc_40344_n1032), .B(_abc_40344_n1251), .C(_abc_40344_n1820), .Y(_abc_40344_n1821) );
  AOI21X1 AOI21X1_83 ( .A(_abc_40344_n1005), .B(_abc_40344_n1819), .C(_abc_40344_n1822), .Y(_abc_40344_n1823) );
  AOI21X1 AOI21X1_84 ( .A(_abc_40344_n1267), .B(_abc_40344_n1313), .C(_abc_40344_n1825), .Y(_abc_40344_n1826) );
  AOI21X1 AOI21X1_85 ( .A(_abc_40344_n1571), .B(_abc_40344_n1831), .C(_abc_40344_n1590), .Y(_abc_40344_n1832) );
  AOI21X1 AOI21X1_86 ( .A(_abc_40344_n1032), .B(_abc_40344_n1100), .C(_abc_40344_n1835), .Y(_abc_40344_n1836) );
  AOI21X1 AOI21X1_87 ( .A(_abc_40344_n1005), .B(_abc_40344_n1834), .C(_abc_40344_n1837), .Y(_abc_40344_n1838) );
  AOI21X1 AOI21X1_88 ( .A(_abc_40344_n1032), .B(_abc_40344_n1273), .C(_abc_40344_n1842), .Y(_abc_40344_n1843) );
  AOI21X1 AOI21X1_89 ( .A(_abc_40344_n1005), .B(_abc_40344_n1841), .C(_abc_40344_n1844), .Y(_abc_40344_n1845) );
  AOI21X1 AOI21X1_9 ( .A(_abc_40344_n661), .B(_abc_40344_n664), .C(_abc_40344_n559_1), .Y(_abc_40344_n752) );
  AOI21X1 AOI21X1_90 ( .A(_abc_40344_n1032), .B(_abc_40344_n825), .C(_abc_40344_n1855), .Y(_abc_40344_n1856) );
  AOI21X1 AOI21X1_91 ( .A(_abc_40344_n1005), .B(_abc_40344_n1853), .C(_abc_40344_n1857), .Y(_abc_40344_n1858) );
  AOI21X1 AOI21X1_92 ( .A(_abc_40344_n1616), .B(_abc_40344_n1860), .C(_abc_40344_n1590), .Y(_abc_40344_n1861) );
  AOI21X1 AOI21X1_93 ( .A(_abc_40344_n1032), .B(_abc_40344_n1124), .C(_abc_40344_n1864), .Y(_abc_40344_n1865) );
  AOI21X1 AOI21X1_94 ( .A(_abc_40344_n1005), .B(_abc_40344_n1863), .C(_abc_40344_n1866), .Y(_abc_40344_n1867) );
  AOI21X1 AOI21X1_95 ( .A(_abc_40344_n1032), .B(_abc_40344_n714), .C(_abc_40344_n1873), .Y(_abc_40344_n1874) );
  AOI21X1 AOI21X1_96 ( .A(_abc_40344_n1005), .B(_abc_40344_n1871), .C(_abc_40344_n1875), .Y(_abc_40344_n1876) );
  AOI21X1 AOI21X1_97 ( .A(_abc_40344_n1717), .B(_abc_40344_n1878), .C(_abc_40344_n1880), .Y(_abc_40344_n1881) );
  AOI21X1 AOI21X1_98 ( .A(_abc_40344_n1032), .B(_abc_40344_n1495), .C(_abc_40344_n1889), .Y(_abc_40344_n1890) );
  AOI21X1 AOI21X1_99 ( .A(_abc_40344_n1886), .B(_abc_40344_n1005), .C(_abc_40344_n1891), .Y(_abc_40344_n1892) );
  AOI22X1 AOI22X1_1 ( .A(_abc_40344_n574), .B(_abc_40344_n596_1), .C(IR_REG_28_), .D(_abc_40344_n598), .Y(_abc_40344_n599) );
  AOI22X1 AOI22X1_10 ( .A(_abc_40344_n601), .B(_abc_40344_n704), .C(_abc_40344_n605), .D(_abc_40344_n609), .Y(_abc_40344_n705_1) );
  AOI22X1 AOI22X1_100 ( .A(_abc_40344_n1418), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1414), .Y(_abc_40344_n2331_1) );
  AOI22X1 AOI22X1_101 ( .A(_abc_40344_n1421_1), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1429), .Y(_abc_40344_n2338) );
  AOI22X1 AOI22X1_102 ( .A(_abc_40344_n1433), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1440), .Y(_abc_40344_n2342) );
  AOI22X1 AOI22X1_103 ( .A(_abc_40344_n2162), .B(_abc_40344_n1434), .C(_abc_40344_n2165), .D(_abc_40344_n1441), .Y(_abc_40344_n2344) );
  AOI22X1 AOI22X1_104 ( .A(_abc_40344_n1099), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1110), .Y(_abc_40344_n2352) );
  AOI22X1 AOI22X1_105 ( .A(_abc_40344_n2343), .B(_abc_40344_n2345), .C(_abc_40344_n2351), .D(_abc_40344_n2353), .Y(_abc_40344_n2354) );
  AOI22X1 AOI22X1_106 ( .A(_abc_40344_n1083), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1090_1), .Y(_abc_40344_n2359) );
  AOI22X1 AOI22X1_107 ( .A(_abc_40344_n2162), .B(_abc_40344_n1463), .C(_abc_40344_n586), .D(_abc_40344_n1091), .Y(_abc_40344_n2364) );
  AOI22X1 AOI22X1_108 ( .A(_abc_40344_n1462), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1577), .Y(_abc_40344_n2367) );
  AOI22X1 AOI22X1_109 ( .A(_abc_40344_n2162), .B(_abc_40344_n1491), .C(_abc_40344_n586), .D(_abc_40344_n1471), .Y(_abc_40344_n2370) );
  AOI22X1 AOI22X1_11 ( .A(_abc_40344_n650), .B(_abc_40344_n698), .C(_abc_40344_n700), .D(_abc_40344_n714), .Y(_abc_40344_n715) );
  AOI22X1 AOI22X1_110 ( .A(_abc_40344_n2162), .B(_abc_40344_n1495), .C(_abc_40344_n586), .D(_abc_40344_n1488), .Y(_abc_40344_n2376) );
  AOI22X1 AOI22X1_111 ( .A(_abc_40344_n1494), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1506), .Y(_abc_40344_n2378) );
  AOI22X1 AOI22X1_112 ( .A(_abc_40344_n2371), .B(_abc_40344_n2372), .C(_abc_40344_n2377), .D(_abc_40344_n2379), .Y(_abc_40344_n2380_1) );
  AOI22X1 AOI22X1_113 ( .A(_abc_40344_n1040), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1074), .Y(_abc_40344_n2382) );
  AOI22X1 AOI22X1_114 ( .A(_abc_40344_n2162), .B(_abc_40344_n1076), .C(_abc_40344_n2165), .D(_abc_40344_n1073), .Y(_abc_40344_n2384) );
  AOI22X1 AOI22X1_115 ( .A(_abc_40344_n2162), .B(_abc_40344_n1649), .C(_abc_40344_n586), .D(_abc_40344_n1073), .Y(_abc_40344_n2389_1) );
  AOI22X1 AOI22X1_116 ( .A(_abc_40344_n2383), .B(_abc_40344_n2385), .C(_abc_40344_n2390), .D(_abc_40344_n2392), .Y(_abc_40344_n2393) );
  AOI22X1 AOI22X1_117 ( .A(_abc_40344_n2162), .B(_abc_40344_n2394), .C(_abc_40344_n2165), .D(_abc_40344_n1645), .Y(_abc_40344_n2395) );
  AOI22X1 AOI22X1_118 ( .A(_abc_40344_n2165), .B(_abc_40344_n1926), .C(_abc_40344_n2173), .D(_abc_40344_n1646), .Y(_abc_40344_n2397) );
  AOI22X1 AOI22X1_119 ( .A(_abc_40344_n2096), .B(_abc_40344_n2165), .C(_abc_40344_n2162), .D(_abc_40344_n2401), .Y(_abc_40344_n2402) );
  AOI22X1 AOI22X1_12 ( .A(_abc_40344_n637), .B(_abc_40344_n633_1), .C(_abc_40344_n647), .D(_abc_40344_n721), .Y(_abc_40344_n722) );
  AOI22X1 AOI22X1_120 ( .A(_abc_40344_n2165), .B(_abc_40344_n2401), .C(_abc_40344_n2096), .D(_abc_40344_n2404), .Y(_abc_40344_n2405) );
  AOI22X1 AOI22X1_121 ( .A(_abc_40344_n2403), .B(_abc_40344_n2405), .C(_abc_40344_n2398), .D(_abc_40344_n2396), .Y(_abc_40344_n2406) );
  AOI22X1 AOI22X1_122 ( .A(_abc_40344_n2101), .B(_abc_40344_n2162), .C(_abc_40344_n2165), .D(_abc_40344_n1917), .Y(_abc_40344_n2413) );
  AOI22X1 AOI22X1_123 ( .A(_abc_40344_n1021), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1994), .Y(_abc_40344_n2422) );
  AOI22X1 AOI22X1_124 ( .A(_abc_40344_n2421), .B(_abc_40344_n2422), .C(_abc_40344_n2424), .D(_abc_40344_n2423), .Y(_abc_40344_n2425) );
  AOI22X1 AOI22X1_125 ( .A(_abc_40344_n2426), .B(_abc_40344_n2427), .C(_abc_40344_n2235), .D(_abc_40344_n2236), .Y(_abc_40344_n2428_1) );
  AOI22X1 AOI22X1_126 ( .A(_abc_40344_n863), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n869), .Y(_abc_40344_n2434) );
  AOI22X1 AOI22X1_127 ( .A(_abc_40344_n2435_1), .B(_abc_40344_n2224), .C(_abc_40344_n2434), .D(_abc_40344_n2433), .Y(_abc_40344_n2436) );
  AOI22X1 AOI22X1_128 ( .A(_abc_40344_n2416_1), .B(_abc_40344_n645), .C(_abc_40344_n2562), .D(_abc_40344_n2468), .Y(_abc_40344_n2563) );
  AOI22X1 AOI22X1_129 ( .A(_abc_40344_n602), .B(_abc_40344_n712), .C(_abc_40344_n2666_1), .D(_abc_40344_n2789), .Y(_abc_40344_n2790) );
  AOI22X1 AOI22X1_13 ( .A(_abc_40344_n698), .B(_abc_40344_n700), .C(_abc_40344_n722), .D(_abc_40344_n714), .Y(_abc_40344_n723) );
  AOI22X1 AOI22X1_130 ( .A(ADDR_REG_6_), .B(_abc_40344_n2673), .C(_abc_40344_n2792), .D(_abc_40344_n2791), .Y(_abc_40344_n2793) );
  AOI22X1 AOI22X1_131 ( .A(_abc_40344_n602), .B(_abc_40344_n1372), .C(_abc_40344_n2666_1), .D(_abc_40344_n2824), .Y(_abc_40344_n2825) );
  AOI22X1 AOI22X1_132 ( .A(_abc_40344_n3040), .B(_abc_40344_n3045), .C(_abc_40344_n3043), .D(_abc_40344_n3038), .Y(_abc_40344_n3046) );
  AOI22X1 AOI22X1_133 ( .A(_abc_40344_n3124), .B(_abc_40344_n3131), .C(_abc_40344_n3127), .D(_abc_40344_n3134), .Y(_abc_40344_n3135) );
  AOI22X1 AOI22X1_134 ( .A(_abc_40344_n3188), .B(_abc_40344_n3190), .C(_abc_40344_n3177), .D(_abc_40344_n3186), .Y(_abc_40344_n3191) );
  AOI22X1 AOI22X1_135 ( .A(_abc_40344_n1030_1), .B(_abc_40344_n1541), .C(_abc_40344_n3068), .D(_abc_40344_n3239), .Y(_abc_40344_n3240) );
  AOI22X1 AOI22X1_136 ( .A(_abc_40344_n1507_1), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3246), .Y(_abc_40344_n3247) );
  AOI22X1 AOI22X1_137 ( .A(_abc_40344_n1488), .B(_abc_40344_n3220), .C(_abc_40344_n3227), .D(_abc_40344_n3268), .Y(_abc_40344_n3269_1) );
  AOI22X1 AOI22X1_138 ( .A(_abc_40344_n1471), .B(_abc_40344_n3220), .C(_abc_40344_n3284), .D(_abc_40344_n3285), .Y(_abc_40344_n3286) );
  AOI22X1 AOI22X1_139 ( .A(_abc_40344_n1030_1), .B(_abc_40344_n1726), .C(_abc_40344_n3068), .D(_abc_40344_n3291), .Y(_abc_40344_n3292) );
  AOI22X1 AOI22X1_14 ( .A(REG2_REG_5_), .B(_abc_40344_n695), .C(REG0_REG_5_), .D(_abc_40344_n673), .Y(_abc_40344_n735) );
  AOI22X1 AOI22X1_140 ( .A(_abc_40344_n1091), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3296), .Y(_abc_40344_n3297) );
  AOI22X1 AOI22X1_141 ( .A(_abc_40344_n995), .B(_abc_40344_n1463), .C(_abc_40344_n3103), .D(_abc_40344_n1488), .Y(_abc_40344_n3343) );
  AOI22X1 AOI22X1_142 ( .A(_abc_40344_n1111), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3351), .Y(_abc_40344_n3352) );
  AOI22X1 AOI22X1_143 ( .A(_abc_40344_n1186), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3459), .Y(_abc_40344_n3463) );
  AOI22X1 AOI22X1_144 ( .A(REG2_REG_17_), .B(_abc_40344_n3067), .C(_abc_40344_n1178), .D(_abc_40344_n3110), .Y(_abc_40344_n3496) );
  AOI22X1 AOI22X1_145 ( .A(_abc_40344_n1210), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3500), .Y(_abc_40344_n3501) );
  AOI22X1 AOI22X1_146 ( .A(_abc_40344_n1234), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3520), .Y(_abc_40344_n3521) );
  AOI22X1 AOI22X1_147 ( .A(_abc_40344_n1260), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3541), .Y(_abc_40344_n3542) );
  AOI22X1 AOI22X1_148 ( .A(_abc_40344_n1309), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3564), .Y(_abc_40344_n3565) );
  AOI22X1 AOI22X1_149 ( .A(_abc_40344_n1030_1), .B(_abc_40344_n1256), .C(_abc_40344_n1234), .D(_abc_40344_n3233), .Y(_abc_40344_n3568) );
  AOI22X1 AOI22X1_15 ( .A(_abc_40344_n650), .B(_abc_40344_n742), .C(_abc_40344_n700), .D(_abc_40344_n734), .Y(_abc_40344_n743) );
  AOI22X1 AOI22X1_150 ( .A(_abc_40344_n1285), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3581_1), .Y(_abc_40344_n3582) );
  AOI22X1 AOI22X1_151 ( .A(_abc_40344_n1335), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3594), .Y(_abc_40344_n3595) );
  AOI22X1 AOI22X1_152 ( .A(_abc_40344_n1030_1), .B(_abc_40344_n1278), .C(_abc_40344_n3602), .D(_abc_40344_n3066), .Y(_abc_40344_n3603) );
  AOI22X1 AOI22X1_153 ( .A(_abc_40344_n1273), .B(_abc_40344_n3110), .C(_abc_40344_n3068), .D(_abc_40344_n3605), .Y(_abc_40344_n3606) );
  AOI22X1 AOI22X1_154 ( .A(_abc_40344_n1362), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3619), .Y(_abc_40344_n3620) );
  AOI22X1 AOI22X1_155 ( .A(_abc_40344_n1285), .B(_abc_40344_n3103), .C(_abc_40344_n995), .D(_abc_40344_n1327), .Y(_abc_40344_n3627) );
  AOI22X1 AOI22X1_156 ( .A(_abc_40344_n1019), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3640), .Y(_abc_40344_n3641) );
  AOI22X1 AOI22X1_157 ( .A(_abc_40344_n915_1), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3655), .Y(_abc_40344_n3656) );
  AOI22X1 AOI22X1_158 ( .A(_abc_40344_n1362), .B(_abc_40344_n3233), .C(_abc_40344_n3068), .D(_abc_40344_n3665), .Y(_abc_40344_n3666) );
  AOI22X1 AOI22X1_159 ( .A(_abc_40344_n698), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3675), .Y(_abc_40344_n3676) );
  AOI22X1 AOI22X1_16 ( .A(_abc_40344_n685_1), .B(_abc_40344_n779), .C(REG2_REG_4_), .D(_abc_40344_n695), .Y(_abc_40344_n780_1) );
  AOI22X1 AOI22X1_160 ( .A(_abc_40344_n742), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3689), .Y(_abc_40344_n3690) );
  AOI22X1 AOI22X1_161 ( .A(_abc_40344_n785), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3707), .Y(_abc_40344_n3708) );
  AOI22X1 AOI22X1_162 ( .A(_abc_40344_n3103), .B(_abc_40344_n698), .C(_abc_40344_n995), .D(_abc_40344_n734), .Y(_abc_40344_n3713) );
  AOI22X1 AOI22X1_163 ( .A(_abc_40344_n779), .B(_abc_40344_n1030_1), .C(REG2_REG_4_), .D(_abc_40344_n3067), .Y(_abc_40344_n3737) );
  AOI22X1 AOI22X1_164 ( .A(_abc_40344_n3103), .B(_abc_40344_n785), .C(_abc_40344_n995), .D(_abc_40344_n813), .Y(_abc_40344_n3739) );
  AOI22X1 AOI22X1_165 ( .A(_abc_40344_n829_1), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3745), .Y(_abc_40344_n3746) );
  AOI22X1 AOI22X1_166 ( .A(_abc_40344_n688_1), .B(_abc_40344_n1030_1), .C(REG2_REG_3_), .D(_abc_40344_n3067), .Y(_abc_40344_n3754) );
  AOI22X1 AOI22X1_167 ( .A(_abc_40344_n864), .B(_abc_40344_n3220), .C(_abc_40344_n3223), .D(_abc_40344_n3759), .Y(_abc_40344_n3760) );
  AOI22X1 AOI22X1_168 ( .A(_abc_40344_n3103), .B(_abc_40344_n808), .C(_abc_40344_n995), .D(_abc_40344_n825), .Y(_abc_40344_n3762) );
  AOI22X1 AOI22X1_169 ( .A(_abc_40344_n3103), .B(_abc_40344_n829_1), .C(_abc_40344_n995), .D(_abc_40344_n856), .Y(_abc_40344_n3775_1) );
  AOI22X1 AOI22X1_17 ( .A(_abc_40344_n650), .B(_abc_40344_n785), .C(_abc_40344_n700), .D(_abc_40344_n777_1), .Y(_abc_40344_n786) );
  AOI22X1 AOI22X1_170 ( .A(REG3_REG_0_), .B(_abc_40344_n1030_1), .C(REG2_REG_0_), .D(_abc_40344_n3067), .Y(_abc_40344_n3792_1) );
  AOI22X1 AOI22X1_171 ( .A(DATAI_28_), .B(n1336), .C(IR_REG_28_), .D(_abc_40344_n3860), .Y(_abc_40344_n3872) );
  AOI22X1 AOI22X1_172 ( .A(DATAI_19_), .B(n1336), .C(IR_REG_19_), .D(_abc_40344_n3860), .Y(_abc_40344_n3912) );
  AOI22X1 AOI22X1_173 ( .A(DATAI_12_), .B(n1336), .C(IR_REG_12_), .D(_abc_40344_n3860), .Y(_abc_40344_n3945) );
  AOI22X1 AOI22X1_174 ( .A(_abc_40344_n4016), .B(_abc_40344_n4017), .C(_abc_40344_n4015), .D(_abc_40344_n2650_1), .Y(_abc_40344_n4018) );
  AOI22X1 AOI22X1_175 ( .A(_abc_40344_n3725), .B(_abc_40344_n3718), .C(_abc_40344_n4048), .D(_abc_40344_n3707), .Y(_abc_40344_n4070_1) );
  AOI22X1 AOI22X1_176 ( .A(_abc_40344_n1234), .B(_abc_40344_n3103), .C(_abc_40344_n995), .D(_abc_40344_n1251), .Y(_abc_40344_n4117) );
  AOI22X1 AOI22X1_177 ( .A(_abc_40344_n995), .B(_abc_40344_n1201), .C(_abc_40344_n3725), .D(_abc_40344_n3530), .Y(_abc_40344_n4132) );
  AOI22X1 AOI22X1_178 ( .A(_abc_40344_n995), .B(_abc_40344_n1153), .C(_abc_40344_n3725), .D(_abc_40344_n3510), .Y(_abc_40344_n4139) );
  AOI22X1 AOI22X1_179 ( .A(_abc_40344_n995), .B(_abc_40344_n1100), .C(_abc_40344_n3103), .D(_abc_40344_n1091), .Y(_abc_40344_n4176) );
  AOI22X1 AOI22X1_18 ( .A(_abc_40344_n798), .B(_abc_40344_n803), .C(_abc_40344_n793), .D(_abc_40344_n792), .Y(_abc_40344_n804) );
  AOI22X1 AOI22X1_180 ( .A(_abc_40344_n995), .B(_abc_40344_n1084), .C(_abc_40344_n3103), .D(_abc_40344_n1471), .Y(_abc_40344_n4184) );
  AOI22X1 AOI22X1_19 ( .A(_abc_40344_n685_1), .B(_abc_40344_n688_1), .C(REG2_REG_3_), .D(_abc_40344_n695), .Y(_abc_40344_n807_1) );
  AOI22X1 AOI22X1_2 ( .A(_abc_40344_n562), .B(_abc_40344_n564), .C(_abc_40344_n636), .D(_abc_40344_n635), .Y(_abc_40344_n637) );
  AOI22X1 AOI22X1_20 ( .A(_abc_40344_n700), .B(_abc_40344_n808), .C(_abc_40344_n722), .D(_abc_40344_n813), .Y(_abc_40344_n814) );
  AOI22X1 AOI22X1_21 ( .A(_abc_40344_n650), .B(_abc_40344_n808), .C(_abc_40344_n700), .D(_abc_40344_n813), .Y(_abc_40344_n818_1) );
  AOI22X1 AOI22X1_22 ( .A(REG3_REG_2_), .B(_abc_40344_n685_1), .C(REG0_REG_2_), .D(_abc_40344_n673), .Y(_abc_40344_n828) );
  AOI22X1 AOI22X1_23 ( .A(_abc_40344_n650), .B(_abc_40344_n829_1), .C(_abc_40344_n700), .D(_abc_40344_n825), .Y(_abc_40344_n830) );
  AOI22X1 AOI22X1_24 ( .A(_abc_40344_n700), .B(_abc_40344_n829_1), .C(_abc_40344_n722), .D(_abc_40344_n825), .Y(_abc_40344_n832) );
  AOI22X1 AOI22X1_25 ( .A(_abc_40344_n834), .B(_abc_40344_n824_1), .C(_abc_40344_n793), .D(_abc_40344_n792), .Y(_abc_40344_n835_1) );
  AOI22X1 AOI22X1_26 ( .A(_abc_40344_n864), .B(_abc_40344_n650), .C(_abc_40344_n700), .D(_abc_40344_n856), .Y(_abc_40344_n865) );
  AOI22X1 AOI22X1_27 ( .A(_abc_40344_n864), .B(_abc_40344_n700), .C(_abc_40344_n722), .D(_abc_40344_n856), .Y(_abc_40344_n866_1) );
  AOI22X1 AOI22X1_28 ( .A(_abc_40344_n581), .B(REG1_REG_0_), .C(_abc_40344_n700), .D(_abc_40344_n887), .Y(_abc_40344_n888) );
  AOI22X1 AOI22X1_29 ( .A(_abc_40344_n581), .B(IR_REG_0_), .C(_abc_40344_n887), .D(_abc_40344_n650), .Y(_abc_40344_n891) );
  AOI22X1 AOI22X1_3 ( .A(_abc_40344_n637), .B(_abc_40344_n633_1), .C(_abc_40344_n647), .D(_abc_40344_n649_1), .Y(_abc_40344_n650) );
  AOI22X1 AOI22X1_30 ( .A(_abc_40344_n880), .B(_abc_40344_n888), .C(_abc_40344_n890), .D(_abc_40344_n891), .Y(_abc_40344_n892) );
  AOI22X1 AOI22X1_31 ( .A(_abc_40344_n895), .B(_abc_40344_n830), .C(_abc_40344_n816), .D(_abc_40344_n818_1), .Y(_abc_40344_n896) );
  AOI22X1 AOI22X1_32 ( .A(_abc_40344_n685_1), .B(_abc_40344_n912), .C(REG0_REG_7_), .D(_abc_40344_n673), .Y(_abc_40344_n913) );
  AOI22X1 AOI22X1_33 ( .A(REG2_REG_7_), .B(_abc_40344_n695), .C(REG1_REG_7_), .D(_abc_40344_n696), .Y(_abc_40344_n914) );
  AOI22X1 AOI22X1_34 ( .A(_abc_40344_n650), .B(_abc_40344_n915_1), .C(_abc_40344_n700), .D(_abc_40344_n908), .Y(_abc_40344_n916) );
  AOI22X1 AOI22X1_35 ( .A(_abc_40344_n700), .B(_abc_40344_n915_1), .C(_abc_40344_n722), .D(_abc_40344_n908), .Y(_abc_40344_n930) );
  AOI22X1 AOI22X1_36 ( .A(STATE_REG), .B(_abc_40344_n999), .C(_abc_40344_n997), .D(_abc_40344_n983), .Y(_abc_40344_n1000) );
  AOI22X1 AOI22X1_37 ( .A(_abc_40344_n722), .B(_abc_40344_n1076), .C(_abc_40344_n700), .D(_abc_40344_n1073), .Y(_abc_40344_n1077) );
  AOI22X1 AOI22X1_38 ( .A(_abc_40344_n673), .B(REG0_REG_23_), .C(REG1_REG_23_), .D(_abc_40344_n696), .Y(_abc_40344_n1088) );
  AOI22X1 AOI22X1_39 ( .A(_abc_40344_n700), .B(_abc_40344_n1084), .C(_abc_40344_n650), .D(_abc_40344_n1091), .Y(_abc_40344_n1092) );
  AOI22X1 AOI22X1_4 ( .A(_abc_40344_n668_1), .B(_abc_40344_n672), .C(_abc_40344_n652_1), .D(_abc_40344_n666_1), .Y(_abc_40344_n673) );
  AOI22X1 AOI22X1_40 ( .A(_abc_40344_n700), .B(_abc_40344_n1100), .C(_abc_40344_n650), .D(_abc_40344_n1111), .Y(_abc_40344_n1112) );
  AOI22X1 AOI22X1_41 ( .A(_abc_40344_n700), .B(_abc_40344_n1124), .C(_abc_40344_n650), .D(_abc_40344_n1134), .Y(_abc_40344_n1135_1) );
  AOI22X1 AOI22X1_42 ( .A(_abc_40344_n700), .B(_abc_40344_n1153), .C(_abc_40344_n650), .D(_abc_40344_n1168), .Y(_abc_40344_n1169) );
  AOI22X1 AOI22X1_43 ( .A(_abc_40344_n700), .B(_abc_40344_n1178), .C(_abc_40344_n650), .D(_abc_40344_n1186), .Y(_abc_40344_n1187) );
  AOI22X1 AOI22X1_44 ( .A(_abc_40344_n722), .B(_abc_40344_n1178), .C(_abc_40344_n700), .D(_abc_40344_n1186), .Y(_abc_40344_n1189) );
  AOI22X1 AOI22X1_45 ( .A(_abc_40344_n650), .B(_abc_40344_n1210), .C(_abc_40344_n700), .D(_abc_40344_n1201), .Y(_abc_40344_n1211) );
  AOI22X1 AOI22X1_46 ( .A(_abc_40344_n650), .B(_abc_40344_n1234), .C(_abc_40344_n700), .D(_abc_40344_n1224), .Y(_abc_40344_n1235) );
  AOI22X1 AOI22X1_47 ( .A(_abc_40344_n700), .B(_abc_40344_n1234), .C(_abc_40344_n722), .D(_abc_40344_n1224), .Y(_abc_40344_n1236) );
  AOI22X1 AOI22X1_48 ( .A(_abc_40344_n650), .B(_abc_40344_n1260), .C(_abc_40344_n700), .D(_abc_40344_n1251), .Y(_abc_40344_n1261) );
  AOI22X1 AOI22X1_49 ( .A(_abc_40344_n650), .B(_abc_40344_n1285), .C(_abc_40344_n700), .D(_abc_40344_n1273), .Y(_abc_40344_n1286) );
  AOI22X1 AOI22X1_5 ( .A(_abc_40344_n683_1), .B(_abc_40344_n684), .C(_abc_40344_n675), .D(_abc_40344_n674_1), .Y(_abc_40344_n685_1) );
  AOI22X1 AOI22X1_50 ( .A(_abc_40344_n700), .B(_abc_40344_n1285), .C(_abc_40344_n722), .D(_abc_40344_n1273), .Y(_abc_40344_n1287) );
  AOI22X1 AOI22X1_51 ( .A(_abc_40344_n700), .B(_abc_40344_n1309), .C(_abc_40344_n722), .D(_abc_40344_n1308), .Y(_abc_40344_n1310) );
  AOI22X1 AOI22X1_52 ( .A(_abc_40344_n650), .B(_abc_40344_n1335), .C(_abc_40344_n700), .D(_abc_40344_n1327), .Y(_abc_40344_n1336) );
  AOI22X1 AOI22X1_53 ( .A(_abc_40344_n700), .B(_abc_40344_n1335), .C(_abc_40344_n722), .D(_abc_40344_n1327), .Y(_abc_40344_n1337) );
  AOI22X1 AOI22X1_54 ( .A(_abc_40344_n1320), .B(_abc_40344_n1339), .C(_abc_40344_n1267), .D(_abc_40344_n1316), .Y(_abc_40344_n1340) );
  AOI22X1 AOI22X1_55 ( .A(_abc_40344_n1362), .B(_abc_40344_n650), .C(_abc_40344_n700), .D(_abc_40344_n1350), .Y(_abc_40344_n1363) );
  AOI22X1 AOI22X1_56 ( .A(_abc_40344_n1362), .B(_abc_40344_n700), .C(_abc_40344_n722), .D(_abc_40344_n1350), .Y(_abc_40344_n1365) );
  AOI22X1 AOI22X1_57 ( .A(_abc_40344_n700), .B(_abc_40344_n1404), .C(_abc_40344_n650), .D(_abc_40344_n1415), .Y(_abc_40344_n1416) );
  AOI22X1 AOI22X1_58 ( .A(REG2_REG_21_), .B(_abc_40344_n695), .C(REG1_REG_21_), .D(_abc_40344_n696), .Y(_abc_40344_n1438) );
  AOI22X1 AOI22X1_59 ( .A(_abc_40344_n700), .B(_abc_40344_n1434), .C(_abc_40344_n650), .D(_abc_40344_n1441), .Y(_abc_40344_n1442) );
  AOI22X1 AOI22X1_6 ( .A(_abc_40344_n685_1), .B(_abc_40344_n693), .C(REG0_REG_6_), .D(_abc_40344_n673), .Y(_abc_40344_n694_1) );
  AOI22X1 AOI22X1_60 ( .A(_abc_40344_n700), .B(_abc_40344_n1463), .C(_abc_40344_n650), .D(_abc_40344_n1471), .Y(_abc_40344_n1472) );
  AOI22X1 AOI22X1_61 ( .A(_abc_40344_n722), .B(_abc_40344_n1463), .C(_abc_40344_n700), .D(_abc_40344_n1471), .Y(_abc_40344_n1474) );
  AOI22X1 AOI22X1_62 ( .A(_abc_40344_n722), .B(_abc_40344_n1491), .C(_abc_40344_n700), .D(_abc_40344_n1488), .Y(_abc_40344_n1492) );
  AOI22X1 AOI22X1_63 ( .A(_abc_40344_n700), .B(_abc_40344_n1495), .C(_abc_40344_n650), .D(_abc_40344_n1507_1), .Y(_abc_40344_n1508_1) );
  AOI22X1 AOI22X1_64 ( .A(_abc_40344_n1629), .B(_abc_40344_n1635), .C(_abc_40344_n1638), .D(_abc_40344_n1637), .Y(_abc_40344_n1639) );
  AOI22X1 AOI22X1_65 ( .A(REG3_REG_1_), .B(_abc_40344_n983), .C(_abc_40344_n829_1), .D(_abc_40344_n1020), .Y(_abc_40344_n1676) );
  AOI22X1 AOI22X1_66 ( .A(_abc_40344_n1020), .B(_abc_40344_n742), .C(_abc_40344_n808), .D(_abc_40344_n1022), .Y(_abc_40344_n1778) );
  AOI22X1 AOI22X1_67 ( .A(_abc_40344_n983), .B(_abc_40344_n1278), .C(_abc_40344_n1309), .D(_abc_40344_n1020), .Y(_abc_40344_n1840) );
  AOI22X1 AOI22X1_68 ( .A(_abc_40344_n2034), .B(_abc_40344_n2070), .C(_abc_40344_n2047), .D(_abc_40344_n2067), .Y(_abc_40344_n2071) );
  AOI22X1 AOI22X1_69 ( .A(_abc_40344_n2115), .B(_abc_40344_n2120), .C(_abc_40344_n2012), .D(_abc_40344_n2123), .Y(_abc_40344_n2124) );
  AOI22X1 AOI22X1_7 ( .A(_abc_40344_n674_1), .B(_abc_40344_n675), .C(_abc_40344_n668_1), .D(_abc_40344_n672), .Y(_abc_40344_n695) );
  AOI22X1 AOI22X1_70 ( .A(_abc_40344_n2086), .B(_abc_40344_n2150), .C(_abc_40344_n1978), .D(_abc_40344_n2153), .Y(_abc_40344_n2154) );
  AOI22X1 AOI22X1_71 ( .A(_abc_40344_n624), .B(_abc_40344_n2159), .C(_abc_40344_n2160), .D(_abc_40344_n639_1), .Y(_abc_40344_n2161) );
  AOI22X1 AOI22X1_72 ( .A(_abc_40344_n808), .B(_abc_40344_n2165), .C(_abc_40344_n586), .D(_abc_40344_n829_1), .Y(_abc_40344_n2166) );
  AOI22X1 AOI22X1_73 ( .A(_abc_40344_n785), .B(_abc_40344_n2165), .C(_abc_40344_n586), .D(_abc_40344_n808), .Y(_abc_40344_n2171) );
  AOI22X1 AOI22X1_74 ( .A(_abc_40344_n2170), .B(_abc_40344_n2171), .C(_abc_40344_n2174), .D(_abc_40344_n2177), .Y(_abc_40344_n2178) );
  AOI22X1 AOI22X1_75 ( .A(_abc_40344_n698), .B(_abc_40344_n2165), .C(_abc_40344_n586), .D(_abc_40344_n742), .Y(_abc_40344_n2182) );
  AOI22X1 AOI22X1_76 ( .A(_abc_40344_n586), .B(_abc_40344_n785), .C(_abc_40344_n2165), .D(_abc_40344_n742), .Y(_abc_40344_n2185) );
  AOI22X1 AOI22X1_77 ( .A(_abc_40344_n915_1), .B(_abc_40344_n2165), .C(_abc_40344_n586), .D(_abc_40344_n698), .Y(_abc_40344_n2193) );
  AOI22X1 AOI22X1_78 ( .A(_abc_40344_n809), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1609), .Y(_abc_40344_n2210) );
  AOI22X1 AOI22X1_79 ( .A(_abc_40344_n841), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n2022), .Y(_abc_40344_n2216) );
  AOI22X1 AOI22X1_8 ( .A(_abc_40344_n683_1), .B(_abc_40344_n684), .C(_abc_40344_n652_1), .D(_abc_40344_n666_1), .Y(_abc_40344_n696) );
  AOI22X1 AOI22X1_80 ( .A(_abc_40344_n2228), .B(_abc_40344_n2229), .C(_abc_40344_n2220), .D(_abc_40344_n2221), .Y(_abc_40344_n2230) );
  AOI22X1 AOI22X1_81 ( .A(_abc_40344_n2215), .B(_abc_40344_n2216), .C(_abc_40344_n2230), .D(_abc_40344_n2226), .Y(_abc_40344_n2231) );
  AOI22X1 AOI22X1_82 ( .A(_abc_40344_n927_1), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n919), .Y(_abc_40344_n2236) );
  AOI22X1 AOI22X1_83 ( .A(_abc_40344_n1787), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1969), .Y(_abc_40344_n2242) );
  AOI22X1 AOI22X1_84 ( .A(_abc_40344_n1361), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1906), .Y(_abc_40344_n2247) );
  AOI22X1 AOI22X1_85 ( .A(_abc_40344_n1018), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1375), .Y(_abc_40344_n2252) );
  AOI22X1 AOI22X1_86 ( .A(_abc_40344_n2188), .B(_abc_40344_n2257), .C(_abc_40344_n2185), .D(_abc_40344_n2256), .Y(_abc_40344_n2258) );
  AOI22X1 AOI22X1_87 ( .A(_abc_40344_n1259), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1264), .Y(_abc_40344_n2276) );
  AOI22X1 AOI22X1_88 ( .A(_abc_40344_n1305), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1295), .Y(_abc_40344_n2277_1) );
  AOI22X1 AOI22X1_89 ( .A(_abc_40344_n2275), .B(_abc_40344_n2276), .C(_abc_40344_n2279), .D(_abc_40344_n2277_1), .Y(_abc_40344_n2280) );
  AOI22X1 AOI22X1_9 ( .A(REG2_REG_6_), .B(_abc_40344_n695), .C(REG1_REG_6_), .D(_abc_40344_n696), .Y(_abc_40344_n697) );
  AOI22X1 AOI22X1_90 ( .A(_abc_40344_n1284), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1973), .Y(_abc_40344_n2281) );
  AOI22X1 AOI22X1_91 ( .A(_abc_40344_n2241), .B(_abc_40344_n2242), .C(_abc_40344_n2283), .D(_abc_40344_n2281), .Y(_abc_40344_n2284) );
  AOI22X1 AOI22X1_92 ( .A(_abc_40344_n586), .B(_abc_40344_n1260), .C(_abc_40344_n2165), .D(_abc_40344_n1234), .Y(_abc_40344_n2294) );
  AOI22X1 AOI22X1_93 ( .A(_abc_40344_n2290), .B(_abc_40344_n2291), .C(_abc_40344_n2296), .D(_abc_40344_n2295), .Y(_abc_40344_n2297) );
  AOI22X1 AOI22X1_94 ( .A(_abc_40344_n1209_1), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1200), .Y(_abc_40344_n2304) );
  AOI22X1 AOI22X1_95 ( .A(_abc_40344_n1152_1), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1167), .Y(_abc_40344_n2313) );
  AOI22X1 AOI22X1_96 ( .A(_abc_40344_n2303), .B(_abc_40344_n2305), .C(_abc_40344_n2314_1), .D(_abc_40344_n2312), .Y(_abc_40344_n2315) );
  AOI22X1 AOI22X1_97 ( .A(_abc_40344_n1185), .B(_abc_40344_n2173), .C(_abc_40344_n2165), .D(_abc_40344_n1949), .Y(_abc_40344_n2319) );
  AOI22X1 AOI22X1_98 ( .A(_abc_40344_n2311), .B(_abc_40344_n2313), .C(_abc_40344_n2319), .D(_abc_40344_n2318), .Y(_abc_40344_n2320) );
  AOI22X1 AOI22X1_99 ( .A(_abc_40344_n1137), .B(_abc_40344_n2165), .C(_abc_40344_n2173), .D(_abc_40344_n1138), .Y(_abc_40344_n2326) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n978), .Q(ADDR_REG_19_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n1014), .Q(ADDR_REG_10_) );
  DFFPOSX1 DFFPOSX1_100 ( .CLK(clock), .D(n403), .Q(D_REG_13_) );
  DFFPOSX1 DFFPOSX1_101 ( .CLK(clock), .D(n408), .Q(D_REG_14_) );
  DFFPOSX1 DFFPOSX1_102 ( .CLK(clock), .D(n413), .Q(D_REG_15_) );
  DFFPOSX1 DFFPOSX1_103 ( .CLK(clock), .D(n418), .Q(D_REG_16_) );
  DFFPOSX1 DFFPOSX1_104 ( .CLK(clock), .D(n423), .Q(D_REG_17_) );
  DFFPOSX1 DFFPOSX1_105 ( .CLK(clock), .D(n428), .Q(D_REG_18_) );
  DFFPOSX1 DFFPOSX1_106 ( .CLK(clock), .D(n433), .Q(D_REG_19_) );
  DFFPOSX1 DFFPOSX1_107 ( .CLK(clock), .D(n438), .Q(D_REG_20_) );
  DFFPOSX1 DFFPOSX1_108 ( .CLK(clock), .D(n443), .Q(D_REG_21_) );
  DFFPOSX1 DFFPOSX1_109 ( .CLK(clock), .D(n448), .Q(D_REG_22_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n1018), .Q(ADDR_REG_9_) );
  DFFPOSX1 DFFPOSX1_110 ( .CLK(clock), .D(n453), .Q(D_REG_23_) );
  DFFPOSX1 DFFPOSX1_111 ( .CLK(clock), .D(n458), .Q(D_REG_24_) );
  DFFPOSX1 DFFPOSX1_112 ( .CLK(clock), .D(n463), .Q(D_REG_25_) );
  DFFPOSX1 DFFPOSX1_113 ( .CLK(clock), .D(n468), .Q(D_REG_26_) );
  DFFPOSX1 DFFPOSX1_114 ( .CLK(clock), .D(n473), .Q(D_REG_27_) );
  DFFPOSX1 DFFPOSX1_115 ( .CLK(clock), .D(n478), .Q(D_REG_28_) );
  DFFPOSX1 DFFPOSX1_116 ( .CLK(clock), .D(n483), .Q(D_REG_29_) );
  DFFPOSX1 DFFPOSX1_117 ( .CLK(clock), .D(n488), .Q(D_REG_30_) );
  DFFPOSX1 DFFPOSX1_118 ( .CLK(clock), .D(n493), .Q(D_REG_31_) );
  DFFPOSX1 DFFPOSX1_119 ( .CLK(clock), .D(n498), .Q(REG0_REG_0_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n1022), .Q(ADDR_REG_8_) );
  DFFPOSX1 DFFPOSX1_120 ( .CLK(clock), .D(n503), .Q(REG0_REG_1_) );
  DFFPOSX1 DFFPOSX1_121 ( .CLK(clock), .D(n508), .Q(REG0_REG_2_) );
  DFFPOSX1 DFFPOSX1_122 ( .CLK(clock), .D(n513), .Q(REG0_REG_3_) );
  DFFPOSX1 DFFPOSX1_123 ( .CLK(clock), .D(n518), .Q(REG0_REG_4_) );
  DFFPOSX1 DFFPOSX1_124 ( .CLK(clock), .D(n523), .Q(REG0_REG_5_) );
  DFFPOSX1 DFFPOSX1_125 ( .CLK(clock), .D(n528), .Q(REG0_REG_6_) );
  DFFPOSX1 DFFPOSX1_126 ( .CLK(clock), .D(n533), .Q(REG0_REG_7_) );
  DFFPOSX1 DFFPOSX1_127 ( .CLK(clock), .D(n538), .Q(REG0_REG_8_) );
  DFFPOSX1 DFFPOSX1_128 ( .CLK(clock), .D(n543), .Q(REG0_REG_9_) );
  DFFPOSX1 DFFPOSX1_129 ( .CLK(clock), .D(n548), .Q(REG0_REG_10_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n1026), .Q(ADDR_REG_7_) );
  DFFPOSX1 DFFPOSX1_130 ( .CLK(clock), .D(n553), .Q(REG0_REG_11_) );
  DFFPOSX1 DFFPOSX1_131 ( .CLK(clock), .D(n558), .Q(REG0_REG_12_) );
  DFFPOSX1 DFFPOSX1_132 ( .CLK(clock), .D(n563), .Q(REG0_REG_13_) );
  DFFPOSX1 DFFPOSX1_133 ( .CLK(clock), .D(n568), .Q(REG0_REG_14_) );
  DFFPOSX1 DFFPOSX1_134 ( .CLK(clock), .D(n573), .Q(REG0_REG_15_) );
  DFFPOSX1 DFFPOSX1_135 ( .CLK(clock), .D(n578), .Q(REG0_REG_16_) );
  DFFPOSX1 DFFPOSX1_136 ( .CLK(clock), .D(n583), .Q(REG0_REG_17_) );
  DFFPOSX1 DFFPOSX1_137 ( .CLK(clock), .D(n588), .Q(REG0_REG_18_) );
  DFFPOSX1 DFFPOSX1_138 ( .CLK(clock), .D(n593), .Q(REG0_REG_19_) );
  DFFPOSX1 DFFPOSX1_139 ( .CLK(clock), .D(n598), .Q(REG0_REG_20_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n1030), .Q(ADDR_REG_6_) );
  DFFPOSX1 DFFPOSX1_140 ( .CLK(clock), .D(n603), .Q(REG0_REG_21_) );
  DFFPOSX1 DFFPOSX1_141 ( .CLK(clock), .D(n608), .Q(REG0_REG_22_) );
  DFFPOSX1 DFFPOSX1_142 ( .CLK(clock), .D(n613), .Q(REG0_REG_23_) );
  DFFPOSX1 DFFPOSX1_143 ( .CLK(clock), .D(n618), .Q(REG0_REG_24_) );
  DFFPOSX1 DFFPOSX1_144 ( .CLK(clock), .D(n623), .Q(REG0_REG_25_) );
  DFFPOSX1 DFFPOSX1_145 ( .CLK(clock), .D(n628), .Q(REG0_REG_26_) );
  DFFPOSX1 DFFPOSX1_146 ( .CLK(clock), .D(n633), .Q(REG0_REG_27_) );
  DFFPOSX1 DFFPOSX1_147 ( .CLK(clock), .D(n638), .Q(REG0_REG_28_) );
  DFFPOSX1 DFFPOSX1_148 ( .CLK(clock), .D(n643), .Q(REG0_REG_29_) );
  DFFPOSX1 DFFPOSX1_149 ( .CLK(clock), .D(n648), .Q(REG0_REG_30_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n1034), .Q(ADDR_REG_5_) );
  DFFPOSX1 DFFPOSX1_150 ( .CLK(clock), .D(n653), .Q(REG0_REG_31_) );
  DFFPOSX1 DFFPOSX1_151 ( .CLK(clock), .D(n658), .Q(REG1_REG_0_) );
  DFFPOSX1 DFFPOSX1_152 ( .CLK(clock), .D(n663), .Q(REG1_REG_1_) );
  DFFPOSX1 DFFPOSX1_153 ( .CLK(clock), .D(n668), .Q(REG1_REG_2_) );
  DFFPOSX1 DFFPOSX1_154 ( .CLK(clock), .D(n673), .Q(REG1_REG_3_) );
  DFFPOSX1 DFFPOSX1_155 ( .CLK(clock), .D(n678), .Q(REG1_REG_4_) );
  DFFPOSX1 DFFPOSX1_156 ( .CLK(clock), .D(n683), .Q(REG1_REG_5_) );
  DFFPOSX1 DFFPOSX1_157 ( .CLK(clock), .D(n688), .Q(REG1_REG_6_) );
  DFFPOSX1 DFFPOSX1_158 ( .CLK(clock), .D(n693), .Q(REG1_REG_7_) );
  DFFPOSX1 DFFPOSX1_159 ( .CLK(clock), .D(n698), .Q(REG1_REG_8_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n1038), .Q(ADDR_REG_4_) );
  DFFPOSX1 DFFPOSX1_160 ( .CLK(clock), .D(n703), .Q(REG1_REG_9_) );
  DFFPOSX1 DFFPOSX1_161 ( .CLK(clock), .D(n708), .Q(REG1_REG_10_) );
  DFFPOSX1 DFFPOSX1_162 ( .CLK(clock), .D(n713), .Q(REG1_REG_11_) );
  DFFPOSX1 DFFPOSX1_163 ( .CLK(clock), .D(n718), .Q(REG1_REG_12_) );
  DFFPOSX1 DFFPOSX1_164 ( .CLK(clock), .D(n723), .Q(REG1_REG_13_) );
  DFFPOSX1 DFFPOSX1_165 ( .CLK(clock), .D(n728), .Q(REG1_REG_14_) );
  DFFPOSX1 DFFPOSX1_166 ( .CLK(clock), .D(n733), .Q(REG1_REG_15_) );
  DFFPOSX1 DFFPOSX1_167 ( .CLK(clock), .D(n738), .Q(REG1_REG_16_) );
  DFFPOSX1 DFFPOSX1_168 ( .CLK(clock), .D(n743), .Q(REG1_REG_17_) );
  DFFPOSX1 DFFPOSX1_169 ( .CLK(clock), .D(n748), .Q(REG1_REG_18_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n1042), .Q(ADDR_REG_3_) );
  DFFPOSX1 DFFPOSX1_170 ( .CLK(clock), .D(n753), .Q(REG1_REG_19_) );
  DFFPOSX1 DFFPOSX1_171 ( .CLK(clock), .D(n758), .Q(REG1_REG_20_) );
  DFFPOSX1 DFFPOSX1_172 ( .CLK(clock), .D(n763), .Q(REG1_REG_21_) );
  DFFPOSX1 DFFPOSX1_173 ( .CLK(clock), .D(n768), .Q(REG1_REG_22_) );
  DFFPOSX1 DFFPOSX1_174 ( .CLK(clock), .D(n773), .Q(REG1_REG_23_) );
  DFFPOSX1 DFFPOSX1_175 ( .CLK(clock), .D(n778), .Q(REG1_REG_24_) );
  DFFPOSX1 DFFPOSX1_176 ( .CLK(clock), .D(n783), .Q(REG1_REG_25_) );
  DFFPOSX1 DFFPOSX1_177 ( .CLK(clock), .D(n788), .Q(REG1_REG_26_) );
  DFFPOSX1 DFFPOSX1_178 ( .CLK(clock), .D(n793), .Q(REG1_REG_27_) );
  DFFPOSX1 DFFPOSX1_179 ( .CLK(clock), .D(n798), .Q(REG1_REG_28_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n1046), .Q(ADDR_REG_2_) );
  DFFPOSX1 DFFPOSX1_180 ( .CLK(clock), .D(n803), .Q(REG1_REG_29_) );
  DFFPOSX1 DFFPOSX1_181 ( .CLK(clock), .D(n808), .Q(REG1_REG_30_) );
  DFFPOSX1 DFFPOSX1_182 ( .CLK(clock), .D(n813), .Q(REG1_REG_31_) );
  DFFPOSX1 DFFPOSX1_183 ( .CLK(clock), .D(n818), .Q(REG2_REG_0_) );
  DFFPOSX1 DFFPOSX1_184 ( .CLK(clock), .D(n823), .Q(REG2_REG_1_) );
  DFFPOSX1 DFFPOSX1_185 ( .CLK(clock), .D(n828), .Q(REG2_REG_2_) );
  DFFPOSX1 DFFPOSX1_186 ( .CLK(clock), .D(n833), .Q(REG2_REG_3_) );
  DFFPOSX1 DFFPOSX1_187 ( .CLK(clock), .D(n838), .Q(REG2_REG_4_) );
  DFFPOSX1 DFFPOSX1_188 ( .CLK(clock), .D(n843), .Q(REG2_REG_5_) );
  DFFPOSX1 DFFPOSX1_189 ( .CLK(clock), .D(n848), .Q(REG2_REG_6_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n1050), .Q(ADDR_REG_1_) );
  DFFPOSX1 DFFPOSX1_190 ( .CLK(clock), .D(n853), .Q(REG2_REG_7_) );
  DFFPOSX1 DFFPOSX1_191 ( .CLK(clock), .D(n858), .Q(REG2_REG_8_) );
  DFFPOSX1 DFFPOSX1_192 ( .CLK(clock), .D(n863), .Q(REG2_REG_9_) );
  DFFPOSX1 DFFPOSX1_193 ( .CLK(clock), .D(n868), .Q(REG2_REG_10_) );
  DFFPOSX1 DFFPOSX1_194 ( .CLK(clock), .D(n873), .Q(REG2_REG_11_) );
  DFFPOSX1 DFFPOSX1_195 ( .CLK(clock), .D(n878), .Q(REG2_REG_12_) );
  DFFPOSX1 DFFPOSX1_196 ( .CLK(clock), .D(n883), .Q(REG2_REG_13_) );
  DFFPOSX1 DFFPOSX1_197 ( .CLK(clock), .D(n888), .Q(REG2_REG_14_) );
  DFFPOSX1 DFFPOSX1_198 ( .CLK(clock), .D(n893), .Q(REG2_REG_15_) );
  DFFPOSX1 DFFPOSX1_199 ( .CLK(clock), .D(n898), .Q(REG2_REG_16_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n982), .Q(ADDR_REG_18_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n1054), .Q(ADDR_REG_0_) );
  DFFPOSX1 DFFPOSX1_200 ( .CLK(clock), .D(n903), .Q(REG2_REG_17_) );
  DFFPOSX1 DFFPOSX1_201 ( .CLK(clock), .D(n908), .Q(REG2_REG_18_) );
  DFFPOSX1 DFFPOSX1_202 ( .CLK(clock), .D(n913), .Q(REG2_REG_19_) );
  DFFPOSX1 DFFPOSX1_203 ( .CLK(clock), .D(n918), .Q(REG2_REG_20_) );
  DFFPOSX1 DFFPOSX1_204 ( .CLK(clock), .D(n923), .Q(REG2_REG_21_) );
  DFFPOSX1 DFFPOSX1_205 ( .CLK(clock), .D(n928), .Q(REG2_REG_22_) );
  DFFPOSX1 DFFPOSX1_206 ( .CLK(clock), .D(n933), .Q(REG2_REG_23_) );
  DFFPOSX1 DFFPOSX1_207 ( .CLK(clock), .D(n938), .Q(REG2_REG_24_) );
  DFFPOSX1 DFFPOSX1_208 ( .CLK(clock), .D(n943), .Q(REG2_REG_25_) );
  DFFPOSX1 DFFPOSX1_209 ( .CLK(clock), .D(n948), .Q(REG2_REG_26_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n1182), .Q(DATAO_REG_31_) );
  DFFPOSX1 DFFPOSX1_210 ( .CLK(clock), .D(n953), .Q(REG2_REG_27_) );
  DFFPOSX1 DFFPOSX1_211 ( .CLK(clock), .D(n958), .Q(REG2_REG_28_) );
  DFFPOSX1 DFFPOSX1_212 ( .CLK(clock), .D(n963), .Q(REG2_REG_29_) );
  DFFPOSX1 DFFPOSX1_213 ( .CLK(clock), .D(n968), .Q(REG2_REG_30_) );
  DFFPOSX1 DFFPOSX1_214 ( .CLK(clock), .D(n973), .Q(REG2_REG_31_) );
  DFFPOSX1 DFFPOSX1_215 ( .CLK(clock), .D(n1186), .Q(B_REG) );
  DFFPOSX1 DFFPOSX1_216 ( .CLK(clock), .D(n1191), .Q(REG3_REG_15_) );
  DFFPOSX1 DFFPOSX1_217 ( .CLK(clock), .D(n1196), .Q(REG3_REG_26_) );
  DFFPOSX1 DFFPOSX1_218 ( .CLK(clock), .D(n1201), .Q(REG3_REG_6_) );
  DFFPOSX1 DFFPOSX1_219 ( .CLK(clock), .D(n1206), .Q(REG3_REG_18_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(n1178), .Q(DATAO_REG_30_) );
  DFFPOSX1 DFFPOSX1_220 ( .CLK(clock), .D(n1211), .Q(REG3_REG_2_) );
  DFFPOSX1 DFFPOSX1_221 ( .CLK(clock), .D(n1216), .Q(REG3_REG_11_) );
  DFFPOSX1 DFFPOSX1_222 ( .CLK(clock), .D(n1221), .Q(REG3_REG_22_) );
  DFFPOSX1 DFFPOSX1_223 ( .CLK(clock), .D(n1226), .Q(REG3_REG_13_) );
  DFFPOSX1 DFFPOSX1_224 ( .CLK(clock), .D(n1231), .Q(REG3_REG_20_) );
  DFFPOSX1 DFFPOSX1_225 ( .CLK(clock), .D(n1236), .Q(REG3_REG_0_) );
  DFFPOSX1 DFFPOSX1_226 ( .CLK(clock), .D(n1241), .Q(REG3_REG_9_) );
  DFFPOSX1 DFFPOSX1_227 ( .CLK(clock), .D(n1246), .Q(REG3_REG_4_) );
  DFFPOSX1 DFFPOSX1_228 ( .CLK(clock), .D(n1251), .Q(REG3_REG_24_) );
  DFFPOSX1 DFFPOSX1_229 ( .CLK(clock), .D(n1256), .Q(REG3_REG_17_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(n1174), .Q(DATAO_REG_29_) );
  DFFPOSX1 DFFPOSX1_230 ( .CLK(clock), .D(n1261), .Q(REG3_REG_5_) );
  DFFPOSX1 DFFPOSX1_231 ( .CLK(clock), .D(n1266), .Q(REG3_REG_16_) );
  DFFPOSX1 DFFPOSX1_232 ( .CLK(clock), .D(n1271), .Q(REG3_REG_25_) );
  DFFPOSX1 DFFPOSX1_233 ( .CLK(clock), .D(n1276), .Q(REG3_REG_12_) );
  DFFPOSX1 DFFPOSX1_234 ( .CLK(clock), .D(n1281), .Q(REG3_REG_21_) );
  DFFPOSX1 DFFPOSX1_235 ( .CLK(clock), .D(n1286), .Q(REG3_REG_1_) );
  DFFPOSX1 DFFPOSX1_236 ( .CLK(clock), .D(n1291), .Q(REG3_REG_8_) );
  DFFPOSX1 DFFPOSX1_237 ( .CLK(clock), .D(n1296), .Q(REG3_REG_28_) );
  DFFPOSX1 DFFPOSX1_238 ( .CLK(clock), .D(n1301), .Q(REG3_REG_19_) );
  DFFPOSX1 DFFPOSX1_239 ( .CLK(clock), .D(n1306), .Q(REG3_REG_3_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(n1170), .Q(DATAO_REG_28_) );
  DFFPOSX1 DFFPOSX1_240 ( .CLK(clock), .D(n1311), .Q(REG3_REG_10_) );
  DFFPOSX1 DFFPOSX1_241 ( .CLK(clock), .D(n1316), .Q(REG3_REG_23_) );
  DFFPOSX1 DFFPOSX1_242 ( .CLK(clock), .D(n1321), .Q(REG3_REG_14_) );
  DFFPOSX1 DFFPOSX1_243 ( .CLK(clock), .D(n1326), .Q(REG3_REG_27_) );
  DFFPOSX1 DFFPOSX1_244 ( .CLK(clock), .D(n1331), .Q(REG3_REG_7_) );
  DFFPOSX1 DFFPOSX1_245 ( .CLK(clock), .D(n1336), .Q(STATE_REG) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(n1166), .Q(DATAO_REG_27_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(n1162), .Q(DATAO_REG_26_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(n1158), .Q(DATAO_REG_25_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(n1154), .Q(DATAO_REG_24_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(n1150), .Q(DATAO_REG_23_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n986), .Q(ADDR_REG_17_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(n1146), .Q(DATAO_REG_22_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(n1142), .Q(DATAO_REG_21_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(n1138), .Q(DATAO_REG_20_) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(n1134), .Q(DATAO_REG_19_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(n1130), .Q(DATAO_REG_18_) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(n1126), .Q(DATAO_REG_17_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(n1122), .Q(DATAO_REG_16_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(n1118), .Q(DATAO_REG_15_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(n1114), .Q(DATAO_REG_14_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(n1110), .Q(DATAO_REG_13_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n990), .Q(ADDR_REG_16_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(n1106), .Q(DATAO_REG_12_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(n1102), .Q(DATAO_REG_11_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(n1098), .Q(DATAO_REG_10_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(n1094), .Q(DATAO_REG_9_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(n1090), .Q(DATAO_REG_8_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(n1086), .Q(DATAO_REG_7_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(n1082), .Q(DATAO_REG_6_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(n1078), .Q(DATAO_REG_5_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(n1074), .Q(DATAO_REG_4_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(n1070), .Q(DATAO_REG_3_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n994), .Q(ADDR_REG_15_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(n1066), .Q(DATAO_REG_2_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(n1062), .Q(DATAO_REG_1_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(n1058), .Q(DATAO_REG_0_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(n1341), .Q(RD_REG) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(n1345), .Q(WR_REG) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(n178), .Q(IR_REG_0_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(n183), .Q(IR_REG_1_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(n188), .Q(IR_REG_2_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(n193), .Q(IR_REG_3_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(n198), .Q(IR_REG_4_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n998), .Q(ADDR_REG_14_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(n203), .Q(IR_REG_5_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(n208), .Q(IR_REG_6_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(n213), .Q(IR_REG_7_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(n218), .Q(IR_REG_8_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(n223), .Q(IR_REG_9_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(n228), .Q(IR_REG_10_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(n233), .Q(IR_REG_11_) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(clock), .D(n238), .Q(IR_REG_12_) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(clock), .D(n243), .Q(IR_REG_13_) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(clock), .D(n248), .Q(IR_REG_14_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n1002), .Q(ADDR_REG_13_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(clock), .D(n253), .Q(IR_REG_15_) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(clock), .D(n258), .Q(IR_REG_16_) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(clock), .D(n263), .Q(IR_REG_17_) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(clock), .D(n268), .Q(IR_REG_18_) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(clock), .D(n273), .Q(IR_REG_19_) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(clock), .D(n278), .Q(IR_REG_20_) );
  DFFPOSX1 DFFPOSX1_76 ( .CLK(clock), .D(n283), .Q(IR_REG_21_) );
  DFFPOSX1 DFFPOSX1_77 ( .CLK(clock), .D(n288), .Q(IR_REG_22_) );
  DFFPOSX1 DFFPOSX1_78 ( .CLK(clock), .D(n293), .Q(IR_REG_23_) );
  DFFPOSX1 DFFPOSX1_79 ( .CLK(clock), .D(n298), .Q(IR_REG_24_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n1006), .Q(ADDR_REG_12_) );
  DFFPOSX1 DFFPOSX1_80 ( .CLK(clock), .D(n303), .Q(IR_REG_25_) );
  DFFPOSX1 DFFPOSX1_81 ( .CLK(clock), .D(n308), .Q(IR_REG_26_) );
  DFFPOSX1 DFFPOSX1_82 ( .CLK(clock), .D(n313), .Q(IR_REG_27_) );
  DFFPOSX1 DFFPOSX1_83 ( .CLK(clock), .D(n318), .Q(IR_REG_28_) );
  DFFPOSX1 DFFPOSX1_84 ( .CLK(clock), .D(n323), .Q(IR_REG_29_) );
  DFFPOSX1 DFFPOSX1_85 ( .CLK(clock), .D(n328), .Q(IR_REG_30_) );
  DFFPOSX1 DFFPOSX1_86 ( .CLK(clock), .D(n333), .Q(IR_REG_31_) );
  DFFPOSX1 DFFPOSX1_87 ( .CLK(clock), .D(n338), .Q(D_REG_0_) );
  DFFPOSX1 DFFPOSX1_88 ( .CLK(clock), .D(n343), .Q(D_REG_1_) );
  DFFPOSX1 DFFPOSX1_89 ( .CLK(clock), .D(n348), .Q(D_REG_2_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n1010), .Q(ADDR_REG_11_) );
  DFFPOSX1 DFFPOSX1_90 ( .CLK(clock), .D(n353), .Q(D_REG_3_) );
  DFFPOSX1 DFFPOSX1_91 ( .CLK(clock), .D(n358), .Q(D_REG_4_) );
  DFFPOSX1 DFFPOSX1_92 ( .CLK(clock), .D(n363), .Q(D_REG_5_) );
  DFFPOSX1 DFFPOSX1_93 ( .CLK(clock), .D(n368), .Q(D_REG_6_) );
  DFFPOSX1 DFFPOSX1_94 ( .CLK(clock), .D(n373), .Q(D_REG_7_) );
  DFFPOSX1 DFFPOSX1_95 ( .CLK(clock), .D(n378), .Q(D_REG_8_) );
  DFFPOSX1 DFFPOSX1_96 ( .CLK(clock), .D(n383), .Q(D_REG_9_) );
  DFFPOSX1 DFFPOSX1_97 ( .CLK(clock), .D(n388), .Q(D_REG_10_) );
  DFFPOSX1 DFFPOSX1_98 ( .CLK(clock), .D(n393), .Q(D_REG_11_) );
  DFFPOSX1 DFFPOSX1_99 ( .CLK(clock), .D(n398), .Q(D_REG_12_) );
  INVX1 INVX1_1 ( .A(_abc_40344_n526), .Y(_abc_40344_n527) );
  INVX1 INVX1_10 ( .A(_abc_40344_n568), .Y(_abc_40344_n569_1) );
  INVX1 INVX1_100 ( .A(DATAI_15_), .Y(_abc_40344_n1198) );
  INVX1 INVX1_101 ( .A(_abc_40344_n1202), .Y(_abc_40344_n1203) );
  INVX1 INVX1_102 ( .A(REG2_REG_15_), .Y(_abc_40344_n1207) );
  INVX1 INVX1_103 ( .A(_abc_40344_n1213), .Y(_abc_40344_n1214) );
  INVX1 INVX1_104 ( .A(_abc_40344_n1215), .Y(_abc_40344_n1216) );
  INVX1 INVX1_105 ( .A(_abc_40344_n1218), .Y(_abc_40344_n1219) );
  INVX1 INVX1_106 ( .A(REG3_REG_14_), .Y(_abc_40344_n1225_1) );
  INVX1 INVX1_107 ( .A(_abc_40344_n1227), .Y(_abc_40344_n1228) );
  INVX1 INVX1_108 ( .A(REG2_REG_14_), .Y(_abc_40344_n1231) );
  INVX1 INVX1_109 ( .A(_abc_40344_n1237), .Y(_abc_40344_n1238) );
  INVX1 INVX1_11 ( .A(_abc_40344_n547), .Y(_abc_40344_n575_1) );
  INVX1 INVX1_110 ( .A(_abc_40344_n1240_1), .Y(_abc_40344_n1241) );
  INVX1 INVX1_111 ( .A(IR_REG_10_), .Y(_abc_40344_n1243) );
  INVX1 INVX1_112 ( .A(REG1_REG_13_), .Y(_abc_40344_n1252) );
  INVX1 INVX1_113 ( .A(REG0_REG_13_), .Y(_abc_40344_n1253) );
  INVX1 INVX1_114 ( .A(REG2_REG_13_), .Y(_abc_40344_n1255) );
  INVX1 INVX1_115 ( .A(_abc_40344_n1256), .Y(_abc_40344_n1257) );
  INVX1 INVX1_116 ( .A(_abc_40344_n1261), .Y(_abc_40344_n1262) );
  INVX1 INVX1_117 ( .A(REG2_REG_11_), .Y(_abc_40344_n1274) );
  INVX1 INVX1_118 ( .A(_abc_40344_n1275), .Y(_abc_40344_n1276) );
  INVX1 INVX1_119 ( .A(_abc_40344_n1278), .Y(_abc_40344_n1279) );
  INVX1 INVX1_12 ( .A(_abc_40344_n595_1), .Y(_abc_40344_n597) );
  INVX1 INVX1_120 ( .A(REG1_REG_11_), .Y(_abc_40344_n1281) );
  INVX1 INVX1_121 ( .A(REG0_REG_11_), .Y(_abc_40344_n1282_1) );
  INVX1 INVX1_122 ( .A(REG0_REG_12_), .Y(_abc_40344_n1297) );
  INVX1 INVX1_123 ( .A(REG3_REG_12_), .Y(_abc_40344_n1299) );
  INVX1 INVX1_124 ( .A(_abc_40344_n1301), .Y(_abc_40344_n1302) );
  INVX1 INVX1_125 ( .A(_abc_40344_n1319), .Y(_abc_40344_n1320) );
  INVX1 INVX1_126 ( .A(DATAI_10_), .Y(_abc_40344_n1321) );
  INVX1 INVX1_127 ( .A(REG0_REG_10_), .Y(_abc_40344_n1328) );
  INVX1 INVX1_128 ( .A(_abc_40344_n1329), .Y(_abc_40344_n1330) );
  INVX1 INVX1_129 ( .A(REG1_REG_10_), .Y(_abc_40344_n1332) );
  INVX1 INVX1_13 ( .A(IR_REG_28_), .Y(_abc_40344_n600_1) );
  INVX1 INVX1_130 ( .A(DATAI_9_), .Y(_abc_40344_n1341) );
  INVX1 INVX1_131 ( .A(_abc_40344_n1246), .Y(_abc_40344_n1342) );
  INVX1 INVX1_132 ( .A(IR_REG_9_), .Y(_abc_40344_n1345) );
  INVX1 INVX1_133 ( .A(REG1_REG_9_), .Y(_abc_40344_n1351) );
  INVX1 INVX1_134 ( .A(REG0_REG_9_), .Y(_abc_40344_n1352) );
  INVX1 INVX1_135 ( .A(_abc_40344_n1051_1), .Y(_abc_40344_n1355) );
  INVX1 INVX1_136 ( .A(REG3_REG_9_), .Y(_abc_40344_n1356) );
  INVX1 INVX1_137 ( .A(_abc_40344_n1358), .Y(_abc_40344_n1359_1) );
  INVX1 INVX1_138 ( .A(_abc_40344_n1363), .Y(_abc_40344_n1364) );
  INVX1 INVX1_139 ( .A(_abc_40344_n1367), .Y(_abc_40344_n1368) );
  INVX1 INVX1_14 ( .A(IR_REG_27_), .Y(_abc_40344_n604) );
  INVX1 INVX1_140 ( .A(_abc_40344_n1372), .Y(_abc_40344_n1373) );
  INVX1 INVX1_141 ( .A(_abc_40344_n1379), .Y(_abc_40344_n1380) );
  INVX1 INVX1_142 ( .A(_abc_40344_n1376), .Y(_abc_40344_n1381) );
  INVX1 INVX1_143 ( .A(_abc_40344_n1378), .Y(_abc_40344_n1382) );
  INVX1 INVX1_144 ( .A(_abc_40344_n1398), .Y(_abc_40344_n1399) );
  INVX1 INVX1_145 ( .A(REG3_REG_19_), .Y(_abc_40344_n1405) );
  INVX1 INVX1_146 ( .A(_abc_40344_n1407), .Y(_abc_40344_n1408) );
  INVX1 INVX1_147 ( .A(REG2_REG_19_), .Y(_abc_40344_n1411) );
  INVX1 INVX1_148 ( .A(REG1_REG_19_), .Y(_abc_40344_n1412) );
  INVX1 INVX1_149 ( .A(_abc_40344_n1414), .Y(_abc_40344_n1415) );
  INVX1 INVX1_15 ( .A(IR_REG_21_), .Y(_abc_40344_n612) );
  INVX1 INVX1_150 ( .A(_abc_40344_n1416), .Y(_abc_40344_n1417) );
  INVX1 INVX1_151 ( .A(_abc_40344_n1446), .Y(_abc_40344_n1447) );
  INVX1 INVX1_152 ( .A(_abc_40344_n1420), .Y(_abc_40344_n1450) );
  INVX1 INVX1_153 ( .A(_abc_40344_n1451_1), .Y(_abc_40344_n1452) );
  INVX1 INVX1_154 ( .A(_abc_40344_n1457), .Y(_abc_40344_n1458) );
  INVX1 INVX1_155 ( .A(REG1_REG_24_), .Y(_abc_40344_n1467) );
  INVX1 INVX1_156 ( .A(_abc_40344_n1472), .Y(_abc_40344_n1473) );
  INVX1 INVX1_157 ( .A(_abc_40344_n1482), .Y(_abc_40344_n1483) );
  INVX1 INVX1_158 ( .A(REG1_REG_25_), .Y(_abc_40344_n1484) );
  INVX1 INVX1_159 ( .A(_abc_40344_n1499), .Y(_abc_40344_n1500) );
  INVX1 INVX1_16 ( .A(IR_REG_20_), .Y(_abc_40344_n613) );
  INVX1 INVX1_160 ( .A(REG1_REG_26_), .Y(_abc_40344_n1501) );
  INVX1 INVX1_161 ( .A(_abc_40344_n1504), .Y(_abc_40344_n1505_1) );
  INVX1 INVX1_162 ( .A(_abc_40344_n1513), .Y(_abc_40344_n1514_1) );
  INVX1 INVX1_163 ( .A(_abc_40344_n1517_1), .Y(_abc_40344_n1518) );
  INVX1 INVX1_164 ( .A(_abc_40344_n1191), .Y(_abc_40344_n1524) );
  INVX1 INVX1_165 ( .A(_abc_40344_n1401), .Y(_abc_40344_n1527) );
  INVX1 INVX1_166 ( .A(_abc_40344_n1448), .Y(_abc_40344_n1529) );
  INVX1 INVX1_167 ( .A(_abc_40344_n1521), .Y(_abc_40344_n1534) );
  INVX1 INVX1_168 ( .A(_abc_40344_n1543), .Y(_abc_40344_n1544) );
  INVX1 INVX1_169 ( .A(REG1_REG_28_), .Y(_abc_40344_n1545) );
  INVX1 INVX1_17 ( .A(IR_REG_22_), .Y(_abc_40344_n620) );
  INVX1 INVX1_170 ( .A(_abc_40344_n1559), .Y(_abc_40344_n1560) );
  INVX1 INVX1_171 ( .A(_abc_40344_n1339), .Y(_abc_40344_n1588) );
  INVX1 INVX1_172 ( .A(_abc_40344_n844), .Y(_abc_40344_n1602) );
  INVX1 INVX1_173 ( .A(_abc_40344_n1610), .Y(_abc_40344_n1611) );
  INVX1 INVX1_174 ( .A(_abc_40344_n1081), .Y(_abc_40344_n1636) );
  INVX1 INVX1_175 ( .A(REG1_REG_29_), .Y(_abc_40344_n1641) );
  INVX1 INVX1_176 ( .A(_abc_40344_n1541), .Y(_abc_40344_n1648) );
  INVX1 INVX1_177 ( .A(DATAI_8_), .Y(_abc_40344_n1663) );
  INVX1 INVX1_178 ( .A(_abc_40344_n893), .Y(_abc_40344_n1671) );
  INVX1 INVX1_179 ( .A(REG3_REG_1_), .Y(_abc_40344_n1678) );
  INVX1 INVX1_18 ( .A(_abc_40344_n651_1), .Y(_abc_40344_n652_1) );
  INVX1 INVX1_180 ( .A(_abc_40344_n1454), .Y(_abc_40344_n1689) );
  INVX1 INVX1_181 ( .A(_abc_40344_n1436), .Y(_abc_40344_n1693) );
  INVX1 INVX1_182 ( .A(_abc_40344_n1703), .Y(_abc_40344_n1704) );
  INVX1 INVX1_183 ( .A(_abc_40344_n1515), .Y(_abc_40344_n1719) );
  INVX1 INVX1_184 ( .A(_abc_40344_n1481), .Y(_abc_40344_n1726) );
  INVX1 INVX1_185 ( .A(_abc_40344_n1172), .Y(_abc_40344_n1732) );
  INVX1 INVX1_186 ( .A(_abc_40344_n1400), .Y(_abc_40344_n1750) );
  INVX1 INVX1_187 ( .A(REG3_REG_17_), .Y(_abc_40344_n1757) );
  INVX1 INVX1_188 ( .A(_abc_40344_n1763), .Y(_abc_40344_n1765) );
  INVX1 INVX1_189 ( .A(REG3_REG_0_), .Y(_abc_40344_n1794) );
  INVX1 INVX1_19 ( .A(_abc_40344_n655), .Y(_abc_40344_n656) );
  INVX1 INVX1_190 ( .A(_abc_40344_n1421_1), .Y(_abc_40344_n1812) );
  INVX1 INVX1_191 ( .A(REG3_REG_2_), .Y(_abc_40344_n1854) );
  INVX1 INVX1_192 ( .A(_abc_40344_n693), .Y(_abc_40344_n1872) );
  INVX1 INVX1_193 ( .A(_abc_40344_n1715), .Y(_abc_40344_n1878) );
  INVX1 INVX1_194 ( .A(_abc_40344_n1511_1), .Y(_abc_40344_n1879) );
  INVX1 INVX1_195 ( .A(_abc_40344_n1887), .Y(_abc_40344_n1888) );
  INVX1 INVX1_196 ( .A(REG1_REG_31_), .Y(_abc_40344_n1911) );
  INVX1 INVX1_197 ( .A(_abc_40344_n1914), .Y(_abc_40344_n1915) );
  INVX1 INVX1_198 ( .A(REG1_REG_30_), .Y(_abc_40344_n1919) );
  INVX1 INVX1_199 ( .A(_abc_40344_n1923), .Y(_abc_40344_n1924) );
  INVX1 INVX1_2 ( .A(IR_REG_8_), .Y(_abc_40344_n528) );
  INVX1 INVX1_20 ( .A(_abc_40344_n658_1), .Y(_abc_40344_n659) );
  INVX1 INVX1_200 ( .A(DATAI_25_), .Y(_abc_40344_n1931) );
  INVX1 INVX1_201 ( .A(_abc_40344_n1939), .Y(_abc_40344_n1940) );
  INVX1 INVX1_202 ( .A(_abc_40344_n1943), .Y(_abc_40344_n1944) );
  INVX1 INVX1_203 ( .A(_abc_40344_n1957), .Y(_abc_40344_n1958) );
  INVX1 INVX1_204 ( .A(_abc_40344_n1962), .Y(_abc_40344_n1963) );
  INVX1 INVX1_205 ( .A(_abc_40344_n1325), .Y(_abc_40344_n1967) );
  INVX1 INVX1_206 ( .A(_abc_40344_n1975), .Y(_abc_40344_n1976) );
  INVX1 INVX1_207 ( .A(_abc_40344_n1978), .Y(_abc_40344_n1979) );
  INVX1 INVX1_208 ( .A(_abc_40344_n1983), .Y(_abc_40344_n1984) );
  INVX1 INVX1_209 ( .A(REG0_REG_6_), .Y(_abc_40344_n1987) );
  INVX1 INVX1_21 ( .A(IR_REG_30_), .Y(_abc_40344_n662) );
  INVX1 INVX1_210 ( .A(REG1_REG_6_), .Y(_abc_40344_n1989) );
  INVX1 INVX1_211 ( .A(_abc_40344_n712), .Y(_abc_40344_n1992) );
  INVX1 INVX1_212 ( .A(_abc_40344_n1995), .Y(_abc_40344_n1996) );
  INVX1 INVX1_213 ( .A(_abc_40344_n1934), .Y(_abc_40344_n2002) );
  INVX1 INVX1_214 ( .A(_abc_40344_n2005), .Y(_abc_40344_n2006) );
  INVX1 INVX1_215 ( .A(DATAI_27_), .Y(_abc_40344_n2009) );
  INVX1 INVX1_216 ( .A(REG1_REG_3_), .Y(_abc_40344_n2014) );
  INVX1 INVX1_217 ( .A(REG0_REG_3_), .Y(_abc_40344_n2015) );
  INVX1 INVX1_218 ( .A(_abc_40344_n807_1), .Y(_abc_40344_n2017) );
  INVX1 INVX1_219 ( .A(_abc_40344_n2023), .Y(_abc_40344_n2024) );
  INVX1 INVX1_22 ( .A(_abc_40344_n667), .Y(_abc_40344_n668_1) );
  INVX1 INVX1_220 ( .A(_abc_40344_n1946), .Y(_abc_40344_n2033) );
  INVX1 INVX1_221 ( .A(_abc_40344_n2034), .Y(_abc_40344_n2055) );
  INVX1 INVX1_222 ( .A(_abc_40344_n2059), .Y(_abc_40344_n2060) );
  INVX1 INVX1_223 ( .A(_abc_40344_n2064), .Y(_abc_40344_n2065) );
  INVX1 INVX1_224 ( .A(_abc_40344_n2073), .Y(_abc_40344_n2074) );
  INVX1 INVX1_225 ( .A(_abc_40344_n2077), .Y(_abc_40344_n2078) );
  INVX1 INVX1_226 ( .A(_abc_40344_n2082), .Y(_abc_40344_n2083) );
  INVX1 INVX1_227 ( .A(_abc_40344_n1997), .Y(_abc_40344_n2085) );
  INVX1 INVX1_228 ( .A(_abc_40344_n2088), .Y(_abc_40344_n2089) );
  INVX1 INVX1_229 ( .A(_abc_40344_n1917), .Y(_abc_40344_n2102) );
  INVX1 INVX1_23 ( .A(IR_REG_29_), .Y(_abc_40344_n670) );
  INVX1 INVX1_230 ( .A(_abc_40344_n2001), .Y(_abc_40344_n2116) );
  INVX1 INVX1_231 ( .A(_abc_40344_n2118), .Y(_abc_40344_n2119) );
  INVX1 INVX1_232 ( .A(_abc_40344_n2134), .Y(_abc_40344_n2135) );
  INVX1 INVX1_233 ( .A(_abc_40344_n2137), .Y(_abc_40344_n2138) );
  INVX1 INVX1_234 ( .A(_abc_40344_n2143), .Y(_abc_40344_n2146) );
  INVX1 INVX1_235 ( .A(DATAI_4_), .Y(_abc_40344_n2168) );
  INVX1 INVX1_236 ( .A(_abc_40344_n779), .Y(_abc_40344_n2201) );
  INVX1 INVX1_237 ( .A(REG2_REG_4_), .Y(_abc_40344_n2203) );
  INVX1 INVX1_238 ( .A(_abc_40344_n2275), .Y(_abc_40344_n2290) );
  INVX1 INVX1_239 ( .A(_abc_40344_n2276), .Y(_abc_40344_n2291) );
  INVX1 INVX1_24 ( .A(REG3_REG_6_), .Y(_abc_40344_n686) );
  INVX1 INVX1_240 ( .A(_abc_40344_n2279), .Y(_abc_40344_n2292) );
  INVX1 INVX1_241 ( .A(_abc_40344_n2302), .Y(_abc_40344_n2303) );
  INVX1 INVX1_242 ( .A(_abc_40344_n2304), .Y(_abc_40344_n2305) );
  INVX1 INVX1_243 ( .A(_abc_40344_n2306), .Y(_abc_40344_n2307) );
  INVX1 INVX1_244 ( .A(_abc_40344_n2311), .Y(_abc_40344_n2312) );
  INVX1 INVX1_245 ( .A(_abc_40344_n2313), .Y(_abc_40344_n2314_1) );
  INVX1 INVX1_246 ( .A(_abc_40344_n2320), .Y(_abc_40344_n2321) );
  INVX1 INVX1_247 ( .A(_abc_40344_n2339), .Y(_abc_40344_n2340_1) );
  INVX1 INVX1_248 ( .A(_abc_40344_n2342), .Y(_abc_40344_n2343) );
  INVX1 INVX1_249 ( .A(_abc_40344_n2352), .Y(_abc_40344_n2353) );
  INVX1 INVX1_25 ( .A(REG3_REG_4_), .Y(_abc_40344_n687) );
  INVX1 INVX1_250 ( .A(_abc_40344_n2354), .Y(_abc_40344_n2355) );
  INVX1 INVX1_251 ( .A(_abc_40344_n2361), .Y(_abc_40344_n2362_1) );
  INVX1 INVX1_252 ( .A(_abc_40344_n2365), .Y(_abc_40344_n2366) );
  INVX1 INVX1_253 ( .A(_abc_40344_n2368), .Y(_abc_40344_n2369_1) );
  INVX1 INVX1_254 ( .A(_abc_40344_n2378), .Y(_abc_40344_n2379) );
  INVX1 INVX1_255 ( .A(_abc_40344_n2380_1), .Y(_abc_40344_n2381) );
  INVX1 INVX1_256 ( .A(_abc_40344_n2382), .Y(_abc_40344_n2383) );
  INVX1 INVX1_257 ( .A(_abc_40344_n2386), .Y(_abc_40344_n2387) );
  INVX1 INVX1_258 ( .A(_abc_40344_n1550), .Y(_abc_40344_n2391) );
  INVX1 INVX1_259 ( .A(_abc_40344_n2397), .Y(_abc_40344_n2398) );
  INVX1 INVX1_26 ( .A(DATAI_6_), .Y(_abc_40344_n701) );
  INVX1 INVX1_260 ( .A(_abc_40344_n2402), .Y(_abc_40344_n2403) );
  INVX1 INVX1_261 ( .A(_abc_40344_n2406), .Y(_abc_40344_n2407) );
  INVX1 INVX1_262 ( .A(_abc_40344_n2410), .Y(_abc_40344_n2411) );
  INVX1 INVX1_263 ( .A(_abc_40344_n2211), .Y(_abc_40344_n2430) );
  INVX1 INVX1_264 ( .A(_abc_40344_n2315), .Y(_abc_40344_n2452) );
  INVX1 INVX1_265 ( .A(_abc_40344_n2327), .Y(_abc_40344_n2454) );
  INVX1 INVX1_266 ( .A(_abc_40344_n2334), .Y(_abc_40344_n2455) );
  INVX1 INVX1_267 ( .A(_abc_40344_n2346), .Y(_abc_40344_n2457) );
  INVX1 INVX1_268 ( .A(_abc_40344_n2374), .Y(_abc_40344_n2460) );
  INVX1 INVX1_269 ( .A(_abc_40344_n2393), .Y(_abc_40344_n2463) );
  INVX1 INVX1_27 ( .A(_abc_40344_n718), .Y(_abc_40344_n721) );
  INVX1 INVX1_270 ( .A(_abc_40344_n2399), .Y(_abc_40344_n2464) );
  INVX1 INVX1_271 ( .A(_abc_40344_n2413), .Y(_abc_40344_n2467) );
  INVX1 INVX1_272 ( .A(_abc_40344_n1956), .Y(_abc_40344_n2471) );
  INVX1 INVX1_273 ( .A(_abc_40344_n2472), .Y(_abc_40344_n2473) );
  INVX1 INVX1_274 ( .A(_abc_40344_n2049), .Y(_abc_40344_n2478_1) );
  INVX1 INVX1_275 ( .A(_abc_40344_n2482), .Y(_abc_40344_n2483) );
  INVX1 INVX1_276 ( .A(_abc_40344_n2130), .Y(_abc_40344_n2486) );
  INVX1 INVX1_277 ( .A(_abc_40344_n1980), .Y(_abc_40344_n2498) );
  INVX1 INVX1_278 ( .A(_abc_40344_n2042), .Y(_abc_40344_n2502_1) );
  INVX1 INVX1_279 ( .A(_abc_40344_n2516), .Y(_abc_40344_n2517) );
  INVX1 INVX1_28 ( .A(_abc_40344_n726), .Y(_abc_40344_n727_1) );
  INVX1 INVX1_280 ( .A(_abc_40344_n1908), .Y(_abc_40344_n2531) );
  INVX1 INVX1_281 ( .A(_abc_40344_n2056), .Y(_abc_40344_n2537) );
  INVX1 INVX1_282 ( .A(_abc_40344_n2541), .Y(_abc_40344_n2542) );
  INVX1 INVX1_283 ( .A(_abc_40344_n2068), .Y(_abc_40344_n2544) );
  INVX1 INVX1_284 ( .A(_abc_40344_n1927), .Y(_abc_40344_n2557) );
  INVX1 INVX1_285 ( .A(_abc_40344_n1916), .Y(_abc_40344_n2566) );
  INVX1 INVX1_286 ( .A(_abc_40344_n2569), .Y(_abc_40344_n2570) );
  INVX1 INVX1_287 ( .A(_abc_40344_n2571), .Y(_abc_40344_n2572) );
  INVX1 INVX1_288 ( .A(DATAI_28_), .Y(_abc_40344_n2573_1) );
  INVX1 INVX1_289 ( .A(_abc_40344_n2511), .Y(_abc_40344_n2577) );
  INVX1 INVX1_29 ( .A(DATAI_5_), .Y(_abc_40344_n728) );
  INVX1 INVX1_290 ( .A(_abc_40344_n2117), .Y(_abc_40344_n2582) );
  INVX1 INVX1_291 ( .A(_abc_40344_n2587), .Y(_abc_40344_n2588) );
  INVX1 INVX1_292 ( .A(_abc_40344_n1950), .Y(_abc_40344_n2589) );
  INVX1 INVX1_293 ( .A(_abc_40344_n2599_1), .Y(_abc_40344_n2604) );
  INVX1 INVX1_294 ( .A(_abc_40344_n2617), .Y(_abc_40344_n2618) );
  INVX1 INVX1_295 ( .A(_abc_40344_n2619_1), .Y(_abc_40344_n2620) );
  INVX1 INVX1_296 ( .A(_abc_40344_n2609), .Y(_abc_40344_n2623) );
  INVX1 INVX1_297 ( .A(_abc_40344_n2615), .Y(_abc_40344_n2625_1) );
  INVX1 INVX1_298 ( .A(_abc_40344_n2018), .Y(_abc_40344_n2628) );
  INVX1 INVX1_299 ( .A(_abc_40344_n2223), .Y(_abc_40344_n2631) );
  INVX1 INVX1_3 ( .A(IR_REG_3_), .Y(_abc_40344_n529) );
  INVX1 INVX1_30 ( .A(REG3_REG_5_), .Y(_abc_40344_n736) );
  INVX1 INVX1_300 ( .A(_abc_40344_n2635), .Y(_abc_40344_n2636) );
  INVX1 INVX1_301 ( .A(_abc_40344_n717), .Y(_abc_40344_n2643) );
  INVX1 INVX1_302 ( .A(_abc_40344_n2648), .Y(_abc_40344_n2649) );
  INVX1 INVX1_303 ( .A(_abc_40344_n2652), .Y(_abc_40344_n2653) );
  INVX1 INVX1_304 ( .A(_abc_40344_n2664), .Y(_abc_40344_n2665) );
  INVX1 INVX1_305 ( .A(_abc_40344_n2680), .Y(_abc_40344_n2681) );
  INVX1 INVX1_306 ( .A(_abc_40344_n2695), .Y(_abc_40344_n2696) );
  INVX1 INVX1_307 ( .A(_abc_40344_n2677), .Y(_abc_40344_n2704) );
  INVX1 INVX1_308 ( .A(REG2_REG_2_), .Y(_abc_40344_n2712) );
  INVX1 INVX1_309 ( .A(_abc_40344_n2728), .Y(_abc_40344_n2729) );
  INVX1 INVX1_31 ( .A(_abc_40344_n738_1), .Y(_abc_40344_n739) );
  INVX1 INVX1_310 ( .A(_abc_40344_n2737), .Y(_abc_40344_n2738) );
  INVX1 INVX1_311 ( .A(_abc_40344_n587), .Y(_abc_40344_n2774) );
  INVX1 INVX1_312 ( .A(_abc_40344_n1873), .Y(_abc_40344_n2775) );
  INVX1 INVX1_313 ( .A(_abc_40344_n2783), .Y(_abc_40344_n2784) );
  INVX1 INVX1_314 ( .A(_abc_40344_n2802), .Y(_abc_40344_n2803) );
  INVX1 INVX1_315 ( .A(_abc_40344_n2814), .Y(_abc_40344_n2815) );
  INVX1 INVX1_316 ( .A(_abc_40344_n2817), .Y(_abc_40344_n2818) );
  INVX1 INVX1_317 ( .A(ADDR_REG_9_), .Y(_abc_40344_n2828) );
  INVX1 INVX1_318 ( .A(_abc_40344_n2836), .Y(_abc_40344_n2844) );
  INVX1 INVX1_319 ( .A(_abc_40344_n2846), .Y(_abc_40344_n2847) );
  INVX1 INVX1_32 ( .A(_abc_40344_n699), .Y(_abc_40344_n744) );
  INVX1 INVX1_320 ( .A(_abc_40344_n2848), .Y(_abc_40344_n2849) );
  INVX1 INVX1_321 ( .A(_abc_40344_n2854), .Y(_abc_40344_n2855) );
  INVX1 INVX1_322 ( .A(_abc_40344_n2865), .Y(_abc_40344_n2866) );
  INVX1 INVX1_323 ( .A(_abc_40344_n1293_1), .Y(_abc_40344_n2883) );
  INVX1 INVX1_324 ( .A(_abc_40344_n2890), .Y(_abc_40344_n2891) );
  INVX1 INVX1_325 ( .A(_abc_40344_n1249), .Y(_abc_40344_n2911) );
  INVX1 INVX1_326 ( .A(_abc_40344_n2872), .Y(_abc_40344_n2914) );
  INVX1 INVX1_327 ( .A(_abc_40344_n2934), .Y(_abc_40344_n2935) );
  INVX1 INVX1_328 ( .A(_abc_40344_n2936), .Y(_abc_40344_n2937) );
  INVX1 INVX1_329 ( .A(_abc_40344_n2910), .Y(_abc_40344_n2939) );
  INVX1 INVX1_33 ( .A(REG0_REG_5_), .Y(_abc_40344_n751_1) );
  INVX1 INVX1_330 ( .A(_abc_40344_n2912), .Y(_abc_40344_n2940) );
  INVX1 INVX1_331 ( .A(_abc_40344_n2951), .Y(_abc_40344_n2952) );
  INVX1 INVX1_332 ( .A(ADDR_REG_15_), .Y(_abc_40344_n2956) );
  INVX1 INVX1_333 ( .A(_abc_40344_n1899), .Y(_abc_40344_n2957) );
  INVX1 INVX1_334 ( .A(_abc_40344_n2959), .Y(_abc_40344_n2960) );
  INVX1 INVX1_335 ( .A(_abc_40344_n2961), .Y(_abc_40344_n2962) );
  INVX1 INVX1_336 ( .A(_abc_40344_n2970), .Y(_abc_40344_n2971) );
  INVX1 INVX1_337 ( .A(_abc_40344_n2972), .Y(_abc_40344_n2973) );
  INVX1 INVX1_338 ( .A(_abc_40344_n2979), .Y(_abc_40344_n2980) );
  INVX1 INVX1_339 ( .A(_abc_40344_n2985), .Y(_abc_40344_n2986) );
  INVX1 INVX1_34 ( .A(REG2_REG_5_), .Y(_abc_40344_n756) );
  INVX1 INVX1_340 ( .A(_abc_40344_n1176), .Y(_abc_40344_n2991) );
  INVX1 INVX1_341 ( .A(_abc_40344_n2994), .Y(_abc_40344_n2995) );
  INVX1 INVX1_342 ( .A(_abc_40344_n3003), .Y(_abc_40344_n3004) );
  INVX1 INVX1_343 ( .A(_abc_40344_n2878), .Y(_abc_40344_n3008) );
  INVX1 INVX1_344 ( .A(ADDR_REG_17_), .Y(_abc_40344_n3009) );
  INVX1 INVX1_345 ( .A(_abc_40344_n1758), .Y(_abc_40344_n3010) );
  INVX1 INVX1_346 ( .A(_abc_40344_n3016), .Y(_abc_40344_n3039) );
  INVX1 INVX1_347 ( .A(_abc_40344_n3026), .Y(_abc_40344_n3053) );
  INVX1 INVX1_348 ( .A(_abc_40344_n3061), .Y(_abc_40344_n3062) );
  INVX1 INVX1_349 ( .A(_abc_40344_n3084), .Y(_abc_40344_n3085) );
  INVX1 INVX1_35 ( .A(REG1_REG_5_), .Y(_abc_40344_n757) );
  INVX1 INVX1_350 ( .A(DATAI_20_), .Y(_abc_40344_n3087) );
  INVX1 INVX1_351 ( .A(_abc_40344_n3088), .Y(_abc_40344_n3089) );
  INVX1 INVX1_352 ( .A(_abc_40344_n3093), .Y(_abc_40344_n3094) );
  INVX1 INVX1_353 ( .A(_abc_40344_n3104), .Y(_abc_40344_n3105) );
  INVX1 INVX1_354 ( .A(_abc_40344_n2523_1), .Y(_abc_40344_n3123) );
  INVX1 INVX1_355 ( .A(_abc_40344_n2492), .Y(_abc_40344_n3124) );
  INVX1 INVX1_356 ( .A(_abc_40344_n2476), .Y(_abc_40344_n3125_1) );
  INVX1 INVX1_357 ( .A(_abc_40344_n3129), .Y(_abc_40344_n3132) );
  INVX1 INVX1_358 ( .A(_abc_40344_n3133), .Y(_abc_40344_n3134) );
  INVX1 INVX1_359 ( .A(_abc_40344_n2500), .Y(_abc_40344_n3163) );
  INVX1 INVX1_36 ( .A(_abc_40344_n767), .Y(_abc_40344_n768) );
  INVX1 INVX1_360 ( .A(_abc_40344_n3164), .Y(_abc_40344_n3171) );
  INVX1 INVX1_361 ( .A(_abc_40344_n3172_1), .Y(_abc_40344_n3173) );
  INVX1 INVX1_362 ( .A(_abc_40344_n3200), .Y(_abc_40344_n3201) );
  INVX1 INVX1_363 ( .A(_abc_40344_n1487), .Y(_abc_40344_n3204) );
  INVX1 INVX1_364 ( .A(_abc_40344_n3205), .Y(_abc_40344_n3206) );
  INVX1 INVX1_365 ( .A(_abc_40344_n3209), .Y(_abc_40344_n3210) );
  INVX1 INVX1_366 ( .A(_abc_40344_n3216), .Y(_abc_40344_n3217) );
  INVX1 INVX1_367 ( .A(_abc_40344_n3095), .Y(_abc_40344_n3237) );
  INVX1 INVX1_368 ( .A(_abc_40344_n3245), .Y(_abc_40344_n3246) );
  INVX1 INVX1_369 ( .A(_abc_40344_n2518), .Y(_abc_40344_n3262) );
  INVX1 INVX1_37 ( .A(DATAI_3_), .Y(_abc_40344_n812) );
  INVX1 INVX1_370 ( .A(_abc_40344_n2525), .Y(_abc_40344_n3298) );
  INVX1 INVX1_371 ( .A(_abc_40344_n3304), .Y(_abc_40344_n3305) );
  INVX1 INVX1_372 ( .A(_abc_40344_n1971), .Y(_abc_40344_n3306) );
  INVX1 INVX1_373 ( .A(_abc_40344_n2614), .Y(_abc_40344_n3311) );
  INVX1 INVX1_374 ( .A(_abc_40344_n1952), .Y(_abc_40344_n3331) );
  INVX1 INVX1_375 ( .A(_abc_40344_n3343), .Y(_abc_40344_n3344) );
  INVX1 INVX1_376 ( .A(_abc_40344_n3326), .Y(_abc_40344_n3355) );
  INVX1 INVX1_377 ( .A(_abc_40344_n3329), .Y(_abc_40344_n3358) );
  INVX1 INVX1_378 ( .A(_abc_40344_n3359_1), .Y(_abc_40344_n3360) );
  INVX1 INVX1_379 ( .A(_abc_40344_n2515), .Y(_abc_40344_n3363) );
  INVX1 INVX1_38 ( .A(_abc_40344_n816), .Y(_abc_40344_n817) );
  INVX1 INVX1_380 ( .A(_abc_40344_n2470), .Y(_abc_40344_n3398) );
  INVX1 INVX1_381 ( .A(_abc_40344_n3184), .Y(_abc_40344_n3403) );
  INVX1 INVX1_382 ( .A(_abc_40344_n3190), .Y(_abc_40344_n3404) );
  INVX1 INVX1_383 ( .A(_abc_40344_n3193), .Y(_abc_40344_n3405) );
  INVX1 INVX1_384 ( .A(_abc_40344_n3406), .Y(_abc_40344_n3407) );
  INVX1 INVX1_385 ( .A(_abc_40344_n3086), .Y(_abc_40344_n3423) );
  INVX1 INVX1_386 ( .A(_abc_40344_n3433), .Y(_abc_40344_n3434) );
  INVX1 INVX1_387 ( .A(_abc_40344_n3445), .Y(_abc_40344_n3455) );
  INVX1 INVX1_388 ( .A(_abc_40344_n3459), .Y(_abc_40344_n3460) );
  INVX1 INVX1_389 ( .A(_abc_40344_n3465), .Y(_abc_40344_n3466) );
  INVX1 INVX1_39 ( .A(DATAI_2_), .Y(_abc_40344_n819) );
  INVX1 INVX1_390 ( .A(_abc_40344_n3473), .Y(_abc_40344_n3474) );
  INVX1 INVX1_391 ( .A(_abc_40344_n3488), .Y(_abc_40344_n3489) );
  INVX1 INVX1_392 ( .A(_abc_40344_n3492), .Y(_abc_40344_n3493) );
  INVX1 INVX1_393 ( .A(_abc_40344_n3511), .Y(_abc_40344_n3512) );
  INVX1 INVX1_394 ( .A(_abc_40344_n3159), .Y(_abc_40344_n3518) );
  INVX1 INVX1_395 ( .A(_abc_40344_n3508), .Y(_abc_40344_n3525) );
  INVX1 INVX1_396 ( .A(_abc_40344_n3530), .Y(_abc_40344_n3531) );
  INVX1 INVX1_397 ( .A(_abc_40344_n3527), .Y(_abc_40344_n3545) );
  INVX1 INVX1_398 ( .A(_abc_40344_n3547), .Y(_abc_40344_n3548) );
  INVX1 INVX1_399 ( .A(_abc_40344_n3079), .Y(_abc_40344_n3574) );
  INVX1 INVX1_4 ( .A(IR_REG_13_), .Y(_abc_40344_n530) );
  INVX1 INVX1_40 ( .A(_abc_40344_n830), .Y(_abc_40344_n831) );
  INVX1 INVX1_400 ( .A(_abc_40344_n3581_1), .Y(_abc_40344_n3584) );
  INVX1 INVX1_401 ( .A(_abc_40344_n3593), .Y(_abc_40344_n3594) );
  INVX1 INVX1_402 ( .A(_abc_40344_n3596), .Y(_abc_40344_n3597) );
  INVX1 INVX1_403 ( .A(_abc_40344_n2475), .Y(_abc_40344_n3612) );
  INVX1 INVX1_404 ( .A(_abc_40344_n3621), .Y(_abc_40344_n3622) );
  INVX1 INVX1_405 ( .A(_abc_40344_n3077), .Y(_abc_40344_n3623) );
  INVX1 INVX1_406 ( .A(_abc_40344_n3630), .Y(_abc_40344_n3631) );
  INVX1 INVX1_407 ( .A(_abc_40344_n3636), .Y(_abc_40344_n3637) );
  INVX1 INVX1_408 ( .A(_abc_40344_n3639), .Y(_abc_40344_n3640) );
  INVX1 INVX1_409 ( .A(_abc_40344_n1985), .Y(_abc_40344_n3651) );
  INVX1 INVX1_41 ( .A(REG1_REG_2_), .Y(_abc_40344_n836) );
  INVX1 INVX1_410 ( .A(_abc_40344_n3654), .Y(_abc_40344_n3655) );
  INVX1 INVX1_411 ( .A(_abc_40344_n3660), .Y(_abc_40344_n3661) );
  INVX1 INVX1_412 ( .A(_abc_40344_n3075), .Y(_abc_40344_n3663) );
  INVX1 INVX1_413 ( .A(_abc_40344_n3671), .Y(_abc_40344_n3672) );
  INVX1 INVX1_414 ( .A(_abc_40344_n3674), .Y(_abc_40344_n3675) );
  INVX1 INVX1_415 ( .A(_abc_40344_n3688), .Y(_abc_40344_n3689) );
  INVX1 INVX1_416 ( .A(_abc_40344_n3146), .Y(_abc_40344_n3703) );
  INVX1 INVX1_417 ( .A(_abc_40344_n3711), .Y(_abc_40344_n3712) );
  INVX1 INVX1_418 ( .A(_abc_40344_n3719), .Y(_abc_40344_n3720) );
  INVX1 INVX1_419 ( .A(_abc_40344_n3307), .Y(_abc_40344_n3741) );
  INVX1 INVX1_42 ( .A(REG0_REG_2_), .Y(_abc_40344_n837) );
  INVX1 INVX1_420 ( .A(_abc_40344_n3744), .Y(_abc_40344_n3745) );
  INVX1 INVX1_421 ( .A(_abc_40344_n2529_1), .Y(_abc_40344_n3784_1) );
  INVX1 INVX1_422 ( .A(_abc_40344_n3786_1), .Y(_abc_40344_n3787_1) );
  INVX1 INVX1_423 ( .A(_abc_40344_n3796_1), .Y(n493) );
  INVX1 INVX1_424 ( .A(_abc_40344_n3798_1), .Y(n488) );
  INVX1 INVX1_425 ( .A(_abc_40344_n3800), .Y(n483) );
  INVX1 INVX1_426 ( .A(_abc_40344_n3802), .Y(n478) );
  INVX1 INVX1_427 ( .A(_abc_40344_n3804), .Y(n473) );
  INVX1 INVX1_428 ( .A(_abc_40344_n3806), .Y(n468) );
  INVX1 INVX1_429 ( .A(_abc_40344_n3808), .Y(n463) );
  INVX1 INVX1_43 ( .A(DATAI_1_), .Y(_abc_40344_n848) );
  INVX1 INVX1_430 ( .A(_abc_40344_n3810_1), .Y(n458) );
  INVX1 INVX1_431 ( .A(_abc_40344_n3812), .Y(n453) );
  INVX1 INVX1_432 ( .A(_abc_40344_n3814), .Y(n448) );
  INVX1 INVX1_433 ( .A(_abc_40344_n3816), .Y(n443) );
  INVX1 INVX1_434 ( .A(_abc_40344_n3818), .Y(n438) );
  INVX1 INVX1_435 ( .A(_abc_40344_n3820), .Y(n433) );
  INVX1 INVX1_436 ( .A(_abc_40344_n3822), .Y(n428) );
  INVX1 INVX1_437 ( .A(_abc_40344_n3824_1), .Y(n423) );
  INVX1 INVX1_438 ( .A(_abc_40344_n3826), .Y(n418) );
  INVX1 INVX1_439 ( .A(_abc_40344_n3828), .Y(n413) );
  INVX1 INVX1_44 ( .A(_abc_40344_n849_1), .Y(_abc_40344_n850_1) );
  INVX1 INVX1_440 ( .A(_abc_40344_n3830_1), .Y(n408) );
  INVX1 INVX1_441 ( .A(_abc_40344_n3832), .Y(n403) );
  INVX1 INVX1_442 ( .A(_abc_40344_n3834), .Y(n398) );
  INVX1 INVX1_443 ( .A(_abc_40344_n3836_1), .Y(n393) );
  INVX1 INVX1_444 ( .A(_abc_40344_n3838), .Y(n388) );
  INVX1 INVX1_445 ( .A(_abc_40344_n3840), .Y(n383) );
  INVX1 INVX1_446 ( .A(_abc_40344_n3842_1), .Y(n378) );
  INVX1 INVX1_447 ( .A(_abc_40344_n3844), .Y(n373) );
  INVX1 INVX1_448 ( .A(_abc_40344_n3846_1), .Y(n368) );
  INVX1 INVX1_449 ( .A(_abc_40344_n3848), .Y(n363) );
  INVX1 INVX1_45 ( .A(_abc_40344_n853), .Y(_abc_40344_n854_1) );
  INVX1 INVX1_450 ( .A(_abc_40344_n3850), .Y(n358) );
  INVX1 INVX1_451 ( .A(_abc_40344_n3852_1), .Y(n353) );
  INVX1 INVX1_452 ( .A(_abc_40344_n3854), .Y(n348) );
  INVX1 INVX1_453 ( .A(_abc_40344_n3863), .Y(_abc_40344_n3864_1) );
  INVX1 INVX1_454 ( .A(_abc_40344_n3868_1), .Y(_abc_40344_n3869) );
  INVX1 INVX1_455 ( .A(_abc_40344_n3876), .Y(_abc_40344_n3877_1) );
  INVX1 INVX1_456 ( .A(_abc_40344_n3881), .Y(_abc_40344_n3882) );
  INVX1 INVX1_457 ( .A(_abc_40344_n3886_1), .Y(_abc_40344_n3887) );
  INVX1 INVX1_458 ( .A(_abc_40344_n3892), .Y(_abc_40344_n3893_1) );
  INVX1 INVX1_459 ( .A(_abc_40344_n3899), .Y(_abc_40344_n3900_1) );
  INVX1 INVX1_46 ( .A(REG0_REG_1_), .Y(_abc_40344_n857) );
  INVX1 INVX1_460 ( .A(_abc_40344_n3903), .Y(_abc_40344_n3904) );
  INVX1 INVX1_461 ( .A(_abc_40344_n638), .Y(_abc_40344_n3906) );
  INVX1 INVX1_462 ( .A(_abc_40344_n3909), .Y(_abc_40344_n3910) );
  INVX1 INVX1_463 ( .A(_abc_40344_n3913), .Y(_abc_40344_n3914) );
  INVX1 INVX1_464 ( .A(_abc_40344_n1120), .Y(_abc_40344_n3916) );
  INVX1 INVX1_465 ( .A(_abc_40344_n3918), .Y(_abc_40344_n3919) );
  INVX1 INVX1_466 ( .A(IR_REG_17_), .Y(_abc_40344_n3921) );
  INVX1 INVX1_467 ( .A(_abc_40344_n3923), .Y(_abc_40344_n3924) );
  INVX1 INVX1_468 ( .A(_abc_40344_n1146), .Y(_abc_40344_n3926) );
  INVX1 INVX1_469 ( .A(_abc_40344_n3928), .Y(_abc_40344_n3929) );
  INVX1 INVX1_47 ( .A(REG1_REG_1_), .Y(_abc_40344_n860) );
  INVX1 INVX1_470 ( .A(_abc_40344_n3932), .Y(_abc_40344_n3933) );
  INVX1 INVX1_471 ( .A(IR_REG_14_), .Y(_abc_40344_n3935) );
  INVX1 INVX1_472 ( .A(_abc_40344_n3937), .Y(_abc_40344_n3938) );
  INVX1 INVX1_473 ( .A(_abc_40344_n1248), .Y(_abc_40344_n3940) );
  INVX1 INVX1_474 ( .A(_abc_40344_n3942), .Y(_abc_40344_n3943) );
  INVX1 INVX1_475 ( .A(_abc_40344_n3946), .Y(_abc_40344_n3947) );
  INVX1 INVX1_476 ( .A(IR_REG_11_), .Y(_abc_40344_n3949) );
  INVX1 INVX1_477 ( .A(_abc_40344_n3951_1), .Y(_abc_40344_n3952) );
  INVX1 INVX1_478 ( .A(_abc_40344_n3955), .Y(_abc_40344_n3956_1) );
  INVX1 INVX1_479 ( .A(_abc_40344_n1344), .Y(_abc_40344_n3958_1) );
  INVX1 INVX1_48 ( .A(_abc_40344_n865), .Y(_abc_40344_n875) );
  INVX1 INVX1_480 ( .A(_abc_40344_n3960), .Y(_abc_40344_n3961) );
  INVX1 INVX1_481 ( .A(_abc_40344_n3964), .Y(_abc_40344_n3965) );
  INVX1 INVX1_482 ( .A(_abc_40344_n3968), .Y(_abc_40344_n3969) );
  INVX1 INVX1_483 ( .A(_abc_40344_n3972_1), .Y(_abc_40344_n3973) );
  INVX1 INVX1_484 ( .A(_abc_40344_n3976), .Y(_abc_40344_n3977) );
  INVX1 INVX1_485 ( .A(_abc_40344_n3980), .Y(_abc_40344_n3981) );
  INVX1 INVX1_486 ( .A(_abc_40344_n3984), .Y(_abc_40344_n3985_1) );
  INVX1 INVX1_487 ( .A(_abc_40344_n3988), .Y(_abc_40344_n3989) );
  INVX1 INVX1_488 ( .A(_abc_40344_n3992_1), .Y(_abc_40344_n3993) );
  INVX1 INVX1_489 ( .A(_abc_40344_n3997), .Y(_abc_40344_n3998) );
  INVX1 INVX1_49 ( .A(DATAI_0_), .Y(_abc_40344_n877_1) );
  INVX1 INVX1_490 ( .A(_abc_40344_n2558), .Y(_abc_40344_n4000) );
  INVX1 INVX1_491 ( .A(_abc_40344_n3122), .Y(_abc_40344_n4002) );
  INVX1 INVX1_492 ( .A(_abc_40344_n2651), .Y(_abc_40344_n4011) );
  INVX1 INVX1_493 ( .A(D_REG_0_), .Y(_abc_40344_n4031) );
  INVX1 INVX1_494 ( .A(D_REG_1_), .Y(_abc_40344_n4035) );
  INVX1 INVX1_495 ( .A(REG0_REG_17_), .Y(_abc_40344_n4144) );
  INVX1 INVX1_496 ( .A(_abc_40344_n3446), .Y(_abc_40344_n4157) );
  INVX1 INVX1_497 ( .A(_abc_40344_n3425), .Y(_abc_40344_n4164) );
  INVX1 INVX1_5 ( .A(IR_REG_2_), .Y(_abc_40344_n536) );
  INVX1 INVX1_50 ( .A(REG0_REG_0_), .Y(_abc_40344_n884) );
  INVX1 INVX1_51 ( .A(_abc_40344_n900), .Y(_abc_40344_n901) );
  INVX1 INVX1_52 ( .A(DATAI_7_), .Y(_abc_40344_n902_1) );
  INVX1 INVX1_53 ( .A(REG3_REG_7_), .Y(_abc_40344_n910) );
  INVX1 INVX1_54 ( .A(REG2_REG_7_), .Y(_abc_40344_n920) );
  INVX1 INVX1_55 ( .A(_abc_40344_n912), .Y(_abc_40344_n922_1) );
  INVX1 INVX1_56 ( .A(REG1_REG_7_), .Y(_abc_40344_n924) );
  INVX1 INVX1_57 ( .A(REG0_REG_7_), .Y(_abc_40344_n925) );
  INVX1 INVX1_58 ( .A(_abc_40344_n934), .Y(_abc_40344_n938) );
  INVX1 INVX1_59 ( .A(_abc_40344_n933), .Y(_abc_40344_n940) );
  INVX1 INVX1_6 ( .A(IR_REG_1_), .Y(_abc_40344_n537_1) );
  INVX1 INVX1_60 ( .A(_abc_40344_n943_1), .Y(_abc_40344_n944) );
  INVX1 INVX1_61 ( .A(B_REG), .Y(_abc_40344_n945_1) );
  INVX1 INVX1_62 ( .A(_abc_40344_n565_1), .Y(_abc_40344_n947) );
  INVX1 INVX1_63 ( .A(_abc_40344_n942), .Y(_abc_40344_n948_1) );
  INVX1 INVX1_64 ( .A(_abc_40344_n950), .Y(_abc_40344_n952) );
  INVX1 INVX1_65 ( .A(_abc_40344_n989), .Y(_abc_40344_n998) );
  INVX1 INVX1_66 ( .A(_abc_40344_n1000), .Y(_abc_40344_n1001) );
  INVX1 INVX1_67 ( .A(_abc_40344_n987), .Y(_abc_40344_n1002) );
  INVX1 INVX1_68 ( .A(_abc_40344_n1003), .Y(_abc_40344_n1004) );
  INVX1 INVX1_69 ( .A(REG0_REG_8_), .Y(_abc_40344_n1008) );
  INVX1 INVX1_7 ( .A(_abc_40344_n551), .Y(_abc_40344_n552) );
  INVX1 INVX1_70 ( .A(_abc_40344_n1015), .Y(_abc_40344_n1016) );
  INVX1 INVX1_71 ( .A(_abc_40344_n1026), .Y(_abc_40344_n1027_1) );
  INVX1 INVX1_72 ( .A(REG3_REG_26_), .Y(_abc_40344_n1041) );
  INVX1 INVX1_73 ( .A(REG3_REG_27_), .Y(_abc_40344_n1042) );
  INVX1 INVX1_74 ( .A(REG3_REG_25_), .Y(_abc_40344_n1044) );
  INVX1 INVX1_75 ( .A(REG3_REG_21_), .Y(_abc_40344_n1045_1) );
  INVX1 INVX1_76 ( .A(REG3_REG_13_), .Y(_abc_40344_n1049_1) );
  INVX1 INVX1_77 ( .A(REG3_REG_11_), .Y(_abc_40344_n1053) );
  INVX1 INVX1_78 ( .A(_abc_40344_n1064), .Y(_abc_40344_n1065) );
  INVX1 INVX1_79 ( .A(REG1_REG_27_), .Y(_abc_40344_n1069) );
  INVX1 INVX1_8 ( .A(IR_REG_26_), .Y(_abc_40344_n554_1) );
  INVX1 INVX1_80 ( .A(_abc_40344_n1079), .Y(_abc_40344_n1080) );
  INVX1 INVX1_81 ( .A(REG2_REG_23_), .Y(_abc_40344_n1087) );
  INVX1 INVX1_82 ( .A(_abc_40344_n1094), .Y(_abc_40344_n1095) );
  INVX1 INVX1_83 ( .A(REG3_REG_22_), .Y(_abc_40344_n1101) );
  INVX1 INVX1_84 ( .A(_abc_40344_n1112), .Y(_abc_40344_n1113) );
  INVX1 INVX1_85 ( .A(_abc_40344_n1117), .Y(_abc_40344_n1118_1) );
  INVX1 INVX1_86 ( .A(_abc_40344_n1127), .Y(_abc_40344_n1128) );
  INVX1 INVX1_87 ( .A(REG1_REG_18_), .Y(_abc_40344_n1132_1) );
  INVX1 INVX1_88 ( .A(_abc_40344_n1135_1), .Y(_abc_40344_n1136) );
  INVX1 INVX1_89 ( .A(_abc_40344_n1142), .Y(_abc_40344_n1143) );
  INVX1 INVX1_9 ( .A(IR_REG_24_), .Y(_abc_40344_n563_1) );
  INVX1 INVX1_90 ( .A(DATAI_16_), .Y(_abc_40344_n1150) );
  INVX1 INVX1_91 ( .A(REG3_REG_15_), .Y(_abc_40344_n1154_1) );
  INVX1 INVX1_92 ( .A(REG3_REG_16_), .Y(_abc_40344_n1155_1) );
  INVX1 INVX1_93 ( .A(_abc_40344_n1158), .Y(_abc_40344_n1159) );
  INVX1 INVX1_94 ( .A(_abc_40344_n1160), .Y(_abc_40344_n1161) );
  INVX1 INVX1_95 ( .A(REG2_REG_16_), .Y(_abc_40344_n1164) );
  INVX1 INVX1_96 ( .A(REG2_REG_17_), .Y(_abc_40344_n1182) );
  INVX1 INVX1_97 ( .A(REG1_REG_17_), .Y(_abc_40344_n1183) );
  INVX1 INVX1_98 ( .A(_abc_40344_n1187), .Y(_abc_40344_n1188) );
  INVX1 INVX1_99 ( .A(_abc_40344_n1193_1), .Y(_abc_40344_n1194) );
  INVX2 INVX2_1 ( .A(IR_REG_0_), .Y(_abc_40344_n538_1) );
  INVX2 INVX2_10 ( .A(_abc_40344_n773), .Y(_abc_40344_n774) );
  INVX2 INVX2_11 ( .A(_abc_40344_n808), .Y(_abc_40344_n809) );
  INVX2 INVX2_12 ( .A(_abc_40344_n863), .Y(_abc_40344_n864) );
  INVX2 INVX2_13 ( .A(REG1_REG_0_), .Y(_abc_40344_n885) );
  INVX2 INVX2_14 ( .A(_abc_40344_n906_1), .Y(_abc_40344_n917) );
  INVX2 INVX2_15 ( .A(_abc_40344_n982), .Y(_abc_40344_n983) );
  INVX2 INVX2_16 ( .A(_abc_40344_n985), .Y(_abc_40344_n986) );
  INVX2 INVX2_17 ( .A(_abc_40344_n990), .Y(_abc_40344_n991) );
  INVX2 INVX2_18 ( .A(_abc_40344_n1005), .Y(_abc_40344_n1006) );
  INVX2 INVX2_19 ( .A(REG1_REG_8_), .Y(_abc_40344_n1007) );
  INVX2 INVX2_2 ( .A(_abc_40344_n549_1), .Y(_abc_40344_n555) );
  INVX2 INVX2_20 ( .A(REG2_REG_8_), .Y(_abc_40344_n1010) );
  INVX2 INVX2_21 ( .A(REG3_REG_8_), .Y(_abc_40344_n1011) );
  INVX2 INVX2_22 ( .A(_abc_40344_n1018), .Y(_abc_40344_n1019) );
  INVX2 INVX2_23 ( .A(_abc_40344_n698), .Y(_abc_40344_n1021) );
  INVX2 INVX2_24 ( .A(_abc_40344_n1028), .Y(_abc_40344_n1029_1) );
  INVX2 INVX2_25 ( .A(_abc_40344_n650), .Y(_abc_40344_n1039) );
  INVX2 INVX2_26 ( .A(REG3_REG_24_), .Y(_abc_40344_n1043) );
  INVX2 INVX2_27 ( .A(REG3_REG_20_), .Y(_abc_40344_n1046) );
  INVX2 INVX2_28 ( .A(REG3_REG_18_), .Y(_abc_40344_n1047) );
  INVX2 INVX2_29 ( .A(REG3_REG_10_), .Y(_abc_40344_n1052_1) );
  INVX2 INVX2_3 ( .A(IR_REG_25_), .Y(_abc_40344_n566) );
  INVX2 INVX2_30 ( .A(_abc_40344_n1083), .Y(_abc_40344_n1084) );
  INVX2 INVX2_31 ( .A(_abc_40344_n1090_1), .Y(_abc_40344_n1091) );
  INVX2 INVX2_32 ( .A(_abc_40344_n1097), .Y(_abc_40344_n1098) );
  INVX2 INVX2_33 ( .A(_abc_40344_n1110), .Y(_abc_40344_n1111) );
  INVX2 INVX2_34 ( .A(IR_REG_18_), .Y(_abc_40344_n1119) );
  INVX2 INVX2_35 ( .A(REG2_REG_18_), .Y(_abc_40344_n1131) );
  INVX2 INVX2_36 ( .A(_abc_40344_n1124), .Y(_abc_40344_n1137) );
  INVX2 INVX2_37 ( .A(IR_REG_16_), .Y(_abc_40344_n1144) );
  INVX2 INVX2_38 ( .A(_abc_40344_n1148), .Y(_abc_40344_n1149) );
  INVX2 INVX2_39 ( .A(_abc_40344_n1152_1), .Y(_abc_40344_n1153) );
  INVX2 INVX2_4 ( .A(_abc_40344_n618), .Y(_abc_40344_n619) );
  INVX2 INVX2_40 ( .A(REG1_REG_16_), .Y(_abc_40344_n1165) );
  INVX2 INVX2_41 ( .A(_abc_40344_n1167), .Y(_abc_40344_n1168) );
  INVX2 INVX2_42 ( .A(_abc_40344_n1185), .Y(_abc_40344_n1186) );
  INVX2 INVX2_43 ( .A(_abc_40344_n1196), .Y(_abc_40344_n1197) );
  INVX2 INVX2_44 ( .A(REG1_REG_15_), .Y(_abc_40344_n1206) );
  INVX2 INVX2_45 ( .A(_abc_40344_n1209_1), .Y(_abc_40344_n1210) );
  INVX2 INVX2_46 ( .A(_abc_40344_n1221), .Y(_abc_40344_n1222) );
  INVX2 INVX2_47 ( .A(REG1_REG_14_), .Y(_abc_40344_n1232) );
  INVX2 INVX2_48 ( .A(REG1_REG_12_), .Y(_abc_40344_n1296) );
  INVX2 INVX2_49 ( .A(_abc_40344_n1305), .Y(_abc_40344_n1309) );
  INVX2 INVX2_5 ( .A(_abc_40344_n625), .Y(_abc_40344_n626) );
  INVX2 INVX2_50 ( .A(_abc_40344_n1347), .Y(_abc_40344_n1348) );
  INVX2 INVX2_51 ( .A(REG2_REG_9_), .Y(_abc_40344_n1354) );
  INVX2 INVX2_52 ( .A(_abc_40344_n1440), .Y(_abc_40344_n1441) );
  INVX2 INVX2_53 ( .A(_abc_40344_n1506), .Y(_abc_40344_n1507_1) );
  INVX2 INVX2_54 ( .A(REG3_REG_28_), .Y(_abc_40344_n1538) );
  INVX2 INVX2_55 ( .A(_abc_40344_n1548), .Y(_abc_40344_n1549) );
  INVX2 INVX2_56 ( .A(_abc_40344_n1471), .Y(_abc_40344_n1577) );
  INVX2 INVX2_57 ( .A(_abc_40344_n1032), .Y(_abc_40344_n1580) );
  INVX2 INVX2_58 ( .A(_abc_40344_n797), .Y(_abc_40344_n1607) );
  INVX2 INVX2_59 ( .A(_abc_40344_n1645), .Y(_abc_40344_n1646) );
  INVX2 INVX2_6 ( .A(_abc_40344_n640), .Y(_abc_40344_n641) );
  INVX2 INVX2_60 ( .A(_abc_40344_n1234), .Y(_abc_40344_n1818) );
  INVX2 INVX2_61 ( .A(DATAI_24_), .Y(_abc_40344_n1933) );
  INVX2 INVX2_62 ( .A(_abc_40344_n1178), .Y(_abc_40344_n1949) );
  INVX2 INVX2_63 ( .A(_abc_40344_n1953), .Y(_abc_40344_n1954) );
  INVX2 INVX2_64 ( .A(_abc_40344_n1224), .Y(_abc_40344_n1961) );
  INVX2 INVX2_65 ( .A(_abc_40344_n823), .Y(_abc_40344_n2020) );
  INVX2 INVX2_66 ( .A(_abc_40344_n2095), .Y(_abc_40344_n2096) );
  INVX2 INVX2_67 ( .A(_abc_40344_n2100), .Y(_abc_40344_n2101) );
  INVX2 INVX2_68 ( .A(_abc_40344_n2121), .Y(_abc_40344_n2122) );
  INVX2 INVX2_69 ( .A(_abc_40344_n1926), .Y(_abc_40344_n2394) );
  INVX2 INVX2_7 ( .A(REG3_REG_3_), .Y(_abc_40344_n688_1) );
  INVX2 INVX2_70 ( .A(_abc_40344_n1922), .Y(_abc_40344_n2401) );
  INVX2 INVX2_71 ( .A(_abc_40344_n1932), .Y(_abc_40344_n2513) );
  INVX2 INVX2_72 ( .A(_abc_40344_n2520), .Y(_abc_40344_n2521) );
  INVX2 INVX2_73 ( .A(_abc_40344_n2666_1), .Y(_abc_40344_n2667) );
  INVX2 INVX2_74 ( .A(n1341), .Y(_abc_40344_n2673) );
  INVX2 INVX2_75 ( .A(_abc_40344_n2705), .Y(_abc_40344_n2706) );
  INVX2 INVX2_76 ( .A(REG1_REG_4_), .Y(_abc_40344_n2748) );
  INVX2 INVX2_77 ( .A(_abc_40344_n1271), .Y(_abc_40344_n2863) );
  INVX2 INVX2_78 ( .A(_abc_40344_n2870), .Y(_abc_40344_n2871) );
  INVX2 INVX2_79 ( .A(_abc_40344_n1122), .Y(_abc_40344_n3017) );
  INVX2 INVX2_8 ( .A(_abc_40344_n708), .Y(_abc_40344_n709) );
  INVX2 INVX2_80 ( .A(_abc_40344_n2556), .Y(_abc_40344_n3120) );
  INVX2 INVX2_81 ( .A(_abc_40344_n3220), .Y(_abc_40344_n3379) );
  INVX2 INVX2_82 ( .A(_abc_40344_n2543_1), .Y(_abc_40344_n3478_1) );
  INVX2 INVX2_9 ( .A(_abc_40344_n732_1), .Y(_abc_40344_n748) );
  INVX4 INVX4_1 ( .A(STATE_REG), .Y(_abc_40344_n523) );
  INVX4 INVX4_10 ( .A(_abc_40344_n1200), .Y(_abc_40344_n1201) );
  INVX4 INVX4_11 ( .A(_abc_40344_n1259), .Y(_abc_40344_n1260) );
  INVX4 INVX4_12 ( .A(_abc_40344_n1284), .Y(_abc_40344_n1285) );
  INVX4 INVX4_13 ( .A(_abc_40344_n1361), .Y(_abc_40344_n1362) );
  INVX4 INVX4_14 ( .A(_abc_40344_n1404), .Y(_abc_40344_n1418) );
  INVX4 INVX4_15 ( .A(_abc_40344_n1433), .Y(_abc_40344_n1434) );
  INVX4 INVX4_16 ( .A(_abc_40344_n1462), .Y(_abc_40344_n1463) );
  INVX4 INVX4_17 ( .A(_abc_40344_n1488), .Y(_abc_40344_n1489) );
  INVX4 INVX4_18 ( .A(_abc_40344_n1477), .Y(_abc_40344_n1491) );
  INVX4 INVX4_19 ( .A(_abc_40344_n1494), .Y(_abc_40344_n1495) );
  INVX4 INVX4_2 ( .A(_abc_40344_n646), .Y(_abc_40344_n648) );
  INVX4 INVX4_20 ( .A(_abc_40344_n993), .Y(_abc_40344_n1590) );
  INVX4 INVX4_21 ( .A(_abc_40344_n1630), .Y(_abc_40344_n1649) );
  INVX4 INVX4_22 ( .A(_abc_40344_n3068), .Y(_abc_40344_n3069) );
  INVX4 INVX4_23 ( .A(_abc_40344_n3110), .Y(_abc_40344_n3111) );
  INVX4 INVX4_24 ( .A(_abc_40344_n3233), .Y(_abc_40344_n3244) );
  INVX4 INVX4_25 ( .A(_abc_40344_n3223), .Y(_abc_40344_n3261) );
  INVX4 INVX4_26 ( .A(_abc_40344_n3725), .Y(_abc_40344_n3726) );
  INVX4 INVX4_27 ( .A(_abc_40344_n4040_1), .Y(_abc_40344_n4041) );
  INVX4 INVX4_28 ( .A(_abc_40344_n4237), .Y(_abc_40344_n4238_1) );
  INVX4 INVX4_3 ( .A(_abc_40344_n776), .Y(_abc_40344_n777_1) );
  INVX4 INVX4_4 ( .A(_abc_40344_n785), .Y(_abc_40344_n787_1) );
  INVX4 INVX4_5 ( .A(_abc_40344_n979), .Y(_abc_40344_n980) );
  INVX4 INVX4_6 ( .A(_abc_40344_n627), .Y(_abc_40344_n984) );
  INVX4 INVX4_7 ( .A(_abc_40344_n1073), .Y(_abc_40344_n1074) );
  INVX4 INVX4_8 ( .A(_abc_40344_n1040), .Y(_abc_40344_n1076) );
  INVX4 INVX4_9 ( .A(_abc_40344_n1099), .Y(_abc_40344_n1100) );
  INVX8 INVX8_1 ( .A(IR_REG_31_), .Y(_abc_40344_n559_1) );
  INVX8 INVX8_10 ( .A(n1336), .Y(_abc_40344_n1033) );
  INVX8 INVX8_11 ( .A(_abc_40344_n1020), .Y(_abc_40344_n1537) );
  INVX8 INVX8_12 ( .A(_abc_40344_n1554), .Y(_abc_40344_n1555) );
  INVX8 INVX8_13 ( .A(_abc_40344_n2161), .Y(_abc_40344_n2162) );
  INVX8 INVX8_14 ( .A(_abc_40344_n2172), .Y(_abc_40344_n2173) );
  INVX8 INVX8_15 ( .A(_abc_40344_n2165), .Y(_abc_40344_n2179) );
  INVX8 INVX8_16 ( .A(_abc_40344_n2674), .Y(_abc_40344_n2675) );
  INVX8 INVX8_17 ( .A(_abc_40344_n3066), .Y(_abc_40344_n3067) );
  INVX8 INVX8_18 ( .A(_abc_40344_n995), .Y(_abc_40344_n3109) );
  INVX8 INVX8_19 ( .A(_abc_40344_n3218), .Y(_abc_40344_n3219) );
  INVX8 INVX8_2 ( .A(_abc_40344_n585), .Y(_abc_40344_n586) );
  INVX8 INVX8_20 ( .A(_abc_40344_n3227), .Y(_abc_40344_n3228) );
  INVX8 INVX8_21 ( .A(_abc_40344_n3103), .Y(_abc_40344_n3232) );
  INVX8 INVX8_22 ( .A(_abc_40344_n3856), .Y(_abc_40344_n3857) );
  INVX8 INVX8_23 ( .A(_abc_40344_n3860), .Y(_abc_40344_n3861_1) );
  INVX8 INVX8_24 ( .A(_abc_40344_n4042), .Y(_abc_40344_n4043) );
  INVX8 INVX8_25 ( .A(_abc_40344_n4048), .Y(_abc_40344_n4049) );
  INVX8 INVX8_26 ( .A(n1345), .Y(_abc_40344_n4329_1) );
  INVX8 INVX8_3 ( .A(_abc_40344_n588), .Y(_abc_40344_n589) );
  INVX8 INVX8_4 ( .A(_abc_40344_n602), .Y(_abc_40344_n603) );
  INVX8 INVX8_5 ( .A(_abc_40344_n610_1), .Y(_abc_40344_n611_1) );
  INVX8 INVX8_6 ( .A(nRESET_G), .Y(_abc_40344_n630_1) );
  INVX8 INVX8_7 ( .A(_abc_40344_n719), .Y(_abc_40344_n720) );
  INVX8 INVX8_8 ( .A(_abc_40344_n1022), .Y(_abc_40344_n1023_1) );
  INVX8 INVX8_9 ( .A(_abc_40344_n1030_1), .Y(_abc_40344_n1031) );
  NAND2X1 NAND2X1_1 ( .A(_abc_40344_n524), .B(_abc_40344_n525), .Y(_abc_40344_n526) );
  NAND2X1 NAND2X1_10 ( .A(IR_REG_23_), .B(_abc_40344_n559_1), .Y(_abc_40344_n584_1) );
  NAND2X1 NAND2X1_100 ( .A(REG3_REG_8_), .B(REG3_REG_9_), .Y(_abc_40344_n1050) );
  NAND2X1 NAND2X1_101 ( .A(REG3_REG_19_), .B(_abc_40344_n1059), .Y(_abc_40344_n1060) );
  NAND2X1 NAND2X1_102 ( .A(_abc_40344_n1067), .B(_abc_40344_n1066_1), .Y(_abc_40344_n1068) );
  NAND2X1 NAND2X1_103 ( .A(REG2_REG_27_), .B(_abc_40344_n695), .Y(_abc_40344_n1070) );
  NAND2X1 NAND2X1_104 ( .A(_abc_40344_n1075), .B(_abc_40344_n1078_1), .Y(_abc_40344_n1079) );
  NAND2X1 NAND2X1_105 ( .A(REG3_REG_22_), .B(_abc_40344_n1062), .Y(_abc_40344_n1085) );
  NAND2X1 NAND2X1_106 ( .A(_abc_40344_n1092), .B(_abc_40344_n1095), .Y(_abc_40344_n1096) );
  NAND2X1 NAND2X1_107 ( .A(REG3_REG_21_), .B(_abc_40344_n1102), .Y(_abc_40344_n1103_1) );
  NAND2X1 NAND2X1_108 ( .A(REG0_REG_22_), .B(_abc_40344_n673), .Y(_abc_40344_n1106) );
  NAND2X1 NAND2X1_109 ( .A(REG2_REG_22_), .B(_abc_40344_n695), .Y(_abc_40344_n1107) );
  NAND2X1 NAND2X1_11 ( .A(_abc_40344_n586), .B(_abc_40344_n581), .Y(_abc_40344_n587) );
  NAND2X1 NAND2X1_110 ( .A(REG1_REG_22_), .B(_abc_40344_n696), .Y(_abc_40344_n1108) );
  NAND2X1 NAND2X1_111 ( .A(_abc_40344_n1113), .B(_abc_40344_n1115), .Y(_abc_40344_n1116) );
  NAND2X1 NAND2X1_112 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1119), .Y(_abc_40344_n1121) );
  NAND2X1 NAND2X1_113 ( .A(REG0_REG_18_), .B(_abc_40344_n673), .Y(_abc_40344_n1129) );
  NAND2X1 NAND2X1_114 ( .A(_abc_40344_n1136), .B(_abc_40344_n1140), .Y(_abc_40344_n1141) );
  NAND2X1 NAND2X1_115 ( .A(_abc_40344_n525), .B(_abc_40344_n574), .Y(_abc_40344_n1145) );
  NAND2X1 NAND2X1_116 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1144), .Y(_abc_40344_n1147) );
  NAND2X1 NAND2X1_117 ( .A(REG3_REG_14_), .B(_abc_40344_n1056), .Y(_abc_40344_n1156) );
  NAND2X1 NAND2X1_118 ( .A(REG0_REG_16_), .B(_abc_40344_n673), .Y(_abc_40344_n1162) );
  NAND2X1 NAND2X1_119 ( .A(_abc_40344_n1169), .B(_abc_40344_n1171), .Y(_abc_40344_n1172) );
  NAND2X1 NAND2X1_12 ( .A(_abc_40344_n551), .B(_abc_40344_n594), .Y(_abc_40344_n595_1) );
  NAND2X1 NAND2X1_120 ( .A(IR_REG_31_), .B(_abc_40344_n1174), .Y(_abc_40344_n1175) );
  NAND2X1 NAND2X1_121 ( .A(REG0_REG_17_), .B(_abc_40344_n673), .Y(_abc_40344_n1180_1) );
  NAND2X1 NAND2X1_122 ( .A(IR_REG_31_), .B(_abc_40344_n1194), .Y(_abc_40344_n1195) );
  NAND2X1 NAND2X1_123 ( .A(REG0_REG_15_), .B(_abc_40344_n673), .Y(_abc_40344_n1204) );
  NAND2X1 NAND2X1_124 ( .A(_abc_40344_n1211), .B(_abc_40344_n1214), .Y(_abc_40344_n1217) );
  NAND2X1 NAND2X1_125 ( .A(IR_REG_14_), .B(_abc_40344_n559_1), .Y(_abc_40344_n1220) );
  NAND2X1 NAND2X1_126 ( .A(REG0_REG_14_), .B(_abc_40344_n673), .Y(_abc_40344_n1229) );
  NAND2X1 NAND2X1_127 ( .A(_abc_40344_n1235), .B(_abc_40344_n1238), .Y(_abc_40344_n1239) );
  NAND2X1 NAND2X1_128 ( .A(_abc_40344_n559_1), .B(_abc_40344_n530), .Y(_abc_40344_n1242) );
  NAND2X1 NAND2X1_129 ( .A(_abc_40344_n528), .B(_abc_40344_n1244), .Y(_abc_40344_n1245) );
  NAND2X1 NAND2X1_13 ( .A(_abc_40344_n559_1), .B(_abc_40344_n600_1), .Y(_abc_40344_n601) );
  NAND2X1 NAND2X1_130 ( .A(_abc_40344_n1249), .B(_abc_40344_n705_1), .Y(_abc_40344_n1263) );
  NAND2X1 NAND2X1_131 ( .A(_abc_40344_n1243), .B(_abc_40344_n1246), .Y(_abc_40344_n1268) );
  NAND2X1 NAND2X1_132 ( .A(IR_REG_31_), .B(_abc_40344_n1269), .Y(_abc_40344_n1270) );
  NAND2X1 NAND2X1_133 ( .A(_abc_40344_n1054), .B(_abc_40344_n1051_1), .Y(_abc_40344_n1275) );
  NAND2X1 NAND2X1_134 ( .A(_abc_40344_n1247), .B(_abc_40344_n1290), .Y(_abc_40344_n1291) );
  NAND2X1 NAND2X1_135 ( .A(IR_REG_31_), .B(_abc_40344_n1291), .Y(_abc_40344_n1292) );
  NAND2X1 NAND2X1_136 ( .A(_abc_40344_n705_1), .B(_abc_40344_n1293_1), .Y(_abc_40344_n1294) );
  NAND2X1 NAND2X1_137 ( .A(_abc_40344_n1299), .B(_abc_40344_n1275), .Y(_abc_40344_n1300) );
  NAND2X1 NAND2X1_138 ( .A(REG2_REG_12_), .B(_abc_40344_n695), .Y(_abc_40344_n1303) );
  NAND2X1 NAND2X1_139 ( .A(_abc_40344_n1262), .B(_abc_40344_n1266), .Y(_abc_40344_n1313) );
  NAND2X1 NAND2X1_14 ( .A(_abc_40344_n559_1), .B(_abc_40344_n604), .Y(_abc_40344_n605) );
  NAND2X1 NAND2X1_140 ( .A(_abc_40344_n1306), .B(_abc_40344_n1311), .Y(_abc_40344_n1314) );
  NAND2X1 NAND2X1_141 ( .A(_abc_40344_n1286), .B(_abc_40344_n1288), .Y(_abc_40344_n1318) );
  NAND2X1 NAND2X1_142 ( .A(_abc_40344_n1322), .B(_abc_40344_n1268), .Y(_abc_40344_n1323) );
  NAND2X1 NAND2X1_143 ( .A(IR_REG_10_), .B(_abc_40344_n559_1), .Y(_abc_40344_n1324) );
  NAND2X1 NAND2X1_144 ( .A(_abc_40344_n1325), .B(_abc_40344_n705_1), .Y(_abc_40344_n1326) );
  NAND2X1 NAND2X1_145 ( .A(REG2_REG_10_), .B(_abc_40344_n695), .Y(_abc_40344_n1333) );
  NAND2X1 NAND2X1_146 ( .A(IR_REG_9_), .B(_abc_40344_n1245), .Y(_abc_40344_n1343_1) );
  NAND2X1 NAND2X1_147 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1345), .Y(_abc_40344_n1346) );
  NAND2X1 NAND2X1_148 ( .A(_abc_40344_n1348), .B(_abc_40344_n705_1), .Y(_abc_40344_n1349) );
  NAND2X1 NAND2X1_149 ( .A(_abc_40344_n1369), .B(_abc_40344_n1245), .Y(_abc_40344_n1370) );
  NAND2X1 NAND2X1_15 ( .A(_abc_40344_n604), .B(_abc_40344_n557_1), .Y(_abc_40344_n606) );
  NAND2X1 NAND2X1_150 ( .A(IR_REG_8_), .B(_abc_40344_n559_1), .Y(_abc_40344_n1371_1) );
  NAND2X1 NAND2X1_151 ( .A(_abc_40344_n1373), .B(_abc_40344_n705_1), .Y(_abc_40344_n1374) );
  NAND2X1 NAND2X1_152 ( .A(_abc_40344_n1364), .B(_abc_40344_n1366), .Y(_abc_40344_n1390) );
  NAND2X1 NAND2X1_153 ( .A(_abc_40344_n1188), .B(_abc_40344_n1190), .Y(_abc_40344_n1400) );
  NAND2X1 NAND2X1_154 ( .A(REG0_REG_19_), .B(_abc_40344_n673), .Y(_abc_40344_n1409_1) );
  NAND2X1 NAND2X1_155 ( .A(_abc_40344_n1422), .B(_abc_40344_n1061), .Y(_abc_40344_n1423) );
  NAND2X1 NAND2X1_156 ( .A(REG0_REG_20_), .B(_abc_40344_n673), .Y(_abc_40344_n1425) );
  NAND2X1 NAND2X1_157 ( .A(REG2_REG_20_), .B(_abc_40344_n695), .Y(_abc_40344_n1426) );
  NAND2X1 NAND2X1_158 ( .A(REG1_REG_20_), .B(_abc_40344_n696), .Y(_abc_40344_n1427) );
  NAND2X1 NAND2X1_159 ( .A(REG0_REG_21_), .B(_abc_40344_n673), .Y(_abc_40344_n1437) );
  NAND2X1 NAND2X1_16 ( .A(_abc_40344_n605), .B(_abc_40344_n609), .Y(_abc_40344_n610_1) );
  NAND2X1 NAND2X1_160 ( .A(_abc_40344_n1437), .B(_abc_40344_n1438), .Y(_abc_40344_n1439_1) );
  NAND2X1 NAND2X1_161 ( .A(_abc_40344_n1442), .B(_abc_40344_n1444), .Y(_abc_40344_n1445) );
  NAND2X1 NAND2X1_162 ( .A(_abc_40344_n1430), .B(_abc_40344_n1432), .Y(_abc_40344_n1454) );
  NAND2X1 NAND2X1_163 ( .A(_abc_40344_n1445), .B(_abc_40344_n1456), .Y(_abc_40344_n1457) );
  NAND2X1 NAND2X1_164 ( .A(_abc_40344_n1096), .B(_abc_40344_n1460), .Y(_abc_40344_n1461) );
  NAND2X1 NAND2X1_165 ( .A(_abc_40344_n1043), .B(_abc_40344_n1063), .Y(_abc_40344_n1465) );
  NAND2X1 NAND2X1_166 ( .A(_abc_40344_n1465), .B(_abc_40344_n1464), .Y(_abc_40344_n1466) );
  NAND2X1 NAND2X1_167 ( .A(REG2_REG_24_), .B(_abc_40344_n695), .Y(_abc_40344_n1468) );
  NAND2X1 NAND2X1_168 ( .A(_abc_40344_n1044), .B(_abc_40344_n1479), .Y(_abc_40344_n1480) );
  NAND2X1 NAND2X1_169 ( .A(REG0_REG_25_), .B(_abc_40344_n673), .Y(_abc_40344_n1482) );
  NAND2X1 NAND2X1_17 ( .A(_abc_40344_n613), .B(_abc_40344_n546_1), .Y(_abc_40344_n614) );
  NAND2X1 NAND2X1_170 ( .A(REG2_REG_25_), .B(_abc_40344_n695), .Y(_abc_40344_n1485) );
  NAND2X1 NAND2X1_171 ( .A(_abc_40344_n1041), .B(_abc_40344_n1064), .Y(_abc_40344_n1497) );
  NAND2X1 NAND2X1_172 ( .A(REG0_REG_26_), .B(_abc_40344_n673), .Y(_abc_40344_n1499) );
  NAND2X1 NAND2X1_173 ( .A(REG2_REG_26_), .B(_abc_40344_n695), .Y(_abc_40344_n1502) );
  NAND2X1 NAND2X1_174 ( .A(_abc_40344_n1508_1), .B(_abc_40344_n1510), .Y(_abc_40344_n1511_1) );
  NAND2X1 NAND2X1_175 ( .A(_abc_40344_n1473), .B(_abc_40344_n1475), .Y(_abc_40344_n1515) );
  NAND2X1 NAND2X1_176 ( .A(_abc_40344_n1490), .B(_abc_40344_n1493), .Y(_abc_40344_n1517_1) );
  NAND2X1 NAND2X1_177 ( .A(_abc_40344_n1511_1), .B(_abc_40344_n1520_1), .Y(_abc_40344_n1521) );
  NAND2X1 NAND2X1_178 ( .A(_abc_40344_n1524), .B(_abc_40344_n1525), .Y(_abc_40344_n1526) );
  NAND2X1 NAND2X1_179 ( .A(_abc_40344_n993), .B(_abc_40344_n1535), .Y(_abc_40344_n1536) );
  NAND2X1 NAND2X1_18 ( .A(IR_REG_21_), .B(_abc_40344_n559_1), .Y(_abc_40344_n617_1) );
  NAND2X1 NAND2X1_180 ( .A(REG0_REG_28_), .B(_abc_40344_n673), .Y(_abc_40344_n1543) );
  NAND2X1 NAND2X1_181 ( .A(REG2_REG_28_), .B(_abc_40344_n695), .Y(_abc_40344_n1546) );
  NAND2X1 NAND2X1_182 ( .A(_abc_40344_n1340), .B(_abc_40344_n1393), .Y(_abc_40344_n1559) );
  NAND2X1 NAND2X1_183 ( .A(_abc_40344_n1239), .B(_abc_40344_n1241), .Y(_abc_40344_n1561) );
  NAND2X1 NAND2X1_184 ( .A(_abc_40344_n1561), .B(_abc_40344_n1560), .Y(_abc_40344_n1563) );
  NAND2X1 NAND2X1_185 ( .A(_abc_40344_n993), .B(_abc_40344_n1563), .Y(_abc_40344_n1564) );
  NAND2X1 NAND2X1_186 ( .A(_abc_40344_n1336), .B(_abc_40344_n1338), .Y(_abc_40344_n1587) );
  NAND2X1 NAND2X1_187 ( .A(_abc_40344_n1587), .B(_abc_40344_n1588), .Y(_abc_40344_n1589) );
  NAND2X1 NAND2X1_188 ( .A(_abc_40344_n1597), .B(_abc_40344_n1592), .Y(n1311) );
  NAND2X1 NAND2X1_189 ( .A(_abc_40344_n830), .B(_abc_40344_n895), .Y(_abc_40344_n1601) );
  NAND2X1 NAND2X1_19 ( .A(_abc_40344_n631), .B(_abc_40344_n629), .Y(n1341) );
  NAND2X1 NAND2X1_190 ( .A(_abc_40344_n1005), .B(_abc_40344_n1605), .Y(_abc_40344_n1606) );
  NAND2X1 NAND2X1_191 ( .A(_abc_40344_n1607), .B(_abc_40344_n705_1), .Y(_abc_40344_n1608) );
  NAND2X1 NAND2X1_192 ( .A(_abc_40344_n1416), .B(_abc_40344_n1450), .Y(_abc_40344_n1618) );
  NAND2X1 NAND2X1_193 ( .A(REG2_REG_29_), .B(_abc_40344_n695), .Y(_abc_40344_n1642) );
  NAND2X1 NAND2X1_194 ( .A(_abc_40344_n790), .B(_abc_40344_n898), .Y(_abc_40344_n1656) );
  NAND2X1 NAND2X1_195 ( .A(_abc_40344_n993), .B(_abc_40344_n1660), .Y(_abc_40344_n1661) );
  NAND2X1 NAND2X1_196 ( .A(_abc_40344_n1372), .B(_abc_40344_n705_1), .Y(_abc_40344_n1664) );
  NAND2X1 NAND2X1_197 ( .A(_abc_40344_n1454), .B(_abc_40344_n1686), .Y(_abc_40344_n1687) );
  NAND2X1 NAND2X1_198 ( .A(_abc_40344_n1314), .B(_abc_40344_n1317_1), .Y(_abc_40344_n1701) );
  NAND2X1 NAND2X1_199 ( .A(_abc_40344_n1318), .B(_abc_40344_n1705), .Y(_abc_40344_n1706) );
  NAND2X1 NAND2X1_2 ( .A(_abc_40344_n532), .B(_abc_40344_n533), .Y(_abc_40344_n534) );
  NAND2X1 NAND2X1_20 ( .A(IR_REG_25_), .B(_abc_40344_n559_1), .Y(_abc_40344_n636) );
  NAND2X1 NAND2X1_200 ( .A(_abc_40344_n993), .B(_abc_40344_n1721), .Y(_abc_40344_n1722) );
  NAND2X1 NAND2X1_201 ( .A(_abc_40344_n769), .B(_abc_40344_n768), .Y(_abc_40344_n1742) );
  NAND2X1 NAND2X1_202 ( .A(_abc_40344_n847), .B(_abc_40344_n897), .Y(_abc_40344_n1773) );
  NAND2X1 NAND2X1_203 ( .A(_abc_40344_n790), .B(_abc_40344_n791), .Y(_abc_40344_n1774) );
  NAND2X1 NAND2X1_204 ( .A(_abc_40344_n1390), .B(_abc_40344_n1368), .Y(_abc_40344_n1783) );
  NAND2X1 NAND2X1_205 ( .A(_abc_40344_n1783), .B(_abc_40344_n1782), .Y(_abc_40344_n1785) );
  NAND2X1 NAND2X1_206 ( .A(_abc_40344_n993), .B(_abc_40344_n1785), .Y(_abc_40344_n1786) );
  NAND2X1 NAND2X1_207 ( .A(_abc_40344_n1116), .B(_abc_40344_n1118_1), .Y(_abc_40344_n1831) );
  NAND2X1 NAND2X1_208 ( .A(_abc_40344_n1838), .B(_abc_40344_n1833), .Y(n1221) );
  NAND2X1 NAND2X1_209 ( .A(_abc_40344_n1318), .B(_abc_40344_n1289), .Y(_abc_40344_n1846) );
  NAND2X1 NAND2X1_21 ( .A(_abc_40344_n546_1), .B(_abc_40344_n621), .Y(_abc_40344_n642) );
  NAND2X1 NAND2X1_210 ( .A(_abc_40344_n1846), .B(_abc_40344_n1704), .Y(_abc_40344_n1848) );
  NAND2X1 NAND2X1_211 ( .A(_abc_40344_n993), .B(_abc_40344_n1848), .Y(_abc_40344_n1849) );
  NAND2X1 NAND2X1_212 ( .A(_abc_40344_n844), .B(_abc_40344_n1601), .Y(_abc_40344_n1851) );
  NAND2X1 NAND2X1_213 ( .A(_abc_40344_n1141), .B(_abc_40344_n1143), .Y(_abc_40344_n1860) );
  NAND2X1 NAND2X1_214 ( .A(_abc_40344_n1867), .B(_abc_40344_n1862), .Y(n1206) );
  NAND2X1 NAND2X1_215 ( .A(_abc_40344_n1515), .B(_abc_40344_n1517_1), .Y(_abc_40344_n1882) );
  NAND2X1 NAND2X1_216 ( .A(_abc_40344_n993), .B(_abc_40344_n1884), .Y(_abc_40344_n1885) );
  NAND2X1 NAND2X1_217 ( .A(_abc_40344_n1497), .B(_abc_40344_n1496), .Y(_abc_40344_n1887) );
  NAND2X1 NAND2X1_218 ( .A(_abc_40344_n1239), .B(_abc_40344_n1394), .Y(_abc_40344_n1894) );
  NAND2X1 NAND2X1_219 ( .A(_abc_40344_n1217), .B(_abc_40344_n1216), .Y(_abc_40344_n1895) );
  NAND2X1 NAND2X1_22 ( .A(_abc_40344_n642), .B(_abc_40344_n643), .Y(_abc_40344_n644) );
  NAND2X1 NAND2X1_220 ( .A(_abc_40344_n1902), .B(_abc_40344_n1897), .Y(n1191) );
  NAND2X1 NAND2X1_221 ( .A(_abc_40344_n1347), .B(_abc_40344_n705_1), .Y(_abc_40344_n1905) );
  NAND2X1 NAND2X1_222 ( .A(REG0_REG_31_), .B(_abc_40344_n673), .Y(_abc_40344_n1912) );
  NAND2X1 NAND2X1_223 ( .A(REG0_REG_30_), .B(_abc_40344_n673), .Y(_abc_40344_n1920) );
  NAND2X1 NAND2X1_224 ( .A(_abc_40344_n1926), .B(_abc_40344_n1645), .Y(_abc_40344_n1927) );
  NAND2X1 NAND2X1_225 ( .A(_abc_40344_n1925), .B(_abc_40344_n1927), .Y(_abc_40344_n1928) );
  NAND2X1 NAND2X1_226 ( .A(_abc_40344_n1084), .B(_abc_40344_n1090_1), .Y(_abc_40344_n1945) );
  NAND2X1 NAND2X1_227 ( .A(_abc_40344_n1958), .B(_abc_40344_n1955), .Y(_abc_40344_n1959) );
  NAND2X1 NAND2X1_228 ( .A(_abc_40344_n1967), .B(_abc_40344_n705_1), .Y(_abc_40344_n1968) );
  NAND2X1 NAND2X1_229 ( .A(_abc_40344_n705_1), .B(_abc_40344_n1271), .Y(_abc_40344_n1972) );
  NAND2X1 NAND2X1_23 ( .A(IR_REG_31_), .B(_abc_40344_n644), .Y(_abc_40344_n645) );
  NAND2X1 NAND2X1_230 ( .A(_abc_40344_n1940), .B(_abc_40344_n1965), .Y(_abc_40344_n1982) );
  NAND2X1 NAND2X1_231 ( .A(REG2_REG_6_), .B(_abc_40344_n695), .Y(_abc_40344_n1990) );
  NAND2X1 NAND2X1_232 ( .A(_abc_40344_n1992), .B(_abc_40344_n705_1), .Y(_abc_40344_n1993) );
  NAND2X1 NAND2X1_233 ( .A(_abc_40344_n2008), .B(_abc_40344_n2012), .Y(_abc_40344_n2013) );
  NAND2X1 NAND2X1_234 ( .A(_abc_40344_n685_1), .B(_abc_40344_n1541), .Y(_abc_40344_n2027) );
  NAND2X1 NAND2X1_235 ( .A(_abc_40344_n2056), .B(_abc_40344_n1960), .Y(_abc_40344_n2057) );
  NAND2X1 NAND2X1_236 ( .A(_abc_40344_n1404), .B(_abc_40344_n1414), .Y(_abc_40344_n2064) );
  NAND2X1 NAND2X1_237 ( .A(_abc_40344_n2065), .B(_abc_40344_n1904), .Y(_abc_40344_n2066) );
  NAND2X1 NAND2X1_238 ( .A(_abc_40344_n2068), .B(_abc_40344_n1965), .Y(_abc_40344_n2069) );
  NAND2X1 NAND2X1_239 ( .A(_abc_40344_n2074), .B(_abc_40344_n1904), .Y(_abc_40344_n2075) );
  NAND2X1 NAND2X1_24 ( .A(_abc_40344_n619), .B(_abc_40344_n648), .Y(_abc_40344_n649_1) );
  NAND2X1 NAND2X1_240 ( .A(_abc_40344_n2076), .B(_abc_40344_n1958), .Y(_abc_40344_n2077) );
  NAND2X1 NAND2X1_241 ( .A(_abc_40344_n2078), .B(_abc_40344_n1904), .Y(_abc_40344_n2079) );
  NAND2X1 NAND2X1_242 ( .A(_abc_40344_n2047), .B(_abc_40344_n2080), .Y(_abc_40344_n2081) );
  NAND2X1 NAND2X1_243 ( .A(_abc_40344_n1964), .B(_abc_40344_n1960), .Y(_abc_40344_n2110) );
  NAND2X1 NAND2X1_244 ( .A(_abc_40344_n1495), .B(_abc_40344_n1506), .Y(_abc_40344_n2117) );
  NAND2X1 NAND2X1_245 ( .A(_abc_40344_n2130), .B(_abc_40344_n1984), .Y(_abc_40344_n2131) );
  NAND2X1 NAND2X1_246 ( .A(_abc_40344_n863), .B(_abc_40344_n856), .Y(_abc_40344_n2137) );
  NAND2X1 NAND2X1_247 ( .A(_abc_40344_n2005), .B(_abc_40344_n2140), .Y(_abc_40344_n2141) );
  NAND2X1 NAND2X1_248 ( .A(_abc_40344_n2151), .B(_abc_40344_n1904), .Y(_abc_40344_n2152) );
  NAND2X1 NAND2X1_249 ( .A(IR_REG_22_), .B(_abc_40344_n559_1), .Y(_abc_40344_n2159) );
  NAND2X1 NAND2X1_25 ( .A(_abc_40344_n545_1), .B(_abc_40344_n549_1), .Y(_abc_40344_n654) );
  NAND2X1 NAND2X1_250 ( .A(_abc_40344_n559_1), .B(_abc_40344_n613), .Y(_abc_40344_n2160) );
  NAND2X1 NAND2X1_251 ( .A(_abc_40344_n812), .B(_abc_40344_n802), .Y(_abc_40344_n2163) );
  NAND2X1 NAND2X1_252 ( .A(_abc_40344_n2164), .B(_abc_40344_n2166), .Y(_abc_40344_n2167) );
  NAND2X1 NAND2X1_253 ( .A(_abc_40344_n2168), .B(_abc_40344_n802), .Y(_abc_40344_n2169) );
  NAND2X1 NAND2X1_254 ( .A(_abc_40344_n2173), .B(_abc_40344_n787_1), .Y(_abc_40344_n2174) );
  NAND2X1 NAND2X1_255 ( .A(_abc_40344_n773), .B(_abc_40344_n705_1), .Y(_abc_40344_n2175) );
  NAND2X1 NAND2X1_256 ( .A(DATAI_4_), .B(_abc_40344_n802), .Y(_abc_40344_n2176) );
  NAND2X1 NAND2X1_257 ( .A(DATAI_5_), .B(_abc_40344_n802), .Y(_abc_40344_n2187) );
  NAND2X1 NAND2X1_258 ( .A(_abc_40344_n2205), .B(_abc_40344_n2200), .Y(_abc_40344_n2206) );
  NAND2X1 NAND2X1_259 ( .A(_abc_40344_n2213), .B(_abc_40344_n2212), .Y(_abc_40344_n2214) );
  NAND2X1 NAND2X1_26 ( .A(_abc_40344_n664), .B(_abc_40344_n661), .Y(_abc_40344_n665) );
  NAND2X1 NAND2X1_260 ( .A(_abc_40344_n877_1), .B(_abc_40344_n802), .Y(_abc_40344_n2222) );
  NAND2X1 NAND2X1_261 ( .A(_abc_40344_n2236), .B(_abc_40344_n2235), .Y(_abc_40344_n2237) );
  NAND2X1 NAND2X1_262 ( .A(_abc_40344_n2238), .B(_abc_40344_n2239), .Y(_abc_40344_n2240) );
  NAND2X1 NAND2X1_263 ( .A(_abc_40344_n2243), .B(_abc_40344_n2244), .Y(_abc_40344_n2245) );
  NAND2X1 NAND2X1_264 ( .A(_abc_40344_n728), .B(_abc_40344_n802), .Y(_abc_40344_n2255) );
  NAND2X1 NAND2X1_265 ( .A(_abc_40344_n2173), .B(_abc_40344_n763), .Y(_abc_40344_n2257) );
  NAND2X1 NAND2X1_266 ( .A(_abc_40344_n2195), .B(_abc_40344_n2194), .Y(_abc_40344_n2260) );
  NAND2X1 NAND2X1_267 ( .A(_abc_40344_n2184), .B(_abc_40344_n2183), .Y(_abc_40344_n2261) );
  NAND2X1 NAND2X1_268 ( .A(DATAI_10_), .B(_abc_40344_n802), .Y(_abc_40344_n2264) );
  NAND2X1 NAND2X1_269 ( .A(_abc_40344_n1321), .B(_abc_40344_n802), .Y(_abc_40344_n2267) );
  NAND2X1 NAND2X1_27 ( .A(IR_REG_31_), .B(_abc_40344_n665), .Y(_abc_40344_n666_1) );
  NAND2X1 NAND2X1_270 ( .A(_abc_40344_n2331_1), .B(_abc_40344_n2330), .Y(_abc_40344_n2332) );
  NAND2X1 NAND2X1_271 ( .A(_abc_40344_n2326), .B(_abc_40344_n2325), .Y(_abc_40344_n2333) );
  NAND2X1 NAND2X1_272 ( .A(_abc_40344_n2338), .B(_abc_40344_n2337), .Y(_abc_40344_n2341) );
  NAND2X1 NAND2X1_273 ( .A(_abc_40344_n586), .B(_abc_40344_n1441), .Y(_abc_40344_n2350) );
  NAND2X1 NAND2X1_274 ( .A(_abc_40344_n2359), .B(_abc_40344_n2358), .Y(_abc_40344_n2360) );
  NAND2X1 NAND2X1_275 ( .A(_abc_40344_n2367), .B(_abc_40344_n2366), .Y(_abc_40344_n2373) );
  NAND2X1 NAND2X1_276 ( .A(_abc_40344_n2418), .B(_abc_40344_n2419), .Y(_abc_40344_n2420) );
  NAND2X1 NAND2X1_277 ( .A(_abc_40344_n2216), .B(_abc_40344_n2215), .Y(_abc_40344_n2431) );
  NAND2X1 NAND2X1_278 ( .A(_abc_40344_n2217), .B(_abc_40344_n2218), .Y(_abc_40344_n2432) );
  NAND2X1 NAND2X1_279 ( .A(_abc_40344_n2422), .B(_abc_40344_n2421), .Y(_abc_40344_n2443) );
  NAND2X1 NAND2X1_28 ( .A(IR_REG_30_), .B(_abc_40344_n559_1), .Y(_abc_40344_n675) );
  NAND2X1 NAND2X1_280 ( .A(_abc_40344_n2001), .B(_abc_40344_n2117), .Y(_abc_40344_n2469) );
  NAND2X1 NAND2X1_281 ( .A(_abc_40344_n2479), .B(_abc_40344_n2478_1), .Y(_abc_40344_n2480) );
  NAND2X1 NAND2X1_282 ( .A(_abc_40344_n1974), .B(_abc_40344_n2122), .Y(_abc_40344_n2484_1) );
  NAND2X1 NAND2X1_283 ( .A(_abc_40344_n1985), .B(_abc_40344_n2486), .Y(_abc_40344_n2487) );
  NAND2X1 NAND2X1_284 ( .A(_abc_40344_n2137), .B(_abc_40344_n2142), .Y(_abc_40344_n2488) );
  NAND2X1 NAND2X1_285 ( .A(_abc_40344_n809), .B(_abc_40344_n813), .Y(_abc_40344_n2490) );
  NAND2X1 NAND2X1_286 ( .A(_abc_40344_n2490), .B(_abc_40344_n2018), .Y(_abc_40344_n2491) );
  NAND2X1 NAND2X1_287 ( .A(_abc_40344_n2498), .B(_abc_40344_n2089), .Y(_abc_40344_n2499) );
  NAND2X1 NAND2X1_288 ( .A(_abc_40344_n1947), .B(_abc_40344_n2502_1), .Y(_abc_40344_n2503) );
  NAND2X1 NAND2X1_289 ( .A(_abc_40344_n1076), .B(_abc_40344_n1074), .Y(_abc_40344_n2511) );
  NAND2X1 NAND2X1_29 ( .A(_abc_40344_n535), .B(_abc_40344_n543), .Y(_abc_40344_n677) );
  NAND2X1 NAND2X1_290 ( .A(_abc_40344_n2010), .B(_abc_40344_n2511), .Y(_abc_40344_n2512) );
  NAND2X1 NAND2X1_291 ( .A(_abc_40344_n1100), .B(_abc_40344_n1110), .Y(_abc_40344_n2515) );
  NAND2X1 NAND2X1_292 ( .A(_abc_40344_n1943), .B(_abc_40344_n2515), .Y(_abc_40344_n2516) );
  NAND2X1 NAND2X1_293 ( .A(_abc_40344_n1463), .B(_abc_40344_n1471), .Y(_abc_40344_n2519) );
  NAND2X1 NAND2X1_294 ( .A(_abc_40344_n2519), .B(_abc_40344_n2518), .Y(_abc_40344_n2520) );
  NAND2X1 NAND2X1_295 ( .A(_abc_40344_n1083), .B(_abc_40344_n1090_1), .Y(_abc_40344_n2522) );
  NAND2X1 NAND2X1_296 ( .A(_abc_40344_n1084), .B(_abc_40344_n1091), .Y(_abc_40344_n2523_1) );
  NAND2X1 NAND2X1_297 ( .A(_abc_40344_n2522), .B(_abc_40344_n2523_1), .Y(_abc_40344_n2524) );
  NAND2X1 NAND2X1_298 ( .A(_abc_40344_n2223), .B(_abc_40344_n2528), .Y(_abc_40344_n2529_1) );
  NAND2X1 NAND2X1_299 ( .A(_abc_40344_n2530), .B(_abc_40344_n2531), .Y(_abc_40344_n2532) );
  NAND2X1 NAND2X1_3 ( .A(_abc_40344_n540), .B(_abc_40344_n541_1), .Y(_abc_40344_n542_1) );
  NAND2X1 NAND2X1_30 ( .A(_abc_40344_n600_1), .B(_abc_40344_n549_1), .Y(_abc_40344_n678) );
  NAND2X1 NAND2X1_300 ( .A(_abc_40344_n1962), .B(_abc_40344_n2537), .Y(_abc_40344_n2538) );
  NAND2X1 NAND2X1_301 ( .A(_abc_40344_n1938), .B(_abc_40344_n2544), .Y(_abc_40344_n2545) );
  NAND2X1 NAND2X1_302 ( .A(_abc_40344_n2134), .B(_abc_40344_n2024), .Y(_abc_40344_n2546) );
  NAND2X1 NAND2X1_303 ( .A(_abc_40344_n1649), .B(_abc_40344_n1550), .Y(_abc_40344_n2555) );
  NAND2X1 NAND2X1_304 ( .A(_abc_40344_n1904), .B(_abc_40344_n2555), .Y(_abc_40344_n2556) );
  NAND2X1 NAND2X1_305 ( .A(_abc_40344_n2413), .B(_abc_40344_n2412), .Y(_abc_40344_n2564) );
  NAND2X1 NAND2X1_306 ( .A(_abc_40344_n2030), .B(_abc_40344_n2591), .Y(_abc_40344_n2592) );
  NAND2X1 NAND2X1_307 ( .A(_abc_40344_n1954), .B(_abc_40344_n2030), .Y(_abc_40344_n2596) );
  NAND2X1 NAND2X1_308 ( .A(_abc_40344_n2602), .B(_abc_40344_n2593_1), .Y(_abc_40344_n2609) );
  NAND2X1 NAND2X1_309 ( .A(_abc_40344_n2628), .B(_abc_40344_n2626), .Y(_abc_40344_n2629) );
  NAND2X1 NAND2X1_31 ( .A(_abc_40344_n679), .B(_abc_40344_n680), .Y(_abc_40344_n681) );
  NAND2X1 NAND2X1_310 ( .A(_abc_40344_n1489), .B(_abc_40344_n2637), .Y(_abc_40344_n2638) );
  NAND2X1 NAND2X1_311 ( .A(_abc_40344_n1491), .B(_abc_40344_n2637), .Y(_abc_40344_n2639) );
  NAND2X1 NAND2X1_312 ( .A(_abc_40344_n648), .B(_abc_40344_n717), .Y(_abc_40344_n2641) );
  NAND2X1 NAND2X1_313 ( .A(_abc_40344_n646), .B(_abc_40344_n626), .Y(_abc_40344_n2644_1) );
  NAND2X1 NAND2X1_314 ( .A(IR_REG_0_), .B(REG2_REG_0_), .Y(_abc_40344_n2680) );
  NAND2X1 NAND2X1_315 ( .A(_abc_40344_n2685), .B(_abc_40344_n2676), .Y(n1054) );
  NAND2X1 NAND2X1_316 ( .A(REG2_REG_1_), .B(_abc_40344_n2688), .Y(_abc_40344_n2689) );
  NAND2X1 NAND2X1_317 ( .A(_abc_40344_n2680), .B(_abc_40344_n853), .Y(_abc_40344_n2690) );
  NAND2X1 NAND2X1_318 ( .A(_abc_40344_n2689), .B(_abc_40344_n2692_1), .Y(_abc_40344_n2693) );
  NAND2X1 NAND2X1_319 ( .A(REG1_REG_1_), .B(_abc_40344_n2694), .Y(_abc_40344_n2695) );
  NAND2X1 NAND2X1_32 ( .A(IR_REG_29_), .B(_abc_40344_n559_1), .Y(_abc_40344_n684) );
  NAND2X1 NAND2X1_320 ( .A(_abc_40344_n2715), .B(_abc_40344_n2717), .Y(_abc_40344_n2718) );
  NAND2X1 NAND2X1_321 ( .A(_abc_40344_n2722_1), .B(_abc_40344_n610_1), .Y(_abc_40344_n2723) );
  NAND2X1 NAND2X1_322 ( .A(REG2_REG_3_), .B(_abc_40344_n797), .Y(_abc_40344_n2730_1) );
  NAND2X1 NAND2X1_323 ( .A(_abc_40344_n2730_1), .B(_abc_40344_n2729), .Y(_abc_40344_n2731) );
  NAND2X1 NAND2X1_324 ( .A(REG1_REG_3_), .B(_abc_40344_n2735), .Y(_abc_40344_n2736) );
  NAND2X1 NAND2X1_325 ( .A(_abc_40344_n2736), .B(_abc_40344_n2738), .Y(_abc_40344_n2739) );
  NAND2X1 NAND2X1_326 ( .A(REG2_REG_4_), .B(_abc_40344_n773), .Y(_abc_40344_n2752) );
  NAND2X1 NAND2X1_327 ( .A(_abc_40344_n2203), .B(_abc_40344_n774), .Y(_abc_40344_n2753) );
  NAND2X1 NAND2X1_328 ( .A(_abc_40344_n2752), .B(_abc_40344_n2753), .Y(_abc_40344_n2754) );
  NAND2X1 NAND2X1_329 ( .A(_abc_40344_n2760_1), .B(_abc_40344_n2772), .Y(n1034) );
  NAND2X1 NAND2X1_33 ( .A(REG3_REG_5_), .B(_abc_40344_n689), .Y(_abc_40344_n690) );
  NAND2X1 NAND2X1_330 ( .A(REG1_REG_5_), .B(_abc_40344_n2762), .Y(_abc_40344_n2776) );
  NAND2X1 NAND2X1_331 ( .A(_abc_40344_n2776), .B(_abc_40344_n2777), .Y(_abc_40344_n2778) );
  NAND2X1 NAND2X1_332 ( .A(REG1_REG_6_), .B(_abc_40344_n712), .Y(_abc_40344_n2779) );
  NAND2X1 NAND2X1_333 ( .A(_abc_40344_n1989), .B(_abc_40344_n1992), .Y(_abc_40344_n2780) );
  NAND2X1 NAND2X1_334 ( .A(_abc_40344_n2779), .B(_abc_40344_n2780), .Y(_abc_40344_n2781) );
  NAND2X1 NAND2X1_335 ( .A(REG2_REG_6_), .B(_abc_40344_n712), .Y(_abc_40344_n2785) );
  NAND2X1 NAND2X1_336 ( .A(_abc_40344_n2785), .B(_abc_40344_n2784), .Y(_abc_40344_n2786) );
  NAND2X1 NAND2X1_337 ( .A(REG1_REG_7_), .B(_abc_40344_n906_1), .Y(_abc_40344_n2798) );
  NAND2X1 NAND2X1_338 ( .A(_abc_40344_n924), .B(_abc_40344_n917), .Y(_abc_40344_n2799) );
  NAND2X1 NAND2X1_339 ( .A(_abc_40344_n2798), .B(_abc_40344_n2799), .Y(_abc_40344_n2800) );
  NAND2X1 NAND2X1_34 ( .A(_abc_40344_n694_1), .B(_abc_40344_n697), .Y(_abc_40344_n698) );
  NAND2X1 NAND2X1_340 ( .A(_abc_40344_n920), .B(_abc_40344_n917), .Y(_abc_40344_n2805) );
  NAND2X1 NAND2X1_341 ( .A(REG1_REG_9_), .B(_abc_40344_n1348), .Y(_abc_40344_n2835) );
  NAND2X1 NAND2X1_342 ( .A(_abc_40344_n1351), .B(_abc_40344_n1347), .Y(_abc_40344_n2836) );
  NAND2X1 NAND2X1_343 ( .A(_abc_40344_n2836), .B(_abc_40344_n2835), .Y(_abc_40344_n2837) );
  NAND2X1 NAND2X1_344 ( .A(REG1_REG_10_), .B(_abc_40344_n2845), .Y(_abc_40344_n2848) );
  NAND2X1 NAND2X1_345 ( .A(_abc_40344_n1967), .B(_abc_40344_n2848), .Y(_abc_40344_n2851) );
  NAND2X1 NAND2X1_346 ( .A(REG2_REG_10_), .B(_abc_40344_n1325), .Y(_abc_40344_n2853) );
  NAND2X1 NAND2X1_347 ( .A(_abc_40344_n2853), .B(_abc_40344_n2855), .Y(_abc_40344_n2856) );
  NAND2X1 NAND2X1_348 ( .A(REG1_REG_11_), .B(_abc_40344_n2863), .Y(_abc_40344_n2864) );
  NAND2X1 NAND2X1_349 ( .A(_abc_40344_n2864), .B(_abc_40344_n2866), .Y(_abc_40344_n2867) );
  NAND2X1 NAND2X1_35 ( .A(_abc_40344_n618), .B(_abc_40344_n640), .Y(_abc_40344_n699) );
  NAND2X1 NAND2X1_350 ( .A(_abc_40344_n1296), .B(_abc_40344_n1293_1), .Y(_abc_40344_n2882) );
  NAND2X1 NAND2X1_351 ( .A(REG1_REG_12_), .B(_abc_40344_n2883), .Y(_abc_40344_n2884) );
  NAND2X1 NAND2X1_352 ( .A(_abc_40344_n2882), .B(_abc_40344_n2884), .Y(_abc_40344_n2885) );
  NAND2X1 NAND2X1_353 ( .A(REG2_REG_12_), .B(_abc_40344_n2883), .Y(_abc_40344_n2892) );
  NAND2X1 NAND2X1_354 ( .A(_abc_40344_n2892), .B(_abc_40344_n2891), .Y(_abc_40344_n2893) );
  NAND2X1 NAND2X1_355 ( .A(_abc_40344_n2897), .B(_abc_40344_n2684), .Y(_abc_40344_n2898) );
  NAND2X1 NAND2X1_356 ( .A(_abc_40344_n2897), .B(_abc_40344_n2677), .Y(_abc_40344_n2900) );
  NAND2X1 NAND2X1_357 ( .A(REG1_REG_13_), .B(_abc_40344_n2905), .Y(_abc_40344_n2906) );
  NAND2X1 NAND2X1_358 ( .A(_abc_40344_n2907), .B(_abc_40344_n2906), .Y(_abc_40344_n2908) );
  NAND2X1 NAND2X1_359 ( .A(_abc_40344_n2918), .B(_abc_40344_n2684), .Y(_abc_40344_n2919) );
  NAND2X1 NAND2X1_36 ( .A(_abc_40344_n529), .B(_abc_40344_n572), .Y(_abc_40344_n706) );
  NAND2X1 NAND2X1_360 ( .A(ADDR_REG_13_), .B(_abc_40344_n2675), .Y(_abc_40344_n2920) );
  NAND2X1 NAND2X1_361 ( .A(_abc_40344_n2911), .B(_abc_40344_n2907), .Y(_abc_40344_n2925) );
  NAND2X1 NAND2X1_362 ( .A(_abc_40344_n1232), .B(_abc_40344_n2926), .Y(_abc_40344_n2927) );
  NAND2X1 NAND2X1_363 ( .A(_abc_40344_n2906), .B(_abc_40344_n2925), .Y(_abc_40344_n2928) );
  NAND2X1 NAND2X1_364 ( .A(REG1_REG_14_), .B(_abc_40344_n2928), .Y(_abc_40344_n2929) );
  NAND2X1 NAND2X1_365 ( .A(_abc_40344_n2937), .B(_abc_40344_n2935), .Y(_abc_40344_n2938) );
  NAND2X1 NAND2X1_366 ( .A(_abc_40344_n2933), .B(_abc_40344_n2947), .Y(n998) );
  NAND2X1 NAND2X1_367 ( .A(_abc_40344_n2960), .B(_abc_40344_n2962), .Y(_abc_40344_n2963) );
  NAND2X1 NAND2X1_368 ( .A(_abc_40344_n2971), .B(_abc_40344_n2973), .Y(_abc_40344_n2974) );
  NAND2X1 NAND2X1_369 ( .A(REG2_REG_16_), .B(_abc_40344_n1149), .Y(_abc_40344_n2978) );
  NAND2X1 NAND2X1_37 ( .A(IR_REG_6_), .B(_abc_40344_n559_1), .Y(_abc_40344_n711) );
  NAND2X1 NAND2X1_370 ( .A(_abc_40344_n2978), .B(_abc_40344_n2980), .Y(_abc_40344_n2981) );
  NAND2X1 NAND2X1_371 ( .A(REG1_REG_17_), .B(_abc_40344_n2991), .Y(_abc_40344_n2992) );
  NAND2X1 NAND2X1_372 ( .A(_abc_40344_n1183), .B(_abc_40344_n1176), .Y(_abc_40344_n2993) );
  NAND2X1 NAND2X1_373 ( .A(_abc_40344_n2993), .B(_abc_40344_n2992), .Y(_abc_40344_n2994) );
  NAND2X1 NAND2X1_374 ( .A(_abc_40344_n1196), .B(_abc_40344_n2975), .Y(_abc_40344_n2996) );
  NAND2X1 NAND2X1_375 ( .A(REG2_REG_17_), .B(_abc_40344_n2991), .Y(_abc_40344_n3001) );
  NAND2X1 NAND2X1_376 ( .A(_abc_40344_n1182), .B(_abc_40344_n1176), .Y(_abc_40344_n3002) );
  NAND2X1 NAND2X1_377 ( .A(_abc_40344_n3002), .B(_abc_40344_n3001), .Y(_abc_40344_n3003) );
  NAND2X1 NAND2X1_378 ( .A(_abc_40344_n2818), .B(_abc_40344_n3031), .Y(_abc_40344_n3032) );
  NAND2X1 NAND2X1_379 ( .A(REG2_REG_19_), .B(_abc_40344_n646), .Y(_abc_40344_n3041_1) );
  NAND2X1 NAND2X1_38 ( .A(_abc_40344_n633_1), .B(_abc_40344_n637), .Y(_abc_40344_n716) );
  NAND2X1 NAND2X1_380 ( .A(_abc_40344_n1411), .B(_abc_40344_n648), .Y(_abc_40344_n3044) );
  NAND2X1 NAND2X1_381 ( .A(REG1_REG_19_), .B(_abc_40344_n646), .Y(_abc_40344_n3054) );
  NAND2X1 NAND2X1_382 ( .A(_abc_40344_n1412), .B(_abc_40344_n648), .Y(_abc_40344_n3055) );
  NAND2X1 NAND2X1_383 ( .A(_abc_40344_n3054), .B(_abc_40344_n3055), .Y(_abc_40344_n3057) );
  NAND2X1 NAND2X1_384 ( .A(_abc_40344_n869), .B(_abc_40344_n1797), .Y(_abc_40344_n3070) );
  NAND2X1 NAND2X1_385 ( .A(_abc_40344_n1609), .B(_abc_40344_n3071), .Y(_abc_40344_n3072) );
  NAND2X1 NAND2X1_386 ( .A(_abc_40344_n750), .B(_abc_40344_n3073), .Y(_abc_40344_n3074) );
  NAND2X1 NAND2X1_387 ( .A(_abc_40344_n919), .B(_abc_40344_n3075), .Y(_abc_40344_n3076) );
  NAND2X1 NAND2X1_388 ( .A(_abc_40344_n1906), .B(_abc_40344_n3077), .Y(_abc_40344_n3078) );
  NAND2X1 NAND2X1_389 ( .A(_abc_40344_n1152_1), .B(_abc_40344_n1200), .Y(_abc_40344_n3083) );
  NAND2X1 NAND2X1_39 ( .A(_abc_40344_n720), .B(_abc_40344_n723), .Y(_abc_40344_n724) );
  NAND2X1 NAND2X1_390 ( .A(_abc_40344_n3096), .B(_abc_40344_n3095), .Y(_abc_40344_n3097) );
  NAND2X1 NAND2X1_391 ( .A(_abc_40344_n1922), .B(_abc_40344_n3098), .Y(_abc_40344_n3099) );
  NAND2X1 NAND2X1_392 ( .A(_abc_40344_n1916), .B(_abc_40344_n3099), .Y(_abc_40344_n3100) );
  NAND2X1 NAND2X1_393 ( .A(_abc_40344_n2401), .B(_abc_40344_n3098), .Y(_abc_40344_n3115) );
  NAND2X1 NAND2X1_394 ( .A(_abc_40344_n787_1), .B(_abc_40344_n776), .Y(_abc_40344_n3139) );
  NAND2X1 NAND2X1_395 ( .A(_abc_40344_n841), .B(_abc_40344_n2022), .Y(_abc_40344_n3141) );
  NAND2X1 NAND2X1_396 ( .A(_abc_40344_n763), .B(_abc_40344_n750), .Y(_abc_40344_n3148) );
  NAND2X1 NAND2X1_397 ( .A(_abc_40344_n3135), .B(_abc_40344_n3158), .Y(_abc_40344_n3159) );
  NAND2X1 NAND2X1_398 ( .A(_abc_40344_n1433), .B(_abc_40344_n1440), .Y(_abc_40344_n3177) );
  NAND2X1 NAND2X1_399 ( .A(_abc_40344_n3193), .B(_abc_40344_n3188), .Y(_abc_40344_n3194) );
  NAND2X1 NAND2X1_4 ( .A(_abc_40344_n545_1), .B(_abc_40344_n546_1), .Y(_abc_40344_n547) );
  NAND2X1 NAND2X1_40 ( .A(_abc_40344_n729_1), .B(_abc_40344_n709), .Y(_abc_40344_n730) );
  NAND2X1 NAND2X1_400 ( .A(_abc_40344_n1494), .B(_abc_40344_n1506), .Y(_abc_40344_n3199) );
  NAND2X1 NAND2X1_401 ( .A(_abc_40344_n3120), .B(_abc_40344_n3212), .Y(_abc_40344_n3213) );
  NAND2X1 NAND2X1_402 ( .A(_abc_40344_n3213), .B(_abc_40344_n3214), .Y(_abc_40344_n3215) );
  NAND2X1 NAND2X1_403 ( .A(_abc_40344_n3220), .B(_abc_40344_n1073), .Y(_abc_40344_n3221_1) );
  NAND2X1 NAND2X1_404 ( .A(_abc_40344_n3236), .B(_abc_40344_n3240), .Y(_abc_40344_n3241) );
  NAND2X1 NAND2X1_405 ( .A(_abc_40344_n3250), .B(_abc_40344_n3247), .Y(_abc_40344_n3251) );
  NAND2X1 NAND2X1_406 ( .A(_abc_40344_n3290), .B(_abc_40344_n3292), .Y(_abc_40344_n3293) );
  NAND2X1 NAND2X1_407 ( .A(_abc_40344_n3323), .B(_abc_40344_n3321), .Y(_abc_40344_n3324) );
  NAND2X1 NAND2X1_408 ( .A(_abc_40344_n3066), .B(_abc_40344_n3339), .Y(_abc_40344_n3340) );
  NAND2X1 NAND2X1_409 ( .A(_abc_40344_n3349), .B(_abc_40344_n3340), .Y(n938) );
  NAND2X1 NAND2X1_41 ( .A(IR_REG_5_), .B(_abc_40344_n559_1), .Y(_abc_40344_n731) );
  NAND2X1 NAND2X1_410 ( .A(_abc_40344_n3356), .B(_abc_40344_n3355), .Y(_abc_40344_n3357) );
  NAND2X1 NAND2X1_411 ( .A(_abc_40344_n3360), .B(_abc_40344_n3357), .Y(_abc_40344_n3361) );
  NAND2X1 NAND2X1_412 ( .A(_abc_40344_n3352), .B(_abc_40344_n3368), .Y(_abc_40344_n3369) );
  NAND2X1 NAND2X1_413 ( .A(_abc_40344_n3066), .B(_abc_40344_n3369), .Y(_abc_40344_n3370) );
  NAND2X1 NAND2X1_414 ( .A(_abc_40344_n3218), .B(_abc_40344_n3351), .Y(_abc_40344_n3371) );
  NAND2X1 NAND2X1_415 ( .A(_abc_40344_n3089), .B(_abc_40344_n3086), .Y(_abc_40344_n3386) );
  NAND2X1 NAND2X1_416 ( .A(_abc_40344_n3068), .B(_abc_40344_n3396), .Y(_abc_40344_n3397) );
  NAND2X1 NAND2X1_417 ( .A(_abc_40344_n3411_1), .B(_abc_40344_n3412), .Y(_abc_40344_n3413) );
  NAND2X1 NAND2X1_418 ( .A(_abc_40344_n3397), .B(_abc_40344_n3421), .Y(n923) );
  NAND2X1 NAND2X1_419 ( .A(_abc_40344_n3432), .B(_abc_40344_n3431_1), .Y(_abc_40344_n3433) );
  NAND2X1 NAND2X1_42 ( .A(_abc_40344_n732_1), .B(_abc_40344_n705_1), .Y(_abc_40344_n733) );
  NAND2X1 NAND2X1_420 ( .A(_abc_40344_n3223), .B(_abc_40344_n3434), .Y(_abc_40344_n3435) );
  NAND2X1 NAND2X1_421 ( .A(_abc_40344_n3437), .B(_abc_40344_n3066), .Y(_abc_40344_n3438) );
  NAND2X1 NAND2X1_422 ( .A(_abc_40344_n3452), .B(_abc_40344_n3457_1), .Y(n913) );
  NAND2X1 NAND2X1_423 ( .A(_abc_40344_n3303), .B(_abc_40344_n3324), .Y(_abc_40344_n3461) );
  NAND2X1 NAND2X1_424 ( .A(_abc_40344_n3068), .B(_abc_40344_n3468), .Y(_abc_40344_n3469) );
  NAND2X1 NAND2X1_425 ( .A(_abc_40344_n1131), .B(_abc_40344_n3067), .Y(_abc_40344_n3471) );
  NAND2X1 NAND2X1_426 ( .A(_abc_40344_n3068), .B(_abc_40344_n3490), .Y(_abc_40344_n3491) );
  NAND2X1 NAND2X1_427 ( .A(_abc_40344_n3066), .B(_abc_40344_n3505), .Y(_abc_40344_n3506_1) );
  NAND2X1 NAND2X1_428 ( .A(_abc_40344_n3218), .B(_abc_40344_n3500), .Y(_abc_40344_n3507) );
  NAND2X1 NAND2X1_429 ( .A(_abc_40344_n3066), .B(_abc_40344_n3523), .Y(_abc_40344_n3524) );
  NAND2X1 NAND2X1_43 ( .A(_abc_40344_n737), .B(_abc_40344_n690), .Y(_abc_40344_n738_1) );
  NAND2X1 NAND2X1_430 ( .A(_abc_40344_n1973), .B(_abc_40344_n3079), .Y(_abc_40344_n3526) );
  NAND2X1 NAND2X1_431 ( .A(_abc_40344_n1264), .B(_abc_40344_n3527), .Y(_abc_40344_n3528) );
  NAND2X1 NAND2X1_432 ( .A(_abc_40344_n3524), .B(_abc_40344_n3537), .Y(n893) );
  NAND2X1 NAND2X1_433 ( .A(_abc_40344_n3066), .B(_abc_40344_n3543), .Y(_abc_40344_n3544) );
  NAND2X1 NAND2X1_434 ( .A(_abc_40344_n3544), .B(_abc_40344_n3555_1), .Y(n888) );
  NAND2X1 NAND2X1_435 ( .A(_abc_40344_n3557), .B(_abc_40344_n3528), .Y(_abc_40344_n3558) );
  NAND2X1 NAND2X1_436 ( .A(_abc_40344_n3218), .B(_abc_40344_n3564), .Y(_abc_40344_n3567) );
  NAND2X1 NAND2X1_437 ( .A(_abc_40344_n3575), .B(_abc_40344_n3545), .Y(_abc_40344_n3576) );
  NAND2X1 NAND2X1_438 ( .A(_abc_40344_n3227), .B(_abc_40344_n3578), .Y(_abc_40344_n3579) );
  NAND2X1 NAND2X1_439 ( .A(_abc_40344_n995), .B(_abc_40344_n1308), .Y(_abc_40344_n3585) );
  NAND2X1 NAND2X1_44 ( .A(_abc_40344_n739), .B(_abc_40344_n685_1), .Y(_abc_40344_n740) );
  NAND2X1 NAND2X1_440 ( .A(_abc_40344_n3068), .B(_abc_40344_n3625), .Y(_abc_40344_n3626) );
  NAND2X1 NAND2X1_441 ( .A(_abc_40344_n3627), .B(_abc_40344_n3066), .Y(_abc_40344_n3628) );
  NAND2X1 NAND2X1_442 ( .A(_abc_40344_n3066), .B(_abc_40344_n3657), .Y(_abc_40344_n3658) );
  NAND2X1 NAND2X1_443 ( .A(_abc_40344_n3668), .B(_abc_40344_n3658), .Y(n858) );
  NAND2X1 NAND2X1_444 ( .A(_abc_40344_n714), .B(_abc_40344_n3074), .Y(_abc_40344_n3686) );
  NAND2X1 NAND2X1_445 ( .A(_abc_40344_n3686), .B(_abc_40344_n3663), .Y(_abc_40344_n3687) );
  NAND2X1 NAND2X1_446 ( .A(_abc_40344_n3713), .B(_abc_40344_n3712), .Y(_abc_40344_n3714) );
  NAND2X1 NAND2X1_447 ( .A(_abc_40344_n3066), .B(_abc_40344_n3714), .Y(_abc_40344_n3715) );
  NAND2X1 NAND2X1_448 ( .A(_abc_40344_n3218), .B(_abc_40344_n3707), .Y(_abc_40344_n3716) );
  NAND2X1 NAND2X1_449 ( .A(_abc_40344_n3739), .B(_abc_40344_n3751), .Y(_abc_40344_n3752) );
  NAND2X1 NAND2X1_45 ( .A(REG1_REG_5_), .B(_abc_40344_n696), .Y(_abc_40344_n741) );
  NAND2X1 NAND2X1_450 ( .A(_abc_40344_n3066), .B(_abc_40344_n3752), .Y(_abc_40344_n3753) );
  NAND2X1 NAND2X1_451 ( .A(_abc_40344_n3759), .B(_abc_40344_n3218), .Y(_abc_40344_n3766_1) );
  NAND2X1 NAND2X1_452 ( .A(_abc_40344_n3791_1), .B(_abc_40344_n3792_1), .Y(n818) );
  NAND2X1 NAND2X1_453 ( .A(D_REG_31_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3796_1) );
  NAND2X1 NAND2X1_454 ( .A(D_REG_30_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3798_1) );
  NAND2X1 NAND2X1_455 ( .A(D_REG_29_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3800) );
  NAND2X1 NAND2X1_456 ( .A(D_REG_28_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3802) );
  NAND2X1 NAND2X1_457 ( .A(D_REG_27_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3804) );
  NAND2X1 NAND2X1_458 ( .A(D_REG_26_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3806) );
  NAND2X1 NAND2X1_459 ( .A(D_REG_25_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3808) );
  NAND2X1 NAND2X1_46 ( .A(_abc_40344_n748), .B(_abc_40344_n705_1), .Y(_abc_40344_n749_1) );
  NAND2X1 NAND2X1_460 ( .A(D_REG_24_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3810_1) );
  NAND2X1 NAND2X1_461 ( .A(D_REG_23_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3812) );
  NAND2X1 NAND2X1_462 ( .A(D_REG_22_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3814) );
  NAND2X1 NAND2X1_463 ( .A(D_REG_21_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3816) );
  NAND2X1 NAND2X1_464 ( .A(D_REG_20_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3818) );
  NAND2X1 NAND2X1_465 ( .A(D_REG_19_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3820) );
  NAND2X1 NAND2X1_466 ( .A(D_REG_18_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3822) );
  NAND2X1 NAND2X1_467 ( .A(D_REG_17_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3824_1) );
  NAND2X1 NAND2X1_468 ( .A(D_REG_16_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3826) );
  NAND2X1 NAND2X1_469 ( .A(D_REG_15_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3828) );
  NAND2X1 NAND2X1_47 ( .A(_abc_40344_n684), .B(_abc_40344_n683_1), .Y(_abc_40344_n760) );
  NAND2X1 NAND2X1_470 ( .A(D_REG_14_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3830_1) );
  NAND2X1 NAND2X1_471 ( .A(D_REG_13_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3832) );
  NAND2X1 NAND2X1_472 ( .A(D_REG_12_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3834) );
  NAND2X1 NAND2X1_473 ( .A(D_REG_11_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3836_1) );
  NAND2X1 NAND2X1_474 ( .A(D_REG_10_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3838) );
  NAND2X1 NAND2X1_475 ( .A(D_REG_9_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3840) );
  NAND2X1 NAND2X1_476 ( .A(D_REG_8_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3842_1) );
  NAND2X1 NAND2X1_477 ( .A(D_REG_7_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3844) );
  NAND2X1 NAND2X1_478 ( .A(D_REG_6_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3846_1) );
  NAND2X1 NAND2X1_479 ( .A(D_REG_5_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3848) );
  NAND2X1 NAND2X1_48 ( .A(_abc_40344_n719), .B(_abc_40344_n764), .Y(_abc_40344_n766) );
  NAND2X1 NAND2X1_480 ( .A(D_REG_4_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3850) );
  NAND2X1 NAND2X1_481 ( .A(D_REG_3_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3852_1) );
  NAND2X1 NAND2X1_482 ( .A(D_REG_2_), .B(_abc_40344_n3795_1), .Y(_abc_40344_n3854) );
  NAND2X1 NAND2X1_483 ( .A(_abc_40344_n3856), .B(_abc_40344_n599), .Y(_abc_40344_n3871_1) );
  NAND2X1 NAND2X1_484 ( .A(_abc_40344_n557_1), .B(_abc_40344_n553_1), .Y(_abc_40344_n3879) );
  NAND2X1 NAND2X1_485 ( .A(_abc_40344_n622), .B(_abc_40344_n623), .Y(_abc_40344_n3897_1) );
  NAND2X1 NAND2X1_486 ( .A(nRESET_G), .B(_abc_40344_n3912), .Y(_abc_40344_n3913) );
  NAND2X1 NAND2X1_487 ( .A(nRESET_G), .B(_abc_40344_n3945), .Y(_abc_40344_n3946) );
  NAND2X1 NAND2X1_488 ( .A(_abc_40344_n3999_1), .B(_abc_40344_n3212), .Y(_abc_40344_n4007) );
  NAND2X1 NAND2X1_489 ( .A(_abc_40344_n3998), .B(_abc_40344_n4009), .Y(_abc_40344_n4010) );
  NAND2X1 NAND2X1_49 ( .A(_abc_40344_n770), .B(_abc_40344_n707_1), .Y(_abc_40344_n771) );
  NAND2X1 NAND2X1_490 ( .A(_abc_40344_n1926), .B(_abc_40344_n3097), .Y(_abc_40344_n4021) );
  NAND2X1 NAND2X1_491 ( .A(_abc_40344_n4022), .B(_abc_40344_n4021), .Y(_abc_40344_n4023) );
  NAND2X1 NAND2X1_492 ( .A(_abc_40344_n4008), .B(_abc_40344_n4006_1), .Y(_abc_40344_n4024) );
  NAND2X1 NAND2X1_493 ( .A(_abc_40344_n4020_1), .B(_abc_40344_n4029), .Y(n963) );
  NAND2X1 NAND2X1_494 ( .A(_abc_40344_n4048), .B(_abc_40344_n3759), .Y(_abc_40344_n4055) );
  NAND2X1 NAND2X1_495 ( .A(_abc_40344_n3624), .B(_abc_40344_n3574), .Y(_abc_40344_n4098) );
  NAND2X1 NAND2X1_496 ( .A(_abc_40344_n4100), .B(_abc_40344_n3622), .Y(_abc_40344_n4101_1) );
  NAND2X1 NAND2X1_497 ( .A(_abc_40344_n4048), .B(_abc_40344_n3541), .Y(_abc_40344_n4123) );
  NAND2X1 NAND2X1_498 ( .A(_abc_40344_n4048), .B(_abc_40344_n3520), .Y(_abc_40344_n4131_1) );
  NAND2X1 NAND2X1_499 ( .A(_abc_40344_n4048), .B(_abc_40344_n3500), .Y(_abc_40344_n4138) );
  NAND2X1 NAND2X1_5 ( .A(_abc_40344_n549_1), .B(_abc_40344_n548), .Y(_abc_40344_n550_1) );
  NAND2X1 NAND2X1_50 ( .A(IR_REG_4_), .B(_abc_40344_n559_1), .Y(_abc_40344_n772) );
  NAND2X1 NAND2X1_500 ( .A(_abc_40344_n4048), .B(_abc_40344_n3480), .Y(_abc_40344_n4145) );
  NAND2X1 NAND2X1_501 ( .A(_abc_40344_n4168), .B(_abc_40344_n4167_1), .Y(n598) );
  NAND2X1 NAND2X1_502 ( .A(_abc_40344_n4174), .B(_abc_40344_n4173_1), .Y(n603) );
  NAND2X1 NAND2X1_503 ( .A(_abc_40344_n4048), .B(_abc_40344_n3351), .Y(_abc_40344_n4182) );
  NAND2X1 NAND2X1_504 ( .A(_abc_40344_n3725), .B(_abc_40344_n3372), .Y(_abc_40344_n4183_1) );
  NAND2X1 NAND2X1_505 ( .A(_abc_40344_n4187_1), .B(_abc_40344_n4186), .Y(n613) );
  NAND2X1 NAND2X1_506 ( .A(_abc_40344_n4193_1), .B(_abc_40344_n4192), .Y(n618) );
  NAND2X1 NAND2X1_507 ( .A(_abc_40344_n4199_1), .B(_abc_40344_n4198), .Y(n623) );
  NAND2X1 NAND2X1_508 ( .A(_abc_40344_n4205_1), .B(_abc_40344_n4204), .Y(n628) );
  NAND2X1 NAND2X1_509 ( .A(_abc_40344_n4211_1), .B(_abc_40344_n4210), .Y(n633) );
  NAND2X1 NAND2X1_51 ( .A(_abc_40344_n668_1), .B(_abc_40344_n672), .Y(_abc_40344_n782) );
  NAND2X1 NAND2X1_510 ( .A(_abc_40344_n4217_1), .B(_abc_40344_n4216), .Y(n638) );
  NAND2X1 NAND2X1_511 ( .A(_abc_40344_n4222), .B(_abc_40344_n4219_1), .Y(_abc_40344_n4223_1) );
  NAND2X1 NAND2X1_512 ( .A(_abc_40344_n4225_1), .B(_abc_40344_n4224), .Y(n643) );
  NAND2X1 NAND2X1_513 ( .A(_abc_40344_n4230), .B(_abc_40344_n4229_1), .Y(n648) );
  NAND2X1 NAND2X1_514 ( .A(_abc_40344_n4295_1), .B(_abc_40344_n4294), .Y(n758) );
  NAND2X1 NAND2X1_515 ( .A(_abc_40344_n4298_1), .B(_abc_40344_n4297), .Y(n763) );
  NAND2X1 NAND2X1_516 ( .A(_abc_40344_n4303), .B(_abc_40344_n4302_1), .Y(n773) );
  NAND2X1 NAND2X1_517 ( .A(_abc_40344_n4306), .B(_abc_40344_n4305_1), .Y(n778) );
  NAND2X1 NAND2X1_518 ( .A(_abc_40344_n4309), .B(_abc_40344_n4308_1), .Y(n783) );
  NAND2X1 NAND2X1_519 ( .A(_abc_40344_n4312), .B(_abc_40344_n4311_1), .Y(n788) );
  NAND2X1 NAND2X1_52 ( .A(_abc_40344_n786), .B(_abc_40344_n789), .Y(_abc_40344_n790) );
  NAND2X1 NAND2X1_520 ( .A(_abc_40344_n4315), .B(_abc_40344_n4314_1), .Y(n793) );
  NAND2X1 NAND2X1_521 ( .A(_abc_40344_n4318), .B(_abc_40344_n4317_1), .Y(n798) );
  NAND2X1 NAND2X1_522 ( .A(_abc_40344_n4321), .B(_abc_40344_n4320_1), .Y(n803) );
  NAND2X1 NAND2X1_53 ( .A(IR_REG_3_), .B(_abc_40344_n539), .Y(_abc_40344_n794) );
  NAND2X1 NAND2X1_54 ( .A(_abc_40344_n706), .B(_abc_40344_n794), .Y(_abc_40344_n795) );
  NAND2X1 NAND2X1_55 ( .A(IR_REG_3_), .B(_abc_40344_n559_1), .Y(_abc_40344_n796) );
  NAND2X1 NAND2X1_56 ( .A(_abc_40344_n797), .B(_abc_40344_n705_1), .Y(_abc_40344_n798) );
  NAND2X1 NAND2X1_57 ( .A(IR_REG_27_), .B(_abc_40344_n557_1), .Y(_abc_40344_n799) );
  NAND2X1 NAND2X1_58 ( .A(IR_REG_27_), .B(_abc_40344_n559_1), .Y(_abc_40344_n801_1) );
  NAND2X1 NAND2X1_59 ( .A(DATAI_3_), .B(_abc_40344_n802), .Y(_abc_40344_n803) );
  NAND2X1 NAND2X1_6 ( .A(IR_REG_26_), .B(_abc_40344_n559_1), .Y(_abc_40344_n560) );
  NAND2X1 NAND2X1_60 ( .A(REG0_REG_3_), .B(_abc_40344_n673), .Y(_abc_40344_n805) );
  NAND2X1 NAND2X1_61 ( .A(REG1_REG_3_), .B(_abc_40344_n696), .Y(_abc_40344_n806) );
  NAND2X1 NAND2X1_62 ( .A(_abc_40344_n719), .B(_abc_40344_n814), .Y(_abc_40344_n815) );
  NAND2X1 NAND2X1_63 ( .A(_abc_40344_n811), .B(_abc_40344_n815), .Y(_abc_40344_n816) );
  NAND2X1 NAND2X1_64 ( .A(_abc_40344_n820), .B(_abc_40344_n539), .Y(_abc_40344_n821) );
  NAND2X1 NAND2X1_65 ( .A(IR_REG_2_), .B(_abc_40344_n559_1), .Y(_abc_40344_n822) );
  NAND2X1 NAND2X1_66 ( .A(REG1_REG_2_), .B(_abc_40344_n696), .Y(_abc_40344_n826_1) );
  NAND2X1 NAND2X1_67 ( .A(_abc_40344_n719), .B(_abc_40344_n832), .Y(_abc_40344_n833) );
  NAND2X1 NAND2X1_68 ( .A(DATAI_2_), .B(_abc_40344_n802), .Y(_abc_40344_n834) );
  NAND2X1 NAND2X1_69 ( .A(REG3_REG_2_), .B(_abc_40344_n685_1), .Y(_abc_40344_n839) );
  NAND2X1 NAND2X1_7 ( .A(_abc_40344_n562), .B(_abc_40344_n564), .Y(_abc_40344_n565_1) );
  NAND2X1 NAND2X1_70 ( .A(_abc_40344_n839), .B(_abc_40344_n827), .Y(_abc_40344_n840) );
  NAND2X1 NAND2X1_71 ( .A(_abc_40344_n818_1), .B(_abc_40344_n844), .Y(_abc_40344_n845) );
  NAND2X1 NAND2X1_72 ( .A(IR_REG_1_), .B(_abc_40344_n559_1), .Y(_abc_40344_n852) );
  NAND2X1 NAND2X1_73 ( .A(_abc_40344_n719), .B(_abc_40344_n866_1), .Y(_abc_40344_n867) );
  NAND2X1 NAND2X1_74 ( .A(_abc_40344_n867), .B(_abc_40344_n872), .Y(_abc_40344_n873) );
  NAND2X1 NAND2X1_75 ( .A(_abc_40344_n865), .B(_abc_40344_n873), .Y(_abc_40344_n874) );
  NAND2X1 NAND2X1_76 ( .A(_abc_40344_n722), .B(_abc_40344_n879), .Y(_abc_40344_n880) );
  NAND2X1 NAND2X1_77 ( .A(REG3_REG_0_), .B(_abc_40344_n685_1), .Y(_abc_40344_n882) );
  NAND2X1 NAND2X1_78 ( .A(_abc_40344_n882), .B(_abc_40344_n881), .Y(_abc_40344_n883) );
  NAND2X1 NAND2X1_79 ( .A(_abc_40344_n700), .B(_abc_40344_n879), .Y(_abc_40344_n890) );
  NAND2X1 NAND2X1_8 ( .A(_abc_40344_n559_1), .B(_abc_40344_n566), .Y(_abc_40344_n567_1) );
  NAND2X1 NAND2X1_80 ( .A(_abc_40344_n893), .B(_abc_40344_n876), .Y(_abc_40344_n894) );
  NAND2X1 NAND2X1_81 ( .A(_abc_40344_n843), .B(_abc_40344_n833), .Y(_abc_40344_n895) );
  NAND2X1 NAND2X1_82 ( .A(_abc_40344_n768), .B(_abc_40344_n899), .Y(_abc_40344_n900) );
  NAND2X1 NAND2X1_83 ( .A(IR_REG_7_), .B(_abc_40344_n559_1), .Y(_abc_40344_n905) );
  NAND2X1 NAND2X1_84 ( .A(_abc_40344_n906_1), .B(_abc_40344_n705_1), .Y(_abc_40344_n907) );
  NAND2X1 NAND2X1_85 ( .A(REG3_REG_7_), .B(_abc_40344_n691), .Y(_abc_40344_n909) );
  NAND2X1 NAND2X1_86 ( .A(_abc_40344_n913), .B(_abc_40344_n914), .Y(_abc_40344_n915_1) );
  NAND2X1 NAND2X1_87 ( .A(_abc_40344_n705_1), .B(_abc_40344_n917), .Y(_abc_40344_n918) );
  NAND2X1 NAND2X1_88 ( .A(_abc_40344_n760), .B(_abc_40344_n758), .Y(_abc_40344_n921) );
  NAND2X1 NAND2X1_89 ( .A(_abc_40344_n719), .B(_abc_40344_n928), .Y(_abc_40344_n929) );
  NAND2X1 NAND2X1_9 ( .A(_abc_40344_n551), .B(_abc_40344_n556), .Y(_abc_40344_n568) );
  NAND2X1 NAND2X1_90 ( .A(_abc_40344_n720), .B(_abc_40344_n930), .Y(_abc_40344_n931) );
  NAND2X1 NAND2X1_91 ( .A(_abc_40344_n933), .B(_abc_40344_n934), .Y(_abc_40344_n935_1) );
  NAND2X1 NAND2X1_92 ( .A(_abc_40344_n946), .B(_abc_40344_n949), .Y(_abc_40344_n950) );
  NAND2X1 NAND2X1_93 ( .A(_abc_40344_n953), .B(_abc_40344_n954), .Y(_abc_40344_n955_1) );
  NAND2X1 NAND2X1_94 ( .A(_abc_40344_n956), .B(_abc_40344_n957), .Y(_abc_40344_n958) );
  NAND2X1 NAND2X1_95 ( .A(_abc_40344_n976), .B(_abc_40344_n975_1), .Y(_abc_40344_n977) );
  NAND2X1 NAND2X1_96 ( .A(_abc_40344_n978), .B(_abc_40344_n980), .Y(_abc_40344_n981_1) );
  NAND2X1 NAND2X1_97 ( .A(_abc_40344_n995), .B(_abc_40344_n990), .Y(_abc_40344_n996) );
  NAND2X1 NAND2X1_98 ( .A(REG3_REG_6_), .B(REG3_REG_7_), .Y(_abc_40344_n1012) );
  NAND2X1 NAND2X1_99 ( .A(REG3_REG_16_), .B(REG3_REG_17_), .Y(_abc_40344_n1048) );
  NAND3X1 NAND3X1_1 ( .A(_abc_40344_n528), .B(_abc_40344_n529), .C(_abc_40344_n530), .Y(_abc_40344_n531) );
  NAND3X1 NAND3X1_10 ( .A(_abc_40344_n565_1), .B(_abc_40344_n567_1), .C(_abc_40344_n579), .Y(_abc_40344_n580) );
  NAND3X1 NAND3X1_100 ( .A(_abc_40344_n1076), .B(_abc_40344_n1923), .C(_abc_40344_n2102), .Y(_abc_40344_n2106) );
  NAND3X1 NAND3X1_101 ( .A(_abc_40344_n1927), .B(_abc_40344_n2107), .C(_abc_40344_n1904), .Y(_abc_40344_n2108) );
  NAND3X1 NAND3X1_102 ( .A(_abc_40344_n2099), .B(_abc_40344_n2108), .C(_abc_40344_n2105), .Y(_abc_40344_n2109) );
  NAND3X1 NAND3X1_103 ( .A(_abc_40344_n1904), .B(_abc_40344_n2127), .C(_abc_40344_n2012), .Y(_abc_40344_n2128) );
  NAND3X1 NAND3X1_104 ( .A(_abc_40344_n2128), .B(_abc_40344_n2124), .C(_abc_40344_n2114), .Y(_abc_40344_n2129) );
  NAND3X1 NAND3X1_105 ( .A(_abc_40344_n1929), .B(_abc_40344_n2132), .C(_abc_40344_n1978), .Y(_abc_40344_n2133) );
  NAND3X1 NAND3X1_106 ( .A(_abc_40344_n2136), .B(_abc_40344_n2138), .C(_abc_40344_n1904), .Y(_abc_40344_n2139) );
  NAND3X1 NAND3X1_107 ( .A(_abc_40344_n2136), .B(_abc_40344_n2148), .C(_abc_40344_n1943), .Y(_abc_40344_n2149) );
  NAND3X1 NAND3X1_108 ( .A(_abc_40344_n2133), .B(_abc_40344_n2141), .C(_abc_40344_n2154), .Y(_abc_40344_n2155) );
  NAND3X1 NAND3X1_109 ( .A(_abc_40344_n2054), .B(_abc_40344_n2094), .C(_abc_40344_n2156), .Y(_abc_40344_n2157) );
  NAND3X1 NAND3X1_11 ( .A(_abc_40344_n524), .B(_abc_40344_n525), .C(_abc_40344_n592), .Y(_abc_40344_n593_1) );
  NAND3X1 NAND3X1_110 ( .A(_abc_40344_n2162), .B(_abc_40344_n1608), .C(_abc_40344_n2163), .Y(_abc_40344_n2164) );
  NAND3X1 NAND3X1_111 ( .A(_abc_40344_n2162), .B(_abc_40344_n775_1), .C(_abc_40344_n2169), .Y(_abc_40344_n2170) );
  NAND3X1 NAND3X1_112 ( .A(_abc_40344_n2165), .B(_abc_40344_n2175), .C(_abc_40344_n2176), .Y(_abc_40344_n2177) );
  NAND3X1 NAND3X1_113 ( .A(_abc_40344_n2165), .B(_abc_40344_n733), .C(_abc_40344_n2187), .Y(_abc_40344_n2188) );
  NAND3X1 NAND3X1_114 ( .A(_abc_40344_n1796), .B(_abc_40344_n1675), .C(_abc_40344_n2222), .Y(_abc_40344_n2223) );
  NAND3X1 NAND3X1_115 ( .A(_abc_40344_n887), .B(_abc_40344_n2165), .C(_abc_40344_n1797), .Y(_abc_40344_n2224) );
  NAND3X1 NAND3X1_116 ( .A(_abc_40344_n2162), .B(_abc_40344_n749_1), .C(_abc_40344_n2255), .Y(_abc_40344_n2256) );
  NAND3X1 NAND3X1_117 ( .A(_abc_40344_n2260), .B(_abc_40344_n2261), .C(_abc_40344_n2259), .Y(_abc_40344_n2262) );
  NAND3X1 NAND3X1_118 ( .A(_abc_40344_n2269), .B(_abc_40344_n2271), .C(_abc_40344_n2270), .Y(_abc_40344_n2272) );
  NAND3X1 NAND3X1_119 ( .A(_abc_40344_n2246), .B(_abc_40344_n2247), .C(_abc_40344_n2269), .Y(_abc_40344_n2273) );
  NAND3X1 NAND3X1_12 ( .A(_abc_40344_n549_1), .B(_abc_40344_n597), .C(_abc_40344_n548), .Y(_abc_40344_n598) );
  NAND3X1 NAND3X1_120 ( .A(_abc_40344_n2272), .B(_abc_40344_n2273), .C(_abc_40344_n2285), .Y(_abc_40344_n2286) );
  NAND3X1 NAND3X1_121 ( .A(_abc_40344_n2349), .B(_abc_40344_n2350), .C(_abc_40344_n2348), .Y(_abc_40344_n2351) );
  NAND3X1 NAND3X1_122 ( .A(_abc_40344_n627), .B(_abc_40344_n2413), .C(_abc_40344_n2412), .Y(_abc_40344_n2414) );
  NAND3X1 NAND3X1_123 ( .A(_abc_40344_n640), .B(_abc_40344_n2158), .C(_abc_40344_n2414), .Y(_abc_40344_n2415) );
  NAND3X1 NAND3X1_124 ( .A(_abc_40344_n2210), .B(_abc_40344_n2198), .C(_abc_40344_n2209), .Y(_abc_40344_n2417) );
  NAND3X1 NAND3X1_125 ( .A(_abc_40344_n2425), .B(_abc_40344_n2428_1), .C(_abc_40344_n2417), .Y(_abc_40344_n2429) );
  NAND3X1 NAND3X1_126 ( .A(_abc_40344_n1675), .B(_abc_40344_n2173), .C(_abc_40344_n879), .Y(_abc_40344_n2435_1) );
  NAND3X1 NAND3X1_127 ( .A(_abc_40344_n2183), .B(_abc_40344_n2184), .C(_abc_40344_n2237), .Y(_abc_40344_n2442) );
  NAND3X1 NAND3X1_128 ( .A(_abc_40344_n2258), .B(_abc_40344_n2443), .C(_abc_40344_n2237), .Y(_abc_40344_n2444) );
  NAND3X1 NAND3X1_129 ( .A(_abc_40344_n2442), .B(_abc_40344_n2444), .C(_abc_40344_n2441), .Y(_abc_40344_n2445) );
  NAND3X1 NAND3X1_13 ( .A(IR_REG_27_), .B(_abc_40344_n607), .C(_abc_40344_n577_1), .Y(_abc_40344_n608_1) );
  NAND3X1 NAND3X1_130 ( .A(_abc_40344_n2284), .B(_abc_40344_n2273), .C(_abc_40344_n2280), .Y(_abc_40344_n2447) );
  NAND3X1 NAND3X1_131 ( .A(_abc_40344_n2485), .B(_abc_40344_n2496_1), .C(_abc_40344_n2481), .Y(_abc_40344_n2497) );
  NAND3X1 NAND3X1_132 ( .A(_abc_40344_n2470), .B(_abc_40344_n2474), .C(_abc_40344_n2508), .Y(_abc_40344_n2509) );
  NAND3X1 NAND3X1_133 ( .A(_abc_40344_n2533), .B(_abc_40344_n2539), .C(_abc_40344_n2548), .Y(_abc_40344_n2549_1) );
  NAND3X1 NAND3X1_134 ( .A(_abc_40344_n2526), .B(_abc_40344_n2550), .C(_abc_40344_n2524), .Y(_abc_40344_n2551) );
  NAND3X1 NAND3X1_135 ( .A(_abc_40344_n2517), .B(_abc_40344_n2514), .C(_abc_40344_n2552), .Y(_abc_40344_n2553) );
  NAND3X1 NAND3X1_136 ( .A(_abc_40344_n2510), .B(_abc_40344_n2554), .C(_abc_40344_n2559), .Y(_abc_40344_n2560) );
  NAND3X1 NAND3X1_137 ( .A(_abc_40344_n1934), .B(_abc_40344_n2596), .C(_abc_40344_n2595), .Y(_abc_40344_n2597) );
  NAND3X1 NAND3X1_138 ( .A(_abc_40344_n2478_1), .B(_abc_40344_n2544), .C(_abc_40344_n2599_1), .Y(_abc_40344_n2600) );
  NAND3X1 NAND3X1_139 ( .A(_abc_40344_n1939), .B(_abc_40344_n2602), .C(_abc_40344_n2593_1), .Y(_abc_40344_n2603) );
  NAND3X1 NAND3X1_14 ( .A(IR_REG_31_), .B(_abc_40344_n608_1), .C(_abc_40344_n606), .Y(_abc_40344_n609) );
  NAND3X1 NAND3X1_140 ( .A(_abc_40344_n2603), .B(_abc_40344_n2607), .C(_abc_40344_n2598), .Y(_abc_40344_n2608) );
  NAND3X1 NAND3X1_141 ( .A(_abc_40344_n2498), .B(_abc_40344_n2060), .C(_abc_40344_n2083), .Y(_abc_40344_n2624) );
  NAND3X1 NAND3X1_142 ( .A(_abc_40344_n2137), .B(_abc_40344_n2024), .C(_abc_40344_n2632), .Y(_abc_40344_n2633) );
  NAND3X1 NAND3X1_143 ( .A(_abc_40344_n2586), .B(_abc_40344_n2638), .C(_abc_40344_n2639), .Y(_abc_40344_n2640) );
  NAND3X1 NAND3X1_144 ( .A(_abc_40344_n648), .B(_abc_40344_n2657), .C(_abc_40344_n2560), .Y(_abc_40344_n2658) );
  NAND3X1 NAND3X1_145 ( .A(_abc_40344_n587), .B(_abc_40344_n2669), .C(_abc_40344_n2668), .Y(_abc_40344_n2670) );
  NAND3X1 NAND3X1_146 ( .A(_abc_40344_n2711), .B(_abc_40344_n2725), .C(_abc_40344_n2710), .Y(n1046) );
  NAND3X1 NAND3X1_147 ( .A(_abc_40344_n2746), .B(_abc_40344_n2758), .C(_abc_40344_n2710), .Y(n1038) );
  NAND3X1 NAND3X1_148 ( .A(_abc_40344_n2776), .B(_abc_40344_n2779), .C(_abc_40344_n2777), .Y(_abc_40344_n2796) );
  NAND3X1 NAND3X1_149 ( .A(_abc_40344_n2780), .B(_abc_40344_n2799), .C(_abc_40344_n2796), .Y(_abc_40344_n2812) );
  NAND3X1 NAND3X1_15 ( .A(_abc_40344_n620), .B(_abc_40344_n575_1), .C(_abc_40344_n621), .Y(_abc_40344_n622) );
  NAND3X1 NAND3X1_150 ( .A(_abc_40344_n1007), .B(_abc_40344_n2798), .C(_abc_40344_n2812), .Y(_abc_40344_n2814) );
  NAND3X1 NAND3X1_151 ( .A(_abc_40344_n2848), .B(_abc_40344_n2864), .C(_abc_40344_n2886), .Y(_abc_40344_n2887) );
  NAND3X1 NAND3X1_152 ( .A(_abc_40344_n2898), .B(_abc_40344_n2900), .C(_abc_40344_n2899), .Y(_abc_40344_n2901) );
  NAND3X1 NAND3X1_153 ( .A(_abc_40344_n2866), .B(_abc_40344_n2882), .C(_abc_40344_n2887), .Y(_abc_40344_n2904) );
  NAND3X1 NAND3X1_154 ( .A(_abc_40344_n1252), .B(_abc_40344_n2884), .C(_abc_40344_n2904), .Y(_abc_40344_n2907) );
  NAND3X1 NAND3X1_155 ( .A(_abc_40344_n2914), .B(_abc_40344_n2892), .C(_abc_40344_n2894), .Y(_abc_40344_n2915) );
  NAND3X1 NAND3X1_156 ( .A(_abc_40344_n2919), .B(_abc_40344_n2921), .C(_abc_40344_n2920), .Y(_abc_40344_n2922) );
  NAND3X1 NAND3X1_157 ( .A(_abc_40344_n2891), .B(_abc_40344_n2940), .C(_abc_40344_n2915), .Y(_abc_40344_n2941) );
  NAND3X1 NAND3X1_158 ( .A(_abc_40344_n1206), .B(_abc_40344_n2929), .C(_abc_40344_n2949), .Y(_abc_40344_n2951) );
  NAND3X1 NAND3X1_159 ( .A(_abc_40344_n2939), .B(_abc_40344_n2935), .C(_abc_40344_n2941), .Y(_abc_40344_n2964) );
  NAND3X1 NAND3X1_16 ( .A(IR_REG_31_), .B(_abc_40344_n622), .C(_abc_40344_n623), .Y(_abc_40344_n624) );
  NAND3X1 NAND3X1_160 ( .A(REG1_REG_15_), .B(_abc_40344_n2927), .C(_abc_40344_n2931), .Y(_abc_40344_n2975) );
  NAND3X1 NAND3X1_161 ( .A(_abc_40344_n2951), .B(_abc_40344_n2973), .C(_abc_40344_n2996), .Y(_abc_40344_n2997) );
  NAND3X1 NAND3X1_162 ( .A(_abc_40344_n3007), .B(_abc_40344_n3012), .C(_abc_40344_n3000), .Y(n986) );
  NAND3X1 NAND3X1_163 ( .A(_abc_40344_n2937), .B(_abc_40344_n2962), .C(_abc_40344_n2964), .Y(_abc_40344_n3020) );
  NAND3X1 NAND3X1_164 ( .A(_abc_40344_n2960), .B(_abc_40344_n2978), .C(_abc_40344_n3020), .Y(_abc_40344_n3021) );
  NAND3X1 NAND3X1_165 ( .A(_abc_40344_n2980), .B(_abc_40344_n3002), .C(_abc_40344_n3021), .Y(_abc_40344_n3022) );
  NAND3X1 NAND3X1_166 ( .A(_abc_40344_n2971), .B(_abc_40344_n2992), .C(_abc_40344_n2997), .Y(_abc_40344_n3029) );
  NAND3X1 NAND3X1_167 ( .A(_abc_40344_n2993), .B(_abc_40344_n3028), .C(_abc_40344_n3029), .Y(_abc_40344_n3031) );
  NAND3X1 NAND3X1_168 ( .A(_abc_40344_n602), .B(_abc_40344_n648), .C(_abc_40344_n2684), .Y(_abc_40344_n3034) );
  NAND3X1 NAND3X1_169 ( .A(_abc_40344_n602), .B(_abc_40344_n648), .C(_abc_40344_n2677), .Y(_abc_40344_n3035) );
  NAND3X1 NAND3X1_17 ( .A(IR_REG_31_), .B(_abc_40344_n568), .C(_abc_40344_n634), .Y(_abc_40344_n635) );
  NAND3X1 NAND3X1_170 ( .A(_abc_40344_n3034), .B(_abc_40344_n3035), .C(_abc_40344_n3036), .Y(_abc_40344_n3037) );
  NAND3X1 NAND3X1_171 ( .A(_abc_40344_n3001), .B(_abc_40344_n3039), .C(_abc_40344_n3022), .Y(_abc_40344_n3040) );
  NAND3X1 NAND3X1_172 ( .A(_abc_40344_n2973), .B(_abc_40344_n2993), .C(_abc_40344_n3049), .Y(_abc_40344_n3050) );
  NAND3X1 NAND3X1_173 ( .A(_abc_40344_n3054), .B(_abc_40344_n3053), .C(_abc_40344_n3055), .Y(_abc_40344_n3056) );
  NAND3X1 NAND3X1_174 ( .A(_abc_40344_n978), .B(_abc_40344_n990), .C(_abc_40344_n3064), .Y(_abc_40344_n3065) );
  NAND3X1 NAND3X1_175 ( .A(_abc_40344_n3080), .B(_abc_40344_n3081_1), .C(_abc_40344_n3079), .Y(_abc_40344_n3082) );
  NAND3X1 NAND3X1_176 ( .A(_abc_40344_n3089), .B(_abc_40344_n3090), .C(_abc_40344_n3086), .Y(_abc_40344_n3091) );
  NAND3X1 NAND3X1_177 ( .A(_abc_40344_n3157), .B(_abc_40344_n3134), .C(_abc_40344_n3155), .Y(_abc_40344_n3158) );
  NAND3X1 NAND3X1_178 ( .A(_abc_40344_n625), .B(_abc_40344_n646), .C(_abc_40344_n699), .Y(_abc_40344_n3222) );
  NAND3X1 NAND3X1_179 ( .A(_abc_40344_n3213), .B(_abc_40344_n3223), .C(_abc_40344_n3214), .Y(_abc_40344_n3224) );
  NAND3X1 NAND3X1_18 ( .A(_abc_40344_n524), .B(_abc_40344_n525), .C(_abc_40344_n546_1), .Y(_abc_40344_n653) );
  NAND3X1 NAND3X1_180 ( .A(_abc_40344_n3221_1), .B(_abc_40344_n3230), .C(_abc_40344_n3224), .Y(_abc_40344_n3231) );
  NAND3X1 NAND3X1_181 ( .A(_abc_40344_n3298), .B(_abc_40344_n3303), .C(_abc_40344_n3324), .Y(_abc_40344_n3325) );
  NAND3X1 NAND3X1_182 ( .A(_abc_40344_n2030), .B(_abc_40344_n1945), .C(_abc_40344_n3327), .Y(_abc_40344_n3328) );
  NAND3X1 NAND3X1_183 ( .A(_abc_40344_n3371), .B(_abc_40344_n3377), .C(_abc_40344_n3370), .Y(n933) );
  NAND3X1 NAND3X1_184 ( .A(_abc_40344_n2517), .B(_abc_40344_n3360), .C(_abc_40344_n3357), .Y(_abc_40344_n3382) );
  NAND3X1 NAND3X1_185 ( .A(_abc_40344_n3429), .B(_abc_40344_n3428), .C(_abc_40344_n3435), .Y(_abc_40344_n3436) );
  NAND3X1 NAND3X1_186 ( .A(_abc_40344_n3472), .B(_abc_40344_n3474), .C(_abc_40344_n3469), .Y(_abc_40344_n3475) );
  NAND3X1 NAND3X1_187 ( .A(_abc_40344_n3495), .B(_abc_40344_n3496), .C(_abc_40344_n3491), .Y(_abc_40344_n3497) );
  NAND3X1 NAND3X1_188 ( .A(_abc_40344_n3507), .B(_abc_40344_n3516), .C(_abc_40344_n3506_1), .Y(n898) );
  NAND3X1 NAND3X1_189 ( .A(_abc_40344_n3568), .B(_abc_40344_n3570), .C(_abc_40344_n3567), .Y(_abc_40344_n3571) );
  NAND3X1 NAND3X1_19 ( .A(_abc_40344_n551), .B(_abc_40344_n594), .C(_abc_40344_n657), .Y(_abc_40344_n658_1) );
  NAND3X1 NAND3X1_190 ( .A(_abc_40344_n3601), .B(_abc_40344_n3603), .C(_abc_40344_n3606), .Y(_abc_40344_n3607) );
  NAND3X1 NAND3X1_191 ( .A(_abc_40344_n3629), .B(_abc_40344_n3631), .C(_abc_40344_n3626), .Y(_abc_40344_n3632_1) );
  NAND3X1 NAND3X1_192 ( .A(_abc_40344_n3716), .B(_abc_40344_n3722), .C(_abc_40344_n3715), .Y(n843) );
  NAND3X1 NAND3X1_193 ( .A(nRESET_G), .B(_abc_40344_n3737), .C(_abc_40344_n3736), .Y(n838) );
  NAND3X1 NAND3X1_194 ( .A(nRESET_G), .B(_abc_40344_n3754), .C(_abc_40344_n3753), .Y(n833) );
  NAND3X1 NAND3X1_195 ( .A(_abc_40344_n3768), .B(_abc_40344_n3765), .C(_abc_40344_n3766_1), .Y(n828) );
  NAND3X1 NAND3X1_196 ( .A(_abc_40344_n3779_1), .B(_abc_40344_n3782_1), .C(_abc_40344_n3780_1), .Y(n823) );
  NAND3X1 NAND3X1_197 ( .A(nRESET_G), .B(_abc_40344_n3872), .C(_abc_40344_n3871_1), .Y(n318) );
  NAND3X1 NAND3X1_198 ( .A(_abc_40344_n4002), .B(_abc_40344_n3210), .C(_abc_40344_n4003), .Y(_abc_40344_n4004) );
  NAND3X1 NAND3X1_199 ( .A(_abc_40344_n4001), .B(_abc_40344_n3121), .C(_abc_40344_n4004), .Y(_abc_40344_n4005) );
  NAND3X1 NAND3X1_2 ( .A(_abc_40344_n536), .B(_abc_40344_n537_1), .C(_abc_40344_n538_1), .Y(_abc_40344_n539) );
  NAND3X1 NAND3X1_20 ( .A(_abc_40344_n659), .B(_abc_40344_n535), .C(_abc_40344_n543), .Y(_abc_40344_n660) );
  NAND3X1 NAND3X1_200 ( .A(_abc_40344_n3999_1), .B(_abc_40344_n4000), .C(_abc_40344_n4005), .Y(_abc_40344_n4006_1) );
  NAND3X1 NAND3X1_201 ( .A(_abc_40344_n4001), .B(_abc_40344_n2558), .C(_abc_40344_n4007), .Y(_abc_40344_n4008) );
  NAND3X1 NAND3X1_202 ( .A(_abc_40344_n3223), .B(_abc_40344_n4008), .C(_abc_40344_n4006_1), .Y(_abc_40344_n4009) );
  NAND3X1 NAND3X1_203 ( .A(_abc_40344_n2394), .B(_abc_40344_n3096), .C(_abc_40344_n3095), .Y(_abc_40344_n4022) );
  NAND3X1 NAND3X1_204 ( .A(_abc_40344_n990), .B(_abc_40344_n1029_1), .C(_abc_40344_n951), .Y(_abc_40344_n4039) );
  NAND3X1 NAND3X1_205 ( .A(_abc_40344_n3762), .B(_abc_40344_n4055), .C(_abc_40344_n4057), .Y(_abc_40344_n4058_1) );
  NAND3X1 NAND3X1_206 ( .A(nRESET_G), .B(_abc_40344_n4068), .C(_abc_40344_n4067), .Y(n518) );
  NAND3X1 NAND3X1_207 ( .A(_abc_40344_n3713), .B(_abc_40344_n4070_1), .C(_abc_40344_n3712), .Y(_abc_40344_n4071) );
  NAND3X1 NAND3X1_208 ( .A(nRESET_G), .B(_abc_40344_n4128), .C(_abc_40344_n4127), .Y(n568) );
  NAND3X1 NAND3X1_209 ( .A(_abc_40344_n4130), .B(_abc_40344_n4131_1), .C(_abc_40344_n4132), .Y(_abc_40344_n4133) );
  NAND3X1 NAND3X1_21 ( .A(_abc_40344_n662), .B(_abc_40344_n655), .C(_abc_40344_n663), .Y(_abc_40344_n664) );
  NAND3X1 NAND3X1_210 ( .A(nRESET_G), .B(_abc_40344_n4135), .C(_abc_40344_n4134), .Y(n573) );
  NAND3X1 NAND3X1_211 ( .A(_abc_40344_n4137_1), .B(_abc_40344_n4138), .C(_abc_40344_n4139), .Y(_abc_40344_n4140) );
  NAND3X1 NAND3X1_212 ( .A(nRESET_G), .B(_abc_40344_n4142), .C(_abc_40344_n4141), .Y(n578) );
  NAND3X1 NAND3X1_213 ( .A(_abc_40344_n4145), .B(_abc_40344_n4147), .C(_abc_40344_n3489), .Y(_abc_40344_n4148) );
  NAND3X1 NAND3X1_214 ( .A(nRESET_G), .B(_abc_40344_n4154), .C(_abc_40344_n4153), .Y(n588) );
  NAND3X1 NAND3X1_215 ( .A(nRESET_G), .B(_abc_40344_n4162), .C(_abc_40344_n4161), .Y(n593) );
  NAND3X1 NAND3X1_216 ( .A(_abc_40344_n4182), .B(_abc_40344_n4184), .C(_abc_40344_n4183_1), .Y(_abc_40344_n4185_1) );
  NAND3X1 NAND3X1_217 ( .A(_abc_40344_n4048), .B(_abc_40344_n4008), .C(_abc_40344_n4006_1), .Y(_abc_40344_n4219_1) );
  NAND3X1 NAND3X1_218 ( .A(nRESET_G), .B(_abc_40344_n4235), .C(_abc_40344_n4234), .Y(n653) );
  NAND3X1 NAND3X1_219 ( .A(nRESET_G), .B(_abc_40344_n4327), .C(_abc_40344_n4326_1), .Y(n813) );
  NAND3X1 NAND3X1_22 ( .A(IR_REG_31_), .B(_abc_40344_n664), .C(_abc_40344_n661), .Y(_abc_40344_n674_1) );
  NAND3X1 NAND3X1_23 ( .A(_abc_40344_n655), .B(_abc_40344_n659), .C(_abc_40344_n574), .Y(_abc_40344_n676) );
  NAND3X1 NAND3X1_24 ( .A(IR_REG_31_), .B(_abc_40344_n676), .C(_abc_40344_n682), .Y(_abc_40344_n683_1) );
  NAND3X1 NAND3X1_25 ( .A(_abc_40344_n602), .B(_abc_40344_n712), .C(_abc_40344_n610_1), .Y(_abc_40344_n713_1) );
  NAND3X1 NAND3X1_26 ( .A(_abc_40344_n740), .B(_abc_40344_n741), .C(_abc_40344_n735), .Y(_abc_40344_n742) );
  NAND3X1 NAND3X1_27 ( .A(_abc_40344_n743), .B(_abc_40344_n766), .C(_abc_40344_n765), .Y(_abc_40344_n769) );
  NAND3X1 NAND3X1_28 ( .A(_abc_40344_n602), .B(_abc_40344_n774), .C(_abc_40344_n610_1), .Y(_abc_40344_n775_1) );
  NAND3X1 NAND3X1_29 ( .A(REG0_REG_4_), .B(_abc_40344_n782), .C(_abc_40344_n781), .Y(_abc_40344_n783) );
  NAND3X1 NAND3X1_3 ( .A(_abc_40344_n527), .B(_abc_40344_n535), .C(_abc_40344_n543), .Y(_abc_40344_n544) );
  NAND3X1 NAND3X1_30 ( .A(REG1_REG_4_), .B(_abc_40344_n760), .C(_abc_40344_n781), .Y(_abc_40344_n784) );
  NAND3X1 NAND3X1_31 ( .A(_abc_40344_n783), .B(_abc_40344_n784), .C(_abc_40344_n780_1), .Y(_abc_40344_n785) );
  NAND3X1 NAND3X1_32 ( .A(IR_REG_31_), .B(_abc_40344_n598), .C(_abc_40344_n799), .Y(_abc_40344_n800_1) );
  NAND3X1 NAND3X1_33 ( .A(_abc_40344_n800_1), .B(_abc_40344_n801_1), .C(_abc_40344_n602), .Y(_abc_40344_n802) );
  NAND3X1 NAND3X1_34 ( .A(_abc_40344_n807_1), .B(_abc_40344_n805), .C(_abc_40344_n806), .Y(_abc_40344_n808) );
  NAND3X1 NAND3X1_35 ( .A(_abc_40344_n602), .B(_abc_40344_n823), .C(_abc_40344_n610_1), .Y(_abc_40344_n824_1) );
  NAND3X1 NAND3X1_36 ( .A(REG2_REG_2_), .B(_abc_40344_n758), .C(_abc_40344_n782), .Y(_abc_40344_n827) );
  NAND3X1 NAND3X1_37 ( .A(_abc_40344_n826_1), .B(_abc_40344_n827), .C(_abc_40344_n828), .Y(_abc_40344_n829_1) );
  NAND3X1 NAND3X1_38 ( .A(_abc_40344_n831), .B(_abc_40344_n843), .C(_abc_40344_n833), .Y(_abc_40344_n844) );
  NAND3X1 NAND3X1_39 ( .A(_abc_40344_n602), .B(_abc_40344_n854_1), .C(_abc_40344_n610_1), .Y(_abc_40344_n855) );
  NAND3X1 NAND3X1_4 ( .A(_abc_40344_n554_1), .B(_abc_40344_n551), .C(_abc_40344_n556), .Y(_abc_40344_n557_1) );
  NAND3X1 NAND3X1_40 ( .A(REG3_REG_1_), .B(_abc_40344_n760), .C(_abc_40344_n758), .Y(_abc_40344_n858) );
  NAND3X1 NAND3X1_41 ( .A(REG2_REG_1_), .B(_abc_40344_n758), .C(_abc_40344_n782), .Y(_abc_40344_n861) );
  NAND3X1 NAND3X1_42 ( .A(_abc_40344_n602), .B(_abc_40344_n853), .C(_abc_40344_n610_1), .Y(_abc_40344_n868) );
  NAND3X1 NAND3X1_43 ( .A(_abc_40344_n875), .B(_abc_40344_n867), .C(_abc_40344_n872), .Y(_abc_40344_n876) );
  NAND3X1 NAND3X1_44 ( .A(IR_REG_0_), .B(_abc_40344_n602), .C(_abc_40344_n610_1), .Y(_abc_40344_n878) );
  NAND3X1 NAND3X1_45 ( .A(REG2_REG_0_), .B(_abc_40344_n758), .C(_abc_40344_n782), .Y(_abc_40344_n881) );
  NAND3X1 NAND3X1_46 ( .A(_abc_40344_n874), .B(_abc_40344_n896), .C(_abc_40344_n894), .Y(_abc_40344_n897) );
  NAND3X1 NAND3X1_47 ( .A(_abc_40344_n791), .B(_abc_40344_n847), .C(_abc_40344_n897), .Y(_abc_40344_n898) );
  NAND3X1 NAND3X1_48 ( .A(_abc_40344_n769), .B(_abc_40344_n790), .C(_abc_40344_n898), .Y(_abc_40344_n899) );
  NAND3X1 NAND3X1_49 ( .A(_abc_40344_n916), .B(_abc_40344_n931), .C(_abc_40344_n929), .Y(_abc_40344_n933) );
  NAND3X1 NAND3X1_5 ( .A(IR_REG_31_), .B(_abc_40344_n557_1), .C(_abc_40344_n553_1), .Y(_abc_40344_n558) );
  NAND3X1 NAND3X1_50 ( .A(_abc_40344_n715), .B(_abc_40344_n724), .C(_abc_40344_n725), .Y(_abc_40344_n934) );
  NAND3X1 NAND3X1_51 ( .A(B_REG), .B(_abc_40344_n947), .C(_abc_40344_n948_1), .Y(_abc_40344_n949) );
  NAND3X1 NAND3X1_52 ( .A(_abc_40344_n962), .B(_abc_40344_n963), .C(_abc_40344_n959), .Y(_abc_40344_n964) );
  NAND3X1 NAND3X1_53 ( .A(_abc_40344_n965), .B(_abc_40344_n966), .C(_abc_40344_n967), .Y(_abc_40344_n968) );
  NAND3X1 NAND3X1_54 ( .A(_abc_40344_n972_1), .B(_abc_40344_n973), .C(_abc_40344_n971), .Y(_abc_40344_n974) );
  NAND3X1 NAND3X1_55 ( .A(REG3_REG_12_), .B(_abc_40344_n1054), .C(_abc_40344_n1051_1), .Y(_abc_40344_n1055) );
  NAND3X1 NAND3X1_56 ( .A(REG3_REG_14_), .B(REG3_REG_15_), .C(_abc_40344_n1056), .Y(_abc_40344_n1057) );
  NAND3X1 NAND3X1_57 ( .A(REG3_REG_22_), .B(REG3_REG_23_), .C(_abc_40344_n1062), .Y(_abc_40344_n1063) );
  NAND3X1 NAND3X1_58 ( .A(REG3_REG_26_), .B(REG3_REG_27_), .C(_abc_40344_n1064), .Y(_abc_40344_n1067) );
  NAND3X1 NAND3X1_59 ( .A(_abc_40344_n1107), .B(_abc_40344_n1106), .C(_abc_40344_n1108), .Y(_abc_40344_n1109) );
  NAND3X1 NAND3X1_6 ( .A(IR_REG_31_), .B(_abc_40344_n563_1), .C(_abc_40344_n550_1), .Y(_abc_40344_n564) );
  NAND3X1 NAND3X1_60 ( .A(_abc_40344_n1243), .B(_abc_40344_n532), .C(_abc_40344_n1246), .Y(_abc_40344_n1247) );
  NAND3X1 NAND3X1_61 ( .A(_abc_40344_n1267), .B(_abc_40344_n1318), .C(_abc_40344_n1317_1), .Y(_abc_40344_n1319) );
  NAND3X1 NAND3X1_62 ( .A(_abc_40344_n933), .B(_abc_40344_n934), .C(_abc_40344_n769), .Y(_abc_40344_n1387) );
  NAND3X1 NAND3X1_63 ( .A(_abc_40344_n790), .B(_abc_40344_n1388), .C(_abc_40344_n898), .Y(_abc_40344_n1389) );
  NAND3X1 NAND3X1_64 ( .A(_abc_40344_n1390), .B(_abc_40344_n1386), .C(_abc_40344_n1389), .Y(_abc_40344_n1391) );
  NAND3X1 NAND3X1_65 ( .A(_abc_40344_n1368), .B(_abc_40344_n1392), .C(_abc_40344_n1391), .Y(_abc_40344_n1393) );
  NAND3X1 NAND3X1_66 ( .A(_abc_40344_n1241), .B(_abc_40344_n1340), .C(_abc_40344_n1393), .Y(_abc_40344_n1394) );
  NAND3X1 NAND3X1_67 ( .A(_abc_40344_n1217), .B(_abc_40344_n1239), .C(_abc_40344_n1394), .Y(_abc_40344_n1395) );
  NAND3X1 NAND3X1_68 ( .A(_abc_40344_n1426), .B(_abc_40344_n1425), .C(_abc_40344_n1427), .Y(_abc_40344_n1428) );
  NAND3X1 NAND3X1_69 ( .A(_abc_40344_n1098), .B(_abc_40344_n1116), .C(_abc_40344_n1459), .Y(_abc_40344_n1460) );
  NAND3X1 NAND3X1_7 ( .A(_abc_40344_n532), .B(_abc_40344_n533), .C(_abc_40344_n570), .Y(_abc_40344_n571_1) );
  NAND3X1 NAND3X1_70 ( .A(_abc_40344_n1141), .B(_abc_40344_n1527), .C(_abc_40344_n1526), .Y(_abc_40344_n1528) );
  NAND3X1 NAND3X1_71 ( .A(_abc_40344_n1143), .B(_abc_40344_n1529), .C(_abc_40344_n1528), .Y(_abc_40344_n1530) );
  NAND3X1 NAND3X1_72 ( .A(_abc_40344_n1116), .B(_abc_40344_n1457), .C(_abc_40344_n1530), .Y(_abc_40344_n1531) );
  NAND3X1 NAND3X1_73 ( .A(_abc_40344_n1096), .B(_abc_40344_n1118_1), .C(_abc_40344_n1531), .Y(_abc_40344_n1532) );
  NAND3X1 NAND3X1_74 ( .A(_abc_40344_n538_1), .B(_abc_40344_n602), .C(_abc_40344_n610_1), .Y(_abc_40344_n1796) );
  NAND3X1 NAND3X1_75 ( .A(_abc_40344_n1267), .B(_abc_40344_n1313), .C(_abc_40344_n1317_1), .Y(_abc_40344_n1828) );
  NAND3X1 NAND3X1_76 ( .A(_abc_40344_n1904), .B(_abc_40344_n1909), .C(_abc_40344_n1929), .Y(_abc_40344_n1930) );
  NAND3X1 NAND3X1_77 ( .A(_abc_40344_n1934), .B(_abc_40344_n1936), .C(_abc_40344_n1932), .Y(_abc_40344_n1937) );
  NAND3X1 NAND3X1_78 ( .A(_abc_40344_n685_1), .B(_abc_40344_n1465), .C(_abc_40344_n1464), .Y(_abc_40344_n1941) );
  NAND3X1 NAND3X1_79 ( .A(_abc_40344_n1463), .B(_abc_40344_n1470), .C(_abc_40344_n1941), .Y(_abc_40344_n1942) );
  NAND3X1 NAND3X1_8 ( .A(_abc_40344_n540), .B(_abc_40344_n541_1), .C(_abc_40344_n572), .Y(_abc_40344_n573_1) );
  NAND3X1 NAND3X1_80 ( .A(_abc_40344_n1942), .B(_abc_40344_n1944), .C(_abc_40344_n1945), .Y(_abc_40344_n1946) );
  NAND3X1 NAND3X1_81 ( .A(_abc_40344_n1940), .B(_abc_40344_n1946), .C(_abc_40344_n1965), .Y(_abc_40344_n1966) );
  NAND3X1 NAND3X1_82 ( .A(_abc_40344_n1904), .B(_abc_40344_n1980), .C(_abc_40344_n1929), .Y(_abc_40344_n1981) );
  NAND3X1 NAND3X1_83 ( .A(_abc_40344_n1984), .B(_abc_40344_n1985), .C(_abc_40344_n1976), .Y(_abc_40344_n1986) );
  NAND3X1 NAND3X1_84 ( .A(_abc_40344_n1997), .B(_abc_40344_n1999), .C(_abc_40344_n1946), .Y(_abc_40344_n2000) );
  NAND3X1 NAND3X1_85 ( .A(_abc_40344_n2001), .B(_abc_40344_n1936), .C(_abc_40344_n2003), .Y(_abc_40344_n2004) );
  NAND3X1 NAND3X1_86 ( .A(_abc_40344_n1925), .B(_abc_40344_n1927), .C(_abc_40344_n2010), .Y(_abc_40344_n2011) );
  NAND3X1 NAND3X1_87 ( .A(_abc_40344_n602), .B(_abc_40344_n2020), .C(_abc_40344_n610_1), .Y(_abc_40344_n2021) );
  NAND3X1 NAND3X1_88 ( .A(_abc_40344_n1929), .B(_abc_40344_n2032), .C(_abc_40344_n2034), .Y(_abc_40344_n2035) );
  NAND3X1 NAND3X1_89 ( .A(_abc_40344_n1929), .B(_abc_40344_n2040), .C(_abc_40344_n2034), .Y(_abc_40344_n2041) );
  NAND3X1 NAND3X1_9 ( .A(_abc_40344_n527), .B(_abc_40344_n575_1), .C(_abc_40344_n574), .Y(_abc_40344_n576) );
  NAND3X1 NAND3X1_90 ( .A(_abc_40344_n1955), .B(_abc_40344_n1946), .C(_abc_40344_n2001), .Y(_abc_40344_n2046) );
  NAND3X1 NAND3X1_91 ( .A(_abc_40344_n2047), .B(_abc_40344_n1929), .C(_abc_40344_n2045), .Y(_abc_40344_n2048) );
  NAND3X1 NAND3X1_92 ( .A(_abc_40344_n1962), .B(_abc_40344_n2049), .C(_abc_40344_n1960), .Y(_abc_40344_n2050) );
  NAND3X1 NAND3X1_93 ( .A(_abc_40344_n1929), .B(_abc_40344_n2051), .C(_abc_40344_n2034), .Y(_abc_40344_n2052) );
  NAND3X1 NAND3X1_94 ( .A(_abc_40344_n2048), .B(_abc_40344_n2041), .C(_abc_40344_n2052), .Y(_abc_40344_n2053) );
  NAND3X1 NAND3X1_95 ( .A(_abc_40344_n1904), .B(_abc_40344_n2084), .C(_abc_40344_n2086), .Y(_abc_40344_n2087) );
  NAND3X1 NAND3X1_96 ( .A(_abc_40344_n813), .B(_abc_40344_n809), .C(_abc_40344_n2089), .Y(_abc_40344_n2090) );
  NAND3X1 NAND3X1_97 ( .A(_abc_40344_n1929), .B(_abc_40344_n2091), .C(_abc_40344_n2005), .Y(_abc_40344_n2092) );
  NAND3X1 NAND3X1_98 ( .A(_abc_40344_n2087), .B(_abc_40344_n2092), .C(_abc_40344_n2081), .Y(_abc_40344_n2093) );
  NAND3X1 NAND3X1_99 ( .A(_abc_40344_n1649), .B(_abc_40344_n1923), .C(_abc_40344_n2102), .Y(_abc_40344_n2103) );
  NOR2X1 NOR2X1_1 ( .A(IR_REG_17_), .B(IR_REG_16_), .Y(_abc_40344_n524) );
  NOR2X1 NOR2X1_10 ( .A(IR_REG_19_), .B(IR_REG_18_), .Y(_abc_40344_n546_1) );
  NOR2X1 NOR2X1_100 ( .A(_abc_40344_n1235), .B(_abc_40344_n1238), .Y(_abc_40344_n1240_1) );
  NOR2X1 NOR2X1_101 ( .A(_abc_40344_n542_1), .B(_abc_40344_n706), .Y(_abc_40344_n1244) );
  NOR2X1 NOR2X1_102 ( .A(IR_REG_9_), .B(_abc_40344_n1245), .Y(_abc_40344_n1246) );
  NOR2X1 NOR2X1_103 ( .A(DATAI_13_), .B(_abc_40344_n705_1), .Y(_abc_40344_n1250) );
  NOR2X1 NOR2X1_104 ( .A(_abc_40344_n1254_1), .B(_abc_40344_n1258), .Y(_abc_40344_n1259) );
  NOR2X1 NOR2X1_105 ( .A(DATAI_11_), .B(_abc_40344_n705_1), .Y(_abc_40344_n1272) );
  NOR2X1 NOR2X1_106 ( .A(_abc_40344_n1277), .B(_abc_40344_n1276), .Y(_abc_40344_n1278) );
  NOR2X1 NOR2X1_107 ( .A(_abc_40344_n1283), .B(_abc_40344_n1280), .Y(_abc_40344_n1284) );
  NOR2X1 NOR2X1_108 ( .A(_abc_40344_n1298), .B(_abc_40344_n1304_1), .Y(_abc_40344_n1305) );
  NOR2X1 NOR2X1_109 ( .A(DATAI_12_), .B(_abc_40344_n705_1), .Y(_abc_40344_n1307) );
  NOR2X1 NOR2X1_11 ( .A(_abc_40344_n547), .B(_abc_40344_n544), .Y(_abc_40344_n548) );
  NOR2X1 NOR2X1_110 ( .A(_abc_40344_n1336), .B(_abc_40344_n1338), .Y(_abc_40344_n1339) );
  NOR2X1 NOR2X1_111 ( .A(_abc_40344_n1353), .B(_abc_40344_n1360), .Y(_abc_40344_n1361) );
  NOR2X1 NOR2X1_112 ( .A(_abc_40344_n1364), .B(_abc_40344_n1366), .Y(_abc_40344_n1367) );
  NOR2X1 NOR2X1_113 ( .A(_abc_40344_n1376), .B(_abc_40344_n1378), .Y(_abc_40344_n1379) );
  NOR2X1 NOR2X1_114 ( .A(_abc_40344_n1381), .B(_abc_40344_n1382), .Y(_abc_40344_n1383_1) );
  NOR2X1 NOR2X1_115 ( .A(_abc_40344_n1379), .B(_abc_40344_n1387), .Y(_abc_40344_n1388) );
  NOR2X1 NOR2X1_116 ( .A(_abc_40344_n1188), .B(_abc_40344_n1190), .Y(_abc_40344_n1397) );
  NOR2X1 NOR2X1_117 ( .A(_abc_40344_n1169), .B(_abc_40344_n1171), .Y(_abc_40344_n1398) );
  NOR2X1 NOR2X1_118 ( .A(_abc_40344_n1413), .B(_abc_40344_n1410), .Y(_abc_40344_n1414) );
  NOR2X1 NOR2X1_119 ( .A(_abc_40344_n921), .B(_abc_40344_n1423), .Y(_abc_40344_n1424) );
  NOR2X1 NOR2X1_12 ( .A(IR_REG_23_), .B(IR_REG_22_), .Y(_abc_40344_n549_1) );
  NOR2X1 NOR2X1_120 ( .A(_abc_40344_n1428), .B(_abc_40344_n1424), .Y(_abc_40344_n1429) );
  NOR2X1 NOR2X1_121 ( .A(_abc_40344_n1416), .B(_abc_40344_n1450), .Y(_abc_40344_n1451_1) );
  NOR2X1 NOR2X1_122 ( .A(_abc_40344_n1473), .B(_abc_40344_n1475), .Y(_abc_40344_n1476) );
  NOR2X1 NOR2X1_123 ( .A(_abc_40344_n1043), .B(_abc_40344_n1063), .Y(_abc_40344_n1479) );
  NOR2X1 NOR2X1_124 ( .A(_abc_40344_n1486), .B(_abc_40344_n1483), .Y(_abc_40344_n1487) );
  NOR2X1 NOR2X1_125 ( .A(_abc_40344_n1503_1), .B(_abc_40344_n1500), .Y(_abc_40344_n1504) );
  NOR2X1 NOR2X1_126 ( .A(_abc_40344_n1505_1), .B(_abc_40344_n1498), .Y(_abc_40344_n1506) );
  NOR2X1 NOR2X1_127 ( .A(_abc_40344_n1476), .B(_abc_40344_n1512), .Y(_abc_40344_n1513) );
  NOR2X1 NOR2X1_128 ( .A(_abc_40344_n1508_1), .B(_abc_40344_n1510), .Y(_abc_40344_n1516_1) );
  NOR2X1 NOR2X1_129 ( .A(_abc_40344_n1518), .B(_abc_40344_n1516_1), .Y(_abc_40344_n1519) );
  NOR2X1 NOR2X1_13 ( .A(IR_REG_25_), .B(IR_REG_24_), .Y(_abc_40344_n551) );
  NOR2X1 NOR2X1_130 ( .A(_abc_40344_n1082), .B(_abc_40344_n1522), .Y(_abc_40344_n1523) );
  NOR2X1 NOR2X1_131 ( .A(_abc_40344_n1538), .B(_abc_40344_n1067), .Y(_abc_40344_n1540) );
  NOR2X1 NOR2X1_132 ( .A(_abc_40344_n1540), .B(_abc_40344_n1539), .Y(_abc_40344_n1541) );
  NOR2X1 NOR2X1_133 ( .A(_abc_40344_n1547), .B(_abc_40344_n1544), .Y(_abc_40344_n1548) );
  NOR2X1 NOR2X1_134 ( .A(_abc_40344_n1549), .B(_abc_40344_n1542), .Y(_abc_40344_n1550) );
  NOR2X1 NOR2X1_135 ( .A(_abc_40344_n1561), .B(_abc_40344_n1560), .Y(_abc_40344_n1562) );
  NOR2X1 NOR2X1_136 ( .A(_abc_40344_n1458), .B(_abc_40344_n1449), .Y(_abc_40344_n1571) );
  NOR2X1 NOR2X1_137 ( .A(_abc_40344_n1110), .B(_abc_40344_n1023_1), .Y(_abc_40344_n1576) );
  NOR2X1 NOR2X1_138 ( .A(_abc_40344_n1577), .B(_abc_40344_n1537), .Y(_abc_40344_n1578) );
  NOR2X1 NOR2X1_139 ( .A(_abc_40344_n1401), .B(_abc_40344_n1396_1), .Y(_abc_40344_n1616) );
  NOR2X1 NOR2X1_14 ( .A(_abc_40344_n571_1), .B(_abc_40344_n573_1), .Y(_abc_40344_n574) );
  NOR2X1 NOR2X1_140 ( .A(_abc_40344_n1080), .B(_abc_40344_n1534), .Y(_abc_40344_n1628) );
  NOR2X1 NOR2X1_141 ( .A(_abc_40344_n1081), .B(_abc_40344_n1634), .Y(_abc_40344_n1635) );
  NOR2X1 NOR2X1_142 ( .A(_abc_40344_n1387), .B(_abc_40344_n1656), .Y(_abc_40344_n1657) );
  NOR2X1 NOR2X1_143 ( .A(_abc_40344_n1385), .B(_abc_40344_n1657), .Y(_abc_40344_n1658) );
  NOR2X1 NOR2X1_144 ( .A(_abc_40344_n1655), .B(_abc_40344_n1658), .Y(_abc_40344_n1659) );
  NOR2X1 NOR2X1_145 ( .A(_abc_40344_n886), .B(_abc_40344_n883), .Y(_abc_40344_n1675) );
  NOR2X1 NOR2X1_146 ( .A(_abc_40344_n1689), .B(_abc_40344_n1685), .Y(_abc_40344_n1690) );
  NOR2X1 NOR2X1_147 ( .A(_abc_40344_n1490), .B(_abc_40344_n1493), .Y(_abc_40344_n1715) );
  NOR2X1 NOR2X1_148 ( .A(_abc_40344_n1715), .B(_abc_40344_n1518), .Y(_abc_40344_n1716) );
  NOR2X1 NOR2X1_149 ( .A(_abc_40344_n1716), .B(_abc_40344_n1717), .Y(_abc_40344_n1718) );
  NOR2X1 NOR2X1_15 ( .A(_abc_40344_n566), .B(_abc_40344_n577_1), .Y(_abc_40344_n578_1) );
  NOR2X1 NOR2X1_150 ( .A(_abc_40344_n1577), .B(_abc_40344_n1023_1), .Y(_abc_40344_n1723) );
  NOR2X1 NOR2X1_151 ( .A(_abc_40344_n1537), .B(_abc_40344_n1506), .Y(_abc_40344_n1724) );
  NOR2X1 NOR2X1_152 ( .A(_abc_40344_n1398), .B(_abc_40344_n1732), .Y(_abc_40344_n1733) );
  NOR2X1 NOR2X1_153 ( .A(_abc_40344_n1750), .B(_abc_40344_n1751), .Y(_abc_40344_n1752) );
  NOR2X1 NOR2X1_154 ( .A(_abc_40344_n1476), .B(_abc_40344_n1719), .Y(_abc_40344_n1763) );
  NOR2X1 NOR2X1_155 ( .A(_abc_40344_n1783), .B(_abc_40344_n1782), .Y(_abc_40344_n1784) );
  NOR2X1 NOR2X1_156 ( .A(_abc_40344_n1331_1), .B(_abc_40344_n1334), .Y(_abc_40344_n1787) );
  NOR2X1 NOR2X1_157 ( .A(_abc_40344_n863), .B(_abc_40344_n1006), .Y(_abc_40344_n1801) );
  NOR2X1 NOR2X1_158 ( .A(_abc_40344_n1430), .B(_abc_40344_n1432), .Y(_abc_40344_n1807) );
  NOR2X1 NOR2X1_159 ( .A(_abc_40344_n1807), .B(_abc_40344_n1689), .Y(_abc_40344_n1808) );
  NOR2X1 NOR2X1_16 ( .A(_abc_40344_n561_1), .B(_abc_40344_n580), .Y(_abc_40344_n581) );
  NOR2X1 NOR2X1_160 ( .A(_abc_40344_n1306), .B(_abc_40344_n1311), .Y(_abc_40344_n1824) );
  NOR2X1 NOR2X1_161 ( .A(_abc_40344_n1846), .B(_abc_40344_n1704), .Y(_abc_40344_n1847) );
  NOR2X1 NOR2X1_162 ( .A(_abc_40344_n726), .B(_abc_40344_n938), .Y(_abc_40344_n1869) );
  NOR2X1 NOR2X1_163 ( .A(_abc_40344_n1516_1), .B(_abc_40344_n1512), .Y(_abc_40344_n1883) );
  NOR2X1 NOR2X1_164 ( .A(_abc_40344_n1019), .B(_abc_40344_n1375), .Y(_abc_40344_n1908) );
  NOR2X1 NOR2X1_165 ( .A(_abc_40344_n1910), .B(_abc_40344_n1913), .Y(_abc_40344_n1914) );
  NOR2X1 NOR2X1_166 ( .A(_abc_40344_n1916), .B(_abc_40344_n1915), .Y(_abc_40344_n1917) );
  NOR2X1 NOR2X1_167 ( .A(_abc_40344_n1924), .B(_abc_40344_n1917), .Y(_abc_40344_n1925) );
  NOR2X1 NOR2X1_168 ( .A(_abc_40344_n1084), .B(_abc_40344_n1090_1), .Y(_abc_40344_n1935) );
  NOR2X1 NOR2X1_169 ( .A(_abc_40344_n1137), .B(_abc_40344_n1134), .Y(_abc_40344_n1948) );
  NOR2X1 NOR2X1_17 ( .A(_abc_40344_n523), .B(_abc_40344_n587), .Y(_abc_40344_n588) );
  NOR2X1 NOR2X1_170 ( .A(_abc_40344_n1434), .B(_abc_40344_n1440), .Y(_abc_40344_n1952) );
  NOR2X1 NOR2X1_171 ( .A(_abc_40344_n1954), .B(_abc_40344_n1952), .Y(_abc_40344_n1955) );
  NOR2X1 NOR2X1_172 ( .A(_abc_40344_n1951), .B(_abc_40344_n1959), .Y(_abc_40344_n1960) );
  NOR2X1 NOR2X1_173 ( .A(_abc_40344_n1309), .B(_abc_40344_n1295), .Y(_abc_40344_n1971) );
  NOR2X1 NOR2X1_174 ( .A(_abc_40344_n785), .B(_abc_40344_n776), .Y(_abc_40344_n1980) );
  NOR2X1 NOR2X1_175 ( .A(_abc_40344_n1996), .B(_abc_40344_n1986), .Y(_abc_40344_n1997) );
  NOR2X1 NOR2X1_176 ( .A(_abc_40344_n763), .B(_abc_40344_n734), .Y(_abc_40344_n1998) );
  NOR2X1 NOR2X1_177 ( .A(_abc_40344_n2000), .B(_abc_40344_n1982), .Y(_abc_40344_n2008) );
  NOR2X1 NOR2X1_178 ( .A(_abc_40344_n2004), .B(_abc_40344_n2011), .Y(_abc_40344_n2012) );
  NOR2X1 NOR2X1_179 ( .A(_abc_40344_n829_1), .B(_abc_40344_n2022), .Y(_abc_40344_n2023) );
  NOR2X1 NOR2X1_18 ( .A(RESET_G), .B(_abc_40344_n589), .Y(n1345) );
  NOR2X1 NOR2X1_180 ( .A(_abc_40344_n2024), .B(_abc_40344_n2019), .Y(_abc_40344_n2025) );
  NOR2X1 NOR2X1_181 ( .A(_abc_40344_n1433), .B(_abc_40344_n1441), .Y(_abc_40344_n2029) );
  NOR2X1 NOR2X1_182 ( .A(_abc_40344_n2033), .B(_abc_40344_n2004), .Y(_abc_40344_n2034) );
  NOR2X1 NOR2X1_183 ( .A(_abc_40344_n1421_1), .B(_abc_40344_n2037), .Y(_abc_40344_n2038) );
  NOR2X1 NOR2X1_184 ( .A(_abc_40344_n2039), .B(_abc_40344_n2028), .Y(_abc_40344_n2040) );
  NOR2X1 NOR2X1_185 ( .A(_abc_40344_n1152_1), .B(_abc_40344_n1168), .Y(_abc_40344_n2042) );
  NOR2X1 NOR2X1_186 ( .A(_abc_40344_n2044), .B(_abc_40344_n2028), .Y(_abc_40344_n2045) );
  NOR2X1 NOR2X1_187 ( .A(_abc_40344_n2046), .B(_abc_40344_n1937), .Y(_abc_40344_n2047) );
  NOR2X1 NOR2X1_188 ( .A(_abc_40344_n1234), .B(_abc_40344_n1961), .Y(_abc_40344_n2049) );
  NOR2X1 NOR2X1_189 ( .A(_abc_40344_n2050), .B(_abc_40344_n2028), .Y(_abc_40344_n2051) );
  NOR2X1 NOR2X1_19 ( .A(RESET_G), .B(STATE_REG), .Y(n1336) );
  NOR2X1 NOR2X1_190 ( .A(_abc_40344_n1200), .B(_abc_40344_n1210), .Y(_abc_40344_n2056) );
  NOR2X1 NOR2X1_191 ( .A(_abc_40344_n2057), .B(_abc_40344_n2028), .Y(_abc_40344_n2058) );
  NOR2X1 NOR2X1_192 ( .A(_abc_40344_n698), .B(_abc_40344_n1994), .Y(_abc_40344_n2059) );
  NOR2X1 NOR2X1_193 ( .A(_abc_40344_n2011), .B(_abc_40344_n2066), .Y(_abc_40344_n2067) );
  NOR2X1 NOR2X1_194 ( .A(_abc_40344_n1260), .B(_abc_40344_n1264), .Y(_abc_40344_n2068) );
  NOR2X1 NOR2X1_195 ( .A(_abc_40344_n1186), .B(_abc_40344_n1949), .Y(_abc_40344_n2076) );
  NOR2X1 NOR2X1_196 ( .A(_abc_40344_n742), .B(_abc_40344_n750), .Y(_abc_40344_n2082) );
  NOR2X1 NOR2X1_197 ( .A(_abc_40344_n2083), .B(_abc_40344_n1966), .Y(_abc_40344_n2084) );
  NOR2X1 NOR2X1_198 ( .A(_abc_40344_n787_1), .B(_abc_40344_n777_1), .Y(_abc_40344_n2088) );
  NOR2X1 NOR2X1_199 ( .A(_abc_40344_n2090), .B(_abc_40344_n2028), .Y(_abc_40344_n2091) );
  NOR2X1 NOR2X1_2 ( .A(IR_REG_15_), .B(IR_REG_14_), .Y(_abc_40344_n525) );
  NOR2X1 NOR2X1_20 ( .A(IR_REG_26_), .B(IR_REG_27_), .Y(_abc_40344_n594) );
  NOR2X1 NOR2X1_200 ( .A(_abc_40344_n2093), .B(_abc_40344_n2072), .Y(_abc_40344_n2094) );
  NOR2X1 NOR2X1_201 ( .A(_abc_40344_n1918), .B(_abc_40344_n1921), .Y(_abc_40344_n2095) );
  NOR2X1 NOR2X1_202 ( .A(_abc_40344_n1922), .B(_abc_40344_n2096), .Y(_abc_40344_n2097) );
  NOR2X1 NOR2X1_203 ( .A(_abc_40344_n1926), .B(_abc_40344_n1645), .Y(_abc_40344_n2098) );
  NOR2X1 NOR2X1_204 ( .A(_abc_40344_n2106), .B(_abc_40344_n1073), .Y(_abc_40344_n2107) );
  NOR2X1 NOR2X1_205 ( .A(_abc_40344_n2028), .B(_abc_40344_n2011), .Y(_abc_40344_n2115) );
  NOR2X1 NOR2X1_206 ( .A(_abc_40344_n1477), .B(_abc_40344_n1488), .Y(_abc_40344_n2118) );
  NOR2X1 NOR2X1_207 ( .A(_abc_40344_n1285), .B(_abc_40344_n1973), .Y(_abc_40344_n2121) );
  NOR2X1 NOR2X1_208 ( .A(_abc_40344_n1335), .B(_abc_40344_n1969), .Y(_abc_40344_n2125) );
  NOR2X1 NOR2X1_209 ( .A(_abc_40344_n2126), .B(_abc_40344_n1966), .Y(_abc_40344_n2127) );
  NOR2X1 NOR2X1_21 ( .A(IR_REG_26_), .B(IR_REG_25_), .Y(_abc_40344_n607) );
  NOR2X1 NOR2X1_210 ( .A(_abc_40344_n915_1), .B(_abc_40344_n919), .Y(_abc_40344_n2130) );
  NOR2X1 NOR2X1_211 ( .A(_abc_40344_n2131), .B(_abc_40344_n2028), .Y(_abc_40344_n2132) );
  NOR2X1 NOR2X1_212 ( .A(_abc_40344_n2135), .B(_abc_40344_n2019), .Y(_abc_40344_n2136) );
  NOR2X1 NOR2X1_213 ( .A(_abc_40344_n2011), .B(_abc_40344_n2139), .Y(_abc_40344_n2140) );
  NOR2X1 NOR2X1_214 ( .A(_abc_40344_n1362), .B(_abc_40344_n1906), .Y(_abc_40344_n2151) );
  NOR2X1 NOR2X1_215 ( .A(_abc_40344_n2011), .B(_abc_40344_n2152), .Y(_abc_40344_n2153) );
  NOR2X1 NOR2X1_216 ( .A(_abc_40344_n2155), .B(_abc_40344_n2129), .Y(_abc_40344_n2156) );
  NOR2X1 NOR2X1_217 ( .A(_abc_40344_n2172), .B(_abc_40344_n785), .Y(_abc_40344_n2207) );
  NOR2X1 NOR2X1_218 ( .A(_abc_40344_n2252), .B(_abc_40344_n2251), .Y(_abc_40344_n2253_1) );
  NOR2X1 NOR2X1_219 ( .A(_abc_40344_n2172), .B(_abc_40344_n1335), .Y(_abc_40344_n2266) );
  NOR2X1 NOR2X1_22 ( .A(_abc_40344_n614), .B(_abc_40344_n544), .Y(_abc_40344_n615) );
  NOR2X1 NOR2X1_220 ( .A(_abc_40344_n2283), .B(_abc_40344_n2281), .Y(_abc_40344_n2288_1) );
  NOR2X1 NOR2X1_221 ( .A(_abc_40344_n2161), .B(_abc_40344_n1200), .Y(_abc_40344_n2300) );
  NOR2X1 NOR2X1_222 ( .A(_abc_40344_n2300), .B(_abc_40344_n2301), .Y(_abc_40344_n2302) );
  NOR2X1 NOR2X1_223 ( .A(_abc_40344_n2161), .B(_abc_40344_n1152_1), .Y(_abc_40344_n2309) );
  NOR2X1 NOR2X1_224 ( .A(_abc_40344_n2309), .B(_abc_40344_n2310), .Y(_abc_40344_n2311) );
  NOR2X1 NOR2X1_225 ( .A(_abc_40344_n2161), .B(_abc_40344_n1949), .Y(_abc_40344_n2316) );
  NOR2X1 NOR2X1_226 ( .A(_abc_40344_n2316), .B(_abc_40344_n2317), .Y(_abc_40344_n2318) );
  NOR2X1 NOR2X1_227 ( .A(_abc_40344_n2161), .B(_abc_40344_n1137), .Y(_abc_40344_n2323) );
  NOR2X1 NOR2X1_228 ( .A(_abc_40344_n2323), .B(_abc_40344_n2324), .Y(_abc_40344_n2325) );
  NOR2X1 NOR2X1_229 ( .A(_abc_40344_n2161), .B(_abc_40344_n1418), .Y(_abc_40344_n2328) );
  NOR2X1 NOR2X1_23 ( .A(_abc_40344_n626), .B(_abc_40344_n619), .Y(_abc_40344_n627) );
  NOR2X1 NOR2X1_230 ( .A(_abc_40344_n2328), .B(_abc_40344_n2329), .Y(_abc_40344_n2330) );
  NOR2X1 NOR2X1_231 ( .A(_abc_40344_n2179), .B(_abc_40344_n1090_1), .Y(_abc_40344_n2356) );
  NOR2X1 NOR2X1_232 ( .A(_abc_40344_n2357), .B(_abc_40344_n2356), .Y(_abc_40344_n2358) );
  NOR2X1 NOR2X1_233 ( .A(_abc_40344_n2101), .B(_abc_40344_n1917), .Y(_abc_40344_n2408_1) );
  NOR2X1 NOR2X1_234 ( .A(_abc_40344_n585), .B(_abc_40344_n2162), .Y(_abc_40344_n2409) );
  NOR2X1 NOR2X1_235 ( .A(_abc_40344_n2248), .B(_abc_40344_n2440), .Y(_abc_40344_n2441) );
  NOR2X1 NOR2X1_236 ( .A(_abc_40344_n2289), .B(_abc_40344_n2298), .Y(_abc_40344_n2450) );
  NOR2X1 NOR2X1_237 ( .A(_abc_40344_n1952), .B(_abc_40344_n2029), .Y(_abc_40344_n2470) );
  NOR2X1 NOR2X1_238 ( .A(_abc_40344_n2471), .B(_abc_40344_n2065), .Y(_abc_40344_n2472) );
  NOR2X1 NOR2X1_239 ( .A(_abc_40344_n2097), .B(_abc_40344_n2473), .Y(_abc_40344_n2474) );
  NOR2X1 NOR2X1_24 ( .A(_abc_40344_n523), .B(_abc_40344_n630_1), .Y(_abc_40344_n631) );
  NOR2X1 NOR2X1_240 ( .A(_abc_40344_n698), .B(_abc_40344_n714), .Y(_abc_40344_n2475) );
  NOR2X1 NOR2X1_241 ( .A(_abc_40344_n1021), .B(_abc_40344_n1994), .Y(_abc_40344_n2476) );
  NOR2X1 NOR2X1_242 ( .A(_abc_40344_n2475), .B(_abc_40344_n2476), .Y(_abc_40344_n2477) );
  NOR2X1 NOR2X1_243 ( .A(_abc_40344_n2477), .B(_abc_40344_n2480), .Y(_abc_40344_n2481) );
  NOR2X1 NOR2X1_244 ( .A(_abc_40344_n1998), .B(_abc_40344_n2082), .Y(_abc_40344_n2482) );
  NOR2X1 NOR2X1_245 ( .A(_abc_40344_n2483), .B(_abc_40344_n2484_1), .Y(_abc_40344_n2485) );
  NOR2X1 NOR2X1_246 ( .A(_abc_40344_n2488), .B(_abc_40344_n2487), .Y(_abc_40344_n2489) );
  NOR2X1 NOR2X1_247 ( .A(_abc_40344_n1335), .B(_abc_40344_n1327), .Y(_abc_40344_n2492) );
  NOR2X1 NOR2X1_248 ( .A(_abc_40344_n1787), .B(_abc_40344_n1969), .Y(_abc_40344_n2493) );
  NOR2X1 NOR2X1_249 ( .A(_abc_40344_n2492), .B(_abc_40344_n2493), .Y(_abc_40344_n2494) );
  NOR2X1 NOR2X1_25 ( .A(IR_REG_31_), .B(IR_REG_30_), .Y(_abc_40344_n651_1) );
  NOR2X1 NOR2X1_250 ( .A(_abc_40344_n2491), .B(_abc_40344_n2494), .Y(_abc_40344_n2495) );
  NOR2X1 NOR2X1_251 ( .A(_abc_40344_n1309), .B(_abc_40344_n1308), .Y(_abc_40344_n2500) );
  NOR2X1 NOR2X1_252 ( .A(_abc_40344_n1305), .B(_abc_40344_n1295), .Y(_abc_40344_n2501) );
  NOR2X1 NOR2X1_253 ( .A(_abc_40344_n2504), .B(_abc_40344_n2503), .Y(_abc_40344_n2505) );
  NOR2X1 NOR2X1_254 ( .A(_abc_40344_n2497), .B(_abc_40344_n2507), .Y(_abc_40344_n2508) );
  NOR2X1 NOR2X1_255 ( .A(_abc_40344_n2469), .B(_abc_40344_n2509), .Y(_abc_40344_n2510) );
  NOR2X1 NOR2X1_256 ( .A(_abc_40344_n2118), .B(_abc_40344_n2513), .Y(_abc_40344_n2514) );
  NOR2X1 NOR2X1_257 ( .A(_abc_40344_n1124), .B(_abc_40344_n1138), .Y(_abc_40344_n2525) );
  NOR2X1 NOR2X1_258 ( .A(_abc_40344_n2525), .B(_abc_40344_n1948), .Y(_abc_40344_n2526) );
  NOR2X1 NOR2X1_259 ( .A(_abc_40344_n2529_1), .B(_abc_40344_n2532), .Y(_abc_40344_n2533) );
  NOR2X1 NOR2X1_26 ( .A(_abc_40344_n654), .B(_abc_40344_n653), .Y(_abc_40344_n655) );
  NOR2X1 NOR2X1_260 ( .A(_abc_40344_n1362), .B(_abc_40344_n1350), .Y(_abc_40344_n2534) );
  NOR2X1 NOR2X1_261 ( .A(_abc_40344_n1361), .B(_abc_40344_n1906), .Y(_abc_40344_n2535) );
  NOR2X1 NOR2X1_262 ( .A(_abc_40344_n2534), .B(_abc_40344_n2535), .Y(_abc_40344_n2536) );
  NOR2X1 NOR2X1_263 ( .A(_abc_40344_n2536), .B(_abc_40344_n2538), .Y(_abc_40344_n2539) );
  NOR2X1 NOR2X1_264 ( .A(_abc_40344_n1178), .B(_abc_40344_n1186), .Y(_abc_40344_n2540) );
  NOR2X1 NOR2X1_265 ( .A(_abc_40344_n2540), .B(_abc_40344_n2542), .Y(_abc_40344_n2543_1) );
  NOR2X1 NOR2X1_266 ( .A(_abc_40344_n2543_1), .B(_abc_40344_n2547), .Y(_abc_40344_n2548) );
  NOR2X1 NOR2X1_267 ( .A(_abc_40344_n2527), .B(_abc_40344_n2549_1), .Y(_abc_40344_n2550) );
  NOR2X1 NOR2X1_268 ( .A(_abc_40344_n2551), .B(_abc_40344_n2521), .Y(_abc_40344_n2552) );
  NOR2X1 NOR2X1_269 ( .A(_abc_40344_n2512), .B(_abc_40344_n2553), .Y(_abc_40344_n2554) );
  NOR2X1 NOR2X1_27 ( .A(IR_REG_28_), .B(IR_REG_29_), .Y(_abc_40344_n657) );
  NOR2X1 NOR2X1_270 ( .A(_abc_40344_n2558), .B(_abc_40344_n2556), .Y(_abc_40344_n2559) );
  NOR2X1 NOR2X1_271 ( .A(_abc_40344_n618), .B(_abc_40344_n2560), .Y(_abc_40344_n2561) );
  NOR2X1 NOR2X1_272 ( .A(_abc_40344_n640), .B(_abc_40344_n2561), .Y(_abc_40344_n2562) );
  NOR2X1 NOR2X1_273 ( .A(_abc_40344_n2570), .B(_abc_40344_n2098), .Y(_abc_40344_n2574) );
  NOR2X1 NOR2X1_274 ( .A(_abc_40344_n2118), .B(_abc_40344_n2582), .Y(_abc_40344_n2583) );
  NOR2X1 NOR2X1_275 ( .A(_abc_40344_n2590), .B(_abc_40344_n2074), .Y(_abc_40344_n2591) );
  NOR2X1 NOR2X1_276 ( .A(_abc_40344_n2078), .B(_abc_40344_n2592), .Y(_abc_40344_n2593_1) );
  NOR2X1 NOR2X1_277 ( .A(_abc_40344_n2056), .B(_abc_40344_n2042), .Y(_abc_40344_n2599_1) );
  NOR2X1 NOR2X1_278 ( .A(_abc_40344_n2601), .B(_abc_40344_n2600), .Y(_abc_40344_n2602) );
  NOR2X1 NOR2X1_279 ( .A(_abc_40344_n2059), .B(_abc_40344_n2611), .Y(_abc_40344_n2612) );
  NOR2X1 NOR2X1_28 ( .A(IR_REG_31_), .B(IR_REG_29_), .Y(_abc_40344_n667) );
  NOR2X1 NOR2X1_280 ( .A(_abc_40344_n2613), .B(_abc_40344_n2614), .Y(_abc_40344_n2615) );
  NOR2X1 NOR2X1_281 ( .A(_abc_40344_n2624), .B(_abc_40344_n2625_1), .Y(_abc_40344_n2626) );
  NOR2X1 NOR2X1_282 ( .A(_abc_40344_n2633), .B(_abc_40344_n2627), .Y(_abc_40344_n2634) );
  NOR2X1 NOR2X1_283 ( .A(_abc_40344_n2621), .B(_abc_40344_n2608), .Y(_abc_40344_n2646) );
  NOR2X1 NOR2X1_284 ( .A(_abc_40344_n618), .B(_abc_40344_n640), .Y(_abc_40344_n2657) );
  NOR2X1 NOR2X1_285 ( .A(_abc_40344_n523), .B(_abc_40344_n586), .Y(_abc_40344_n2664) );
  NOR2X1 NOR2X1_286 ( .A(_abc_40344_n602), .B(_abc_40344_n610_1), .Y(_abc_40344_n2666_1) );
  NOR2X1 NOR2X1_287 ( .A(_abc_40344_n991), .B(_abc_40344_n2673), .Y(_abc_40344_n2677) );
  NOR2X1 NOR2X1_288 ( .A(_abc_40344_n2665), .B(_abc_40344_n2673), .Y(_abc_40344_n2684) );
  NOR2X1 NOR2X1_289 ( .A(_abc_40344_n2680), .B(_abc_40344_n853), .Y(_abc_40344_n2688) );
  NOR2X1 NOR2X1_29 ( .A(_abc_40344_n656), .B(_abc_40344_n660), .Y(_abc_40344_n669) );
  NOR2X1 NOR2X1_290 ( .A(_abc_40344_n538_1), .B(_abc_40344_n885), .Y(_abc_40344_n2694) );
  NOR2X1 NOR2X1_291 ( .A(REG1_REG_1_), .B(_abc_40344_n2694), .Y(_abc_40344_n2697) );
  NOR2X1 NOR2X1_292 ( .A(_abc_40344_n2697), .B(_abc_40344_n2696), .Y(_abc_40344_n2698_1) );
  NOR2X1 NOR2X1_293 ( .A(_abc_40344_n853), .B(_abc_40344_n2698_1), .Y(_abc_40344_n2699) );
  NOR2X1 NOR2X1_294 ( .A(_abc_40344_n602), .B(_abc_40344_n611_1), .Y(_abc_40344_n2708) );
  NOR2X1 NOR2X1_295 ( .A(_abc_40344_n2712), .B(_abc_40344_n2020), .Y(_abc_40344_n2713) );
  NOR2X1 NOR2X1_296 ( .A(REG2_REG_2_), .B(_abc_40344_n823), .Y(_abc_40344_n2714) );
  NOR2X1 NOR2X1_297 ( .A(_abc_40344_n2714), .B(_abc_40344_n2691), .Y(_abc_40344_n2716) );
  NOR2X1 NOR2X1_298 ( .A(_abc_40344_n2718), .B(_abc_40344_n2667), .Y(_abc_40344_n2719) );
  NOR2X1 NOR2X1_299 ( .A(REG2_REG_3_), .B(_abc_40344_n797), .Y(_abc_40344_n2728) );
  NOR2X1 NOR2X1_3 ( .A(IR_REG_12_), .B(IR_REG_11_), .Y(_abc_40344_n532) );
  NOR2X1 NOR2X1_30 ( .A(_abc_40344_n678), .B(_abc_40344_n526), .Y(_abc_40344_n679) );
  NOR2X1 NOR2X1_300 ( .A(_abc_40344_n2713), .B(_abc_40344_n2716), .Y(_abc_40344_n2732) );
  NOR2X1 NOR2X1_301 ( .A(REG1_REG_3_), .B(_abc_40344_n2735), .Y(_abc_40344_n2737) );
  NOR2X1 NOR2X1_302 ( .A(_abc_40344_n797), .B(_abc_40344_n2739), .Y(_abc_40344_n2740) );
  NOR2X1 NOR2X1_303 ( .A(REG2_REG_6_), .B(_abc_40344_n712), .Y(_abc_40344_n2783) );
  NOR2X1 NOR2X1_304 ( .A(_abc_40344_n523), .B(_abc_40344_n2673), .Y(_abc_40344_n2792) );
  NOR2X1 NOR2X1_305 ( .A(_abc_40344_n920), .B(_abc_40344_n917), .Y(_abc_40344_n2802) );
  NOR2X1 NOR2X1_306 ( .A(_abc_40344_n2813), .B(_abc_40344_n2815), .Y(_abc_40344_n2816_1) );
  NOR2X1 NOR2X1_307 ( .A(REG2_REG_10_), .B(_abc_40344_n1325), .Y(_abc_40344_n2854) );
  NOR2X1 NOR2X1_308 ( .A(REG1_REG_11_), .B(_abc_40344_n2863), .Y(_abc_40344_n2865) );
  NOR2X1 NOR2X1_309 ( .A(_abc_40344_n1274), .B(_abc_40344_n1271), .Y(_abc_40344_n2872) );
  NOR2X1 NOR2X1_31 ( .A(_abc_40344_n547), .B(_abc_40344_n595_1), .Y(_abc_40344_n680) );
  NOR2X1 NOR2X1_310 ( .A(REG2_REG_11_), .B(_abc_40344_n2863), .Y(_abc_40344_n2873) );
  NOR2X1 NOR2X1_311 ( .A(_abc_40344_n2872), .B(_abc_40344_n2873), .Y(_abc_40344_n2874) );
  NOR2X1 NOR2X1_312 ( .A(REG2_REG_12_), .B(_abc_40344_n2883), .Y(_abc_40344_n2890) );
  NOR2X1 NOR2X1_313 ( .A(_abc_40344_n603), .B(_abc_40344_n1293_1), .Y(_abc_40344_n2897) );
  NOR2X1 NOR2X1_314 ( .A(_abc_40344_n1255), .B(_abc_40344_n1249), .Y(_abc_40344_n2910) );
  NOR2X1 NOR2X1_315 ( .A(REG2_REG_13_), .B(_abc_40344_n2911), .Y(_abc_40344_n2912) );
  NOR2X1 NOR2X1_316 ( .A(_abc_40344_n2910), .B(_abc_40344_n2912), .Y(_abc_40344_n2913) );
  NOR2X1 NOR2X1_317 ( .A(_abc_40344_n1249), .B(_abc_40344_n603), .Y(_abc_40344_n2918) );
  NOR2X1 NOR2X1_318 ( .A(_abc_40344_n1231), .B(_abc_40344_n1222), .Y(_abc_40344_n2934) );
  NOR2X1 NOR2X1_319 ( .A(REG2_REG_14_), .B(_abc_40344_n1221), .Y(_abc_40344_n2936) );
  NOR2X1 NOR2X1_32 ( .A(_abc_40344_n687), .B(_abc_40344_n688_1), .Y(_abc_40344_n689) );
  NOR2X1 NOR2X1_320 ( .A(_abc_40344_n2946), .B(_abc_40344_n2944), .Y(_abc_40344_n2947) );
  NOR2X1 NOR2X1_321 ( .A(_abc_40344_n2950), .B(_abc_40344_n2952), .Y(_abc_40344_n2953) );
  NOR2X1 NOR2X1_322 ( .A(_abc_40344_n1207), .B(_abc_40344_n1196), .Y(_abc_40344_n2959) );
  NOR2X1 NOR2X1_323 ( .A(REG2_REG_15_), .B(_abc_40344_n1197), .Y(_abc_40344_n2961) );
  NOR2X1 NOR2X1_324 ( .A(_abc_40344_n1165), .B(_abc_40344_n1148), .Y(_abc_40344_n2970) );
  NOR2X1 NOR2X1_325 ( .A(REG1_REG_16_), .B(_abc_40344_n1149), .Y(_abc_40344_n2972) );
  NOR2X1 NOR2X1_326 ( .A(REG2_REG_16_), .B(_abc_40344_n1149), .Y(_abc_40344_n2979) );
  NOR2X1 NOR2X1_327 ( .A(_abc_40344_n2988), .B(_abc_40344_n2986), .Y(_abc_40344_n2989) );
  NOR2X1 NOR2X1_328 ( .A(_abc_40344_n1131), .B(_abc_40344_n1122), .Y(_abc_40344_n3016) );
  NOR2X1 NOR2X1_329 ( .A(REG2_REG_18_), .B(_abc_40344_n3017), .Y(_abc_40344_n3018) );
  NOR2X1 NOR2X1_33 ( .A(_abc_40344_n686), .B(_abc_40344_n690), .Y(_abc_40344_n691) );
  NOR2X1 NOR2X1_330 ( .A(_abc_40344_n3016), .B(_abc_40344_n3018), .Y(_abc_40344_n3019) );
  NOR2X1 NOR2X1_331 ( .A(_abc_40344_n1132_1), .B(_abc_40344_n1122), .Y(_abc_40344_n3026) );
  NOR2X1 NOR2X1_332 ( .A(REG1_REG_18_), .B(_abc_40344_n3017), .Y(_abc_40344_n3027) );
  NOR2X1 NOR2X1_333 ( .A(_abc_40344_n3026), .B(_abc_40344_n3027), .Y(_abc_40344_n3028) );
  NOR2X1 NOR2X1_334 ( .A(_abc_40344_n1197), .B(_abc_40344_n2950), .Y(_abc_40344_n3048) );
  NOR2X1 NOR2X1_335 ( .A(_abc_40344_n986), .B(_abc_40344_n1002), .Y(_abc_40344_n3061) );
  NOR2X1 NOR2X1_336 ( .A(_abc_40344_n951), .B(_abc_40344_n3063), .Y(_abc_40344_n3064) );
  NOR2X1 NOR2X1_337 ( .A(_abc_40344_n3062), .B(_abc_40344_n3067), .Y(_abc_40344_n3068) );
  NOR2X1 NOR2X1_338 ( .A(_abc_40344_n825), .B(_abc_40344_n3070), .Y(_abc_40344_n3071) );
  NOR2X1 NOR2X1_339 ( .A(_abc_40344_n777_1), .B(_abc_40344_n3072), .Y(_abc_40344_n3073) );
  NOR2X1 NOR2X1_34 ( .A(_abc_40344_n692), .B(_abc_40344_n691), .Y(_abc_40344_n693) );
  NOR2X1 NOR2X1_340 ( .A(_abc_40344_n714), .B(_abc_40344_n3074), .Y(_abc_40344_n3075) );
  NOR2X1 NOR2X1_341 ( .A(_abc_40344_n1665), .B(_abc_40344_n3076), .Y(_abc_40344_n3077) );
  NOR2X1 NOR2X1_342 ( .A(_abc_40344_n1327), .B(_abc_40344_n3078), .Y(_abc_40344_n3079) );
  NOR2X1 NOR2X1_343 ( .A(_abc_40344_n1273), .B(_abc_40344_n1308), .Y(_abc_40344_n3080) );
  NOR2X1 NOR2X1_344 ( .A(_abc_40344_n1251), .B(_abc_40344_n1224), .Y(_abc_40344_n3081_1) );
  NOR2X1 NOR2X1_345 ( .A(_abc_40344_n1124), .B(_abc_40344_n1178), .Y(_abc_40344_n3084) );
  NOR2X1 NOR2X1_346 ( .A(_abc_40344_n2394), .B(_abc_40344_n3097), .Y(_abc_40344_n3098) );
  NOR2X1 NOR2X1_347 ( .A(_abc_40344_n603), .B(_abc_40344_n984), .Y(_abc_40344_n3103) );
  NOR2X1 NOR2X1_348 ( .A(_abc_40344_n3109), .B(_abc_40344_n3067), .Y(_abc_40344_n3110) );
  NOR2X1 NOR2X1_349 ( .A(_abc_40344_n1040), .B(_abc_40344_n1074), .Y(_abc_40344_n3122) );
  NOR2X1 NOR2X1_35 ( .A(_abc_40344_n677), .B(_abc_40344_n681), .Y(_abc_40344_n702) );
  NOR2X1 NOR2X1_350 ( .A(_abc_40344_n2493), .B(_abc_40344_n2535), .Y(_abc_40344_n3130) );
  NOR2X1 NOR2X1_351 ( .A(_abc_40344_n1675), .B(_abc_40344_n1797), .Y(_abc_40344_n3136) );
  NOR2X1 NOR2X1_352 ( .A(_abc_40344_n3140), .B(_abc_40344_n3142), .Y(_abc_40344_n3143) );
  NOR2X1 NOR2X1_353 ( .A(_abc_40344_n763), .B(_abc_40344_n750), .Y(_abc_40344_n3151) );
  NOR2X1 NOR2X1_354 ( .A(_abc_40344_n787_1), .B(_abc_40344_n776), .Y(_abc_40344_n3152) );
  NOR2X1 NOR2X1_355 ( .A(_abc_40344_n915_1), .B(_abc_40344_n908), .Y(_abc_40344_n3156) );
  NOR2X1 NOR2X1_356 ( .A(_abc_40344_n2475), .B(_abc_40344_n3156), .Y(_abc_40344_n3157) );
  NOR2X1 NOR2X1_357 ( .A(_abc_40344_n1210), .B(_abc_40344_n1201), .Y(_abc_40344_n3160) );
  NOR2X1 NOR2X1_358 ( .A(_abc_40344_n3160), .B(_abc_40344_n3174), .Y(_abc_40344_n3175) );
  NOR2X1 NOR2X1_359 ( .A(_abc_40344_n1812), .B(_abc_40344_n2037), .Y(_abc_40344_n3179) );
  NOR2X1 NOR2X1_36 ( .A(IR_REG_5_), .B(_abc_40344_n707_1), .Y(_abc_40344_n708) );
  NOR2X1 NOR2X1_360 ( .A(_abc_40344_n1124), .B(_abc_40344_n1134), .Y(_abc_40344_n3187) );
  NOR2X1 NOR2X1_361 ( .A(_abc_40344_n3187), .B(_abc_40344_n3181), .Y(_abc_40344_n3188) );
  NOR2X1 NOR2X1_362 ( .A(_abc_40344_n1153), .B(_abc_40344_n1168), .Y(_abc_40344_n3192) );
  NOR2X1 NOR2X1_363 ( .A(_abc_40344_n2540), .B(_abc_40344_n3192), .Y(_abc_40344_n3193) );
  NOR2X1 NOR2X1_364 ( .A(_abc_40344_n921), .B(_abc_40344_n1481), .Y(_abc_40344_n3203) );
  NOR2X1 NOR2X1_365 ( .A(_abc_40344_n646), .B(_abc_40344_n699), .Y(_abc_40344_n3216) );
  NOR2X1 NOR2X1_366 ( .A(_abc_40344_n3217), .B(_abc_40344_n3067), .Y(_abc_40344_n3218) );
  NOR2X1 NOR2X1_367 ( .A(_abc_40344_n602), .B(_abc_40344_n984), .Y(_abc_40344_n3220) );
  NOR2X1 NOR2X1_368 ( .A(_abc_40344_n3232), .B(_abc_40344_n3067), .Y(_abc_40344_n3233) );
  NOR2X1 NOR2X1_369 ( .A(_abc_40344_n1031), .B(_abc_40344_n1068), .Y(_abc_40344_n3253) );
  NOR2X1 NOR2X1_37 ( .A(_abc_40344_n640), .B(_abc_40344_n619), .Y(_abc_40344_n717) );
  NOR2X1 NOR2X1_370 ( .A(_abc_40344_n1084), .B(_abc_40344_n3091), .Y(_abc_40344_n3271) );
  NOR2X1 NOR2X1_371 ( .A(_abc_40344_n1031), .B(_abc_40344_n1888), .Y(_abc_40344_n3275) );
  NOR2X1 NOR2X1_372 ( .A(_abc_40344_n2479), .B(_abc_40344_n2604), .Y(_abc_40344_n3299) );
  NOR2X1 NOR2X1_373 ( .A(_abc_40344_n2076), .B(_abc_40344_n3301), .Y(_abc_40344_n3302) );
  NOR2X1 NOR2X1_374 ( .A(_abc_40344_n2589), .B(_abc_40344_n3302), .Y(_abc_40344_n3303) );
  NOR2X1 NOR2X1_375 ( .A(_abc_40344_n1996), .B(_abc_40344_n2612), .Y(_abc_40344_n3309) );
  NOR2X1 NOR2X1_376 ( .A(_abc_40344_n1907), .B(_abc_40344_n2125), .Y(_abc_40344_n3315) );
  NOR2X1 NOR2X1_377 ( .A(_abc_40344_n2125), .B(_abc_40344_n2121), .Y(_abc_40344_n3317) );
  NOR2X1 NOR2X1_378 ( .A(_abc_40344_n2076), .B(_abc_40344_n3322), .Y(_abc_40344_n3323) );
  NOR2X1 NOR2X1_379 ( .A(_abc_40344_n2590), .B(_abc_40344_n3326), .Y(_abc_40344_n3327) );
  NOR2X1 NOR2X1_38 ( .A(_abc_40344_n755), .B(_abc_40344_n762), .Y(_abc_40344_n763) );
  NOR2X1 NOR2X1_380 ( .A(_abc_40344_n1944), .B(_abc_40344_n1935), .Y(_abc_40344_n3333) );
  NOR2X1 NOR2X1_381 ( .A(_abc_40344_n2524), .B(_abc_40344_n3353), .Y(_abc_40344_n3354) );
  NOR2X1 NOR2X1_382 ( .A(_abc_40344_n2590), .B(_abc_40344_n2029), .Y(_abc_40344_n3356) );
  NOR2X1 NOR2X1_383 ( .A(_abc_40344_n3381), .B(_abc_40344_n3384), .Y(_abc_40344_n3385) );
  NOR2X1 NOR2X1_384 ( .A(_abc_40344_n3391), .B(_abc_40344_n3389), .Y(_abc_40344_n3392) );
  NOR2X1 NOR2X1_385 ( .A(_abc_40344_n3329), .B(_abc_40344_n3327), .Y(_abc_40344_n3399) );
  NOR2X1 NOR2X1_386 ( .A(_abc_40344_n3418), .B(_abc_40344_n3416), .Y(_abc_40344_n3419) );
  NOR2X1 NOR2X1_387 ( .A(_abc_40344_n3449), .B(_abc_40344_n3447), .Y(_abc_40344_n3450) );
  NOR2X1 NOR2X1_388 ( .A(_abc_40344_n3083), .B(_abc_40344_n3082), .Y(_abc_40344_n3465) );
  NOR2X1 NOR2X1_389 ( .A(_abc_40344_n1201), .B(_abc_40344_n3082), .Y(_abc_40344_n3508) );
  NOR2X1 NOR2X1_39 ( .A(REG3_REG_4_), .B(REG3_REG_3_), .Y(_abc_40344_n778) );
  NOR2X1 NOR2X1_390 ( .A(_abc_40344_n1152_1), .B(_abc_40344_n3508), .Y(_abc_40344_n3509) );
  NOR2X1 NOR2X1_391 ( .A(_abc_40344_n3465), .B(_abc_40344_n3509), .Y(_abc_40344_n3510) );
  NOR2X1 NOR2X1_392 ( .A(_abc_40344_n1308), .B(_abc_40344_n3526), .Y(_abc_40344_n3527) );
  NOR2X1 NOR2X1_393 ( .A(_abc_40344_n2500), .B(_abc_40344_n2501), .Y(_abc_40344_n3580) );
  NOR2X1 NOR2X1_394 ( .A(_abc_40344_n3588), .B(_abc_40344_n3586), .Y(_abc_40344_n3589) );
  NOR2X1 NOR2X1_395 ( .A(_abc_40344_n1305), .B(_abc_40344_n3232), .Y(_abc_40344_n3602) );
  NOR2X1 NOR2X1_396 ( .A(_abc_40344_n3662_1), .B(_abc_40344_n3667), .Y(_abc_40344_n3668) );
  NOR2X1 NOR2X1_397 ( .A(_abc_40344_n3703), .B(_abc_40344_n3138), .Y(_abc_40344_n3704) );
  NOR2X1 NOR2X1_398 ( .A(_abc_40344_n641), .B(_abc_40344_n986), .Y(_abc_40344_n3725) );
  NOR2X1 NOR2X1_399 ( .A(_abc_40344_n3228), .B(_abc_40344_n3730), .Y(_abc_40344_n3731) );
  NOR2X1 NOR2X1_4 ( .A(IR_REG_10_), .B(IR_REG_9_), .Y(_abc_40344_n533) );
  NOR2X1 NOR2X1_40 ( .A(_abc_40344_n778), .B(_abc_40344_n689), .Y(_abc_40344_n779) );
  NOR2X1 NOR2X1_400 ( .A(_abc_40344_n3750), .B(_abc_40344_n3747), .Y(_abc_40344_n3751) );
  NOR2X1 NOR2X1_401 ( .A(_abc_40344_n952), .B(_abc_40344_n991), .Y(_abc_40344_n3794_1) );
  NOR2X1 NOR2X1_402 ( .A(_abc_40344_n630_1), .B(_abc_40344_n3794_1), .Y(_abc_40344_n3795_1) );
  NOR2X1 NOR2X1_403 ( .A(_abc_40344_n559_1), .B(_abc_40344_n523), .Y(_abc_40344_n3856) );
  NOR2X1 NOR2X1_404 ( .A(IR_REG_31_), .B(_abc_40344_n523), .Y(_abc_40344_n3860) );
  NOR2X1 NOR2X1_405 ( .A(_abc_40344_n563_1), .B(_abc_40344_n556), .Y(_abc_40344_n3889) );
  NOR2X1 NOR2X1_406 ( .A(_abc_40344_n2558), .B(_abc_40344_n2652), .Y(_abc_40344_n4015) );
  NOR2X1 NOR2X1_407 ( .A(_abc_40344_n4039), .B(_abc_40344_n4038), .Y(_abc_40344_n4040_1) );
  NOR2X1 NOR2X1_408 ( .A(_abc_40344_n980), .B(_abc_40344_n4041), .Y(_abc_40344_n4042) );
  NOR2X1 NOR2X1_409 ( .A(_abc_40344_n625), .B(_abc_40344_n1027_1), .Y(_abc_40344_n4048) );
  NOR2X1 NOR2X1_41 ( .A(_abc_40344_n745), .B(_abc_40344_n809), .Y(_abc_40344_n810) );
  NOR2X1 NOR2X1_410 ( .A(_abc_40344_n3726), .B(_abc_40344_n3763), .Y(_abc_40344_n4056) );
  NOR2X1 NOR2X1_411 ( .A(_abc_40344_n4056), .B(_abc_40344_n3761), .Y(_abc_40344_n4057) );
  NOR2X1 NOR2X1_412 ( .A(_abc_40344_n3109), .B(_abc_40344_n1926), .Y(_abc_40344_n4220) );
  NOR2X1 NOR2X1_413 ( .A(_abc_40344_n979), .B(_abc_40344_n4041), .Y(_abc_40344_n4237) );
  NOR2X1 NOR2X1_42 ( .A(_abc_40344_n838), .B(_abc_40344_n840), .Y(_abc_40344_n841) );
  NOR2X1 NOR2X1_43 ( .A(_abc_40344_n841), .B(_abc_40344_n745), .Y(_abc_40344_n842) );
  NOR2X1 NOR2X1_44 ( .A(_abc_40344_n818_1), .B(_abc_40344_n844), .Y(_abc_40344_n846) );
  NOR2X1 NOR2X1_45 ( .A(_abc_40344_n859), .B(_abc_40344_n862), .Y(_abc_40344_n863) );
  NOR2X1 NOR2X1_46 ( .A(_abc_40344_n869), .B(_abc_40344_n747), .Y(_abc_40344_n870) );
  NOR2X1 NOR2X1_47 ( .A(_abc_40344_n863), .B(_abc_40344_n745), .Y(_abc_40344_n871) );
  NOR2X1 NOR2X1_48 ( .A(_abc_40344_n926), .B(_abc_40344_n923_1), .Y(_abc_40344_n927_1) );
  NOR2X1 NOR2X1_49 ( .A(_abc_40344_n938), .B(_abc_40344_n901), .Y(_abc_40344_n939) );
  NOR2X1 NOR2X1_5 ( .A(_abc_40344_n531), .B(_abc_40344_n534), .Y(_abc_40344_n535) );
  NOR2X1 NOR2X1_50 ( .A(_abc_40344_n633_1), .B(_abc_40344_n942), .Y(_abc_40344_n943_1) );
  NOR2X1 NOR2X1_51 ( .A(D_REG_2_), .B(D_REG_29_), .Y(_abc_40344_n953) );
  NOR2X1 NOR2X1_52 ( .A(D_REG_28_), .B(D_REG_27_), .Y(_abc_40344_n954) );
  NOR2X1 NOR2X1_53 ( .A(D_REG_26_), .B(D_REG_25_), .Y(_abc_40344_n956) );
  NOR2X1 NOR2X1_54 ( .A(D_REG_23_), .B(D_REG_22_), .Y(_abc_40344_n957) );
  NOR2X1 NOR2X1_55 ( .A(_abc_40344_n955_1), .B(_abc_40344_n958), .Y(_abc_40344_n959) );
  NOR2X1 NOR2X1_56 ( .A(D_REG_9_), .B(D_REG_8_), .Y(_abc_40344_n960) );
  NOR2X1 NOR2X1_57 ( .A(D_REG_31_), .B(D_REG_30_), .Y(_abc_40344_n961) );
  NOR2X1 NOR2X1_58 ( .A(D_REG_7_), .B(D_REG_4_), .Y(_abc_40344_n963) );
  NOR2X1 NOR2X1_59 ( .A(D_REG_24_), .B(D_REG_16_), .Y(_abc_40344_n965) );
  NOR2X1 NOR2X1_6 ( .A(IR_REG_6_), .B(IR_REG_5_), .Y(_abc_40344_n540) );
  NOR2X1 NOR2X1_60 ( .A(D_REG_21_), .B(D_REG_20_), .Y(_abc_40344_n966) );
  NOR2X1 NOR2X1_61 ( .A(D_REG_13_), .B(D_REG_18_), .Y(_abc_40344_n967) );
  NOR2X1 NOR2X1_62 ( .A(D_REG_14_), .B(D_REG_12_), .Y(_abc_40344_n969) );
  NOR2X1 NOR2X1_63 ( .A(D_REG_17_), .B(D_REG_10_), .Y(_abc_40344_n970_1) );
  NOR2X1 NOR2X1_64 ( .A(D_REG_11_), .B(D_REG_19_), .Y(_abc_40344_n972_1) );
  NOR2X1 NOR2X1_65 ( .A(D_REG_15_), .B(D_REG_5_), .Y(_abc_40344_n973) );
  NOR2X1 NOR2X1_66 ( .A(_abc_40344_n968), .B(_abc_40344_n974), .Y(_abc_40344_n975_1) );
  NOR2X1 NOR2X1_67 ( .A(D_REG_3_), .B(D_REG_6_), .Y(_abc_40344_n976) );
  NOR2X1 NOR2X1_68 ( .A(_abc_40344_n951), .B(_abc_40344_n981_1), .Y(_abc_40344_n982) );
  NOR2X1 NOR2X1_69 ( .A(_abc_40344_n625), .B(_abc_40344_n618), .Y(_abc_40344_n985) );
  NOR2X1 NOR2X1_7 ( .A(IR_REG_7_), .B(IR_REG_4_), .Y(_abc_40344_n541_1) );
  NOR2X1 NOR2X1_70 ( .A(_abc_40344_n641), .B(_abc_40344_n648), .Y(_abc_40344_n987) );
  NOR2X1 NOR2X1_71 ( .A(_abc_40344_n523), .B(_abc_40344_n989), .Y(_abc_40344_n990) );
  NOR2X1 NOR2X1_72 ( .A(_abc_40344_n992), .B(_abc_40344_n983), .Y(_abc_40344_n993) );
  NOR2X1 NOR2X1_73 ( .A(_abc_40344_n640), .B(_abc_40344_n986), .Y(_abc_40344_n995) );
  NOR2X1 NOR2X1_74 ( .A(_abc_40344_n984), .B(_abc_40344_n1002), .Y(_abc_40344_n1003) );
  NOR2X1 NOR2X1_75 ( .A(_abc_40344_n1004), .B(_abc_40344_n991), .Y(_abc_40344_n1005) );
  NOR2X1 NOR2X1_76 ( .A(_abc_40344_n1009), .B(_abc_40344_n1017), .Y(_abc_40344_n1018) );
  NOR2X1 NOR2X1_77 ( .A(_abc_40344_n603), .B(_abc_40344_n983), .Y(_abc_40344_n1020) );
  NOR2X1 NOR2X1_78 ( .A(_abc_40344_n602), .B(_abc_40344_n983), .Y(_abc_40344_n1022) );
  NOR2X1 NOR2X1_79 ( .A(_abc_40344_n646), .B(_abc_40344_n641), .Y(_abc_40344_n1026) );
  NOR2X1 NOR2X1_8 ( .A(_abc_40344_n539), .B(_abc_40344_n542_1), .Y(_abc_40344_n543) );
  NOR2X1 NOR2X1_80 ( .A(_abc_40344_n986), .B(_abc_40344_n1027_1), .Y(_abc_40344_n1028) );
  NOR2X1 NOR2X1_81 ( .A(_abc_40344_n1029_1), .B(_abc_40344_n991), .Y(_abc_40344_n1030_1) );
  NOR2X1 NOR2X1_82 ( .A(_abc_40344_n1052_1), .B(_abc_40344_n1053), .Y(_abc_40344_n1054) );
  NOR2X1 NOR2X1_83 ( .A(_abc_40344_n1049_1), .B(_abc_40344_n1055), .Y(_abc_40344_n1056) );
  NOR2X1 NOR2X1_84 ( .A(_abc_40344_n1047), .B(_abc_40344_n1058), .Y(_abc_40344_n1059) );
  NOR2X1 NOR2X1_85 ( .A(_abc_40344_n1045_1), .B(_abc_40344_n1061), .Y(_abc_40344_n1062) );
  NOR2X1 NOR2X1_86 ( .A(_abc_40344_n1075), .B(_abc_40344_n1078_1), .Y(_abc_40344_n1081) );
  NOR2X1 NOR2X1_87 ( .A(_abc_40344_n1081), .B(_abc_40344_n1080), .Y(_abc_40344_n1082) );
  NOR2X1 NOR2X1_88 ( .A(_abc_40344_n1092), .B(_abc_40344_n1095), .Y(_abc_40344_n1097) );
  NOR2X1 NOR2X1_89 ( .A(_abc_40344_n1046), .B(_abc_40344_n1060), .Y(_abc_40344_n1102) );
  NOR2X1 NOR2X1_9 ( .A(IR_REG_21_), .B(IR_REG_20_), .Y(_abc_40344_n545_1) );
  NOR2X1 NOR2X1_90 ( .A(_abc_40344_n921), .B(_abc_40344_n1104), .Y(_abc_40344_n1105) );
  NOR2X1 NOR2X1_91 ( .A(_abc_40344_n1109), .B(_abc_40344_n1105), .Y(_abc_40344_n1110) );
  NOR2X1 NOR2X1_92 ( .A(_abc_40344_n1113), .B(_abc_40344_n1115), .Y(_abc_40344_n1117) );
  NOR2X1 NOR2X1_93 ( .A(_abc_40344_n1133), .B(_abc_40344_n1130), .Y(_abc_40344_n1138) );
  NOR2X1 NOR2X1_94 ( .A(_abc_40344_n1136), .B(_abc_40344_n1140), .Y(_abc_40344_n1142) );
  NOR2X1 NOR2X1_95 ( .A(_abc_40344_n1155_1), .B(_abc_40344_n1057), .Y(_abc_40344_n1158) );
  NOR2X1 NOR2X1_96 ( .A(_abc_40344_n1166_1), .B(_abc_40344_n1163), .Y(_abc_40344_n1167) );
  NOR2X1 NOR2X1_97 ( .A(_abc_40344_n1184), .B(_abc_40344_n1181), .Y(_abc_40344_n1185) );
  NOR2X1 NOR2X1_98 ( .A(_abc_40344_n1208), .B(_abc_40344_n1205), .Y(_abc_40344_n1209_1) );
  NOR2X1 NOR2X1_99 ( .A(_abc_40344_n1211), .B(_abc_40344_n1214), .Y(_abc_40344_n1215) );
  NOR3X1 NOR3X1_1 ( .A(_abc_40344_n547), .B(_abc_40344_n555), .C(_abc_40344_n544), .Y(_abc_40344_n556) );
  NOR3X1 NOR3X1_10 ( .A(_abc_40344_n1043), .B(_abc_40344_n1044), .C(_abc_40344_n1063), .Y(_abc_40344_n1064) );
  NOR3X1 NOR3X1_11 ( .A(_abc_40344_n1937), .B(_abc_40344_n1977), .C(_abc_40344_n1966), .Y(_abc_40344_n1978) );
  NOR3X1 NOR3X1_12 ( .A(_abc_40344_n2000), .B(_abc_40344_n1982), .C(_abc_40344_n2004), .Y(_abc_40344_n2005) );
  NOR3X1 NOR3X1_13 ( .A(_abc_40344_n2053), .B(_abc_40344_n2036), .C(_abc_40344_n2007), .Y(_abc_40344_n2054) );
  NOR3X1 NOR3X1_14 ( .A(_abc_40344_n2061), .B(_abc_40344_n2028), .C(_abc_40344_n1982), .Y(_abc_40344_n2062) );
  NOR3X1 NOR3X1_15 ( .A(_abc_40344_n2028), .B(_abc_40344_n2069), .C(_abc_40344_n2011), .Y(_abc_40344_n2070) );
  NOR3X1 NOR3X1_16 ( .A(_abc_40344_n2085), .B(_abc_40344_n2004), .C(_abc_40344_n2011), .Y(_abc_40344_n2086) );
  NOR3X1 NOR3X1_17 ( .A(_abc_40344_n2028), .B(_abc_40344_n2112), .C(_abc_40344_n2011), .Y(_abc_40344_n2113) );
  NOR3X1 NOR3X1_18 ( .A(_abc_40344_n2028), .B(_abc_40344_n2122), .C(_abc_40344_n1966), .Y(_abc_40344_n2123) );
  NOR3X1 NOR3X1_19 ( .A(_abc_40344_n2149), .B(_abc_40344_n2028), .C(_abc_40344_n1982), .Y(_abc_40344_n2150) );
  NOR3X1 NOR3X1_2 ( .A(IR_REG_8_), .B(IR_REG_3_), .C(IR_REG_13_), .Y(_abc_40344_n570) );
  NOR3X1 NOR3X1_20 ( .A(_abc_40344_n2167), .B(_abc_40344_n2180), .C(_abc_40344_n2178), .Y(_abc_40344_n2181) );
  NOR3X1 NOR3X1_21 ( .A(_abc_40344_n2190), .B(_abc_40344_n2196), .C(_abc_40344_n2181), .Y(_abc_40344_n2197) );
  NOR3X1 NOR3X1_22 ( .A(_abc_40344_n2645), .B(_abc_40344_n2571), .C(_abc_40344_n2655), .Y(_abc_40344_n2656) );
  NOR3X1 NOR3X1_23 ( .A(_abc_40344_n2642), .B(_abc_40344_n2660), .C(_abc_40344_n2656), .Y(_abc_40344_n2661) );
  NOR3X1 NOR3X1_24 ( .A(_abc_40344_n3083), .B(_abc_40344_n3085), .C(_abc_40344_n3082), .Y(_abc_40344_n3086) );
  NOR3X1 NOR3X1_25 ( .A(_abc_40344_n3092), .B(_abc_40344_n3094), .C(_abc_40344_n3091), .Y(_abc_40344_n3095) );
  NOR3X1 NOR3X1_26 ( .A(_abc_40344_n4220), .B(_abc_40344_n4019), .C(_abc_40344_n4221_1), .Y(_abc_40344_n4222) );
  NOR3X1 NOR3X1_3 ( .A(IR_REG_2_), .B(IR_REG_1_), .C(IR_REG_0_), .Y(_abc_40344_n572) );
  NOR3X1 NOR3X1_4 ( .A(IR_REG_24_), .B(_abc_40344_n555), .C(_abc_40344_n576), .Y(_abc_40344_n577_1) );
  NOR3X1 NOR3X1_5 ( .A(IR_REG_23_), .B(IR_REG_22_), .C(IR_REG_28_), .Y(_abc_40344_n592) );
  NOR3X1 NOR3X1_6 ( .A(_abc_40344_n547), .B(_abc_40344_n595_1), .C(_abc_40344_n593_1), .Y(_abc_40344_n596_1) );
  NOR3X1 NOR3X1_7 ( .A(_abc_40344_n526), .B(_abc_40344_n571_1), .C(_abc_40344_n573_1), .Y(_abc_40344_n621) );
  NOR3X1 NOR3X1_8 ( .A(_abc_40344_n658_1), .B(_abc_40344_n571_1), .C(_abc_40344_n573_1), .Y(_abc_40344_n663) );
  NOR3X1 NOR3X1_9 ( .A(_abc_40344_n1012), .B(_abc_40344_n1050), .C(_abc_40344_n690), .Y(_abc_40344_n1051_1) );
  OAI21X1 OAI21X1_1 ( .A(_abc_40344_n552), .B(_abc_40344_n550_1), .C(IR_REG_26_), .Y(_abc_40344_n553_1) );
  OAI21X1 OAI21X1_10 ( .A(_abc_40344_n547), .B(_abc_40344_n544), .C(IR_REG_22_), .Y(_abc_40344_n623) );
  OAI21X1 OAI21X1_100 ( .A(_abc_40344_n802), .B(_abc_40344_n1176), .C(_abc_40344_n1177), .Y(_abc_40344_n1178) );
  OAI21X1 OAI21X1_1000 ( .A(_abc_40344_n3287), .B(_abc_40344_n4197_1), .C(_abc_40344_n4237), .Y(_abc_40344_n4308_1) );
  OAI21X1 OAI21X1_1001 ( .A(_abc_40344_n3270), .B(_abc_40344_n4203_1), .C(_abc_40344_n4237), .Y(_abc_40344_n4311_1) );
  OAI21X1 OAI21X1_1002 ( .A(_abc_40344_n4209_1), .B(_abc_40344_n3251), .C(_abc_40344_n4237), .Y(_abc_40344_n4314_1) );
  OAI21X1 OAI21X1_1003 ( .A(_abc_40344_n3231), .B(_abc_40344_n4215_1), .C(_abc_40344_n4237), .Y(_abc_40344_n4317_1) );
  OAI21X1 OAI21X1_1004 ( .A(_abc_40344_n4010), .B(_abc_40344_n4223_1), .C(_abc_40344_n4237), .Y(_abc_40344_n4320_1) );
  OAI21X1 OAI21X1_1005 ( .A(_abc_40344_n4228), .B(_abc_40344_n4227_1), .C(_abc_40344_n4237), .Y(_abc_40344_n4323_1) );
  OAI21X1 OAI21X1_1006 ( .A(_abc_40344_n1919), .B(_abc_40344_n4237), .C(_abc_40344_n4324), .Y(n808) );
  OAI21X1 OAI21X1_1007 ( .A(_abc_40344_n4233_1), .B(_abc_40344_n4232), .C(_abc_40344_n4237), .Y(_abc_40344_n4326_1) );
  OAI21X1 OAI21X1_1008 ( .A(_abc_40344_n979), .B(_abc_40344_n4041), .C(REG1_REG_31_), .Y(_abc_40344_n4327) );
  OAI21X1 OAI21X1_1009 ( .A(_abc_40344_n1675), .B(_abc_40344_n4329_1), .C(_abc_40344_n4330), .Y(n1058) );
  OAI21X1 OAI21X1_101 ( .A(REG3_REG_17_), .B(_abc_40344_n1158), .C(_abc_40344_n1058), .Y(_abc_40344_n1179) );
  OAI21X1 OAI21X1_1010 ( .A(_abc_40344_n863), .B(_abc_40344_n4329_1), .C(_abc_40344_n4332), .Y(n1062) );
  OAI21X1 OAI21X1_1011 ( .A(_abc_40344_n841), .B(_abc_40344_n4329_1), .C(_abc_40344_n4334), .Y(n1066) );
  OAI21X1 OAI21X1_1012 ( .A(_abc_40344_n809), .B(_abc_40344_n4329_1), .C(_abc_40344_n4336), .Y(n1070) );
  OAI21X1 OAI21X1_1013 ( .A(_abc_40344_n787_1), .B(_abc_40344_n4329_1), .C(_abc_40344_n4338), .Y(n1074) );
  OAI21X1 OAI21X1_1014 ( .A(_abc_40344_n763), .B(_abc_40344_n4329_1), .C(_abc_40344_n4340), .Y(n1078) );
  OAI21X1 OAI21X1_1015 ( .A(_abc_40344_n1021), .B(_abc_40344_n4329_1), .C(_abc_40344_n4342), .Y(n1082) );
  OAI21X1 OAI21X1_1016 ( .A(_abc_40344_n927_1), .B(_abc_40344_n4329_1), .C(_abc_40344_n4344), .Y(n1086) );
  OAI21X1 OAI21X1_1017 ( .A(_abc_40344_n1018), .B(_abc_40344_n4329_1), .C(_abc_40344_n4346), .Y(n1090) );
  OAI21X1 OAI21X1_1018 ( .A(_abc_40344_n1361), .B(_abc_40344_n4329_1), .C(_abc_40344_n4348), .Y(n1094) );
  OAI21X1 OAI21X1_1019 ( .A(_abc_40344_n1787), .B(_abc_40344_n4329_1), .C(_abc_40344_n4350), .Y(n1098) );
  OAI21X1 OAI21X1_102 ( .A(_abc_40344_n921), .B(_abc_40344_n1179), .C(_abc_40344_n1180_1), .Y(_abc_40344_n1181) );
  OAI21X1 OAI21X1_1020 ( .A(_abc_40344_n1284), .B(_abc_40344_n4329_1), .C(_abc_40344_n4352), .Y(n1102) );
  OAI21X1 OAI21X1_1021 ( .A(_abc_40344_n1305), .B(_abc_40344_n4329_1), .C(_abc_40344_n4354), .Y(n1106) );
  OAI21X1 OAI21X1_1022 ( .A(_abc_40344_n1259), .B(_abc_40344_n4329_1), .C(_abc_40344_n4356), .Y(n1110) );
  OAI21X1 OAI21X1_1023 ( .A(_abc_40344_n1818), .B(_abc_40344_n4329_1), .C(_abc_40344_n4358), .Y(n1114) );
  OAI21X1 OAI21X1_1024 ( .A(_abc_40344_n1209_1), .B(_abc_40344_n4329_1), .C(_abc_40344_n4360), .Y(n1118) );
  OAI21X1 OAI21X1_1025 ( .A(_abc_40344_n1167), .B(_abc_40344_n4329_1), .C(_abc_40344_n4362), .Y(n1122) );
  OAI21X1 OAI21X1_1026 ( .A(_abc_40344_n1185), .B(_abc_40344_n4329_1), .C(_abc_40344_n4364), .Y(n1126) );
  OAI21X1 OAI21X1_1027 ( .A(_abc_40344_n1138), .B(_abc_40344_n4329_1), .C(_abc_40344_n4366), .Y(n1130) );
  OAI21X1 OAI21X1_1028 ( .A(_abc_40344_n1414), .B(_abc_40344_n4329_1), .C(_abc_40344_n4368), .Y(n1134) );
  OAI21X1 OAI21X1_1029 ( .A(_abc_40344_n1429), .B(_abc_40344_n4329_1), .C(_abc_40344_n4370), .Y(n1138) );
  OAI21X1 OAI21X1_103 ( .A(_abc_40344_n1188), .B(_abc_40344_n1190), .C(_abc_40344_n1172), .Y(_abc_40344_n1191) );
  OAI21X1 OAI21X1_1030 ( .A(_abc_40344_n1440), .B(_abc_40344_n4329_1), .C(_abc_40344_n4372), .Y(n1142) );
  OAI21X1 OAI21X1_1031 ( .A(_abc_40344_n4329_1), .B(_abc_40344_n1110), .C(_abc_40344_n4374), .Y(n1146) );
  OAI21X1 OAI21X1_1032 ( .A(_abc_40344_n4329_1), .B(_abc_40344_n1090_1), .C(_abc_40344_n4376), .Y(n1150) );
  OAI21X1 OAI21X1_1033 ( .A(_abc_40344_n4329_1), .B(_abc_40344_n1577), .C(_abc_40344_n4378), .Y(n1154) );
  OAI21X1 OAI21X1_1034 ( .A(_abc_40344_n4329_1), .B(_abc_40344_n1489), .C(_abc_40344_n4380), .Y(n1158) );
  OAI21X1 OAI21X1_1035 ( .A(_abc_40344_n4329_1), .B(_abc_40344_n1506), .C(_abc_40344_n4382), .Y(n1162) );
  OAI21X1 OAI21X1_1036 ( .A(_abc_40344_n4329_1), .B(_abc_40344_n1074), .C(_abc_40344_n4384), .Y(n1166) );
  OAI21X1 OAI21X1_1037 ( .A(_abc_40344_n4329_1), .B(_abc_40344_n1550), .C(_abc_40344_n4386), .Y(n1170) );
  OAI21X1 OAI21X1_1038 ( .A(_abc_40344_n4329_1), .B(_abc_40344_n1646), .C(_abc_40344_n4388), .Y(n1174) );
  OAI21X1 OAI21X1_1039 ( .A(_abc_40344_n2095), .B(_abc_40344_n4329_1), .C(_abc_40344_n4390), .Y(n1178) );
  OAI21X1 OAI21X1_104 ( .A(IR_REG_14_), .B(_abc_40344_n677), .C(IR_REG_15_), .Y(_abc_40344_n1192) );
  OAI21X1 OAI21X1_1040 ( .A(_abc_40344_n1914), .B(_abc_40344_n4329_1), .C(_abc_40344_n4392), .Y(n1182) );
  OAI21X1 OAI21X1_105 ( .A(IR_REG_31_), .B(IR_REG_15_), .C(_abc_40344_n1195), .Y(_abc_40344_n1196) );
  OAI21X1 OAI21X1_106 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(_abc_40344_n1198), .Y(_abc_40344_n1199) );
  OAI21X1 OAI21X1_107 ( .A(_abc_40344_n802), .B(_abc_40344_n1197), .C(_abc_40344_n1199), .Y(_abc_40344_n1200) );
  OAI21X1 OAI21X1_108 ( .A(_abc_40344_n921), .B(_abc_40344_n1203), .C(_abc_40344_n1204), .Y(_abc_40344_n1205) );
  OAI21X1 OAI21X1_109 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1219), .C(_abc_40344_n1220), .Y(_abc_40344_n1221) );
  OAI21X1 OAI21X1_11 ( .A(IR_REG_31_), .B(_abc_40344_n620), .C(_abc_40344_n624), .Y(_abc_40344_n625) );
  OAI21X1 OAI21X1_110 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_14_), .Y(_abc_40344_n1223) );
  OAI21X1 OAI21X1_111 ( .A(_abc_40344_n802), .B(_abc_40344_n1222), .C(_abc_40344_n1223), .Y(_abc_40344_n1224) );
  OAI21X1 OAI21X1_112 ( .A(_abc_40344_n1049_1), .B(_abc_40344_n1055), .C(_abc_40344_n1225_1), .Y(_abc_40344_n1226) );
  OAI21X1 OAI21X1_113 ( .A(_abc_40344_n921), .B(_abc_40344_n1228), .C(_abc_40344_n1229), .Y(_abc_40344_n1230) );
  OAI21X1 OAI21X1_114 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1248), .C(_abc_40344_n1242), .Y(_abc_40344_n1249) );
  OAI21X1 OAI21X1_115 ( .A(DATAI_13_), .B(_abc_40344_n705_1), .C(_abc_40344_n1263), .Y(_abc_40344_n1264) );
  OAI21X1 OAI21X1_116 ( .A(IR_REG_31_), .B(IR_REG_11_), .C(_abc_40344_n1270), .Y(_abc_40344_n1271) );
  OAI21X1 OAI21X1_117 ( .A(IR_REG_11_), .B(_abc_40344_n1268), .C(IR_REG_12_), .Y(_abc_40344_n1290) );
  OAI21X1 OAI21X1_118 ( .A(IR_REG_31_), .B(IR_REG_12_), .C(_abc_40344_n1292), .Y(_abc_40344_n1293_1) );
  OAI21X1 OAI21X1_119 ( .A(DATAI_12_), .B(_abc_40344_n705_1), .C(_abc_40344_n1294), .Y(_abc_40344_n1295) );
  OAI21X1 OAI21X1_12 ( .A(_abc_40344_n627), .B(_abc_40344_n581), .C(_abc_40344_n586), .Y(_abc_40344_n628) );
  OAI21X1 OAI21X1_120 ( .A(_abc_40344_n921), .B(_abc_40344_n1302), .C(_abc_40344_n1303), .Y(_abc_40344_n1304_1) );
  OAI21X1 OAI21X1_121 ( .A(_abc_40344_n1306), .B(_abc_40344_n1311), .C(_abc_40344_n1267), .Y(_abc_40344_n1312) );
  OAI21X1 OAI21X1_122 ( .A(_abc_40344_n1289), .B(_abc_40344_n1312), .C(_abc_40344_n1315), .Y(_abc_40344_n1316) );
  OAI21X1 OAI21X1_123 ( .A(IR_REG_9_), .B(_abc_40344_n1245), .C(IR_REG_10_), .Y(_abc_40344_n1322) );
  OAI21X1 OAI21X1_124 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1323), .C(_abc_40344_n1324), .Y(_abc_40344_n1325) );
  OAI21X1 OAI21X1_125 ( .A(_abc_40344_n1321), .B(_abc_40344_n705_1), .C(_abc_40344_n1326), .Y(_abc_40344_n1327) );
  OAI21X1 OAI21X1_126 ( .A(_abc_40344_n1332), .B(_abc_40344_n761_1), .C(_abc_40344_n1333), .Y(_abc_40344_n1334) );
  OAI21X1 OAI21X1_127 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1344), .C(_abc_40344_n1346), .Y(_abc_40344_n1347) );
  OAI21X1 OAI21X1_128 ( .A(_abc_40344_n1341), .B(_abc_40344_n705_1), .C(_abc_40344_n1349), .Y(_abc_40344_n1350) );
  OAI21X1 OAI21X1_129 ( .A(_abc_40344_n1011), .B(_abc_40344_n909), .C(_abc_40344_n1356), .Y(_abc_40344_n1357) );
  OAI21X1 OAI21X1_13 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(_abc_40344_n628), .Y(_abc_40344_n629) );
  OAI21X1 OAI21X1_130 ( .A(_abc_40344_n542_1), .B(_abc_40344_n706), .C(IR_REG_8_), .Y(_abc_40344_n1369) );
  OAI21X1 OAI21X1_131 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1370), .C(_abc_40344_n1371_1), .Y(_abc_40344_n1372) );
  OAI21X1 OAI21X1_132 ( .A(DATAI_8_), .B(_abc_40344_n705_1), .C(_abc_40344_n1374), .Y(_abc_40344_n1375) );
  OAI21X1 OAI21X1_133 ( .A(_abc_40344_n932), .B(_abc_40344_n726), .C(_abc_40344_n933), .Y(_abc_40344_n1384) );
  OAI21X1 OAI21X1_134 ( .A(_abc_40344_n935_1), .B(_abc_40344_n768), .C(_abc_40344_n1384), .Y(_abc_40344_n1385) );
  OAI21X1 OAI21X1_135 ( .A(_abc_40344_n1401), .B(_abc_40344_n1396_1), .C(_abc_40344_n1143), .Y(_abc_40344_n1402) );
  OAI21X1 OAI21X1_136 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_19_), .Y(_abc_40344_n1403) );
  OAI21X1 OAI21X1_137 ( .A(_abc_40344_n802), .B(_abc_40344_n646), .C(_abc_40344_n1403), .Y(_abc_40344_n1404) );
  OAI21X1 OAI21X1_138 ( .A(_abc_40344_n1047), .B(_abc_40344_n1058), .C(_abc_40344_n1405), .Y(_abc_40344_n1406) );
  OAI21X1 OAI21X1_139 ( .A(_abc_40344_n921), .B(_abc_40344_n1408), .C(_abc_40344_n1409_1), .Y(_abc_40344_n1410) );
  OAI21X1 OAI21X1_14 ( .A(IR_REG_31_), .B(_abc_40344_n554_1), .C(_abc_40344_n558), .Y(_abc_40344_n633_1) );
  OAI21X1 OAI21X1_140 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_20_), .Y(_abc_40344_n1421_1) );
  OAI21X1 OAI21X1_141 ( .A(_abc_40344_n1405), .B(_abc_40344_n1125), .C(_abc_40344_n1046), .Y(_abc_40344_n1422) );
  OAI21X1 OAI21X1_142 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_21_), .Y(_abc_40344_n1433) );
  OAI21X1 OAI21X1_143 ( .A(_abc_40344_n1046), .B(_abc_40344_n1060), .C(_abc_40344_n1045_1), .Y(_abc_40344_n1435) );
  OAI21X1 OAI21X1_144 ( .A(_abc_40344_n1430), .B(_abc_40344_n1432), .C(_abc_40344_n1445), .Y(_abc_40344_n1446) );
  OAI21X1 OAI21X1_145 ( .A(_abc_40344_n1417), .B(_abc_40344_n1420), .C(_abc_40344_n1447), .Y(_abc_40344_n1448) );
  OAI21X1 OAI21X1_146 ( .A(_abc_40344_n1446), .B(_abc_40344_n1452), .C(_abc_40344_n1455), .Y(_abc_40344_n1456) );
  OAI21X1 OAI21X1_147 ( .A(_abc_40344_n1458), .B(_abc_40344_n1449), .C(_abc_40344_n1118_1), .Y(_abc_40344_n1459) );
  OAI21X1 OAI21X1_148 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_24_), .Y(_abc_40344_n1462) );
  OAI21X1 OAI21X1_149 ( .A(_abc_40344_n1467), .B(_abc_40344_n761_1), .C(_abc_40344_n1468), .Y(_abc_40344_n1469) );
  OAI21X1 OAI21X1_15 ( .A(IR_REG_24_), .B(_abc_40344_n550_1), .C(IR_REG_25_), .Y(_abc_40344_n634) );
  OAI21X1 OAI21X1_150 ( .A(_abc_40344_n921), .B(_abc_40344_n1466), .C(_abc_40344_n1470), .Y(_abc_40344_n1471) );
  OAI21X1 OAI21X1_151 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_25_), .Y(_abc_40344_n1477) );
  OAI21X1 OAI21X1_152 ( .A(_abc_40344_n1043), .B(_abc_40344_n1063), .C(REG3_REG_25_), .Y(_abc_40344_n1478) );
  OAI21X1 OAI21X1_153 ( .A(_abc_40344_n1484), .B(_abc_40344_n761_1), .C(_abc_40344_n1485), .Y(_abc_40344_n1486) );
  OAI21X1 OAI21X1_154 ( .A(_abc_40344_n921), .B(_abc_40344_n1481), .C(_abc_40344_n1487), .Y(_abc_40344_n1488) );
  OAI21X1 OAI21X1_155 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_26_), .Y(_abc_40344_n1494) );
  OAI21X1 OAI21X1_156 ( .A(_abc_40344_n1044), .B(_abc_40344_n1464), .C(REG3_REG_26_), .Y(_abc_40344_n1496) );
  OAI21X1 OAI21X1_157 ( .A(_abc_40344_n1501), .B(_abc_40344_n761_1), .C(_abc_40344_n1502), .Y(_abc_40344_n1503_1) );
  OAI21X1 OAI21X1_158 ( .A(_abc_40344_n1490), .B(_abc_40344_n1493), .C(_abc_40344_n1511_1), .Y(_abc_40344_n1512) );
  OAI21X1 OAI21X1_159 ( .A(_abc_40344_n1512), .B(_abc_40344_n1515), .C(_abc_40344_n1519), .Y(_abc_40344_n1520_1) );
  OAI21X1 OAI21X1_16 ( .A(_abc_40344_n615), .B(_abc_40344_n638), .C(IR_REG_31_), .Y(_abc_40344_n639_1) );
  OAI21X1 OAI21X1_160 ( .A(_abc_40344_n1514_1), .B(_abc_40344_n1461), .C(_abc_40344_n1521), .Y(_abc_40344_n1522) );
  OAI21X1 OAI21X1_161 ( .A(_abc_40344_n1211), .B(_abc_40344_n1214), .C(_abc_40344_n1395), .Y(_abc_40344_n1525) );
  OAI21X1 OAI21X1_162 ( .A(_abc_40344_n1534), .B(_abc_40344_n1533), .C(_abc_40344_n1082), .Y(_abc_40344_n1535) );
  OAI21X1 OAI21X1_163 ( .A(_abc_40344_n1545), .B(_abc_40344_n761_1), .C(_abc_40344_n1546), .Y(_abc_40344_n1547) );
  OAI21X1 OAI21X1_164 ( .A(_abc_40344_n1042), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1552) );
  OAI21X1 OAI21X1_165 ( .A(_abc_40344_n982), .B(_abc_40344_n1006), .C(_abc_40344_n1000), .Y(_abc_40344_n1554) );
  OAI21X1 OAI21X1_166 ( .A(_abc_40344_n1068), .B(_abc_40344_n1555), .C(_abc_40344_n1553), .Y(_abc_40344_n1556) );
  OAI21X1 OAI21X1_167 ( .A(_abc_40344_n1523), .B(_abc_40344_n1536), .C(_abc_40344_n1557), .Y(n1326) );
  OAI21X1 OAI21X1_168 ( .A(_abc_40344_n1225_1), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1566) );
  OAI21X1 OAI21X1_169 ( .A(_abc_40344_n1228), .B(_abc_40344_n1555), .C(_abc_40344_n1567), .Y(_abc_40344_n1568) );
  OAI21X1 OAI21X1_17 ( .A(IR_REG_31_), .B(IR_REG_20_), .C(_abc_40344_n639_1), .Y(_abc_40344_n640) );
  OAI21X1 OAI21X1_170 ( .A(_abc_40344_n1562), .B(_abc_40344_n1564), .C(_abc_40344_n1569), .Y(n1321) );
  OAI21X1 OAI21X1_171 ( .A(_abc_40344_n1117), .B(_abc_40344_n1571), .C(_abc_40344_n1116), .Y(_abc_40344_n1572) );
  OAI21X1 OAI21X1_172 ( .A(_abc_40344_n1573), .B(_abc_40344_n1572), .C(_abc_40344_n993), .Y(_abc_40344_n1575) );
  OAI21X1 OAI21X1_173 ( .A(_abc_40344_n1576), .B(_abc_40344_n1578), .C(_abc_40344_n1005), .Y(_abc_40344_n1579) );
  OAI21X1 OAI21X1_174 ( .A(_abc_40344_n1083), .B(_abc_40344_n1580), .C(_abc_40344_n1581), .Y(_abc_40344_n1582) );
  OAI21X1 OAI21X1_175 ( .A(_abc_40344_n1574), .B(_abc_40344_n1575), .C(_abc_40344_n1584), .Y(n1316) );
  OAI21X1 OAI21X1_176 ( .A(_abc_40344_n1364), .B(_abc_40344_n1366), .C(_abc_40344_n1391), .Y(_abc_40344_n1586) );
  OAI21X1 OAI21X1_177 ( .A(_abc_40344_n1586), .B(_abc_40344_n1589), .C(_abc_40344_n1591), .Y(_abc_40344_n1592) );
  OAI21X1 OAI21X1_178 ( .A(_abc_40344_n1052_1), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1594) );
  OAI21X1 OAI21X1_179 ( .A(_abc_40344_n1330), .B(_abc_40344_n1555), .C(_abc_40344_n1595), .Y(_abc_40344_n1596) );
  OAI21X1 OAI21X1_18 ( .A(IR_REG_18_), .B(_abc_40344_n544), .C(IR_REG_19_), .Y(_abc_40344_n643) );
  OAI21X1 OAI21X1_180 ( .A(_abc_40344_n1602), .B(_abc_40344_n1600), .C(_abc_40344_n1601), .Y(_abc_40344_n1603) );
  OAI21X1 OAI21X1_181 ( .A(DATAI_3_), .B(_abc_40344_n705_1), .C(_abc_40344_n1608), .Y(_abc_40344_n1609) );
  OAI21X1 OAI21X1_182 ( .A(_abc_40344_n688_1), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1610) );
  OAI21X1 OAI21X1_183 ( .A(_abc_40344_n1609), .B(_abc_40344_n1580), .C(_abc_40344_n1611), .Y(_abc_40344_n1612) );
  OAI21X1 OAI21X1_184 ( .A(_abc_40344_n1590), .B(_abc_40344_n1604), .C(_abc_40344_n1614), .Y(n1306) );
  OAI21X1 OAI21X1_185 ( .A(_abc_40344_n1142), .B(_abc_40344_n1616), .C(_abc_40344_n1141), .Y(_abc_40344_n1617) );
  OAI21X1 OAI21X1_186 ( .A(_abc_40344_n1619), .B(_abc_40344_n1617), .C(_abc_40344_n993), .Y(_abc_40344_n1621) );
  OAI21X1 OAI21X1_187 ( .A(_abc_40344_n1405), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1623) );
  OAI21X1 OAI21X1_188 ( .A(_abc_40344_n1408), .B(_abc_40344_n1555), .C(_abc_40344_n1624), .Y(_abc_40344_n1625) );
  OAI21X1 OAI21X1_189 ( .A(_abc_40344_n1620), .B(_abc_40344_n1621), .C(_abc_40344_n1626), .Y(n1301) );
  OAI21X1 OAI21X1_19 ( .A(IR_REG_31_), .B(IR_REG_19_), .C(_abc_40344_n645), .Y(_abc_40344_n646) );
  OAI21X1 OAI21X1_190 ( .A(_abc_40344_n1514_1), .B(_abc_40344_n1461), .C(_abc_40344_n1628), .Y(_abc_40344_n1629) );
  OAI21X1 OAI21X1_191 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_28_), .Y(_abc_40344_n1630) );
  OAI21X1 OAI21X1_192 ( .A(_abc_40344_n1534), .B(_abc_40344_n1533), .C(_abc_40344_n1636), .Y(_abc_40344_n1637) );
  OAI21X1 OAI21X1_193 ( .A(_abc_40344_n1641), .B(_abc_40344_n761_1), .C(_abc_40344_n1642), .Y(_abc_40344_n1643) );
  OAI21X1 OAI21X1_194 ( .A(_abc_40344_n921), .B(_abc_40344_n1640), .C(_abc_40344_n1644), .Y(_abc_40344_n1645) );
  OAI21X1 OAI21X1_195 ( .A(_abc_40344_n1538), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1650) );
  OAI21X1 OAI21X1_196 ( .A(_abc_40344_n1555), .B(_abc_40344_n1648), .C(_abc_40344_n1651), .Y(_abc_40344_n1652) );
  OAI21X1 OAI21X1_197 ( .A(_abc_40344_n1590), .B(_abc_40344_n1639), .C(_abc_40344_n1653), .Y(n1296) );
  OAI21X1 OAI21X1_198 ( .A(_abc_40344_n1379), .B(_abc_40344_n1383_1), .C(_abc_40344_n1658), .Y(_abc_40344_n1660) );
  OAI21X1 OAI21X1_199 ( .A(_abc_40344_n1663), .B(_abc_40344_n705_1), .C(_abc_40344_n1664), .Y(_abc_40344_n1665) );
  OAI21X1 OAI21X1_2 ( .A(_abc_40344_n559_1), .B(_abc_40344_n556), .C(IR_REG_24_), .Y(_abc_40344_n562) );
  OAI21X1 OAI21X1_20 ( .A(_abc_40344_n656), .B(_abc_40344_n660), .C(IR_REG_30_), .Y(_abc_40344_n661) );
  OAI21X1 OAI21X1_200 ( .A(_abc_40344_n1011), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1666) );
  OAI21X1 OAI21X1_201 ( .A(_abc_40344_n1016), .B(_abc_40344_n1555), .C(_abc_40344_n1667), .Y(_abc_40344_n1668) );
  OAI21X1 OAI21X1_202 ( .A(_abc_40344_n1659), .B(_abc_40344_n1661), .C(_abc_40344_n1669), .Y(n1291) );
  OAI21X1 OAI21X1_203 ( .A(_abc_40344_n1671), .B(_abc_40344_n1672), .C(_abc_40344_n993), .Y(_abc_40344_n1674) );
  OAI21X1 OAI21X1_204 ( .A(_abc_40344_n1675), .B(_abc_40344_n1023_1), .C(_abc_40344_n1676), .Y(_abc_40344_n1677) );
  OAI21X1 OAI21X1_205 ( .A(_abc_40344_n1678), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1679) );
  OAI21X1 OAI21X1_206 ( .A(_abc_40344_n1678), .B(_abc_40344_n1000), .C(_abc_40344_n1680), .Y(_abc_40344_n1681) );
  OAI21X1 OAI21X1_207 ( .A(_abc_40344_n1673), .B(_abc_40344_n1674), .C(_abc_40344_n1682), .Y(n1286) );
  OAI21X1 OAI21X1_208 ( .A(_abc_40344_n1417), .B(_abc_40344_n1420), .C(_abc_40344_n1617), .Y(_abc_40344_n1684) );
  OAI21X1 OAI21X1_209 ( .A(_abc_40344_n1416), .B(_abc_40344_n1450), .C(_abc_40344_n1684), .Y(_abc_40344_n1685) );
  OAI21X1 OAI21X1_21 ( .A(_abc_40344_n669), .B(_abc_40344_n671_1), .C(IR_REG_31_), .Y(_abc_40344_n672) );
  OAI21X1 OAI21X1_210 ( .A(_abc_40344_n1430), .B(_abc_40344_n1432), .C(_abc_40344_n1685), .Y(_abc_40344_n1686) );
  OAI21X1 OAI21X1_211 ( .A(_abc_40344_n1442), .B(_abc_40344_n1444), .C(_abc_40344_n1447), .Y(_abc_40344_n1691) );
  OAI21X1 OAI21X1_212 ( .A(_abc_40344_n1691), .B(_abc_40344_n1690), .C(_abc_40344_n993), .Y(_abc_40344_n1692) );
  OAI21X1 OAI21X1_213 ( .A(_abc_40344_n1045_1), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1696) );
  OAI21X1 OAI21X1_214 ( .A(_abc_40344_n1006), .B(_abc_40344_n1695), .C(_abc_40344_n1697), .Y(_abc_40344_n1698) );
  OAI21X1 OAI21X1_215 ( .A(_abc_40344_n1692), .B(_abc_40344_n1688), .C(_abc_40344_n1699), .Y(n1281) );
  OAI21X1 OAI21X1_216 ( .A(_abc_40344_n1702), .B(_abc_40344_n1586), .C(_abc_40344_n1588), .Y(_abc_40344_n1703) );
  OAI21X1 OAI21X1_217 ( .A(_abc_40344_n1286), .B(_abc_40344_n1288), .C(_abc_40344_n1704), .Y(_abc_40344_n1705) );
  OAI21X1 OAI21X1_218 ( .A(_abc_40344_n1701), .B(_abc_40344_n1706), .C(_abc_40344_n993), .Y(_abc_40344_n1708) );
  OAI21X1 OAI21X1_219 ( .A(_abc_40344_n1299), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1710) );
  OAI21X1 OAI21X1_22 ( .A(_abc_40344_n677), .B(_abc_40344_n681), .C(IR_REG_29_), .Y(_abc_40344_n682) );
  OAI21X1 OAI21X1_220 ( .A(_abc_40344_n1302), .B(_abc_40344_n1555), .C(_abc_40344_n1711), .Y(_abc_40344_n1712) );
  OAI21X1 OAI21X1_221 ( .A(_abc_40344_n1707), .B(_abc_40344_n1708), .C(_abc_40344_n1713), .Y(n1276) );
  OAI21X1 OAI21X1_222 ( .A(_abc_40344_n1476), .B(_abc_40344_n1461), .C(_abc_40344_n1515), .Y(_abc_40344_n1717) );
  OAI21X1 OAI21X1_223 ( .A(_abc_40344_n1719), .B(_abc_40344_n1720), .C(_abc_40344_n1716), .Y(_abc_40344_n1721) );
  OAI21X1 OAI21X1_224 ( .A(_abc_40344_n1723), .B(_abc_40344_n1724), .C(_abc_40344_n1005), .Y(_abc_40344_n1725) );
  OAI21X1 OAI21X1_225 ( .A(_abc_40344_n1477), .B(_abc_40344_n1580), .C(_abc_40344_n1727), .Y(_abc_40344_n1728) );
  OAI21X1 OAI21X1_226 ( .A(_abc_40344_n1718), .B(_abc_40344_n1722), .C(_abc_40344_n1730), .Y(n1271) );
  OAI21X1 OAI21X1_227 ( .A(_abc_40344_n1733), .B(_abc_40344_n1525), .C(_abc_40344_n993), .Y(_abc_40344_n1735) );
  OAI21X1 OAI21X1_228 ( .A(_abc_40344_n1155_1), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1737) );
  OAI21X1 OAI21X1_229 ( .A(_abc_40344_n1161), .B(_abc_40344_n1555), .C(_abc_40344_n1738), .Y(_abc_40344_n1739) );
  OAI21X1 OAI21X1_23 ( .A(_abc_40344_n702), .B(_abc_40344_n703), .C(IR_REG_31_), .Y(_abc_40344_n704) );
  OAI21X1 OAI21X1_230 ( .A(_abc_40344_n1734), .B(_abc_40344_n1735), .C(_abc_40344_n1740), .Y(n1266) );
  OAI21X1 OAI21X1_231 ( .A(_abc_40344_n736), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1745) );
  OAI21X1 OAI21X1_232 ( .A(_abc_40344_n738_1), .B(_abc_40344_n1555), .C(_abc_40344_n1746), .Y(_abc_40344_n1747) );
  OAI21X1 OAI21X1_233 ( .A(_abc_40344_n1590), .B(_abc_40344_n1743), .C(_abc_40344_n1748), .Y(n1261) );
  OAI21X1 OAI21X1_234 ( .A(_abc_40344_n1398), .B(_abc_40344_n1525), .C(_abc_40344_n1524), .Y(_abc_40344_n1751) );
  OAI21X1 OAI21X1_235 ( .A(_abc_40344_n1750), .B(_abc_40344_n1397), .C(_abc_40344_n1399), .Y(_abc_40344_n1754) );
  OAI21X1 OAI21X1_236 ( .A(_abc_40344_n1754), .B(_abc_40344_n1753), .C(_abc_40344_n993), .Y(_abc_40344_n1755) );
  OAI21X1 OAI21X1_237 ( .A(_abc_40344_n1757), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1758) );
  OAI21X1 OAI21X1_238 ( .A(_abc_40344_n1179), .B(_abc_40344_n1555), .C(_abc_40344_n1759), .Y(_abc_40344_n1760) );
  OAI21X1 OAI21X1_239 ( .A(_abc_40344_n1755), .B(_abc_40344_n1752), .C(_abc_40344_n1761), .Y(n1256) );
  OAI21X1 OAI21X1_24 ( .A(_abc_40344_n559_1), .B(_abc_40344_n710_1), .C(_abc_40344_n711), .Y(_abc_40344_n712) );
  OAI21X1 OAI21X1_240 ( .A(_abc_40344_n1765), .B(_abc_40344_n1461), .C(_abc_40344_n993), .Y(_abc_40344_n1766) );
  OAI21X1 OAI21X1_241 ( .A(_abc_40344_n1043), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1768) );
  OAI21X1 OAI21X1_242 ( .A(_abc_40344_n1466), .B(_abc_40344_n1555), .C(_abc_40344_n1769), .Y(_abc_40344_n1770) );
  OAI21X1 OAI21X1_243 ( .A(_abc_40344_n1764), .B(_abc_40344_n1766), .C(_abc_40344_n1771), .Y(n1251) );
  OAI21X1 OAI21X1_244 ( .A(_abc_40344_n687), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1776) );
  OAI21X1 OAI21X1_245 ( .A(_abc_40344_n1006), .B(_abc_40344_n1778), .C(_abc_40344_n1777), .Y(_abc_40344_n1779) );
  OAI21X1 OAI21X1_246 ( .A(_abc_40344_n1590), .B(_abc_40344_n1775), .C(_abc_40344_n1780), .Y(n1246) );
  OAI21X1 OAI21X1_247 ( .A(_abc_40344_n1356), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1789) );
  OAI21X1 OAI21X1_248 ( .A(_abc_40344_n1359_1), .B(_abc_40344_n1555), .C(_abc_40344_n1790), .Y(_abc_40344_n1791) );
  OAI21X1 OAI21X1_249 ( .A(_abc_40344_n1784), .B(_abc_40344_n1786), .C(_abc_40344_n1792), .Y(n1241) );
  OAI21X1 OAI21X1_25 ( .A(_abc_40344_n701), .B(_abc_40344_n705_1), .C(_abc_40344_n713_1), .Y(_abc_40344_n714) );
  OAI21X1 OAI21X1_250 ( .A(DATAI_0_), .B(_abc_40344_n705_1), .C(_abc_40344_n1796), .Y(_abc_40344_n1797) );
  OAI21X1 OAI21X1_251 ( .A(_abc_40344_n745), .B(_abc_40344_n1797), .C(_abc_40344_n891), .Y(_abc_40344_n1798) );
  OAI21X1 OAI21X1_252 ( .A(_abc_40344_n1794), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1802) );
  OAI21X1 OAI21X1_253 ( .A(_abc_40344_n1797), .B(_abc_40344_n1580), .C(_abc_40344_n1803), .Y(_abc_40344_n1804) );
  OAI21X1 OAI21X1_254 ( .A(_abc_40344_n1794), .B(_abc_40344_n1555), .C(_abc_40344_n1805), .Y(n1236) );
  OAI21X1 OAI21X1_255 ( .A(_abc_40344_n1808), .B(_abc_40344_n1685), .C(_abc_40344_n993), .Y(_abc_40344_n1810) );
  OAI21X1 OAI21X1_256 ( .A(_abc_40344_n1046), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1813) );
  OAI21X1 OAI21X1_257 ( .A(_abc_40344_n1423), .B(_abc_40344_n1555), .C(_abc_40344_n1814), .Y(_abc_40344_n1815) );
  OAI21X1 OAI21X1_258 ( .A(_abc_40344_n1809), .B(_abc_40344_n1810), .C(_abc_40344_n1816), .Y(n1231) );
  OAI21X1 OAI21X1_259 ( .A(_abc_40344_n1049_1), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1820) );
  OAI21X1 OAI21X1_26 ( .A(_abc_40344_n717), .B(_abc_40344_n718), .C(_abc_40344_n716), .Y(_abc_40344_n719) );
  OAI21X1 OAI21X1_260 ( .A(_abc_40344_n1257), .B(_abc_40344_n1555), .C(_abc_40344_n1821), .Y(_abc_40344_n1822) );
  OAI21X1 OAI21X1_261 ( .A(_abc_40344_n1824), .B(_abc_40344_n1706), .C(_abc_40344_n1314), .Y(_abc_40344_n1825) );
  OAI21X1 OAI21X1_262 ( .A(_abc_40344_n1828), .B(_abc_40344_n1827), .C(_abc_40344_n993), .Y(_abc_40344_n1829) );
  OAI21X1 OAI21X1_263 ( .A(_abc_40344_n1826), .B(_abc_40344_n1829), .C(_abc_40344_n1823), .Y(n1226) );
  OAI21X1 OAI21X1_264 ( .A(_abc_40344_n1571), .B(_abc_40344_n1831), .C(_abc_40344_n1832), .Y(_abc_40344_n1833) );
  OAI21X1 OAI21X1_265 ( .A(_abc_40344_n1101), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1835) );
  OAI21X1 OAI21X1_266 ( .A(_abc_40344_n1104), .B(_abc_40344_n1555), .C(_abc_40344_n1836), .Y(_abc_40344_n1837) );
  OAI21X1 OAI21X1_267 ( .A(_abc_40344_n1023_1), .B(_abc_40344_n1787), .C(_abc_40344_n1840), .Y(_abc_40344_n1841) );
  OAI21X1 OAI21X1_268 ( .A(_abc_40344_n1053), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1842) );
  OAI21X1 OAI21X1_269 ( .A(_abc_40344_n1000), .B(_abc_40344_n1279), .C(_abc_40344_n1843), .Y(_abc_40344_n1844) );
  OAI21X1 OAI21X1_27 ( .A(IR_REG_4_), .B(_abc_40344_n706), .C(IR_REG_5_), .Y(_abc_40344_n729_1) );
  OAI21X1 OAI21X1_270 ( .A(_abc_40344_n1847), .B(_abc_40344_n1849), .C(_abc_40344_n1845), .Y(n1216) );
  OAI21X1 OAI21X1_271 ( .A(_abc_40344_n1854), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1855) );
  OAI21X1 OAI21X1_272 ( .A(_abc_40344_n1854), .B(_abc_40344_n1555), .C(_abc_40344_n1856), .Y(_abc_40344_n1857) );
  OAI21X1 OAI21X1_273 ( .A(_abc_40344_n1590), .B(_abc_40344_n1852), .C(_abc_40344_n1858), .Y(n1211) );
  OAI21X1 OAI21X1_274 ( .A(_abc_40344_n1616), .B(_abc_40344_n1860), .C(_abc_40344_n1861), .Y(_abc_40344_n1862) );
  OAI21X1 OAI21X1_275 ( .A(_abc_40344_n1047), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1864) );
  OAI21X1 OAI21X1_276 ( .A(_abc_40344_n1128), .B(_abc_40344_n1555), .C(_abc_40344_n1865), .Y(_abc_40344_n1866) );
  OAI21X1 OAI21X1_277 ( .A(_abc_40344_n686), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1873) );
  OAI21X1 OAI21X1_278 ( .A(_abc_40344_n1872), .B(_abc_40344_n1555), .C(_abc_40344_n1874), .Y(_abc_40344_n1875) );
  OAI21X1 OAI21X1_279 ( .A(_abc_40344_n1590), .B(_abc_40344_n1870), .C(_abc_40344_n1876), .Y(n1201) );
  OAI21X1 OAI21X1_28 ( .A(_abc_40344_n559_1), .B(_abc_40344_n730), .C(_abc_40344_n731), .Y(_abc_40344_n732_1) );
  OAI21X1 OAI21X1_280 ( .A(_abc_40344_n1516_1), .B(_abc_40344_n1879), .C(_abc_40344_n1517_1), .Y(_abc_40344_n1880) );
  OAI21X1 OAI21X1_281 ( .A(_abc_40344_n1882), .B(_abc_40344_n1720), .C(_abc_40344_n1883), .Y(_abc_40344_n1884) );
  OAI21X1 OAI21X1_282 ( .A(_abc_40344_n1041), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1889) );
  OAI21X1 OAI21X1_283 ( .A(_abc_40344_n1888), .B(_abc_40344_n1555), .C(_abc_40344_n1890), .Y(_abc_40344_n1891) );
  OAI21X1 OAI21X1_284 ( .A(_abc_40344_n1885), .B(_abc_40344_n1881), .C(_abc_40344_n1892), .Y(n1196) );
  OAI21X1 OAI21X1_285 ( .A(_abc_40344_n1894), .B(_abc_40344_n1895), .C(_abc_40344_n1896), .Y(_abc_40344_n1897) );
  OAI21X1 OAI21X1_286 ( .A(_abc_40344_n1154_1), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1899) );
  OAI21X1 OAI21X1_287 ( .A(_abc_40344_n1203), .B(_abc_40344_n1555), .C(_abc_40344_n1900), .Y(_abc_40344_n1901) );
  OAI21X1 OAI21X1_288 ( .A(_abc_40344_n1549), .B(_abc_40344_n1542), .C(_abc_40344_n1630), .Y(_abc_40344_n1904) );
  OAI21X1 OAI21X1_289 ( .A(DATAI_9_), .B(_abc_40344_n705_1), .C(_abc_40344_n1905), .Y(_abc_40344_n1906) );
  OAI21X1 OAI21X1_29 ( .A(_abc_40344_n728), .B(_abc_40344_n705_1), .C(_abc_40344_n733), .Y(_abc_40344_n734) );
  OAI21X1 OAI21X1_290 ( .A(_abc_40344_n1353), .B(_abc_40344_n1360), .C(_abc_40344_n1906), .Y(_abc_40344_n1907) );
  OAI21X1 OAI21X1_291 ( .A(_abc_40344_n1911), .B(_abc_40344_n761_1), .C(_abc_40344_n1912), .Y(_abc_40344_n1913) );
  OAI21X1 OAI21X1_292 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_31_), .Y(_abc_40344_n1916) );
  OAI21X1 OAI21X1_293 ( .A(_abc_40344_n1919), .B(_abc_40344_n761_1), .C(_abc_40344_n1920), .Y(_abc_40344_n1921) );
  OAI21X1 OAI21X1_294 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_30_), .Y(_abc_40344_n1922) );
  OAI21X1 OAI21X1_295 ( .A(_abc_40344_n1918), .B(_abc_40344_n1921), .C(_abc_40344_n1922), .Y(_abc_40344_n1923) );
  OAI21X1 OAI21X1_296 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_29_), .Y(_abc_40344_n1926) );
  OAI21X1 OAI21X1_297 ( .A(_abc_40344_n1931), .B(_abc_40344_n705_1), .C(_abc_40344_n1488), .Y(_abc_40344_n1932) );
  OAI21X1 OAI21X1_298 ( .A(_abc_40344_n1933), .B(_abc_40344_n705_1), .C(_abc_40344_n1471), .Y(_abc_40344_n1934) );
  OAI21X1 OAI21X1_299 ( .A(_abc_40344_n1462), .B(_abc_40344_n1471), .C(_abc_40344_n1935), .Y(_abc_40344_n1936) );
  OAI21X1 OAI21X1_3 ( .A(_abc_40344_n569_1), .B(_abc_40344_n578_1), .C(IR_REG_31_), .Y(_abc_40344_n579) );
  OAI21X1 OAI21X1_30 ( .A(_abc_40344_n687), .B(_abc_40344_n688_1), .C(_abc_40344_n736), .Y(_abc_40344_n737) );
  OAI21X1 OAI21X1_300 ( .A(_abc_40344_n1254_1), .B(_abc_40344_n1258), .C(_abc_40344_n1264), .Y(_abc_40344_n1938) );
  OAI21X1 OAI21X1_301 ( .A(_abc_40344_n1308), .B(_abc_40344_n1305), .C(_abc_40344_n1938), .Y(_abc_40344_n1939) );
  OAI21X1 OAI21X1_302 ( .A(_abc_40344_n1109), .B(_abc_40344_n1105), .C(_abc_40344_n1099), .Y(_abc_40344_n1943) );
  OAI21X1 OAI21X1_303 ( .A(_abc_40344_n1166_1), .B(_abc_40344_n1163), .C(_abc_40344_n1152_1), .Y(_abc_40344_n1947) );
  OAI21X1 OAI21X1_304 ( .A(_abc_40344_n1181), .B(_abc_40344_n1184), .C(_abc_40344_n1949), .Y(_abc_40344_n1950) );
  OAI21X1 OAI21X1_305 ( .A(_abc_40344_n1950), .B(_abc_40344_n1948), .C(_abc_40344_n1947), .Y(_abc_40344_n1951) );
  OAI21X1 OAI21X1_306 ( .A(_abc_40344_n1428), .B(_abc_40344_n1424), .C(_abc_40344_n1421_1), .Y(_abc_40344_n1953) );
  OAI21X1 OAI21X1_307 ( .A(_abc_40344_n1413), .B(_abc_40344_n1410), .C(_abc_40344_n1418), .Y(_abc_40344_n1956) );
  OAI21X1 OAI21X1_308 ( .A(_abc_40344_n1124), .B(_abc_40344_n1138), .C(_abc_40344_n1956), .Y(_abc_40344_n1957) );
  OAI21X1 OAI21X1_309 ( .A(_abc_40344_n1205), .B(_abc_40344_n1208), .C(_abc_40344_n1200), .Y(_abc_40344_n1962) );
  OAI21X1 OAI21X1_31 ( .A(_abc_40344_n561_1), .B(_abc_40344_n580), .C(_abc_40344_n744), .Y(_abc_40344_n745) );
  OAI21X1 OAI21X1_310 ( .A(DATAI_10_), .B(_abc_40344_n705_1), .C(_abc_40344_n1968), .Y(_abc_40344_n1969) );
  OAI21X1 OAI21X1_311 ( .A(_abc_40344_n1331_1), .B(_abc_40344_n1334), .C(_abc_40344_n1969), .Y(_abc_40344_n1970) );
  OAI21X1 OAI21X1_312 ( .A(DATAI_11_), .B(_abc_40344_n705_1), .C(_abc_40344_n1972), .Y(_abc_40344_n1973) );
  OAI21X1 OAI21X1_313 ( .A(_abc_40344_n1280), .B(_abc_40344_n1283), .C(_abc_40344_n1973), .Y(_abc_40344_n1974) );
  OAI21X1 OAI21X1_314 ( .A(_abc_40344_n1974), .B(_abc_40344_n1971), .C(_abc_40344_n1970), .Y(_abc_40344_n1975) );
  OAI21X1 OAI21X1_315 ( .A(_abc_40344_n1495), .B(_abc_40344_n1506), .C(_abc_40344_n1976), .Y(_abc_40344_n1977) );
  OAI21X1 OAI21X1_316 ( .A(_abc_40344_n1018), .B(_abc_40344_n1665), .C(_abc_40344_n1907), .Y(_abc_40344_n1983) );
  OAI21X1 OAI21X1_317 ( .A(_abc_40344_n923_1), .B(_abc_40344_n926), .C(_abc_40344_n919), .Y(_abc_40344_n1985) );
  OAI21X1 OAI21X1_318 ( .A(_abc_40344_n1989), .B(_abc_40344_n761_1), .C(_abc_40344_n1990), .Y(_abc_40344_n1991) );
  OAI21X1 OAI21X1_319 ( .A(DATAI_6_), .B(_abc_40344_n705_1), .C(_abc_40344_n1993), .Y(_abc_40344_n1994) );
  OAI21X1 OAI21X1_32 ( .A(_abc_40344_n626), .B(_abc_40344_n648), .C(_abc_40344_n640), .Y(_abc_40344_n746) );
  OAI21X1 OAI21X1_320 ( .A(_abc_40344_n1988), .B(_abc_40344_n1991), .C(_abc_40344_n1994), .Y(_abc_40344_n1995) );
  OAI21X1 OAI21X1_321 ( .A(_abc_40344_n698), .B(_abc_40344_n1994), .C(_abc_40344_n1998), .Y(_abc_40344_n1999) );
  OAI21X1 OAI21X1_322 ( .A(_abc_40344_n1505_1), .B(_abc_40344_n1498), .C(_abc_40344_n1494), .Y(_abc_40344_n2001) );
  OAI21X1 OAI21X1_323 ( .A(_abc_40344_n2009), .B(_abc_40344_n705_1), .C(_abc_40344_n1073), .Y(_abc_40344_n2010) );
  OAI21X1 OAI21X1_324 ( .A(_abc_40344_n2016), .B(_abc_40344_n2017), .C(_abc_40344_n1609), .Y(_abc_40344_n2018) );
  OAI21X1 OAI21X1_325 ( .A(_abc_40344_n777_1), .B(_abc_40344_n787_1), .C(_abc_40344_n2018), .Y(_abc_40344_n2019) );
  OAI21X1 OAI21X1_326 ( .A(DATAI_2_), .B(_abc_40344_n705_1), .C(_abc_40344_n2021), .Y(_abc_40344_n2022) );
  OAI21X1 OAI21X1_327 ( .A(_abc_40344_n1649), .B(_abc_40344_n1550), .C(_abc_40344_n2025), .Y(_abc_40344_n2026) );
  OAI21X1 OAI21X1_328 ( .A(_abc_40344_n2026), .B(_abc_40344_n2013), .C(_abc_40344_n2035), .Y(_abc_40344_n2036) );
  OAI21X1 OAI21X1_329 ( .A(_abc_40344_n1434), .B(_abc_40344_n1440), .C(_abc_40344_n2038), .Y(_abc_40344_n2039) );
  OAI21X1 OAI21X1_33 ( .A(_abc_40344_n746), .B(_abc_40344_n718), .C(_abc_40344_n716), .Y(_abc_40344_n747) );
  OAI21X1 OAI21X1_330 ( .A(_abc_40344_n1950), .B(_abc_40344_n1948), .C(_abc_40344_n2042), .Y(_abc_40344_n2043) );
  OAI21X1 OAI21X1_331 ( .A(_abc_40344_n2058), .B(_abc_40344_n2062), .C(_abc_40344_n1929), .Y(_abc_40344_n2063) );
  OAI21X1 OAI21X1_332 ( .A(_abc_40344_n2055), .B(_abc_40344_n2063), .C(_abc_40344_n2071), .Y(_abc_40344_n2072) );
  OAI21X1 OAI21X1_333 ( .A(_abc_40344_n1404), .B(_abc_40344_n1414), .C(_abc_40344_n1948), .Y(_abc_40344_n2073) );
  OAI21X1 OAI21X1_334 ( .A(_abc_40344_n2097), .B(_abc_40344_n2098), .C(_abc_40344_n1925), .Y(_abc_40344_n2099) );
  OAI21X1 OAI21X1_335 ( .A(_abc_40344_n1910), .B(_abc_40344_n1913), .C(_abc_40344_n1916), .Y(_abc_40344_n2100) );
  OAI21X1 OAI21X1_336 ( .A(_abc_40344_n1251), .B(_abc_40344_n1259), .C(_abc_40344_n1971), .Y(_abc_40344_n2111) );
  OAI21X1 OAI21X1_337 ( .A(_abc_40344_n2116), .B(_abc_40344_n2119), .C(_abc_40344_n2117), .Y(_abc_40344_n2120) );
  OAI21X1 OAI21X1_338 ( .A(_abc_40344_n1974), .B(_abc_40344_n1971), .C(_abc_40344_n2125), .Y(_abc_40344_n2126) );
  OAI21X1 OAI21X1_339 ( .A(_abc_40344_n838), .B(_abc_40344_n840), .C(_abc_40344_n2022), .Y(_abc_40344_n2134) );
  OAI21X1 OAI21X1_34 ( .A(DATAI_5_), .B(_abc_40344_n705_1), .C(_abc_40344_n749_1), .Y(_abc_40344_n750) );
  OAI21X1 OAI21X1_340 ( .A(_abc_40344_n859), .B(_abc_40344_n862), .C(_abc_40344_n869), .Y(_abc_40344_n2142) );
  OAI21X1 OAI21X1_341 ( .A(_abc_40344_n625), .B(_abc_40344_n646), .C(_abc_40344_n619), .Y(_abc_40344_n2143) );
  OAI21X1 OAI21X1_342 ( .A(_abc_40344_n879), .B(_abc_40344_n2143), .C(_abc_40344_n2142), .Y(_abc_40344_n2144) );
  OAI21X1 OAI21X1_343 ( .A(_abc_40344_n2146), .B(_abc_40344_n1797), .C(_abc_40344_n887), .Y(_abc_40344_n2147) );
  OAI21X1 OAI21X1_344 ( .A(_abc_40344_n619), .B(_abc_40344_n626), .C(_abc_40344_n2157), .Y(_abc_40344_n2158) );
  OAI21X1 OAI21X1_345 ( .A(_abc_40344_n626), .B(_abc_40344_n641), .C(_abc_40344_n585), .Y(_abc_40344_n2172) );
  OAI21X1 OAI21X1_346 ( .A(_abc_40344_n2161), .B(_abc_40344_n1994), .C(_abc_40344_n2182), .Y(_abc_40344_n2183) );
  OAI21X1 OAI21X1_347 ( .A(_abc_40344_n2161), .B(_abc_40344_n750), .C(_abc_40344_n2185), .Y(_abc_40344_n2186) );
  OAI21X1 OAI21X1_348 ( .A(_abc_40344_n742), .B(_abc_40344_n2172), .C(_abc_40344_n2188), .Y(_abc_40344_n2189) );
  OAI21X1 OAI21X1_349 ( .A(_abc_40344_n2161), .B(_abc_40344_n776), .C(_abc_40344_n2171), .Y(_abc_40344_n2191) );
  OAI21X1 OAI21X1_35 ( .A(_abc_40344_n751_1), .B(_abc_40344_n754_1), .C(_abc_40344_n740), .Y(_abc_40344_n755) );
  OAI21X1 OAI21X1_350 ( .A(_abc_40344_n785), .B(_abc_40344_n2172), .C(_abc_40344_n2177), .Y(_abc_40344_n2192) );
  OAI21X1 OAI21X1_351 ( .A(_abc_40344_n2161), .B(_abc_40344_n919), .C(_abc_40344_n2193), .Y(_abc_40344_n2194) );
  OAI21X1 OAI21X1_352 ( .A(_abc_40344_n2016), .B(_abc_40344_n2017), .C(_abc_40344_n586), .Y(_abc_40344_n2200) );
  OAI21X1 OAI21X1_353 ( .A(_abc_40344_n921), .B(_abc_40344_n2201), .C(_abc_40344_n783), .Y(_abc_40344_n2202) );
  OAI21X1 OAI21X1_354 ( .A(_abc_40344_n2203), .B(_abc_40344_n759), .C(_abc_40344_n784), .Y(_abc_40344_n2204) );
  OAI21X1 OAI21X1_355 ( .A(_abc_40344_n2202), .B(_abc_40344_n2204), .C(_abc_40344_n2165), .Y(_abc_40344_n2205) );
  OAI21X1 OAI21X1_356 ( .A(_abc_40344_n2210), .B(_abc_40344_n2198), .C(_abc_40344_n2209), .Y(_abc_40344_n2211) );
  OAI21X1 OAI21X1_357 ( .A(_abc_40344_n859), .B(_abc_40344_n862), .C(_abc_40344_n586), .Y(_abc_40344_n2212) );
  OAI21X1 OAI21X1_358 ( .A(_abc_40344_n838), .B(_abc_40344_n840), .C(_abc_40344_n2165), .Y(_abc_40344_n2213) );
  OAI21X1 OAI21X1_359 ( .A(_abc_40344_n886), .B(_abc_40344_n883), .C(_abc_40344_n586), .Y(_abc_40344_n2217) );
  OAI21X1 OAI21X1_36 ( .A(IR_REG_31_), .B(_abc_40344_n662), .C(_abc_40344_n674_1), .Y(_abc_40344_n758) );
  OAI21X1 OAI21X1_360 ( .A(_abc_40344_n859), .B(_abc_40344_n862), .C(_abc_40344_n2165), .Y(_abc_40344_n2218) );
  OAI21X1 OAI21X1_361 ( .A(_abc_40344_n2161), .B(_abc_40344_n869), .C(_abc_40344_n2219), .Y(_abc_40344_n2220) );
  OAI21X1 OAI21X1_362 ( .A(_abc_40344_n2172), .B(_abc_40344_n2223), .C(_abc_40344_n2224), .Y(_abc_40344_n2225) );
  OAI21X1 OAI21X1_363 ( .A(_abc_40344_n2221), .B(_abc_40344_n2220), .C(_abc_40344_n2225), .Y(_abc_40344_n2226) );
  OAI21X1 OAI21X1_364 ( .A(_abc_40344_n2161), .B(_abc_40344_n2022), .C(_abc_40344_n2227), .Y(_abc_40344_n2228) );
  OAI21X1 OAI21X1_365 ( .A(_abc_40344_n2211), .B(_abc_40344_n2231), .C(_abc_40344_n2197), .Y(_abc_40344_n2232) );
  OAI21X1 OAI21X1_366 ( .A(_abc_40344_n1988), .B(_abc_40344_n1991), .C(_abc_40344_n586), .Y(_abc_40344_n2233) );
  OAI21X1 OAI21X1_367 ( .A(_abc_40344_n2179), .B(_abc_40344_n927_1), .C(_abc_40344_n2233), .Y(_abc_40344_n2234) );
  OAI21X1 OAI21X1_368 ( .A(_abc_40344_n1353), .B(_abc_40344_n1360), .C(_abc_40344_n586), .Y(_abc_40344_n2238) );
  OAI21X1 OAI21X1_369 ( .A(_abc_40344_n1331_1), .B(_abc_40344_n1334), .C(_abc_40344_n2165), .Y(_abc_40344_n2239) );
  OAI21X1 OAI21X1_37 ( .A(_abc_40344_n667), .B(_abc_40344_n753), .C(_abc_40344_n758), .Y(_abc_40344_n759) );
  OAI21X1 OAI21X1_370 ( .A(_abc_40344_n1009), .B(_abc_40344_n1017), .C(_abc_40344_n586), .Y(_abc_40344_n2243) );
  OAI21X1 OAI21X1_371 ( .A(_abc_40344_n1353), .B(_abc_40344_n1360), .C(_abc_40344_n2165), .Y(_abc_40344_n2244) );
  OAI21X1 OAI21X1_372 ( .A(_abc_40344_n926), .B(_abc_40344_n923_1), .C(_abc_40344_n586), .Y(_abc_40344_n2249) );
  OAI21X1 OAI21X1_373 ( .A(_abc_40344_n2179), .B(_abc_40344_n1018), .C(_abc_40344_n2249), .Y(_abc_40344_n2250) );
  OAI21X1 OAI21X1_374 ( .A(_abc_40344_n2184), .B(_abc_40344_n2183), .C(_abc_40344_n2258), .Y(_abc_40344_n2259) );
  OAI21X1 OAI21X1_375 ( .A(_abc_40344_n2291), .B(_abc_40344_n2290), .C(_abc_40344_n2292), .Y(_abc_40344_n2293) );
  OAI21X1 OAI21X1_376 ( .A(_abc_40344_n2161), .B(_abc_40344_n1961), .C(_abc_40344_n2294), .Y(_abc_40344_n2295) );
  OAI21X1 OAI21X1_377 ( .A(_abc_40344_n2277_1), .B(_abc_40344_n2293), .C(_abc_40344_n2297), .Y(_abc_40344_n2298) );
  OAI21X1 OAI21X1_378 ( .A(_abc_40344_n2299), .B(_abc_40344_n2287), .C(_abc_40344_n2307), .Y(_abc_40344_n2308_1) );
  OAI21X1 OAI21X1_379 ( .A(_abc_40344_n2327), .B(_abc_40344_n2322), .C(_abc_40344_n2334), .Y(_abc_40344_n2335) );
  OAI21X1 OAI21X1_38 ( .A(_abc_40344_n651_1), .B(_abc_40344_n752), .C(_abc_40344_n760), .Y(_abc_40344_n761_1) );
  OAI21X1 OAI21X1_380 ( .A(_abc_40344_n585), .B(_abc_40344_n1429), .C(_abc_40344_n2344), .Y(_abc_40344_n2345) );
  OAI21X1 OAI21X1_381 ( .A(_abc_40344_n2343), .B(_abc_40344_n2345), .C(_abc_40344_n2341), .Y(_abc_40344_n2346) );
  OAI21X1 OAI21X1_382 ( .A(_abc_40344_n1109), .B(_abc_40344_n1105), .C(_abc_40344_n2165), .Y(_abc_40344_n2348) );
  OAI21X1 OAI21X1_383 ( .A(_abc_40344_n626), .B(_abc_40344_n641), .C(_abc_40344_n1100), .Y(_abc_40344_n2349) );
  OAI21X1 OAI21X1_384 ( .A(_abc_40344_n2351), .B(_abc_40344_n2353), .C(_abc_40344_n2360), .Y(_abc_40344_n2361) );
  OAI21X1 OAI21X1_385 ( .A(_abc_40344_n2355), .B(_abc_40344_n2347), .C(_abc_40344_n2362_1), .Y(_abc_40344_n2363) );
  OAI21X1 OAI21X1_386 ( .A(_abc_40344_n2179), .B(_abc_40344_n1577), .C(_abc_40344_n2364), .Y(_abc_40344_n2365) );
  OAI21X1 OAI21X1_387 ( .A(_abc_40344_n2179), .B(_abc_40344_n1489), .C(_abc_40344_n2370), .Y(_abc_40344_n2371) );
  OAI21X1 OAI21X1_388 ( .A(_abc_40344_n2372), .B(_abc_40344_n2371), .C(_abc_40344_n2373), .Y(_abc_40344_n2374) );
  OAI21X1 OAI21X1_389 ( .A(_abc_40344_n1506), .B(_abc_40344_n2179), .C(_abc_40344_n2376), .Y(_abc_40344_n2377) );
  OAI21X1 OAI21X1_39 ( .A(IR_REG_3_), .B(_abc_40344_n539), .C(IR_REG_4_), .Y(_abc_40344_n770) );
  OAI21X1 OAI21X1_390 ( .A(_abc_40344_n585), .B(_abc_40344_n1506), .C(_abc_40344_n2384), .Y(_abc_40344_n2385) );
  OAI21X1 OAI21X1_391 ( .A(_abc_40344_n2381), .B(_abc_40344_n2375), .C(_abc_40344_n2387), .Y(_abc_40344_n2388) );
  OAI21X1 OAI21X1_392 ( .A(_abc_40344_n2179), .B(_abc_40344_n1550), .C(_abc_40344_n2389_1), .Y(_abc_40344_n2390) );
  OAI21X1 OAI21X1_393 ( .A(_abc_40344_n585), .B(_abc_40344_n1550), .C(_abc_40344_n2395), .Y(_abc_40344_n2396) );
  OAI21X1 OAI21X1_394 ( .A(_abc_40344_n640), .B(_abc_40344_n1914), .C(_abc_40344_n625), .Y(_abc_40344_n2404) );
  OAI21X1 OAI21X1_395 ( .A(_abc_40344_n2407), .B(_abc_40344_n2400), .C(_abc_40344_n2411), .Y(_abc_40344_n2412) );
  OAI21X1 OAI21X1_396 ( .A(_abc_40344_n755), .B(_abc_40344_n762), .C(_abc_40344_n586), .Y(_abc_40344_n2418) );
  OAI21X1 OAI21X1_397 ( .A(_abc_40344_n1988), .B(_abc_40344_n1991), .C(_abc_40344_n2165), .Y(_abc_40344_n2419) );
  OAI21X1 OAI21X1_398 ( .A(_abc_40344_n2436), .B(_abc_40344_n2437), .C(_abc_40344_n2431), .Y(_abc_40344_n2438) );
  OAI21X1 OAI21X1_399 ( .A(_abc_40344_n2445), .B(_abc_40344_n2439), .C(_abc_40344_n2448), .Y(_abc_40344_n2449) );
  OAI21X1 OAI21X1_4 ( .A(IR_REG_22_), .B(_abc_40344_n576), .C(IR_REG_23_), .Y(_abc_40344_n582) );
  OAI21X1 OAI21X1_40 ( .A(_abc_40344_n559_1), .B(_abc_40344_n771), .C(_abc_40344_n772), .Y(_abc_40344_n773) );
  OAI21X1 OAI21X1_400 ( .A(_abc_40344_n2452), .B(_abc_40344_n2451_1), .C(_abc_40344_n2320), .Y(_abc_40344_n2453) );
  OAI21X1 OAI21X1_401 ( .A(_abc_40344_n2339), .B(_abc_40344_n2456), .C(_abc_40344_n2457), .Y(_abc_40344_n2458_1) );
  OAI21X1 OAI21X1_402 ( .A(_abc_40344_n2368), .B(_abc_40344_n2459), .C(_abc_40344_n2460), .Y(_abc_40344_n2461) );
  OAI21X1 OAI21X1_403 ( .A(_abc_40344_n2463), .B(_abc_40344_n2462), .C(_abc_40344_n2464), .Y(_abc_40344_n2465) );
  OAI21X1 OAI21X1_404 ( .A(_abc_40344_n2467), .B(_abc_40344_n2466), .C(_abc_40344_n627), .Y(_abc_40344_n2468) );
  OAI21X1 OAI21X1_405 ( .A(_abc_40344_n1230), .B(_abc_40344_n1233), .C(_abc_40344_n1961), .Y(_abc_40344_n2479) );
  OAI21X1 OAI21X1_406 ( .A(_abc_40344_n2095), .B(_abc_40344_n2401), .C(_abc_40344_n2408_1), .Y(_abc_40344_n2504) );
  OAI21X1 OAI21X1_407 ( .A(_abc_40344_n2500), .B(_abc_40344_n2501), .C(_abc_40344_n2505), .Y(_abc_40344_n2506) );
  OAI21X1 OAI21X1_408 ( .A(_abc_40344_n1933), .B(_abc_40344_n705_1), .C(_abc_40344_n1577), .Y(_abc_40344_n2518) );
  OAI21X1 OAI21X1_409 ( .A(_abc_40344_n883), .B(_abc_40344_n886), .C(_abc_40344_n1797), .Y(_abc_40344_n2528) );
  OAI21X1 OAI21X1_41 ( .A(DATAI_4_), .B(_abc_40344_n705_1), .C(_abc_40344_n775_1), .Y(_abc_40344_n776) );
  OAI21X1 OAI21X1_410 ( .A(_abc_40344_n1009), .B(_abc_40344_n1017), .C(_abc_40344_n1375), .Y(_abc_40344_n2530) );
  OAI21X1 OAI21X1_411 ( .A(_abc_40344_n1181), .B(_abc_40344_n1184), .C(_abc_40344_n1178), .Y(_abc_40344_n2541) );
  OAI21X1 OAI21X1_412 ( .A(_abc_40344_n1495), .B(_abc_40344_n1506), .C(_abc_40344_n2010), .Y(_abc_40344_n2565) );
  OAI21X1 OAI21X1_413 ( .A(_abc_40344_n1914), .B(_abc_40344_n1924), .C(_abc_40344_n2566), .Y(_abc_40344_n2567_1) );
  OAI21X1 OAI21X1_414 ( .A(_abc_40344_n1910), .B(_abc_40344_n1913), .C(_abc_40344_n2096), .Y(_abc_40344_n2568) );
  OAI21X1 OAI21X1_415 ( .A(_abc_40344_n2570), .B(_abc_40344_n1927), .C(_abc_40344_n2567_1), .Y(_abc_40344_n2571) );
  OAI21X1 OAI21X1_416 ( .A(_abc_40344_n2573_1), .B(_abc_40344_n705_1), .C(_abc_40344_n2574), .Y(_abc_40344_n2575) );
  OAI21X1 OAI21X1_417 ( .A(_abc_40344_n1550), .B(_abc_40344_n2575), .C(_abc_40344_n2572), .Y(_abc_40344_n2576) );
  OAI21X1 OAI21X1_418 ( .A(_abc_40344_n1542), .B(_abc_40344_n1549), .C(_abc_40344_n2578), .Y(_abc_40344_n2579) );
  OAI21X1 OAI21X1_419 ( .A(_abc_40344_n2577), .B(_abc_40344_n2575), .C(_abc_40344_n2579), .Y(_abc_40344_n2580) );
  OAI21X1 OAI21X1_42 ( .A(_abc_40344_n561_1), .B(_abc_40344_n580), .C(_abc_40344_n746), .Y(_abc_40344_n792) );
  OAI21X1 OAI21X1_420 ( .A(_abc_40344_n2577), .B(_abc_40344_n2575), .C(_abc_40344_n1550), .Y(_abc_40344_n2585) );
  OAI21X1 OAI21X1_421 ( .A(_abc_40344_n1945), .B(_abc_40344_n2002), .C(_abc_40344_n1942), .Y(_abc_40344_n2587) );
  OAI21X1 OAI21X1_422 ( .A(_abc_40344_n1421_1), .B(_abc_40344_n2037), .C(_abc_40344_n2064), .Y(_abc_40344_n2590) );
  OAI21X1 OAI21X1_423 ( .A(_abc_40344_n1434), .B(_abc_40344_n1440), .C(_abc_40344_n1943), .Y(_abc_40344_n2594) );
  OAI21X1 OAI21X1_424 ( .A(_abc_40344_n1939), .B(_abc_40344_n2122), .C(_abc_40344_n2111), .Y(_abc_40344_n2601) );
  OAI21X1 OAI21X1_425 ( .A(_abc_40344_n2479), .B(_abc_40344_n2604), .C(_abc_40344_n1958), .Y(_abc_40344_n2605) );
  OAI21X1 OAI21X1_426 ( .A(_abc_40344_n1962), .B(_abc_40344_n2042), .C(_abc_40344_n1947), .Y(_abc_40344_n2606) );
  OAI21X1 OAI21X1_427 ( .A(_abc_40344_n2605), .B(_abc_40344_n2606), .C(_abc_40344_n2593_1), .Y(_abc_40344_n2607) );
  OAI21X1 OAI21X1_428 ( .A(_abc_40344_n908), .B(_abc_40344_n927_1), .C(_abc_40344_n1995), .Y(_abc_40344_n2610) );
  OAI21X1 OAI21X1_429 ( .A(_abc_40344_n1998), .B(_abc_40344_n2088), .C(_abc_40344_n2083), .Y(_abc_40344_n2611) );
  OAI21X1 OAI21X1_43 ( .A(_abc_40344_n561_1), .B(_abc_40344_n580), .C(_abc_40344_n718), .Y(_abc_40344_n793) );
  OAI21X1 OAI21X1_430 ( .A(_abc_40344_n919), .B(_abc_40344_n915_1), .C(_abc_40344_n2531), .Y(_abc_40344_n2614) );
  OAI21X1 OAI21X1_431 ( .A(_abc_40344_n2610), .B(_abc_40344_n2612), .C(_abc_40344_n2615), .Y(_abc_40344_n2616) );
  OAI21X1 OAI21X1_432 ( .A(_abc_40344_n1273), .B(_abc_40344_n1284), .C(_abc_40344_n2616), .Y(_abc_40344_n2617) );
  OAI21X1 OAI21X1_433 ( .A(_abc_40344_n2613), .B(_abc_40344_n1984), .C(_abc_40344_n1970), .Y(_abc_40344_n2619_1) );
  OAI21X1 OAI21X1_434 ( .A(_abc_40344_n1609), .B(_abc_40344_n808), .C(_abc_40344_n2626), .Y(_abc_40344_n2627) );
  OAI21X1 OAI21X1_435 ( .A(_abc_40344_n2134), .B(_abc_40344_n2627), .C(_abc_40344_n2629), .Y(_abc_40344_n2630) );
  OAI21X1 OAI21X1_436 ( .A(_abc_40344_n856), .B(_abc_40344_n863), .C(_abc_40344_n2631), .Y(_abc_40344_n2632) );
  OAI21X1 OAI21X1_437 ( .A(_abc_40344_n2630), .B(_abc_40344_n2634), .C(_abc_40344_n2623), .Y(_abc_40344_n2635) );
  OAI21X1 OAI21X1_438 ( .A(_abc_40344_n2636), .B(_abc_40344_n2622), .C(_abc_40344_n2588), .Y(_abc_40344_n2637) );
  OAI21X1 OAI21X1_439 ( .A(_abc_40344_n1040), .B(_abc_40344_n1073), .C(_abc_40344_n2583), .Y(_abc_40344_n2648) );
  OAI21X1 OAI21X1_44 ( .A(_abc_40344_n559_1), .B(_abc_40344_n795), .C(_abc_40344_n796), .Y(_abc_40344_n797) );
  OAI21X1 OAI21X1_440 ( .A(_abc_40344_n2513), .B(_abc_40344_n2647), .C(_abc_40344_n2649), .Y(_abc_40344_n2650_1) );
  OAI21X1 OAI21X1_441 ( .A(_abc_40344_n1040), .B(_abc_40344_n1073), .C(_abc_40344_n2565), .Y(_abc_40344_n2651) );
  OAI21X1 OAI21X1_442 ( .A(_abc_40344_n1550), .B(_abc_40344_n1649), .C(_abc_40344_n2651), .Y(_abc_40344_n2652) );
  OAI21X1 OAI21X1_443 ( .A(_abc_40344_n1630), .B(_abc_40344_n2391), .C(_abc_40344_n2574), .Y(_abc_40344_n2654) );
  OAI21X1 OAI21X1_444 ( .A(_abc_40344_n618), .B(_abc_40344_n625), .C(_abc_40344_n1026), .Y(_abc_40344_n2659) );
  OAI21X1 OAI21X1_445 ( .A(_abc_40344_n2659), .B(_abc_40344_n2157), .C(_abc_40344_n2658), .Y(_abc_40344_n2660) );
  OAI21X1 OAI21X1_446 ( .A(_abc_40344_n1029_1), .B(_abc_40344_n2564), .C(_abc_40344_n2661), .Y(_abc_40344_n2662) );
  OAI21X1 OAI21X1_447 ( .A(_abc_40344_n2667), .B(_abc_40344_n1004), .C(_abc_40344_n586), .Y(_abc_40344_n2668) );
  OAI21X1 OAI21X1_448 ( .A(_abc_40344_n2665), .B(_abc_40344_n2663), .C(_abc_40344_n2671), .Y(n1186) );
  OAI21X1 OAI21X1_449 ( .A(_abc_40344_n716), .B(_abc_40344_n585), .C(_abc_40344_n2673), .Y(_abc_40344_n2674) );
  OAI21X1 OAI21X1_45 ( .A(_abc_40344_n810), .B(_abc_40344_n804), .C(_abc_40344_n720), .Y(_abc_40344_n811) );
  OAI21X1 OAI21X1_450 ( .A(_abc_40344_n538_1), .B(_abc_40344_n885), .C(_abc_40344_n610_1), .Y(_abc_40344_n2678) );
  OAI21X1 OAI21X1_451 ( .A(IR_REG_0_), .B(REG2_REG_0_), .C(_abc_40344_n2666_1), .Y(_abc_40344_n2682) );
  OAI21X1 OAI21X1_452 ( .A(REG2_REG_1_), .B(_abc_40344_n2688), .C(_abc_40344_n2690), .Y(_abc_40344_n2691) );
  OAI21X1 OAI21X1_453 ( .A(REG2_REG_1_), .B(_abc_40344_n2690), .C(_abc_40344_n2691), .Y(_abc_40344_n2692_1) );
  OAI21X1 OAI21X1_454 ( .A(_abc_40344_n2699), .B(_abc_40344_n2700), .C(_abc_40344_n610_1), .Y(_abc_40344_n2701) );
  OAI21X1 OAI21X1_455 ( .A(_abc_40344_n853), .B(_abc_40344_n603), .C(_abc_40344_n2701), .Y(_abc_40344_n2702) );
  OAI21X1 OAI21X1_456 ( .A(_abc_40344_n2673), .B(_abc_40344_n2665), .C(_abc_40344_n2704), .Y(_abc_40344_n2705) );
  OAI21X1 OAI21X1_457 ( .A(_abc_40344_n2703), .B(_abc_40344_n2706), .C(_abc_40344_n2687), .Y(n1050) );
  OAI21X1 OAI21X1_458 ( .A(_abc_40344_n2683), .B(_abc_40344_n2709), .C(n1345), .Y(_abc_40344_n2710) );
  OAI21X1 OAI21X1_459 ( .A(_abc_40344_n2713), .B(_abc_40344_n2714), .C(_abc_40344_n2691), .Y(_abc_40344_n2715) );
  OAI21X1 OAI21X1_46 ( .A(_abc_40344_n812), .B(_abc_40344_n705_1), .C(_abc_40344_n798), .Y(_abc_40344_n813) );
  OAI21X1 OAI21X1_460 ( .A(_abc_40344_n2712), .B(_abc_40344_n2020), .C(_abc_40344_n2716), .Y(_abc_40344_n2717) );
  OAI21X1 OAI21X1_461 ( .A(_abc_40344_n2697), .B(_abc_40344_n853), .C(_abc_40344_n2695), .Y(_abc_40344_n2721) );
  OAI21X1 OAI21X1_462 ( .A(_abc_40344_n2020), .B(_abc_40344_n603), .C(_abc_40344_n2723), .Y(_abc_40344_n2724) );
  OAI21X1 OAI21X1_463 ( .A(_abc_40344_n2719), .B(_abc_40344_n2724), .C(_abc_40344_n2705), .Y(_abc_40344_n2725) );
  OAI21X1 OAI21X1_464 ( .A(REG1_REG_2_), .B(_abc_40344_n823), .C(_abc_40344_n2721), .Y(_abc_40344_n2734) );
  OAI21X1 OAI21X1_465 ( .A(_abc_40344_n836), .B(_abc_40344_n2020), .C(_abc_40344_n2734), .Y(_abc_40344_n2735) );
  OAI21X1 OAI21X1_466 ( .A(_abc_40344_n2741), .B(_abc_40344_n2740), .C(_abc_40344_n610_1), .Y(_abc_40344_n2742) );
  OAI21X1 OAI21X1_467 ( .A(_abc_40344_n603), .B(_abc_40344_n1607), .C(_abc_40344_n2742), .Y(_abc_40344_n2743) );
  OAI21X1 OAI21X1_468 ( .A(_abc_40344_n2744), .B(_abc_40344_n2706), .C(_abc_40344_n2727), .Y(n1042) );
  OAI21X1 OAI21X1_469 ( .A(_abc_40344_n1607), .B(_abc_40344_n2737), .C(_abc_40344_n2736), .Y(_abc_40344_n2747) );
  OAI21X1 OAI21X1_47 ( .A(IR_REG_1_), .B(IR_REG_0_), .C(IR_REG_2_), .Y(_abc_40344_n820) );
  OAI21X1 OAI21X1_470 ( .A(_abc_40344_n2749), .B(_abc_40344_n2747), .C(_abc_40344_n610_1), .Y(_abc_40344_n2750) );
  OAI21X1 OAI21X1_471 ( .A(_abc_40344_n2728), .B(_abc_40344_n2732), .C(_abc_40344_n2730_1), .Y(_abc_40344_n2755) );
  OAI21X1 OAI21X1_472 ( .A(_abc_40344_n2751), .B(_abc_40344_n2757), .C(_abc_40344_n2705), .Y(_abc_40344_n2758) );
  OAI21X1 OAI21X1_473 ( .A(REG1_REG_4_), .B(_abc_40344_n773), .C(_abc_40344_n2747), .Y(_abc_40344_n2761) );
  OAI21X1 OAI21X1_474 ( .A(_abc_40344_n2748), .B(_abc_40344_n774), .C(_abc_40344_n2761), .Y(_abc_40344_n2762) );
  OAI21X1 OAI21X1_475 ( .A(_abc_40344_n748), .B(_abc_40344_n2763), .C(_abc_40344_n610_1), .Y(_abc_40344_n2764) );
  OAI21X1 OAI21X1_476 ( .A(REG2_REG_4_), .B(_abc_40344_n773), .C(_abc_40344_n2755), .Y(_abc_40344_n2767) );
  OAI21X1 OAI21X1_477 ( .A(_abc_40344_n2766), .B(_abc_40344_n2768_1), .C(_abc_40344_n2769), .Y(_abc_40344_n2770) );
  OAI21X1 OAI21X1_478 ( .A(_abc_40344_n603), .B(_abc_40344_n748), .C(_abc_40344_n2770), .Y(_abc_40344_n2771) );
  OAI21X1 OAI21X1_479 ( .A(_abc_40344_n2771), .B(_abc_40344_n2765), .C(_abc_40344_n2705), .Y(_abc_40344_n2772) );
  OAI21X1 OAI21X1_48 ( .A(_abc_40344_n559_1), .B(_abc_40344_n821), .C(_abc_40344_n822), .Y(_abc_40344_n823) );
  OAI21X1 OAI21X1_480 ( .A(REG1_REG_5_), .B(_abc_40344_n2762), .C(_abc_40344_n732_1), .Y(_abc_40344_n2777) );
  OAI21X1 OAI21X1_481 ( .A(_abc_40344_n756), .B(_abc_40344_n748), .C(_abc_40344_n2768_1), .Y(_abc_40344_n2787) );
  OAI21X1 OAI21X1_482 ( .A(REG2_REG_5_), .B(_abc_40344_n732_1), .C(_abc_40344_n2787), .Y(_abc_40344_n2788) );
  OAI21X1 OAI21X1_483 ( .A(_abc_40344_n611_1), .B(_abc_40344_n2782), .C(_abc_40344_n2790), .Y(_abc_40344_n2791) );
  OAI21X1 OAI21X1_484 ( .A(_abc_40344_n2774), .B(_abc_40344_n2793), .C(_abc_40344_n2775), .Y(n1030) );
  OAI21X1 OAI21X1_485 ( .A(REG1_REG_6_), .B(_abc_40344_n712), .C(_abc_40344_n2796), .Y(_abc_40344_n2797) );
  OAI21X1 OAI21X1_486 ( .A(_abc_40344_n2783), .B(_abc_40344_n2788), .C(_abc_40344_n2785), .Y(_abc_40344_n2804) );
  OAI21X1 OAI21X1_487 ( .A(REG2_REG_7_), .B(_abc_40344_n906_1), .C(_abc_40344_n2804), .Y(_abc_40344_n2807) );
  OAI21X1 OAI21X1_488 ( .A(_abc_40344_n2802), .B(_abc_40344_n2807), .C(_abc_40344_n2666_1), .Y(_abc_40344_n2808) );
  OAI21X1 OAI21X1_489 ( .A(_abc_40344_n2706), .B(_abc_40344_n2810), .C(_abc_40344_n2795), .Y(n1026) );
  OAI21X1 OAI21X1_49 ( .A(_abc_40344_n819), .B(_abc_40344_n705_1), .C(_abc_40344_n824_1), .Y(_abc_40344_n825) );
  OAI21X1 OAI21X1_490 ( .A(_abc_40344_n2677), .B(_abc_40344_n2684), .C(_abc_40344_n610_1), .Y(_abc_40344_n2817) );
  OAI21X1 OAI21X1_491 ( .A(_abc_40344_n1372), .B(_abc_40344_n2816_1), .C(_abc_40344_n2818), .Y(_abc_40344_n2819) );
  OAI21X1 OAI21X1_492 ( .A(_abc_40344_n2706), .B(_abc_40344_n2825), .C(_abc_40344_n2821), .Y(_abc_40344_n2826) );
  OAI21X1 OAI21X1_493 ( .A(_abc_40344_n1010), .B(_abc_40344_n1373), .C(_abc_40344_n2823_1), .Y(_abc_40344_n2830) );
  OAI21X1 OAI21X1_494 ( .A(REG2_REG_8_), .B(_abc_40344_n1372), .C(_abc_40344_n2830), .Y(_abc_40344_n2831) );
  OAI21X1 OAI21X1_495 ( .A(_abc_40344_n2829), .B(_abc_40344_n2831), .C(_abc_40344_n2666_1), .Y(_abc_40344_n2832) );
  OAI21X1 OAI21X1_496 ( .A(_abc_40344_n611_1), .B(_abc_40344_n2839), .C(_abc_40344_n2834), .Y(_abc_40344_n2840) );
  OAI21X1 OAI21X1_497 ( .A(_abc_40344_n2828), .B(_abc_40344_n2674), .C(_abc_40344_n2841), .Y(n1018) );
  OAI21X1 OAI21X1_498 ( .A(_abc_40344_n2844), .B(_abc_40344_n2838), .C(_abc_40344_n2835), .Y(_abc_40344_n2845) );
  OAI21X1 OAI21X1_499 ( .A(_abc_40344_n2849), .B(_abc_40344_n2847), .C(_abc_40344_n1325), .Y(_abc_40344_n2850) );
  OAI21X1 OAI21X1_5 ( .A(_abc_40344_n576), .B(_abc_40344_n555), .C(_abc_40344_n582), .Y(_abc_40344_n583) );
  OAI21X1 OAI21X1_50 ( .A(_abc_40344_n842), .B(_abc_40344_n835_1), .C(_abc_40344_n720), .Y(_abc_40344_n843) );
  OAI21X1 OAI21X1_500 ( .A(_abc_40344_n2847), .B(_abc_40344_n2851), .C(_abc_40344_n2850), .Y(_abc_40344_n2852) );
  OAI21X1 OAI21X1_501 ( .A(_abc_40344_n1354), .B(_abc_40344_n1347), .C(_abc_40344_n2831), .Y(_abc_40344_n2857) );
  OAI21X1 OAI21X1_502 ( .A(REG2_REG_9_), .B(_abc_40344_n1348), .C(_abc_40344_n2857), .Y(_abc_40344_n2858) );
  OAI21X1 OAI21X1_503 ( .A(_abc_40344_n2706), .B(_abc_40344_n2861), .C(_abc_40344_n2843), .Y(n1014) );
  OAI21X1 OAI21X1_504 ( .A(REG1_REG_10_), .B(_abc_40344_n2845), .C(_abc_40344_n2851), .Y(_abc_40344_n2868) );
  OAI21X1 OAI21X1_505 ( .A(_abc_40344_n2677), .B(_abc_40344_n2684), .C(_abc_40344_n2666_1), .Y(_abc_40344_n2870) );
  OAI21X1 OAI21X1_506 ( .A(_abc_40344_n2854), .B(_abc_40344_n2858), .C(_abc_40344_n2853), .Y(_abc_40344_n2875) );
  OAI21X1 OAI21X1_507 ( .A(_abc_40344_n2677), .B(_abc_40344_n2684), .C(_abc_40344_n602), .Y(_abc_40344_n2878) );
  OAI21X1 OAI21X1_508 ( .A(_abc_40344_n1271), .B(_abc_40344_n2878), .C(_abc_40344_n2877), .Y(_abc_40344_n2879) );
  OAI21X1 OAI21X1_509 ( .A(_abc_40344_n2817), .B(_abc_40344_n2869), .C(_abc_40344_n2880), .Y(n1010) );
  OAI21X1 OAI21X1_51 ( .A(IR_REG_1_), .B(IR_REG_0_), .C(IR_REG_31_), .Y(_abc_40344_n849_1) );
  OAI21X1 OAI21X1_510 ( .A(REG1_REG_10_), .B(_abc_40344_n2845), .C(_abc_40344_n1325), .Y(_abc_40344_n2886) );
  OAI21X1 OAI21X1_511 ( .A(REG1_REG_11_), .B(_abc_40344_n2863), .C(_abc_40344_n2887), .Y(_abc_40344_n2888) );
  OAI21X1 OAI21X1_512 ( .A(REG2_REG_11_), .B(_abc_40344_n2863), .C(_abc_40344_n2875), .Y(_abc_40344_n2894) );
  OAI21X1 OAI21X1_513 ( .A(_abc_40344_n1274), .B(_abc_40344_n1271), .C(_abc_40344_n2894), .Y(_abc_40344_n2895) );
  OAI21X1 OAI21X1_514 ( .A(_abc_40344_n2817), .B(_abc_40344_n2889), .C(_abc_40344_n2902), .Y(n1006) );
  OAI21X1 OAI21X1_515 ( .A(_abc_40344_n1296), .B(_abc_40344_n1293_1), .C(_abc_40344_n2904), .Y(_abc_40344_n2905) );
  OAI21X1 OAI21X1_516 ( .A(REG2_REG_12_), .B(_abc_40344_n2883), .C(_abc_40344_n2915), .Y(_abc_40344_n2916) );
  OAI21X1 OAI21X1_517 ( .A(_abc_40344_n2817), .B(_abc_40344_n2909), .C(_abc_40344_n2923), .Y(n1002) );
  OAI21X1 OAI21X1_518 ( .A(_abc_40344_n1232), .B(_abc_40344_n2926), .C(_abc_40344_n1222), .Y(_abc_40344_n2931) );
  OAI21X1 OAI21X1_519 ( .A(_abc_40344_n2930), .B(_abc_40344_n2932), .C(_abc_40344_n2818), .Y(_abc_40344_n2933) );
  OAI21X1 OAI21X1_52 ( .A(_abc_40344_n537_1), .B(_abc_40344_n538_1), .C(_abc_40344_n850_1), .Y(_abc_40344_n851) );
  OAI21X1 OAI21X1_520 ( .A(_abc_40344_n2938), .B(_abc_40344_n2942), .C(_abc_40344_n2871), .Y(_abc_40344_n2943) );
  OAI21X1 OAI21X1_521 ( .A(_abc_40344_n1222), .B(_abc_40344_n2878), .C(_abc_40344_n2945), .Y(_abc_40344_n2946) );
  OAI21X1 OAI21X1_522 ( .A(REG1_REG_14_), .B(_abc_40344_n2928), .C(_abc_40344_n1221), .Y(_abc_40344_n2949) );
  OAI21X1 OAI21X1_523 ( .A(_abc_40344_n1197), .B(_abc_40344_n2953), .C(_abc_40344_n2818), .Y(_abc_40344_n2955) );
  OAI21X1 OAI21X1_524 ( .A(_abc_40344_n2956), .B(_abc_40344_n2674), .C(_abc_40344_n2957), .Y(_abc_40344_n2958) );
  OAI21X1 OAI21X1_525 ( .A(REG2_REG_14_), .B(_abc_40344_n1221), .C(_abc_40344_n2964), .Y(_abc_40344_n2965) );
  OAI21X1 OAI21X1_526 ( .A(_abc_40344_n2954), .B(_abc_40344_n2955), .C(_abc_40344_n2968), .Y(n994) );
  OAI21X1 OAI21X1_527 ( .A(_abc_40344_n1196), .B(_abc_40344_n2952), .C(_abc_40344_n2975), .Y(_abc_40344_n2976) );
  OAI21X1 OAI21X1_528 ( .A(_abc_40344_n1207), .B(_abc_40344_n1196), .C(_abc_40344_n2965), .Y(_abc_40344_n2982) );
  OAI21X1 OAI21X1_529 ( .A(REG2_REG_15_), .B(_abc_40344_n1197), .C(_abc_40344_n2982), .Y(_abc_40344_n2983) );
  OAI21X1 OAI21X1_53 ( .A(_abc_40344_n848), .B(_abc_40344_n705_1), .C(_abc_40344_n855), .Y(_abc_40344_n856) );
  OAI21X1 OAI21X1_530 ( .A(_abc_40344_n2981), .B(_abc_40344_n2983), .C(_abc_40344_n2984), .Y(_abc_40344_n2985) );
  OAI21X1 OAI21X1_531 ( .A(_abc_40344_n1148), .B(_abc_40344_n2878), .C(_abc_40344_n2987), .Y(_abc_40344_n2988) );
  OAI21X1 OAI21X1_532 ( .A(_abc_40344_n2817), .B(_abc_40344_n2977), .C(_abc_40344_n2989), .Y(n990) );
  OAI21X1 OAI21X1_533 ( .A(_abc_40344_n1165), .B(_abc_40344_n1148), .C(_abc_40344_n2997), .Y(_abc_40344_n2998) );
  OAI21X1 OAI21X1_534 ( .A(_abc_40344_n2995), .B(_abc_40344_n2998), .C(_abc_40344_n2999), .Y(_abc_40344_n3000) );
  OAI21X1 OAI21X1_535 ( .A(_abc_40344_n2979), .B(_abc_40344_n2983), .C(_abc_40344_n2978), .Y(_abc_40344_n3005) );
  OAI21X1 OAI21X1_536 ( .A(_abc_40344_n3004), .B(_abc_40344_n3005), .C(_abc_40344_n3006), .Y(_abc_40344_n3007) );
  OAI21X1 OAI21X1_537 ( .A(_abc_40344_n3009), .B(_abc_40344_n2674), .C(_abc_40344_n3010), .Y(_abc_40344_n3011) );
  OAI21X1 OAI21X1_538 ( .A(_abc_40344_n1122), .B(_abc_40344_n2878), .C(_abc_40344_n3014), .Y(_abc_40344_n3015) );
  OAI21X1 OAI21X1_539 ( .A(_abc_40344_n1182), .B(_abc_40344_n1176), .C(_abc_40344_n3022), .Y(_abc_40344_n3023) );
  OAI21X1 OAI21X1_54 ( .A(_abc_40344_n857), .B(_abc_40344_n754_1), .C(_abc_40344_n858), .Y(_abc_40344_n859) );
  OAI21X1 OAI21X1_540 ( .A(_abc_40344_n3030), .B(_abc_40344_n3032), .C(_abc_40344_n3025), .Y(n982) );
  OAI21X1 OAI21X1_541 ( .A(REG2_REG_18_), .B(_abc_40344_n3017), .C(_abc_40344_n3023), .Y(_abc_40344_n3038) );
  OAI21X1 OAI21X1_542 ( .A(_abc_40344_n1131), .B(_abc_40344_n1122), .C(_abc_40344_n3041_1), .Y(_abc_40344_n3042) );
  OAI21X1 OAI21X1_543 ( .A(_abc_40344_n2952), .B(_abc_40344_n3048), .C(_abc_40344_n2971), .Y(_abc_40344_n3049) );
  OAI21X1 OAI21X1_544 ( .A(REG1_REG_18_), .B(_abc_40344_n3017), .C(_abc_40344_n3057), .Y(_abc_40344_n3058) );
  OAI21X1 OAI21X1_545 ( .A(_abc_40344_n2817), .B(_abc_40344_n3059), .C(_abc_40344_n3047), .Y(n978) );
  OAI21X1 OAI21X1_546 ( .A(_abc_40344_n984), .B(_abc_40344_n987), .C(_abc_40344_n979), .Y(_abc_40344_n3063) );
  OAI21X1 OAI21X1_547 ( .A(_abc_40344_n991), .B(_abc_40344_n1029_1), .C(_abc_40344_n3065), .Y(_abc_40344_n3066) );
  OAI21X1 OAI21X1_548 ( .A(_abc_40344_n3087), .B(_abc_40344_n705_1), .C(_abc_40344_n1418), .Y(_abc_40344_n3088) );
  OAI21X1 OAI21X1_549 ( .A(DATAI_22_), .B(DATAI_21_), .C(_abc_40344_n802), .Y(_abc_40344_n3090) );
  OAI21X1 OAI21X1_55 ( .A(_abc_40344_n860), .B(_abc_40344_n761_1), .C(_abc_40344_n861), .Y(_abc_40344_n862) );
  OAI21X1 OAI21X1_550 ( .A(_abc_40344_n1933), .B(_abc_40344_n705_1), .C(_abc_40344_n1083), .Y(_abc_40344_n3092) );
  OAI21X1 OAI21X1_551 ( .A(DATAI_26_), .B(DATAI_25_), .C(_abc_40344_n802), .Y(_abc_40344_n3093) );
  OAI21X1 OAI21X1_552 ( .A(DATAI_27_), .B(DATAI_28_), .C(_abc_40344_n802), .Y(_abc_40344_n3096) );
  OAI21X1 OAI21X1_553 ( .A(_abc_40344_n945_1), .B(_abc_40344_n610_1), .C(_abc_40344_n3103), .Y(_abc_40344_n3104) );
  OAI21X1 OAI21X1_554 ( .A(_abc_40344_n1910), .B(_abc_40344_n1913), .C(_abc_40344_n3105), .Y(_abc_40344_n3106) );
  OAI21X1 OAI21X1_555 ( .A(_abc_40344_n3106), .B(_abc_40344_n3067), .C(nRESET_G), .Y(_abc_40344_n3107) );
  OAI21X1 OAI21X1_556 ( .A(_abc_40344_n1916), .B(_abc_40344_n3111), .C(_abc_40344_n3108), .Y(_abc_40344_n3112) );
  OAI21X1 OAI21X1_557 ( .A(_abc_40344_n2394), .B(_abc_40344_n3097), .C(_abc_40344_n1922), .Y(_abc_40344_n3114) );
  OAI21X1 OAI21X1_558 ( .A(_abc_40344_n1922), .B(_abc_40344_n3111), .C(_abc_40344_n3117), .Y(_abc_40344_n3118) );
  OAI21X1 OAI21X1_559 ( .A(_abc_40344_n2009), .B(_abc_40344_n705_1), .C(_abc_40344_n1074), .Y(_abc_40344_n3121) );
  OAI21X1 OAI21X1_56 ( .A(DATAI_1_), .B(_abc_40344_n705_1), .C(_abc_40344_n868), .Y(_abc_40344_n869) );
  OAI21X1 OAI21X1_560 ( .A(_abc_40344_n908), .B(_abc_40344_n2476), .C(_abc_40344_n915_1), .Y(_abc_40344_n3126) );
  OAI21X1 OAI21X1_561 ( .A(_abc_40344_n919), .B(_abc_40344_n3125_1), .C(_abc_40344_n3126), .Y(_abc_40344_n3127) );
  OAI21X1 OAI21X1_562 ( .A(_abc_40344_n1009), .B(_abc_40344_n1017), .C(_abc_40344_n1665), .Y(_abc_40344_n3128) );
  OAI21X1 OAI21X1_563 ( .A(_abc_40344_n1350), .B(_abc_40344_n1362), .C(_abc_40344_n3124), .Y(_abc_40344_n3129) );
  OAI21X1 OAI21X1_564 ( .A(_abc_40344_n3128), .B(_abc_40344_n3129), .C(_abc_40344_n3130), .Y(_abc_40344_n3131) );
  OAI21X1 OAI21X1_565 ( .A(_abc_40344_n1019), .B(_abc_40344_n1665), .C(_abc_40344_n3132), .Y(_abc_40344_n3133) );
  OAI21X1 OAI21X1_566 ( .A(_abc_40344_n856), .B(_abc_40344_n864), .C(_abc_40344_n3136), .Y(_abc_40344_n3137) );
  OAI21X1 OAI21X1_567 ( .A(_abc_40344_n869), .B(_abc_40344_n863), .C(_abc_40344_n3137), .Y(_abc_40344_n3138) );
  OAI21X1 OAI21X1_568 ( .A(_abc_40344_n734), .B(_abc_40344_n742), .C(_abc_40344_n3139), .Y(_abc_40344_n3140) );
  OAI21X1 OAI21X1_569 ( .A(_abc_40344_n813), .B(_abc_40344_n808), .C(_abc_40344_n3141), .Y(_abc_40344_n3142) );
  OAI21X1 OAI21X1_57 ( .A(_abc_40344_n871), .B(_abc_40344_n870), .C(_abc_40344_n720), .Y(_abc_40344_n872) );
  OAI21X1 OAI21X1_570 ( .A(_abc_40344_n2016), .B(_abc_40344_n2017), .C(_abc_40344_n813), .Y(_abc_40344_n3145) );
  OAI21X1 OAI21X1_571 ( .A(_abc_40344_n838), .B(_abc_40344_n840), .C(_abc_40344_n825), .Y(_abc_40344_n3146) );
  OAI21X1 OAI21X1_572 ( .A(_abc_40344_n813), .B(_abc_40344_n808), .C(_abc_40344_n3149), .Y(_abc_40344_n3150) );
  OAI21X1 OAI21X1_573 ( .A(_abc_40344_n3152), .B(_abc_40344_n3151), .C(_abc_40344_n3148), .Y(_abc_40344_n3153) );
  OAI21X1 OAI21X1_574 ( .A(_abc_40344_n3147_1), .B(_abc_40344_n3150), .C(_abc_40344_n3153), .Y(_abc_40344_n3154) );
  OAI21X1 OAI21X1_575 ( .A(_abc_40344_n1205), .B(_abc_40344_n1208), .C(_abc_40344_n1201), .Y(_abc_40344_n3161) );
  OAI21X1 OAI21X1_576 ( .A(_abc_40344_n1280), .B(_abc_40344_n1283), .C(_abc_40344_n1273), .Y(_abc_40344_n3162) );
  OAI21X1 OAI21X1_577 ( .A(_abc_40344_n1251), .B(_abc_40344_n1260), .C(_abc_40344_n3163), .Y(_abc_40344_n3164) );
  OAI21X1 OAI21X1_578 ( .A(_abc_40344_n3162), .B(_abc_40344_n3164), .C(_abc_40344_n3165), .Y(_abc_40344_n3166) );
  OAI21X1 OAI21X1_579 ( .A(_abc_40344_n1251), .B(_abc_40344_n1260), .C(_abc_40344_n3166), .Y(_abc_40344_n3167) );
  OAI21X1 OAI21X1_58 ( .A(_abc_40344_n877_1), .B(_abc_40344_n705_1), .C(_abc_40344_n878), .Y(_abc_40344_n879) );
  OAI21X1 OAI21X1_580 ( .A(_abc_40344_n1961), .B(_abc_40344_n1818), .C(_abc_40344_n3167), .Y(_abc_40344_n3168) );
  OAI21X1 OAI21X1_581 ( .A(_abc_40344_n1224), .B(_abc_40344_n1234), .C(_abc_40344_n3168), .Y(_abc_40344_n3169) );
  OAI21X1 OAI21X1_582 ( .A(_abc_40344_n3160), .B(_abc_40344_n3169), .C(_abc_40344_n3161), .Y(_abc_40344_n3170) );
  OAI21X1 OAI21X1_583 ( .A(_abc_40344_n1273), .B(_abc_40344_n1285), .C(_abc_40344_n3171), .Y(_abc_40344_n3172_1) );
  OAI21X1 OAI21X1_584 ( .A(_abc_40344_n1224), .B(_abc_40344_n1234), .C(_abc_40344_n3173), .Y(_abc_40344_n3174) );
  OAI21X1 OAI21X1_585 ( .A(_abc_40344_n1133), .B(_abc_40344_n1130), .C(_abc_40344_n1124), .Y(_abc_40344_n3178) );
  OAI21X1 OAI21X1_586 ( .A(_abc_40344_n1434), .B(_abc_40344_n1441), .C(_abc_40344_n3180), .Y(_abc_40344_n3181) );
  OAI21X1 OAI21X1_587 ( .A(_abc_40344_n1428), .B(_abc_40344_n1424), .C(_abc_40344_n1812), .Y(_abc_40344_n3182) );
  OAI21X1 OAI21X1_588 ( .A(_abc_40344_n1413), .B(_abc_40344_n1410), .C(_abc_40344_n1404), .Y(_abc_40344_n3183) );
  OAI21X1 OAI21X1_589 ( .A(_abc_40344_n3178), .B(_abc_40344_n3181), .C(_abc_40344_n3185), .Y(_abc_40344_n3186) );
  OAI21X1 OAI21X1_59 ( .A(IR_REG_6_), .B(_abc_40344_n709), .C(IR_REG_7_), .Y(_abc_40344_n903_1) );
  OAI21X1 OAI21X1_590 ( .A(_abc_40344_n1163), .B(_abc_40344_n1166_1), .C(_abc_40344_n1153), .Y(_abc_40344_n3189) );
  OAI21X1 OAI21X1_591 ( .A(_abc_40344_n3194), .B(_abc_40344_n3176), .C(_abc_40344_n3191), .Y(_abc_40344_n3195) );
  OAI21X1 OAI21X1_592 ( .A(_abc_40344_n1100), .B(_abc_40344_n1111), .C(_abc_40344_n3195), .Y(_abc_40344_n3196) );
  OAI21X1 OAI21X1_593 ( .A(_abc_40344_n1099), .B(_abc_40344_n1110), .C(_abc_40344_n3196), .Y(_abc_40344_n3197) );
  OAI21X1 OAI21X1_594 ( .A(_abc_40344_n3123), .B(_abc_40344_n3197), .C(_abc_40344_n2522), .Y(_abc_40344_n3198) );
  OAI21X1 OAI21X1_595 ( .A(_abc_40344_n1491), .B(_abc_40344_n1488), .C(_abc_40344_n3199), .Y(_abc_40344_n3200) );
  OAI21X1 OAI21X1_596 ( .A(_abc_40344_n1463), .B(_abc_40344_n1471), .C(_abc_40344_n3201), .Y(_abc_40344_n3202) );
  OAI21X1 OAI21X1_597 ( .A(_abc_40344_n3204), .B(_abc_40344_n3203), .C(_abc_40344_n1491), .Y(_abc_40344_n3205) );
  OAI21X1 OAI21X1_598 ( .A(_abc_40344_n2519), .B(_abc_40344_n3200), .C(_abc_40344_n3207), .Y(_abc_40344_n3208) );
  OAI21X1 OAI21X1_599 ( .A(_abc_40344_n3202), .B(_abc_40344_n3198), .C(_abc_40344_n3210), .Y(_abc_40344_n3211) );
  OAI21X1 OAI21X1_6 ( .A(_abc_40344_n559_1), .B(_abc_40344_n583), .C(_abc_40344_n584_1), .Y(_abc_40344_n585) );
  OAI21X1 OAI21X1_60 ( .A(_abc_40344_n542_1), .B(_abc_40344_n706), .C(_abc_40344_n903_1), .Y(_abc_40344_n904) );
  OAI21X1 OAI21X1_600 ( .A(_abc_40344_n3122), .B(_abc_40344_n3211), .C(_abc_40344_n3121), .Y(_abc_40344_n3212) );
  OAI21X1 OAI21X1_601 ( .A(_abc_40344_n699), .B(_abc_40344_n2644_1), .C(_abc_40344_n3222), .Y(_abc_40344_n3223) );
  OAI21X1 OAI21X1_602 ( .A(_abc_40344_n2513), .B(_abc_40344_n2647), .C(_abc_40344_n2583), .Y(_abc_40344_n3225) );
  OAI21X1 OAI21X1_603 ( .A(_abc_40344_n2577), .B(_abc_40344_n3225), .C(_abc_40344_n2651), .Y(_abc_40344_n3226) );
  OAI21X1 OAI21X1_604 ( .A(_abc_40344_n626), .B(_abc_40344_n646), .C(_abc_40344_n2643), .Y(_abc_40344_n3227) );
  OAI21X1 OAI21X1_605 ( .A(_abc_40344_n3120), .B(_abc_40344_n3226), .C(_abc_40344_n3229), .Y(_abc_40344_n3230) );
  OAI21X1 OAI21X1_606 ( .A(_abc_40344_n1630), .B(_abc_40344_n3111), .C(_abc_40344_n3234), .Y(_abc_40344_n3235) );
  OAI21X1 OAI21X1_607 ( .A(_abc_40344_n1076), .B(_abc_40344_n3237), .C(_abc_40344_n1649), .Y(_abc_40344_n3238) );
  OAI21X1 OAI21X1_608 ( .A(_abc_40344_n3215), .B(_abc_40344_n3219), .C(_abc_40344_n3242), .Y(n958) );
  OAI21X1 OAI21X1_609 ( .A(_abc_40344_n2512), .B(_abc_40344_n3225), .C(_abc_40344_n3249), .Y(_abc_40344_n3250) );
  OAI21X1 OAI21X1_61 ( .A(_abc_40344_n559_1), .B(_abc_40344_n904), .C(_abc_40344_n905), .Y(_abc_40344_n906_1) );
  OAI21X1 OAI21X1_610 ( .A(_abc_40344_n1040), .B(_abc_40344_n3111), .C(_abc_40344_n3254), .Y(_abc_40344_n3255) );
  OAI21X1 OAI21X1_611 ( .A(_abc_40344_n3219), .B(_abc_40344_n3245), .C(_abc_40344_n3257), .Y(_abc_40344_n3258) );
  OAI21X1 OAI21X1_612 ( .A(_abc_40344_n1550), .B(_abc_40344_n3244), .C(_abc_40344_n3259), .Y(n953) );
  OAI21X1 OAI21X1_613 ( .A(_abc_40344_n3262), .B(_abc_40344_n3198), .C(_abc_40344_n2519), .Y(_abc_40344_n3263) );
  OAI21X1 OAI21X1_614 ( .A(_abc_40344_n1491), .B(_abc_40344_n1488), .C(_abc_40344_n3263), .Y(_abc_40344_n3264) );
  OAI21X1 OAI21X1_615 ( .A(_abc_40344_n1477), .B(_abc_40344_n1489), .C(_abc_40344_n3264), .Y(_abc_40344_n3265) );
  OAI21X1 OAI21X1_616 ( .A(_abc_40344_n2513), .B(_abc_40344_n2647), .C(_abc_40344_n2119), .Y(_abc_40344_n3267) );
  OAI21X1 OAI21X1_617 ( .A(_abc_40344_n3261), .B(_abc_40344_n3266), .C(_abc_40344_n3269_1), .Y(_abc_40344_n3270) );
  OAI21X1 OAI21X1_618 ( .A(_abc_40344_n1933), .B(_abc_40344_n705_1), .C(_abc_40344_n3271), .Y(_abc_40344_n3272) );
  OAI21X1 OAI21X1_619 ( .A(_abc_40344_n1491), .B(_abc_40344_n3272), .C(_abc_40344_n1495), .Y(_abc_40344_n3273) );
  OAI21X1 OAI21X1_62 ( .A(_abc_40344_n902_1), .B(_abc_40344_n705_1), .C(_abc_40344_n907), .Y(_abc_40344_n908) );
  OAI21X1 OAI21X1_620 ( .A(_abc_40344_n1494), .B(_abc_40344_n3111), .C(_abc_40344_n3276), .Y(_abc_40344_n3277) );
  OAI21X1 OAI21X1_621 ( .A(_abc_40344_n3219), .B(_abc_40344_n3266), .C(_abc_40344_n3279), .Y(_abc_40344_n3280) );
  OAI21X1 OAI21X1_622 ( .A(_abc_40344_n1074), .B(_abc_40344_n3244), .C(_abc_40344_n3281), .Y(n948) );
  OAI21X1 OAI21X1_623 ( .A(_abc_40344_n2118), .B(_abc_40344_n2513), .C(_abc_40344_n2637), .Y(_abc_40344_n3284) );
  OAI21X1 OAI21X1_624 ( .A(_abc_40344_n3261), .B(_abc_40344_n3283), .C(_abc_40344_n3286), .Y(_abc_40344_n3287) );
  OAI21X1 OAI21X1_625 ( .A(_abc_40344_n1477), .B(_abc_40344_n3111), .C(_abc_40344_n3288), .Y(_abc_40344_n3289) );
  OAI21X1 OAI21X1_626 ( .A(_abc_40344_n3219), .B(_abc_40344_n3283), .C(_abc_40344_n3294), .Y(n943) );
  OAI21X1 OAI21X1_627 ( .A(_abc_40344_n1201), .B(_abc_40344_n1209_1), .C(_abc_40344_n1947), .Y(_abc_40344_n3300) );
  OAI21X1 OAI21X1_628 ( .A(_abc_40344_n3300), .B(_abc_40344_n3299), .C(_abc_40344_n2502_1), .Y(_abc_40344_n3301) );
  OAI21X1 OAI21X1_629 ( .A(_abc_40344_n1298), .B(_abc_40344_n1304_1), .C(_abc_40344_n1295), .Y(_abc_40344_n3304) );
  OAI21X1 OAI21X1_63 ( .A(_abc_40344_n686), .B(_abc_40344_n690), .C(_abc_40344_n910), .Y(_abc_40344_n911) );
  OAI21X1 OAI21X1_630 ( .A(_abc_40344_n825), .B(_abc_40344_n841), .C(_abc_40344_n2633), .Y(_abc_40344_n3307) );
  OAI21X1 OAI21X1_631 ( .A(_abc_40344_n2624), .B(_abc_40344_n3308), .C(_abc_40344_n3309), .Y(_abc_40344_n3310) );
  OAI21X1 OAI21X1_632 ( .A(_abc_40344_n1985), .B(_abc_40344_n1908), .C(_abc_40344_n2530), .Y(_abc_40344_n3312) );
  OAI21X1 OAI21X1_633 ( .A(_abc_40344_n1273), .B(_abc_40344_n1284), .C(_abc_40344_n1970), .Y(_abc_40344_n3314_1) );
  OAI21X1 OAI21X1_634 ( .A(_abc_40344_n3314_1), .B(_abc_40344_n3315), .C(_abc_40344_n2122), .Y(_abc_40344_n3316) );
  OAI21X1 OAI21X1_635 ( .A(_abc_40344_n1906), .B(_abc_40344_n1362), .C(_abc_40344_n3317), .Y(_abc_40344_n3318) );
  OAI21X1 OAI21X1_636 ( .A(_abc_40344_n3318), .B(_abc_40344_n3313), .C(_abc_40344_n3316), .Y(_abc_40344_n3319) );
  OAI21X1 OAI21X1_637 ( .A(_abc_40344_n3305), .B(_abc_40344_n3319), .C(_abc_40344_n3306), .Y(_abc_40344_n3320) );
  OAI21X1 OAI21X1_638 ( .A(_abc_40344_n1961), .B(_abc_40344_n1234), .C(_abc_40344_n2599_1), .Y(_abc_40344_n3322) );
  OAI21X1 OAI21X1_639 ( .A(_abc_40344_n1137), .B(_abc_40344_n1134), .C(_abc_40344_n3325), .Y(_abc_40344_n3326) );
  OAI21X1 OAI21X1_64 ( .A(DATAI_7_), .B(_abc_40344_n705_1), .C(_abc_40344_n918), .Y(_abc_40344_n919) );
  OAI21X1 OAI21X1_640 ( .A(_abc_40344_n1956), .B(_abc_40344_n2038), .C(_abc_40344_n1953), .Y(_abc_40344_n3329) );
  OAI21X1 OAI21X1_641 ( .A(_abc_40344_n1099), .B(_abc_40344_n1111), .C(_abc_40344_n1945), .Y(_abc_40344_n3332) );
  OAI21X1 OAI21X1_642 ( .A(_abc_40344_n3331), .B(_abc_40344_n3332), .C(_abc_40344_n3333), .Y(_abc_40344_n3334) );
  OAI21X1 OAI21X1_643 ( .A(_abc_40344_n3330), .B(_abc_40344_n3334), .C(_abc_40344_n1945), .Y(_abc_40344_n3335_1) );
  OAI21X1 OAI21X1_644 ( .A(_abc_40344_n2521), .B(_abc_40344_n3336), .C(_abc_40344_n3227), .Y(_abc_40344_n3338) );
  OAI21X1 OAI21X1_645 ( .A(_abc_40344_n3337), .B(_abc_40344_n3338), .C(_abc_40344_n3297), .Y(_abc_40344_n3339) );
  OAI21X1 OAI21X1_646 ( .A(_abc_40344_n1084), .B(_abc_40344_n3091), .C(_abc_40344_n1463), .Y(_abc_40344_n3341) );
  OAI21X1 OAI21X1_647 ( .A(_abc_40344_n3091), .B(_abc_40344_n3092), .C(_abc_40344_n3341), .Y(_abc_40344_n3342) );
  OAI21X1 OAI21X1_648 ( .A(_abc_40344_n1031), .B(_abc_40344_n1466), .C(_abc_40344_n3345), .Y(_abc_40344_n3346) );
  OAI21X1 OAI21X1_649 ( .A(_abc_40344_n3069), .B(_abc_40344_n3342), .C(_abc_40344_n3347), .Y(_abc_40344_n3348) );
  OAI21X1 OAI21X1_65 ( .A(_abc_40344_n932), .B(_abc_40344_n940), .C(_abc_40344_n727_1), .Y(_abc_40344_n941) );
  OAI21X1 OAI21X1_650 ( .A(_abc_40344_n3329), .B(_abc_40344_n3327), .C(_abc_40344_n2030), .Y(_abc_40344_n3353) );
  OAI21X1 OAI21X1_651 ( .A(_abc_40344_n2029), .B(_abc_40344_n3358), .C(_abc_40344_n3331), .Y(_abc_40344_n3359_1) );
  OAI21X1 OAI21X1_652 ( .A(_abc_40344_n1100), .B(_abc_40344_n1110), .C(_abc_40344_n2524), .Y(_abc_40344_n3362) );
  OAI21X1 OAI21X1_653 ( .A(_abc_40344_n3331), .B(_abc_40344_n3363), .C(_abc_40344_n1943), .Y(_abc_40344_n3364) );
  OAI21X1 OAI21X1_654 ( .A(_abc_40344_n1099), .B(_abc_40344_n1111), .C(_abc_40344_n2524), .Y(_abc_40344_n3365) );
  OAI21X1 OAI21X1_655 ( .A(_abc_40344_n2524), .B(_abc_40344_n3364), .C(_abc_40344_n3365), .Y(_abc_40344_n3366) );
  OAI21X1 OAI21X1_656 ( .A(_abc_40344_n3362), .B(_abc_40344_n3361), .C(_abc_40344_n3366), .Y(_abc_40344_n3367) );
  OAI21X1 OAI21X1_657 ( .A(_abc_40344_n3354), .B(_abc_40344_n3367), .C(_abc_40344_n3227), .Y(_abc_40344_n3368) );
  OAI21X1 OAI21X1_658 ( .A(_abc_40344_n1083), .B(_abc_40344_n3111), .C(_abc_40344_n3373), .Y(_abc_40344_n3374) );
  OAI21X1 OAI21X1_659 ( .A(_abc_40344_n1577), .B(_abc_40344_n3244), .C(_abc_40344_n3375), .Y(_abc_40344_n3376) );
  OAI21X1 OAI21X1_66 ( .A(IR_REG_31_), .B(_abc_40344_n566), .C(_abc_40344_n635), .Y(_abc_40344_n942) );
  OAI21X1 OAI21X1_660 ( .A(_abc_40344_n1944), .B(_abc_40344_n3363), .C(_abc_40344_n3361), .Y(_abc_40344_n3383) );
  OAI21X1 OAI21X1_661 ( .A(_abc_40344_n1434), .B(_abc_40344_n3386), .C(_abc_40344_n1100), .Y(_abc_40344_n3387) );
  OAI21X1 OAI21X1_662 ( .A(_abc_40344_n1099), .B(_abc_40344_n3111), .C(_abc_40344_n3390), .Y(_abc_40344_n3391) );
  OAI21X1 OAI21X1_663 ( .A(_abc_40344_n3219), .B(_abc_40344_n3380), .C(_abc_40344_n3392), .Y(_abc_40344_n3393) );
  OAI21X1 OAI21X1_664 ( .A(_abc_40344_n3067), .B(_abc_40344_n3385), .C(_abc_40344_n3394), .Y(n928) );
  OAI21X1 OAI21X1_665 ( .A(_abc_40344_n3398), .B(_abc_40344_n3399), .C(_abc_40344_n3227), .Y(_abc_40344_n3400) );
  OAI21X1 OAI21X1_666 ( .A(_abc_40344_n1428), .B(_abc_40344_n1424), .C(_abc_40344_n3220), .Y(_abc_40344_n3402) );
  OAI21X1 OAI21X1_667 ( .A(_abc_40344_n3405), .B(_abc_40344_n3176), .C(_abc_40344_n3404), .Y(_abc_40344_n3406) );
  OAI21X1 OAI21X1_668 ( .A(_abc_40344_n3187), .B(_abc_40344_n3407), .C(_abc_40344_n3178), .Y(_abc_40344_n3408) );
  OAI21X1 OAI21X1_669 ( .A(_abc_40344_n1404), .B(_abc_40344_n1415), .C(_abc_40344_n3408), .Y(_abc_40344_n3409) );
  OAI21X1 OAI21X1_67 ( .A(D_REG_1_), .B(_abc_40344_n950), .C(_abc_40344_n944), .Y(_abc_40344_n951) );
  OAI21X1 OAI21X1_670 ( .A(_abc_40344_n3179), .B(_abc_40344_n3409), .C(_abc_40344_n3403), .Y(_abc_40344_n3410) );
  OAI21X1 OAI21X1_671 ( .A(_abc_40344_n1952), .B(_abc_40344_n2029), .C(_abc_40344_n3410), .Y(_abc_40344_n3411_1) );
  OAI21X1 OAI21X1_672 ( .A(_abc_40344_n3261), .B(_abc_40344_n3413), .C(_abc_40344_n3402), .Y(_abc_40344_n3414) );
  OAI21X1 OAI21X1_673 ( .A(_abc_40344_n1433), .B(_abc_40344_n3111), .C(_abc_40344_n3417), .Y(_abc_40344_n3418) );
  OAI21X1 OAI21X1_674 ( .A(_abc_40344_n3219), .B(_abc_40344_n3413), .C(_abc_40344_n3419), .Y(_abc_40344_n3420) );
  OAI21X1 OAI21X1_675 ( .A(_abc_40344_n1404), .B(_abc_40344_n3423), .C(_abc_40344_n1812), .Y(_abc_40344_n3424) );
  OAI21X1 OAI21X1_676 ( .A(_abc_40344_n3423), .B(_abc_40344_n3088), .C(_abc_40344_n3424), .Y(_abc_40344_n3425) );
  OAI21X1 OAI21X1_677 ( .A(_abc_40344_n2527), .B(_abc_40344_n3426), .C(_abc_40344_n3427), .Y(_abc_40344_n3428) );
  OAI21X1 OAI21X1_678 ( .A(_abc_40344_n1413), .B(_abc_40344_n1410), .C(_abc_40344_n3220), .Y(_abc_40344_n3429) );
  OAI21X1 OAI21X1_679 ( .A(_abc_40344_n1418), .B(_abc_40344_n1414), .C(_abc_40344_n3409), .Y(_abc_40344_n3430) );
  OAI21X1 OAI21X1_68 ( .A(_abc_40344_n964), .B(_abc_40344_n977), .C(_abc_40344_n952), .Y(_abc_40344_n978) );
  OAI21X1 OAI21X1_680 ( .A(_abc_40344_n1954), .B(_abc_40344_n2038), .C(_abc_40344_n3430), .Y(_abc_40344_n3432) );
  OAI21X1 OAI21X1_681 ( .A(_abc_40344_n1423), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3439) );
  OAI21X1 OAI21X1_682 ( .A(_abc_40344_n3219), .B(_abc_40344_n3433), .C(_abc_40344_n3441), .Y(_abc_40344_n3442) );
  OAI21X1 OAI21X1_683 ( .A(_abc_40344_n3069), .B(_abc_40344_n3425), .C(_abc_40344_n3443), .Y(n918) );
  OAI21X1 OAI21X1_684 ( .A(_abc_40344_n1418), .B(_abc_40344_n3111), .C(_abc_40344_n3448), .Y(_abc_40344_n3449) );
  OAI21X1 OAI21X1_685 ( .A(_abc_40344_n3069), .B(_abc_40344_n3446), .C(_abc_40344_n3450), .Y(_abc_40344_n3451) );
  OAI21X1 OAI21X1_686 ( .A(_abc_40344_n2473), .B(_abc_40344_n3326), .C(_abc_40344_n3227), .Y(_abc_40344_n3453) );
  OAI21X1 OAI21X1_687 ( .A(_abc_40344_n3454), .B(_abc_40344_n3456), .C(_abc_40344_n3066), .Y(_abc_40344_n3457_1) );
  OAI21X1 OAI21X1_688 ( .A(_abc_40344_n3228), .B(_abc_40344_n3462), .C(_abc_40344_n3463), .Y(_abc_40344_n3464) );
  OAI21X1 OAI21X1_689 ( .A(_abc_40344_n1178), .B(_abc_40344_n3466), .C(_abc_40344_n1124), .Y(_abc_40344_n3467) );
  OAI21X1 OAI21X1_69 ( .A(_abc_40344_n986), .B(_abc_40344_n987), .C(_abc_40344_n984), .Y(_abc_40344_n988) );
  OAI21X1 OAI21X1_690 ( .A(_abc_40344_n3067), .B(_abc_40344_n3470), .C(_abc_40344_n3471), .Y(_abc_40344_n3472) );
  OAI21X1 OAI21X1_691 ( .A(_abc_40344_n1128), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3473) );
  OAI21X1 OAI21X1_692 ( .A(_abc_40344_n3219), .B(_abc_40344_n3460), .C(_abc_40344_n3476), .Y(n908) );
  OAI21X1 OAI21X1_693 ( .A(_abc_40344_n3192), .B(_abc_40344_n3176), .C(_abc_40344_n3189), .Y(_abc_40344_n3479) );
  OAI21X1 OAI21X1_694 ( .A(_abc_40344_n1939), .B(_abc_40344_n3482), .C(_abc_40344_n2544), .Y(_abc_40344_n3483) );
  OAI21X1 OAI21X1_695 ( .A(_abc_40344_n3322), .B(_abc_40344_n3483), .C(_abc_40344_n3301), .Y(_abc_40344_n3484) );
  OAI21X1 OAI21X1_696 ( .A(_abc_40344_n3478_1), .B(_abc_40344_n3484), .C(_abc_40344_n3485), .Y(_abc_40344_n3486) );
  OAI21X1 OAI21X1_697 ( .A(_abc_40344_n1167), .B(_abc_40344_n3379), .C(_abc_40344_n3486), .Y(_abc_40344_n3487) );
  OAI21X1 OAI21X1_698 ( .A(_abc_40344_n1133), .B(_abc_40344_n1130), .C(_abc_40344_n3103), .Y(_abc_40344_n3492) );
  OAI21X1 OAI21X1_699 ( .A(_abc_40344_n1179), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3494) );
  OAI21X1 OAI21X1_7 ( .A(_abc_40344_n559_1), .B(_abc_40344_n599), .C(_abc_40344_n601), .Y(_abc_40344_n602) );
  OAI21X1 OAI21X1_70 ( .A(_abc_40344_n561_1), .B(_abc_40344_n580), .C(_abc_40344_n586), .Y(_abc_40344_n989) );
  OAI21X1 OAI21X1_700 ( .A(_abc_40344_n3067), .B(_abc_40344_n3489), .C(_abc_40344_n3498), .Y(n903) );
  OAI21X1 OAI21X1_701 ( .A(_abc_40344_n2049), .B(_abc_40344_n3483), .C(_abc_40344_n2479), .Y(_abc_40344_n3502) );
  OAI21X1 OAI21X1_702 ( .A(_abc_40344_n3228), .B(_abc_40344_n3504), .C(_abc_40344_n3501), .Y(_abc_40344_n3505) );
  OAI21X1 OAI21X1_703 ( .A(_abc_40344_n1161), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3511) );
  OAI21X1 OAI21X1_704 ( .A(_abc_40344_n1164), .B(_abc_40344_n3066), .C(_abc_40344_n3512), .Y(_abc_40344_n3513) );
  OAI21X1 OAI21X1_705 ( .A(_abc_40344_n1185), .B(_abc_40344_n3244), .C(_abc_40344_n3514), .Y(_abc_40344_n3515) );
  OAI21X1 OAI21X1_706 ( .A(_abc_40344_n3174), .B(_abc_40344_n3518), .C(_abc_40344_n3169), .Y(_abc_40344_n3519) );
  OAI21X1 OAI21X1_707 ( .A(_abc_40344_n3228), .B(_abc_40344_n3522), .C(_abc_40344_n3521), .Y(_abc_40344_n3523) );
  OAI21X1 OAI21X1_708 ( .A(_abc_40344_n1224), .B(_abc_40344_n3528), .C(_abc_40344_n1201), .Y(_abc_40344_n3529) );
  OAI21X1 OAI21X1_709 ( .A(_abc_40344_n1203), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3532) );
  OAI21X1 OAI21X1_71 ( .A(_abc_40344_n941), .B(_abc_40344_n939), .C(_abc_40344_n993), .Y(_abc_40344_n994) );
  OAI21X1 OAI21X1_710 ( .A(_abc_40344_n1200), .B(_abc_40344_n3111), .C(_abc_40344_n3533), .Y(_abc_40344_n3534) );
  OAI21X1 OAI21X1_711 ( .A(_abc_40344_n3069), .B(_abc_40344_n3531), .C(_abc_40344_n3535_1), .Y(_abc_40344_n3536) );
  OAI21X1 OAI21X1_712 ( .A(_abc_40344_n3172_1), .B(_abc_40344_n3518), .C(_abc_40344_n3167), .Y(_abc_40344_n3540) );
  OAI21X1 OAI21X1_713 ( .A(_abc_40344_n3228), .B(_abc_40344_n3539), .C(_abc_40344_n3542), .Y(_abc_40344_n3543) );
  OAI21X1 OAI21X1_714 ( .A(_abc_40344_n1251), .B(_abc_40344_n3545), .C(_abc_40344_n1224), .Y(_abc_40344_n3546) );
  OAI21X1 OAI21X1_715 ( .A(_abc_40344_n1209_1), .B(_abc_40344_n3232), .C(_abc_40344_n3066), .Y(_abc_40344_n3549) );
  OAI21X1 OAI21X1_716 ( .A(REG2_REG_14_), .B(_abc_40344_n3066), .C(_abc_40344_n3549), .Y(_abc_40344_n3550) );
  OAI21X1 OAI21X1_717 ( .A(_abc_40344_n1228), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3551) );
  OAI21X1 OAI21X1_718 ( .A(_abc_40344_n3069), .B(_abc_40344_n3548), .C(_abc_40344_n3553), .Y(_abc_40344_n3554) );
  OAI21X1 OAI21X1_719 ( .A(_abc_40344_n1308), .B(_abc_40344_n3526), .C(_abc_40344_n1251), .Y(_abc_40344_n3557) );
  OAI21X1 OAI21X1_72 ( .A(_abc_40344_n523), .B(_abc_40344_n988), .C(_abc_40344_n996), .Y(_abc_40344_n997) );
  OAI21X1 OAI21X1_720 ( .A(_abc_40344_n2545), .B(_abc_40344_n3320), .C(_abc_40344_n3227), .Y(_abc_40344_n3560) );
  OAI21X1 OAI21X1_721 ( .A(_abc_40344_n1273), .B(_abc_40344_n1285), .C(_abc_40344_n3159), .Y(_abc_40344_n3561) );
  OAI21X1 OAI21X1_722 ( .A(_abc_40344_n1973), .B(_abc_40344_n1284), .C(_abc_40344_n3561), .Y(_abc_40344_n3562) );
  OAI21X1 OAI21X1_723 ( .A(_abc_40344_n2501), .B(_abc_40344_n3562), .C(_abc_40344_n3163), .Y(_abc_40344_n3563) );
  OAI21X1 OAI21X1_724 ( .A(_abc_40344_n3559), .B(_abc_40344_n3560), .C(_abc_40344_n3565), .Y(_abc_40344_n3566) );
  OAI21X1 OAI21X1_725 ( .A(_abc_40344_n1255), .B(_abc_40344_n3066), .C(nRESET_G), .Y(_abc_40344_n3569) );
  OAI21X1 OAI21X1_726 ( .A(_abc_40344_n3069), .B(_abc_40344_n3558), .C(_abc_40344_n3572), .Y(n883) );
  OAI21X1 OAI21X1_727 ( .A(_abc_40344_n1273), .B(_abc_40344_n3574), .C(_abc_40344_n1308), .Y(_abc_40344_n3575) );
  OAI21X1 OAI21X1_728 ( .A(_abc_40344_n2500), .B(_abc_40344_n2501), .C(_abc_40344_n3319), .Y(_abc_40344_n3578) );
  OAI21X1 OAI21X1_729 ( .A(_abc_40344_n3577), .B(_abc_40344_n3579), .C(_abc_40344_n3582), .Y(_abc_40344_n3583) );
  OAI21X1 OAI21X1_73 ( .A(_abc_40344_n984), .B(_abc_40344_n987), .C(_abc_40344_n998), .Y(_abc_40344_n999) );
  OAI21X1 OAI21X1_730 ( .A(_abc_40344_n1031), .B(_abc_40344_n1302), .C(_abc_40344_n3587), .Y(_abc_40344_n3588) );
  OAI21X1 OAI21X1_731 ( .A(_abc_40344_n3219), .B(_abc_40344_n3584), .C(_abc_40344_n3589), .Y(_abc_40344_n3590) );
  OAI21X1 OAI21X1_732 ( .A(_abc_40344_n3069), .B(_abc_40344_n3576), .C(_abc_40344_n3591), .Y(n878) );
  OAI21X1 OAI21X1_733 ( .A(_abc_40344_n2151), .B(_abc_40344_n3313), .C(_abc_40344_n1907), .Y(_abc_40344_n3596) );
  OAI21X1 OAI21X1_734 ( .A(_abc_40344_n2125), .B(_abc_40344_n3597), .C(_abc_40344_n1970), .Y(_abc_40344_n3598) );
  OAI21X1 OAI21X1_735 ( .A(_abc_40344_n3228), .B(_abc_40344_n3599), .C(_abc_40344_n3595), .Y(_abc_40344_n3600) );
  OAI21X1 OAI21X1_736 ( .A(_abc_40344_n1327), .B(_abc_40344_n3078), .C(_abc_40344_n1273), .Y(_abc_40344_n3604_1) );
  OAI21X1 OAI21X1_737 ( .A(_abc_40344_n3219), .B(_abc_40344_n3593), .C(_abc_40344_n3608), .Y(n873) );
  OAI21X1 OAI21X1_738 ( .A(_abc_40344_n923_1), .B(_abc_40344_n926), .C(_abc_40344_n908), .Y(_abc_40344_n3611) );
  OAI21X1 OAI21X1_739 ( .A(_abc_40344_n2476), .B(_abc_40344_n3155), .C(_abc_40344_n3612), .Y(_abc_40344_n3613) );
  OAI21X1 OAI21X1_74 ( .A(_abc_40344_n1012), .B(_abc_40344_n690), .C(_abc_40344_n1011), .Y(_abc_40344_n1013) );
  OAI21X1 OAI21X1_740 ( .A(_abc_40344_n3156), .B(_abc_40344_n3613), .C(_abc_40344_n3611), .Y(_abc_40344_n3614) );
  OAI21X1 OAI21X1_741 ( .A(_abc_40344_n1019), .B(_abc_40344_n1665), .C(_abc_40344_n3614), .Y(_abc_40344_n3615) );
  OAI21X1 OAI21X1_742 ( .A(_abc_40344_n1018), .B(_abc_40344_n1375), .C(_abc_40344_n3615), .Y(_abc_40344_n3616) );
  OAI21X1 OAI21X1_743 ( .A(_abc_40344_n1350), .B(_abc_40344_n1362), .C(_abc_40344_n3616), .Y(_abc_40344_n3617) );
  OAI21X1 OAI21X1_744 ( .A(_abc_40344_n1906), .B(_abc_40344_n1361), .C(_abc_40344_n3617), .Y(_abc_40344_n3618) );
  OAI21X1 OAI21X1_745 ( .A(_abc_40344_n3228), .B(_abc_40344_n3610), .C(_abc_40344_n3620), .Y(_abc_40344_n3621) );
  OAI21X1 OAI21X1_746 ( .A(_abc_40344_n1350), .B(_abc_40344_n3623), .C(_abc_40344_n1327), .Y(_abc_40344_n3624) );
  OAI21X1 OAI21X1_747 ( .A(REG2_REG_10_), .B(_abc_40344_n3066), .C(_abc_40344_n3628), .Y(_abc_40344_n3629) );
  OAI21X1 OAI21X1_748 ( .A(_abc_40344_n1330), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3630) );
  OAI21X1 OAI21X1_749 ( .A(_abc_40344_n3067), .B(_abc_40344_n3622), .C(_abc_40344_n3633), .Y(n868) );
  OAI21X1 OAI21X1_75 ( .A(_abc_40344_n996), .B(_abc_40344_n983), .C(_abc_40344_n1031), .Y(_abc_40344_n1032) );
  OAI21X1 OAI21X1_750 ( .A(_abc_40344_n1665), .B(_abc_40344_n3076), .C(_abc_40344_n1350), .Y(_abc_40344_n3635) );
  OAI21X1 OAI21X1_751 ( .A(_abc_40344_n3228), .B(_abc_40344_n3638), .C(_abc_40344_n3641), .Y(_abc_40344_n3642) );
  OAI21X1 OAI21X1_752 ( .A(_abc_40344_n3109), .B(_abc_40344_n1906), .C(_abc_40344_n3066), .Y(_abc_40344_n3643) );
  OAI21X1 OAI21X1_753 ( .A(REG2_REG_9_), .B(_abc_40344_n3066), .C(_abc_40344_n3643), .Y(_abc_40344_n3644) );
  OAI21X1 OAI21X1_754 ( .A(_abc_40344_n1359_1), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3645) );
  OAI21X1 OAI21X1_755 ( .A(_abc_40344_n3219), .B(_abc_40344_n3639), .C(_abc_40344_n3647), .Y(_abc_40344_n3648) );
  OAI21X1 OAI21X1_756 ( .A(_abc_40344_n3069), .B(_abc_40344_n3637), .C(_abc_40344_n3649), .Y(n863) );
  OAI21X1 OAI21X1_757 ( .A(_abc_40344_n3651), .B(_abc_40344_n3310), .C(_abc_40344_n2486), .Y(_abc_40344_n3652) );
  OAI21X1 OAI21X1_758 ( .A(_abc_40344_n3228), .B(_abc_40344_n3653), .C(_abc_40344_n3656), .Y(_abc_40344_n3657) );
  OAI21X1 OAI21X1_759 ( .A(_abc_40344_n1016), .B(_abc_40344_n1031), .C(_abc_40344_n3659), .Y(_abc_40344_n3660) );
  OAI21X1 OAI21X1_76 ( .A(_abc_40344_n910), .B(_abc_40344_n1033), .C(nRESET_G), .Y(_abc_40344_n1034_1) );
  OAI21X1 OAI21X1_760 ( .A(_abc_40344_n3219), .B(_abc_40344_n3654), .C(_abc_40344_n3661), .Y(_abc_40344_n3662_1) );
  OAI21X1 OAI21X1_761 ( .A(_abc_40344_n908), .B(_abc_40344_n3663), .C(_abc_40344_n1665), .Y(_abc_40344_n3664) );
  OAI21X1 OAI21X1_762 ( .A(_abc_40344_n1375), .B(_abc_40344_n3111), .C(_abc_40344_n3666), .Y(_abc_40344_n3667) );
  OAI21X1 OAI21X1_763 ( .A(_abc_40344_n714), .B(_abc_40344_n3074), .C(_abc_40344_n908), .Y(_abc_40344_n3670) );
  OAI21X1 OAI21X1_764 ( .A(_abc_40344_n3228), .B(_abc_40344_n3673), .C(_abc_40344_n3676), .Y(_abc_40344_n3677) );
  OAI21X1 OAI21X1_765 ( .A(_abc_40344_n1009), .B(_abc_40344_n1017), .C(_abc_40344_n3103), .Y(_abc_40344_n3678) );
  OAI21X1 OAI21X1_766 ( .A(_abc_40344_n922_1), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3679) );
  OAI21X1 OAI21X1_767 ( .A(_abc_40344_n3067), .B(_abc_40344_n3678), .C(_abc_40344_n3680), .Y(_abc_40344_n3681) );
  OAI21X1 OAI21X1_768 ( .A(_abc_40344_n3219), .B(_abc_40344_n3674), .C(_abc_40344_n3682_1), .Y(_abc_40344_n3683) );
  OAI21X1 OAI21X1_769 ( .A(_abc_40344_n3069), .B(_abc_40344_n3672), .C(_abc_40344_n3684), .Y(n853) );
  OAI21X1 OAI21X1_77 ( .A(_abc_40344_n1006), .B(_abc_40344_n1025), .C(_abc_40344_n1035), .Y(_abc_40344_n1036) );
  OAI21X1 OAI21X1_770 ( .A(_abc_40344_n1980), .B(_abc_40344_n3308), .C(_abc_40344_n2089), .Y(_abc_40344_n3691) );
  OAI21X1 OAI21X1_771 ( .A(_abc_40344_n1998), .B(_abc_40344_n3691), .C(_abc_40344_n2083), .Y(_abc_40344_n3692) );
  OAI21X1 OAI21X1_772 ( .A(_abc_40344_n3228), .B(_abc_40344_n3693), .C(_abc_40344_n3690), .Y(_abc_40344_n3694) );
  OAI21X1 OAI21X1_773 ( .A(_abc_40344_n923_1), .B(_abc_40344_n926), .C(_abc_40344_n3103), .Y(_abc_40344_n3695) );
  OAI21X1 OAI21X1_774 ( .A(_abc_40344_n1872), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3696) );
  OAI21X1 OAI21X1_775 ( .A(_abc_40344_n3067), .B(_abc_40344_n3695), .C(_abc_40344_n3697), .Y(_abc_40344_n3698) );
  OAI21X1 OAI21X1_776 ( .A(_abc_40344_n3219), .B(_abc_40344_n3688), .C(_abc_40344_n3699), .Y(_abc_40344_n3700) );
  OAI21X1 OAI21X1_777 ( .A(_abc_40344_n3069), .B(_abc_40344_n3687), .C(_abc_40344_n3701), .Y(n848) );
  OAI21X1 OAI21X1_778 ( .A(_abc_40344_n3142), .B(_abc_40344_n3704), .C(_abc_40344_n3145), .Y(_abc_40344_n3705) );
  OAI21X1 OAI21X1_779 ( .A(_abc_40344_n2482), .B(_abc_40344_n3691), .C(_abc_40344_n3227), .Y(_abc_40344_n3710) );
  OAI21X1 OAI21X1_78 ( .A(_abc_40344_n937), .B(_abc_40344_n994), .C(_abc_40344_n1037), .Y(n1331) );
  OAI21X1 OAI21X1_780 ( .A(_abc_40344_n3709), .B(_abc_40344_n3710), .C(_abc_40344_n3708), .Y(_abc_40344_n3711) );
  OAI21X1 OAI21X1_781 ( .A(_abc_40344_n777_1), .B(_abc_40344_n3072), .C(_abc_40344_n734), .Y(_abc_40344_n3717) );
  OAI21X1 OAI21X1_782 ( .A(_abc_40344_n738_1), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3719) );
  OAI21X1 OAI21X1_783 ( .A(_abc_40344_n756), .B(_abc_40344_n3066), .C(_abc_40344_n3720), .Y(_abc_40344_n3721) );
  OAI21X1 OAI21X1_784 ( .A(_abc_40344_n777_1), .B(_abc_40344_n3072), .C(_abc_40344_n3727_1), .Y(_abc_40344_n3728) );
  OAI21X1 OAI21X1_785 ( .A(_abc_40344_n3261), .B(_abc_40344_n3724), .C(_abc_40344_n3733), .Y(_abc_40344_n3734) );
  OAI21X1 OAI21X1_786 ( .A(_abc_40344_n3729), .B(_abc_40344_n3735), .C(_abc_40344_n3066), .Y(_abc_40344_n3736) );
  OAI21X1 OAI21X1_787 ( .A(_abc_40344_n2491), .B(_abc_40344_n3741), .C(_abc_40344_n3227), .Y(_abc_40344_n3742) );
  OAI21X1 OAI21X1_788 ( .A(_abc_40344_n3703), .B(_abc_40344_n3138), .C(_abc_40344_n3141), .Y(_abc_40344_n3743) );
  OAI21X1 OAI21X1_789 ( .A(_abc_40344_n3740), .B(_abc_40344_n3742), .C(_abc_40344_n3746), .Y(_abc_40344_n3747) );
  OAI21X1 OAI21X1_79 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_27_), .Y(_abc_40344_n1040) );
  OAI21X1 OAI21X1_790 ( .A(_abc_40344_n1609), .B(_abc_40344_n3071), .C(_abc_40344_n3748), .Y(_abc_40344_n3749_1) );
  OAI21X1 OAI21X1_791 ( .A(_abc_40344_n869), .B(_abc_40344_n864), .C(_abc_40344_n2632), .Y(_abc_40344_n3756) );
  OAI21X1 OAI21X1_792 ( .A(_abc_40344_n2546), .B(_abc_40344_n3756), .C(_abc_40344_n3227), .Y(_abc_40344_n3758) );
  OAI21X1 OAI21X1_793 ( .A(_abc_40344_n3757), .B(_abc_40344_n3758), .C(_abc_40344_n3760), .Y(_abc_40344_n3761) );
  OAI21X1 OAI21X1_794 ( .A(_abc_40344_n3062), .B(_abc_40344_n3763), .C(_abc_40344_n3762), .Y(_abc_40344_n3764) );
  OAI21X1 OAI21X1_795 ( .A(_abc_40344_n3764), .B(_abc_40344_n3761), .C(_abc_40344_n3066), .Y(_abc_40344_n3765) );
  OAI21X1 OAI21X1_796 ( .A(_abc_40344_n1854), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3767) );
  OAI21X1 OAI21X1_797 ( .A(_abc_40344_n2631), .B(_abc_40344_n2488), .C(_abc_40344_n3227), .Y(_abc_40344_n3771_1) );
  OAI21X1 OAI21X1_798 ( .A(_abc_40344_n3261), .B(_abc_40344_n3770_1), .C(_abc_40344_n3773_1), .Y(_abc_40344_n3774_1) );
  OAI21X1 OAI21X1_799 ( .A(_abc_40344_n869), .B(_abc_40344_n1797), .C(_abc_40344_n3776_1), .Y(_abc_40344_n3777_1) );
  OAI21X1 OAI21X1_8 ( .A(_abc_40344_n612), .B(_abc_40344_n615), .C(_abc_40344_n576), .Y(_abc_40344_n616) );
  OAI21X1 OAI21X1_80 ( .A(_abc_40344_n1041), .B(_abc_40344_n1065), .C(_abc_40344_n1042), .Y(_abc_40344_n1066_1) );
  OAI21X1 OAI21X1_800 ( .A(_abc_40344_n648), .B(_abc_40344_n3777_1), .C(_abc_40344_n3775_1), .Y(_abc_40344_n3778_1) );
  OAI21X1 OAI21X1_801 ( .A(_abc_40344_n3778_1), .B(_abc_40344_n3774_1), .C(_abc_40344_n3066), .Y(_abc_40344_n3779_1) );
  OAI21X1 OAI21X1_802 ( .A(_abc_40344_n1678), .B(_abc_40344_n1031), .C(nRESET_G), .Y(_abc_40344_n3781_1) );
  OAI21X1 OAI21X1_803 ( .A(_abc_40344_n984), .B(_abc_40344_n1002), .C(_abc_40344_n986), .Y(_abc_40344_n3785_1) );
  OAI21X1 OAI21X1_804 ( .A(_abc_40344_n859), .B(_abc_40344_n862), .C(_abc_40344_n3103), .Y(_abc_40344_n3786_1) );
  OAI21X1 OAI21X1_805 ( .A(_abc_40344_n986), .B(_abc_40344_n1797), .C(_abc_40344_n3786_1), .Y(_abc_40344_n3788_1) );
  OAI21X1 OAI21X1_806 ( .A(_abc_40344_n1027_1), .B(_abc_40344_n3787_1), .C(_abc_40344_n3788_1), .Y(_abc_40344_n3789_1) );
  OAI21X1 OAI21X1_807 ( .A(_abc_40344_n3785_1), .B(_abc_40344_n3784_1), .C(_abc_40344_n3789_1), .Y(_abc_40344_n3790_1) );
  OAI21X1 OAI21X1_808 ( .A(_abc_40344_n3857), .B(_abc_40344_n664), .C(_abc_40344_n3858_1), .Y(n333) );
  OAI21X1 OAI21X1_809 ( .A(_abc_40344_n662), .B(_abc_40344_n3861_1), .C(_abc_40344_n3862), .Y(_abc_40344_n3863) );
  OAI21X1 OAI21X1_81 ( .A(_abc_40344_n1069), .B(_abc_40344_n761_1), .C(_abc_40344_n1070), .Y(_abc_40344_n1071) );
  OAI21X1 OAI21X1_810 ( .A(_abc_40344_n3857), .B(_abc_40344_n665), .C(_abc_40344_n3864_1), .Y(n328) );
  OAI21X1 OAI21X1_811 ( .A(_abc_40344_n656), .B(_abc_40344_n660), .C(_abc_40344_n682), .Y(_abc_40344_n3866) );
  OAI21X1 OAI21X1_812 ( .A(_abc_40344_n670), .B(_abc_40344_n3861_1), .C(_abc_40344_n3867), .Y(_abc_40344_n3868_1) );
  OAI21X1 OAI21X1_813 ( .A(_abc_40344_n3857), .B(_abc_40344_n3866), .C(_abc_40344_n3869), .Y(n323) );
  OAI21X1 OAI21X1_814 ( .A(_abc_40344_n550_1), .B(_abc_40344_n595_1), .C(_abc_40344_n799), .Y(_abc_40344_n3874_1) );
  OAI21X1 OAI21X1_815 ( .A(_abc_40344_n2009), .B(_abc_40344_n1033), .C(_abc_40344_n3875), .Y(_abc_40344_n3876) );
  OAI21X1 OAI21X1_816 ( .A(_abc_40344_n3857), .B(_abc_40344_n3874_1), .C(_abc_40344_n3877_1), .Y(n313) );
  OAI21X1 OAI21X1_817 ( .A(_abc_40344_n554_1), .B(_abc_40344_n3861_1), .C(_abc_40344_n3880_1), .Y(_abc_40344_n3881) );
  OAI21X1 OAI21X1_818 ( .A(_abc_40344_n3857), .B(_abc_40344_n3879), .C(_abc_40344_n3882), .Y(n308) );
  OAI21X1 OAI21X1_819 ( .A(_abc_40344_n550_1), .B(_abc_40344_n552), .C(_abc_40344_n634), .Y(_abc_40344_n3884) );
  OAI21X1 OAI21X1_82 ( .A(_abc_40344_n921), .B(_abc_40344_n1068), .C(_abc_40344_n1072), .Y(_abc_40344_n1073) );
  OAI21X1 OAI21X1_820 ( .A(_abc_40344_n566), .B(_abc_40344_n3861_1), .C(_abc_40344_n3885), .Y(_abc_40344_n3886_1) );
  OAI21X1 OAI21X1_821 ( .A(_abc_40344_n3857), .B(_abc_40344_n3884), .C(_abc_40344_n3887), .Y(n303) );
  OAI21X1 OAI21X1_822 ( .A(IR_REG_24_), .B(_abc_40344_n550_1), .C(_abc_40344_n3856), .Y(_abc_40344_n3890_1) );
  OAI21X1 OAI21X1_823 ( .A(_abc_40344_n563_1), .B(_abc_40344_n3861_1), .C(_abc_40344_n3891), .Y(_abc_40344_n3892) );
  OAI21X1 OAI21X1_824 ( .A(_abc_40344_n3889), .B(_abc_40344_n3890_1), .C(_abc_40344_n3893_1), .Y(n298) );
  OAI21X1 OAI21X1_825 ( .A(_abc_40344_n523), .B(_abc_40344_n586), .C(_abc_40344_n3895), .Y(n293) );
  OAI21X1 OAI21X1_826 ( .A(_abc_40344_n620), .B(_abc_40344_n3861_1), .C(_abc_40344_n3898), .Y(_abc_40344_n3899) );
  OAI21X1 OAI21X1_827 ( .A(_abc_40344_n3857), .B(_abc_40344_n3897_1), .C(_abc_40344_n3900_1), .Y(n288) );
  OAI21X1 OAI21X1_828 ( .A(_abc_40344_n612), .B(_abc_40344_n3861_1), .C(_abc_40344_n3902), .Y(_abc_40344_n3903) );
  OAI21X1 OAI21X1_829 ( .A(_abc_40344_n3857), .B(_abc_40344_n616), .C(_abc_40344_n3904), .Y(n283) );
  OAI21X1 OAI21X1_83 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_23_), .Y(_abc_40344_n1083) );
  OAI21X1 OAI21X1_830 ( .A(_abc_40344_n544), .B(_abc_40344_n614), .C(_abc_40344_n3906), .Y(_abc_40344_n3907) );
  OAI21X1 OAI21X1_831 ( .A(_abc_40344_n613), .B(_abc_40344_n3861_1), .C(_abc_40344_n3908_1), .Y(_abc_40344_n3909) );
  OAI21X1 OAI21X1_832 ( .A(_abc_40344_n3857), .B(_abc_40344_n3907), .C(_abc_40344_n3910), .Y(n278) );
  OAI21X1 OAI21X1_833 ( .A(_abc_40344_n3857), .B(_abc_40344_n644), .C(_abc_40344_n3914), .Y(n273) );
  OAI21X1 OAI21X1_834 ( .A(_abc_40344_n1119), .B(_abc_40344_n3861_1), .C(_abc_40344_n3917), .Y(_abc_40344_n3918) );
  OAI21X1 OAI21X1_835 ( .A(_abc_40344_n3857), .B(_abc_40344_n3916), .C(_abc_40344_n3919), .Y(n268) );
  OAI21X1 OAI21X1_836 ( .A(_abc_40344_n3921), .B(_abc_40344_n3861_1), .C(_abc_40344_n3922), .Y(_abc_40344_n3923) );
  OAI21X1 OAI21X1_837 ( .A(_abc_40344_n3857), .B(_abc_40344_n1174), .C(_abc_40344_n3924), .Y(n263) );
  OAI21X1 OAI21X1_838 ( .A(_abc_40344_n1144), .B(_abc_40344_n3861_1), .C(_abc_40344_n3927), .Y(_abc_40344_n3928) );
  OAI21X1 OAI21X1_839 ( .A(_abc_40344_n3857), .B(_abc_40344_n3926), .C(_abc_40344_n3929), .Y(n258) );
  OAI21X1 OAI21X1_84 ( .A(_abc_40344_n1087), .B(_abc_40344_n759), .C(_abc_40344_n1088), .Y(_abc_40344_n1089) );
  OAI21X1 OAI21X1_840 ( .A(_abc_40344_n1198), .B(_abc_40344_n1033), .C(_abc_40344_n3931), .Y(_abc_40344_n3932) );
  OAI21X1 OAI21X1_841 ( .A(_abc_40344_n3857), .B(_abc_40344_n1194), .C(_abc_40344_n3933), .Y(n253) );
  OAI21X1 OAI21X1_842 ( .A(_abc_40344_n3935), .B(_abc_40344_n3861_1), .C(_abc_40344_n3936), .Y(_abc_40344_n3937) );
  OAI21X1 OAI21X1_843 ( .A(_abc_40344_n3857), .B(_abc_40344_n1219), .C(_abc_40344_n3938), .Y(n248) );
  OAI21X1 OAI21X1_844 ( .A(_abc_40344_n530), .B(_abc_40344_n3861_1), .C(_abc_40344_n3941), .Y(_abc_40344_n3942) );
  OAI21X1 OAI21X1_845 ( .A(_abc_40344_n3857), .B(_abc_40344_n3940), .C(_abc_40344_n3943), .Y(n243) );
  OAI21X1 OAI21X1_846 ( .A(_abc_40344_n3857), .B(_abc_40344_n1291), .C(_abc_40344_n3947), .Y(n238) );
  OAI21X1 OAI21X1_847 ( .A(_abc_40344_n3949), .B(_abc_40344_n3861_1), .C(_abc_40344_n3950), .Y(_abc_40344_n3951_1) );
  OAI21X1 OAI21X1_848 ( .A(_abc_40344_n3857), .B(_abc_40344_n1269), .C(_abc_40344_n3952), .Y(n233) );
  OAI21X1 OAI21X1_849 ( .A(_abc_40344_n1243), .B(_abc_40344_n3861_1), .C(_abc_40344_n3954), .Y(_abc_40344_n3955) );
  OAI21X1 OAI21X1_85 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_22_), .Y(_abc_40344_n1099) );
  OAI21X1 OAI21X1_850 ( .A(_abc_40344_n3857), .B(_abc_40344_n1323), .C(_abc_40344_n3956_1), .Y(n228) );
  OAI21X1 OAI21X1_851 ( .A(_abc_40344_n1345), .B(_abc_40344_n3861_1), .C(_abc_40344_n3959), .Y(_abc_40344_n3960) );
  OAI21X1 OAI21X1_852 ( .A(_abc_40344_n3857), .B(_abc_40344_n3958_1), .C(_abc_40344_n3961), .Y(n223) );
  OAI21X1 OAI21X1_853 ( .A(_abc_40344_n528), .B(_abc_40344_n3861_1), .C(_abc_40344_n3963), .Y(_abc_40344_n3964) );
  OAI21X1 OAI21X1_854 ( .A(_abc_40344_n3857), .B(_abc_40344_n1370), .C(_abc_40344_n3965), .Y(n218) );
  OAI21X1 OAI21X1_855 ( .A(_abc_40344_n902_1), .B(_abc_40344_n1033), .C(_abc_40344_n3967), .Y(_abc_40344_n3968) );
  OAI21X1 OAI21X1_856 ( .A(_abc_40344_n3857), .B(_abc_40344_n904), .C(_abc_40344_n3969), .Y(n213) );
  OAI21X1 OAI21X1_857 ( .A(_abc_40344_n701), .B(_abc_40344_n1033), .C(_abc_40344_n3971), .Y(_abc_40344_n3972_1) );
  OAI21X1 OAI21X1_858 ( .A(_abc_40344_n3857), .B(_abc_40344_n710_1), .C(_abc_40344_n3973), .Y(n208) );
  OAI21X1 OAI21X1_859 ( .A(_abc_40344_n728), .B(_abc_40344_n1033), .C(_abc_40344_n3975), .Y(_abc_40344_n3976) );
  OAI21X1 OAI21X1_86 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1120), .C(_abc_40344_n1121), .Y(_abc_40344_n1122) );
  OAI21X1 OAI21X1_860 ( .A(_abc_40344_n3857), .B(_abc_40344_n730), .C(_abc_40344_n3977), .Y(n203) );
  OAI21X1 OAI21X1_861 ( .A(_abc_40344_n2168), .B(_abc_40344_n1033), .C(_abc_40344_n3979_1), .Y(_abc_40344_n3980) );
  OAI21X1 OAI21X1_862 ( .A(_abc_40344_n3857), .B(_abc_40344_n771), .C(_abc_40344_n3981), .Y(n198) );
  OAI21X1 OAI21X1_863 ( .A(_abc_40344_n812), .B(_abc_40344_n1033), .C(_abc_40344_n3983), .Y(_abc_40344_n3984) );
  OAI21X1 OAI21X1_864 ( .A(_abc_40344_n795), .B(_abc_40344_n3857), .C(_abc_40344_n3985_1), .Y(n193) );
  OAI21X1 OAI21X1_865 ( .A(_abc_40344_n536), .B(_abc_40344_n3861_1), .C(_abc_40344_n3987), .Y(_abc_40344_n3988) );
  OAI21X1 OAI21X1_866 ( .A(_abc_40344_n821), .B(_abc_40344_n3857), .C(_abc_40344_n3989), .Y(n188) );
  OAI21X1 OAI21X1_867 ( .A(_abc_40344_n537_1), .B(_abc_40344_n3861_1), .C(_abc_40344_n3991), .Y(_abc_40344_n3992_1) );
  OAI21X1 OAI21X1_868 ( .A(_abc_40344_n523), .B(_abc_40344_n851), .C(_abc_40344_n3993), .Y(n183) );
  OAI21X1 OAI21X1_869 ( .A(_abc_40344_n877_1), .B(_abc_40344_n1033), .C(_abc_40344_n3995), .Y(n178) );
  OAI21X1 OAI21X1_87 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_18_), .Y(_abc_40344_n1123) );
  OAI21X1 OAI21X1_870 ( .A(_abc_40344_n1549), .B(_abc_40344_n1542), .C(_abc_40344_n1649), .Y(_abc_40344_n3999_1) );
  OAI21X1 OAI21X1_871 ( .A(_abc_40344_n2573_1), .B(_abc_40344_n705_1), .C(_abc_40344_n1550), .Y(_abc_40344_n4001) );
  OAI21X1 OAI21X1_872 ( .A(_abc_40344_n4011), .B(_abc_40344_n4012), .C(_abc_40344_n4013_1), .Y(_abc_40344_n4014) );
  OAI21X1 OAI21X1_873 ( .A(_abc_40344_n2098), .B(_abc_40344_n2557), .C(_abc_40344_n1904), .Y(_abc_40344_n4016) );
  OAI21X1 OAI21X1_874 ( .A(_abc_40344_n2391), .B(_abc_40344_n1630), .C(_abc_40344_n4000), .Y(_abc_40344_n4017) );
  OAI21X1 OAI21X1_875 ( .A(_abc_40344_n4019), .B(_abc_40344_n4010), .C(_abc_40344_n3066), .Y(_abc_40344_n4020_1) );
  OAI21X1 OAI21X1_876 ( .A(_abc_40344_n1031), .B(_abc_40344_n1640), .C(_abc_40344_n4025), .Y(_abc_40344_n4026_1) );
  OAI21X1 OAI21X1_877 ( .A(_abc_40344_n3219), .B(_abc_40344_n4024), .C(_abc_40344_n4027), .Y(_abc_40344_n4028) );
  OAI21X1 OAI21X1_878 ( .A(_abc_40344_n942), .B(_abc_40344_n561_1), .C(_abc_40344_n947), .Y(_abc_40344_n4032) );
  OAI21X1 OAI21X1_879 ( .A(_abc_40344_n4031), .B(_abc_40344_n3794_1), .C(_abc_40344_n4033_1), .Y(n338) );
  OAI21X1 OAI21X1_88 ( .A(_abc_40344_n802), .B(_abc_40344_n1122), .C(_abc_40344_n1123), .Y(_abc_40344_n1124) );
  OAI21X1 OAI21X1_880 ( .A(_abc_40344_n4035), .B(_abc_40344_n3794_1), .C(_abc_40344_n4036), .Y(n343) );
  OAI21X1 OAI21X1_881 ( .A(_abc_40344_n984), .B(_abc_40344_n987), .C(_abc_40344_n978), .Y(_abc_40344_n4038) );
  OAI21X1 OAI21X1_882 ( .A(_abc_40344_n4043), .B(_abc_40344_n4045), .C(_abc_40344_n4046_1), .Y(n498) );
  OAI21X1 OAI21X1_883 ( .A(_abc_40344_n4049), .B(_abc_40344_n3770_1), .C(_abc_40344_n4050), .Y(_abc_40344_n4051) );
  OAI21X1 OAI21X1_884 ( .A(_abc_40344_n4051), .B(_abc_40344_n3774_1), .C(_abc_40344_n4042), .Y(_abc_40344_n4052_1) );
  OAI21X1 OAI21X1_885 ( .A(_abc_40344_n857), .B(_abc_40344_n4042), .C(_abc_40344_n4053), .Y(n503) );
  OAI21X1 OAI21X1_886 ( .A(_abc_40344_n837), .B(_abc_40344_n4042), .C(_abc_40344_n4059), .Y(n508) );
  OAI21X1 OAI21X1_887 ( .A(_abc_40344_n4049), .B(_abc_40344_n3744), .C(_abc_40344_n4061), .Y(_abc_40344_n4062) );
  OAI21X1 OAI21X1_888 ( .A(_abc_40344_n4062), .B(_abc_40344_n3747), .C(_abc_40344_n4042), .Y(_abc_40344_n4063) );
  OAI21X1 OAI21X1_889 ( .A(_abc_40344_n2015), .B(_abc_40344_n4042), .C(_abc_40344_n4064_1), .Y(n513) );
  OAI21X1 OAI21X1_89 ( .A(_abc_40344_n1048), .B(_abc_40344_n1057), .C(_abc_40344_n1047), .Y(_abc_40344_n1126) );
  OAI21X1 OAI21X1_890 ( .A(_abc_40344_n4049), .B(_abc_40344_n3724), .C(_abc_40344_n3728), .Y(_abc_40344_n4066) );
  OAI21X1 OAI21X1_891 ( .A(_abc_40344_n4066), .B(_abc_40344_n3735), .C(_abc_40344_n4042), .Y(_abc_40344_n4067) );
  OAI21X1 OAI21X1_892 ( .A(_abc_40344_n980), .B(_abc_40344_n4041), .C(REG0_REG_4_), .Y(_abc_40344_n4068) );
  OAI21X1 OAI21X1_893 ( .A(_abc_40344_n751_1), .B(_abc_40344_n4042), .C(_abc_40344_n4072), .Y(n523) );
  OAI21X1 OAI21X1_894 ( .A(_abc_40344_n3726), .B(_abc_40344_n3687), .C(_abc_40344_n3695), .Y(_abc_40344_n4074) );
  OAI21X1 OAI21X1_895 ( .A(_abc_40344_n4076), .B(_abc_40344_n3694), .C(_abc_40344_n4042), .Y(_abc_40344_n4077_1) );
  OAI21X1 OAI21X1_896 ( .A(_abc_40344_n1987), .B(_abc_40344_n4042), .C(_abc_40344_n4078), .Y(n528) );
  OAI21X1 OAI21X1_897 ( .A(_abc_40344_n919), .B(_abc_40344_n3109), .C(_abc_40344_n3678), .Y(_abc_40344_n4080) );
  OAI21X1 OAI21X1_898 ( .A(_abc_40344_n4049), .B(_abc_40344_n3674), .C(_abc_40344_n4081), .Y(_abc_40344_n4082) );
  OAI21X1 OAI21X1_899 ( .A(_abc_40344_n4082), .B(_abc_40344_n3677), .C(_abc_40344_n4042), .Y(_abc_40344_n4083_1) );
  OAI21X1 OAI21X1_9 ( .A(_abc_40344_n559_1), .B(_abc_40344_n616), .C(_abc_40344_n617_1), .Y(_abc_40344_n618) );
  OAI21X1 OAI21X1_90 ( .A(_abc_40344_n921), .B(_abc_40344_n1128), .C(_abc_40344_n1129), .Y(_abc_40344_n1130) );
  OAI21X1 OAI21X1_900 ( .A(_abc_40344_n925), .B(_abc_40344_n4042), .C(_abc_40344_n4084), .Y(n533) );
  OAI21X1 OAI21X1_901 ( .A(_abc_40344_n3654), .B(_abc_40344_n4049), .C(_abc_40344_n4087), .Y(_abc_40344_n4088) );
  OAI21X1 OAI21X1_902 ( .A(_abc_40344_n4088), .B(_abc_40344_n3657), .C(_abc_40344_n4042), .Y(_abc_40344_n4089_1) );
  OAI21X1 OAI21X1_903 ( .A(_abc_40344_n1008), .B(_abc_40344_n4042), .C(_abc_40344_n4090), .Y(n538) );
  OAI21X1 OAI21X1_904 ( .A(_abc_40344_n4049), .B(_abc_40344_n3639), .C(_abc_40344_n4093), .Y(_abc_40344_n4094) );
  OAI21X1 OAI21X1_905 ( .A(_abc_40344_n4094), .B(_abc_40344_n3642), .C(_abc_40344_n4042), .Y(_abc_40344_n4095_1) );
  OAI21X1 OAI21X1_906 ( .A(_abc_40344_n1352), .B(_abc_40344_n4042), .C(_abc_40344_n4096), .Y(n543) );
  OAI21X1 OAI21X1_907 ( .A(_abc_40344_n3726), .B(_abc_40344_n4098), .C(_abc_40344_n3627), .Y(_abc_40344_n4099) );
  OAI21X1 OAI21X1_908 ( .A(_abc_40344_n1328), .B(_abc_40344_n4042), .C(_abc_40344_n4102), .Y(n548) );
  OAI21X1 OAI21X1_909 ( .A(_abc_40344_n3593), .B(_abc_40344_n4049), .C(_abc_40344_n4105), .Y(_abc_40344_n4106) );
  OAI21X1 OAI21X1_91 ( .A(_abc_40344_n559_1), .B(_abc_40344_n1146), .C(_abc_40344_n1147), .Y(_abc_40344_n1148) );
  OAI21X1 OAI21X1_910 ( .A(_abc_40344_n4106), .B(_abc_40344_n3600), .C(_abc_40344_n4042), .Y(_abc_40344_n4107_1) );
  OAI21X1 OAI21X1_911 ( .A(_abc_40344_n1282_1), .B(_abc_40344_n4042), .C(_abc_40344_n4108), .Y(n553) );
  OAI21X1 OAI21X1_912 ( .A(_abc_40344_n3726), .B(_abc_40344_n3576), .C(_abc_40344_n3585), .Y(_abc_40344_n4110) );
  OAI21X1 OAI21X1_913 ( .A(_abc_40344_n3584), .B(_abc_40344_n4049), .C(_abc_40344_n4111), .Y(_abc_40344_n4112) );
  OAI21X1 OAI21X1_914 ( .A(_abc_40344_n3583), .B(_abc_40344_n4112), .C(_abc_40344_n4042), .Y(_abc_40344_n4113_1) );
  OAI21X1 OAI21X1_915 ( .A(_abc_40344_n1297), .B(_abc_40344_n4042), .C(_abc_40344_n4114), .Y(n558) );
  OAI21X1 OAI21X1_916 ( .A(_abc_40344_n3726), .B(_abc_40344_n3558), .C(_abc_40344_n4117), .Y(_abc_40344_n4118) );
  OAI21X1 OAI21X1_917 ( .A(_abc_40344_n3566), .B(_abc_40344_n4119_1), .C(_abc_40344_n4042), .Y(_abc_40344_n4120) );
  OAI21X1 OAI21X1_918 ( .A(_abc_40344_n1253), .B(_abc_40344_n4042), .C(_abc_40344_n4121), .Y(n563) );
  OAI21X1 OAI21X1_919 ( .A(_abc_40344_n1209_1), .B(_abc_40344_n3232), .C(_abc_40344_n4123), .Y(_abc_40344_n4124) );
  OAI21X1 OAI21X1_92 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(_abc_40344_n1150), .Y(_abc_40344_n1151) );
  OAI21X1 OAI21X1_920 ( .A(_abc_40344_n3726), .B(_abc_40344_n3548), .C(_abc_40344_n4125_1), .Y(_abc_40344_n4126) );
  OAI21X1 OAI21X1_921 ( .A(_abc_40344_n3543), .B(_abc_40344_n4126), .C(_abc_40344_n4042), .Y(_abc_40344_n4127) );
  OAI21X1 OAI21X1_922 ( .A(_abc_40344_n980), .B(_abc_40344_n4041), .C(REG0_REG_14_), .Y(_abc_40344_n4128) );
  OAI21X1 OAI21X1_923 ( .A(_abc_40344_n1166_1), .B(_abc_40344_n1163), .C(_abc_40344_n3103), .Y(_abc_40344_n4130) );
  OAI21X1 OAI21X1_924 ( .A(_abc_40344_n3523), .B(_abc_40344_n4133), .C(_abc_40344_n4042), .Y(_abc_40344_n4134) );
  OAI21X1 OAI21X1_925 ( .A(_abc_40344_n980), .B(_abc_40344_n4041), .C(REG0_REG_15_), .Y(_abc_40344_n4135) );
  OAI21X1 OAI21X1_926 ( .A(_abc_40344_n1181), .B(_abc_40344_n1184), .C(_abc_40344_n3103), .Y(_abc_40344_n4137_1) );
  OAI21X1 OAI21X1_927 ( .A(_abc_40344_n4140), .B(_abc_40344_n3505), .C(_abc_40344_n4042), .Y(_abc_40344_n4141) );
  OAI21X1 OAI21X1_928 ( .A(_abc_40344_n980), .B(_abc_40344_n4041), .C(REG0_REG_16_), .Y(_abc_40344_n4142) );
  OAI21X1 OAI21X1_929 ( .A(_abc_40344_n3109), .B(_abc_40344_n1949), .C(_abc_40344_n3492), .Y(_abc_40344_n4146) );
  OAI21X1 OAI21X1_93 ( .A(_abc_40344_n802), .B(_abc_40344_n1149), .C(_abc_40344_n1151), .Y(_abc_40344_n1152_1) );
  OAI21X1 OAI21X1_930 ( .A(_abc_40344_n4144), .B(_abc_40344_n4042), .C(_abc_40344_n4149_1), .Y(n583) );
  OAI21X1 OAI21X1_931 ( .A(_abc_40344_n3460), .B(_abc_40344_n4049), .C(_abc_40344_n4151), .Y(_abc_40344_n4152) );
  OAI21X1 OAI21X1_932 ( .A(_abc_40344_n3464), .B(_abc_40344_n4152), .C(_abc_40344_n4042), .Y(_abc_40344_n4153) );
  OAI21X1 OAI21X1_933 ( .A(_abc_40344_n980), .B(_abc_40344_n4041), .C(REG0_REG_18_), .Y(_abc_40344_n4154) );
  OAI21X1 OAI21X1_934 ( .A(_abc_40344_n4049), .B(_abc_40344_n3455), .C(_abc_40344_n4159), .Y(_abc_40344_n4160) );
  OAI21X1 OAI21X1_935 ( .A(_abc_40344_n4160), .B(_abc_40344_n4156), .C(_abc_40344_n4042), .Y(_abc_40344_n4161) );
  OAI21X1 OAI21X1_936 ( .A(_abc_40344_n980), .B(_abc_40344_n4041), .C(REG0_REG_19_), .Y(_abc_40344_n4162) );
  OAI21X1 OAI21X1_937 ( .A(_abc_40344_n4049), .B(_abc_40344_n3433), .C(_abc_40344_n4165), .Y(_abc_40344_n4166) );
  OAI21X1 OAI21X1_938 ( .A(_abc_40344_n4166), .B(_abc_40344_n3436), .C(_abc_40344_n4042), .Y(_abc_40344_n4167_1) );
  OAI21X1 OAI21X1_939 ( .A(_abc_40344_n4049), .B(_abc_40344_n3413), .C(_abc_40344_n4171_1), .Y(_abc_40344_n4172) );
  OAI21X1 OAI21X1_94 ( .A(_abc_40344_n1154_1), .B(_abc_40344_n1156), .C(_abc_40344_n1155_1), .Y(_abc_40344_n1157) );
  OAI21X1 OAI21X1_940 ( .A(_abc_40344_n4172), .B(_abc_40344_n3415), .C(_abc_40344_n4042), .Y(_abc_40344_n4173_1) );
  OAI21X1 OAI21X1_941 ( .A(_abc_40344_n4049), .B(_abc_40344_n3380), .C(_abc_40344_n4176), .Y(_abc_40344_n4177_1) );
  OAI21X1 OAI21X1_942 ( .A(_abc_40344_n4043), .B(_abc_40344_n4179_1), .C(_abc_40344_n4180), .Y(n608) );
  OAI21X1 OAI21X1_943 ( .A(_abc_40344_n4185_1), .B(_abc_40344_n3369), .C(_abc_40344_n4042), .Y(_abc_40344_n4186) );
  OAI21X1 OAI21X1_944 ( .A(_abc_40344_n3726), .B(_abc_40344_n3342), .C(_abc_40344_n3343), .Y(_abc_40344_n4190) );
  OAI21X1 OAI21X1_945 ( .A(_abc_40344_n4191_1), .B(_abc_40344_n3339), .C(_abc_40344_n4042), .Y(_abc_40344_n4192) );
  OAI21X1 OAI21X1_946 ( .A(_abc_40344_n3283), .B(_abc_40344_n4049), .C(_abc_40344_n4196), .Y(_abc_40344_n4197_1) );
  OAI21X1 OAI21X1_947 ( .A(_abc_40344_n3287), .B(_abc_40344_n4197_1), .C(_abc_40344_n4042), .Y(_abc_40344_n4198) );
  OAI21X1 OAI21X1_948 ( .A(_abc_40344_n4049), .B(_abc_40344_n3266), .C(_abc_40344_n4202), .Y(_abc_40344_n4203_1) );
  OAI21X1 OAI21X1_949 ( .A(_abc_40344_n3270), .B(_abc_40344_n4203_1), .C(_abc_40344_n4042), .Y(_abc_40344_n4204) );
  OAI21X1 OAI21X1_95 ( .A(_abc_40344_n921), .B(_abc_40344_n1161), .C(_abc_40344_n1162), .Y(_abc_40344_n1163) );
  OAI21X1 OAI21X1_950 ( .A(_abc_40344_n4049), .B(_abc_40344_n3245), .C(_abc_40344_n4208), .Y(_abc_40344_n4209_1) );
  OAI21X1 OAI21X1_951 ( .A(_abc_40344_n4209_1), .B(_abc_40344_n3251), .C(_abc_40344_n4042), .Y(_abc_40344_n4210) );
  OAI21X1 OAI21X1_952 ( .A(_abc_40344_n4049), .B(_abc_40344_n3215), .C(_abc_40344_n4214), .Y(_abc_40344_n4215_1) );
  OAI21X1 OAI21X1_953 ( .A(_abc_40344_n3231), .B(_abc_40344_n4215_1), .C(_abc_40344_n4042), .Y(_abc_40344_n4216) );
  OAI21X1 OAI21X1_954 ( .A(_abc_40344_n4010), .B(_abc_40344_n4223_1), .C(_abc_40344_n4042), .Y(_abc_40344_n4224) );
  OAI21X1 OAI21X1_955 ( .A(_abc_40344_n3109), .B(_abc_40344_n1922), .C(_abc_40344_n3106), .Y(_abc_40344_n4228) );
  OAI21X1 OAI21X1_956 ( .A(_abc_40344_n4228), .B(_abc_40344_n4227_1), .C(_abc_40344_n4042), .Y(_abc_40344_n4229_1) );
  OAI21X1 OAI21X1_957 ( .A(_abc_40344_n3109), .B(_abc_40344_n1916), .C(_abc_40344_n3106), .Y(_abc_40344_n4233_1) );
  OAI21X1 OAI21X1_958 ( .A(_abc_40344_n4233_1), .B(_abc_40344_n4232), .C(_abc_40344_n4042), .Y(_abc_40344_n4234) );
  OAI21X1 OAI21X1_959 ( .A(_abc_40344_n980), .B(_abc_40344_n4041), .C(REG0_REG_31_), .Y(_abc_40344_n4235) );
  OAI21X1 OAI21X1_96 ( .A(IR_REG_16_), .B(_abc_40344_n1145), .C(IR_REG_17_), .Y(_abc_40344_n1173) );
  OAI21X1 OAI21X1_960 ( .A(_abc_40344_n4045), .B(_abc_40344_n4238_1), .C(_abc_40344_n4239_1), .Y(n658) );
  OAI21X1 OAI21X1_961 ( .A(_abc_40344_n4051), .B(_abc_40344_n3774_1), .C(_abc_40344_n4237), .Y(_abc_40344_n4241_1) );
  OAI21X1 OAI21X1_962 ( .A(_abc_40344_n860), .B(_abc_40344_n4237), .C(_abc_40344_n4242_1), .Y(n663) );
  OAI21X1 OAI21X1_963 ( .A(_abc_40344_n836), .B(_abc_40344_n4237), .C(_abc_40344_n4244_1), .Y(n668) );
  OAI21X1 OAI21X1_964 ( .A(_abc_40344_n4062), .B(_abc_40344_n3747), .C(_abc_40344_n4237), .Y(_abc_40344_n4246) );
  OAI21X1 OAI21X1_965 ( .A(_abc_40344_n2014), .B(_abc_40344_n4237), .C(_abc_40344_n4247_1), .Y(n673) );
  OAI21X1 OAI21X1_966 ( .A(_abc_40344_n4066), .B(_abc_40344_n3735), .C(_abc_40344_n4237), .Y(_abc_40344_n4249) );
  OAI21X1 OAI21X1_967 ( .A(_abc_40344_n2748), .B(_abc_40344_n4237), .C(_abc_40344_n4250_1), .Y(n678) );
  OAI21X1 OAI21X1_968 ( .A(_abc_40344_n757), .B(_abc_40344_n4237), .C(_abc_40344_n4252), .Y(n683) );
  OAI21X1 OAI21X1_969 ( .A(_abc_40344_n4076), .B(_abc_40344_n3694), .C(_abc_40344_n4237), .Y(_abc_40344_n4254_1) );
  OAI21X1 OAI21X1_97 ( .A(_abc_40344_n526), .B(_abc_40344_n677), .C(_abc_40344_n1173), .Y(_abc_40344_n1174) );
  OAI21X1 OAI21X1_970 ( .A(_abc_40344_n1989), .B(_abc_40344_n4237), .C(_abc_40344_n4255), .Y(n688) );
  OAI21X1 OAI21X1_971 ( .A(_abc_40344_n4082), .B(_abc_40344_n3677), .C(_abc_40344_n4237), .Y(_abc_40344_n4257_1) );
  OAI21X1 OAI21X1_972 ( .A(_abc_40344_n924), .B(_abc_40344_n4237), .C(_abc_40344_n4258), .Y(n693) );
  OAI21X1 OAI21X1_973 ( .A(_abc_40344_n4088), .B(_abc_40344_n3657), .C(_abc_40344_n4237), .Y(_abc_40344_n4260_1) );
  OAI21X1 OAI21X1_974 ( .A(_abc_40344_n1007), .B(_abc_40344_n4237), .C(_abc_40344_n4261), .Y(n698) );
  OAI21X1 OAI21X1_975 ( .A(_abc_40344_n4094), .B(_abc_40344_n3642), .C(_abc_40344_n4237), .Y(_abc_40344_n4263_1) );
  OAI21X1 OAI21X1_976 ( .A(_abc_40344_n1351), .B(_abc_40344_n4237), .C(_abc_40344_n4264), .Y(n703) );
  OAI21X1 OAI21X1_977 ( .A(_abc_40344_n1332), .B(_abc_40344_n4237), .C(_abc_40344_n4266_1), .Y(n708) );
  OAI21X1 OAI21X1_978 ( .A(_abc_40344_n4106), .B(_abc_40344_n3600), .C(_abc_40344_n4237), .Y(_abc_40344_n4268_1) );
  OAI21X1 OAI21X1_979 ( .A(_abc_40344_n1281), .B(_abc_40344_n4237), .C(_abc_40344_n4269_1), .Y(n713) );
  OAI21X1 OAI21X1_98 ( .A(IR_REG_31_), .B(IR_REG_17_), .C(_abc_40344_n1175), .Y(_abc_40344_n1176) );
  OAI21X1 OAI21X1_980 ( .A(_abc_40344_n3583), .B(_abc_40344_n4112), .C(_abc_40344_n4237), .Y(_abc_40344_n4271_1) );
  OAI21X1 OAI21X1_981 ( .A(_abc_40344_n1296), .B(_abc_40344_n4237), .C(_abc_40344_n4272_1), .Y(n718) );
  OAI21X1 OAI21X1_982 ( .A(_abc_40344_n3566), .B(_abc_40344_n4119_1), .C(_abc_40344_n4237), .Y(_abc_40344_n4274_1) );
  OAI21X1 OAI21X1_983 ( .A(_abc_40344_n1252), .B(_abc_40344_n4237), .C(_abc_40344_n4275_1), .Y(n723) );
  OAI21X1 OAI21X1_984 ( .A(_abc_40344_n3543), .B(_abc_40344_n4126), .C(_abc_40344_n4237), .Y(_abc_40344_n4277_1) );
  OAI21X1 OAI21X1_985 ( .A(_abc_40344_n1232), .B(_abc_40344_n4237), .C(_abc_40344_n4278_1), .Y(n728) );
  OAI21X1 OAI21X1_986 ( .A(_abc_40344_n3523), .B(_abc_40344_n4133), .C(_abc_40344_n4237), .Y(_abc_40344_n4280_1) );
  OAI21X1 OAI21X1_987 ( .A(_abc_40344_n1206), .B(_abc_40344_n4237), .C(_abc_40344_n4281_1), .Y(n733) );
  OAI21X1 OAI21X1_988 ( .A(_abc_40344_n4140), .B(_abc_40344_n3505), .C(_abc_40344_n4237), .Y(_abc_40344_n4283_1) );
  OAI21X1 OAI21X1_989 ( .A(_abc_40344_n1165), .B(_abc_40344_n4237), .C(_abc_40344_n4284_1), .Y(n738) );
  OAI21X1 OAI21X1_99 ( .A(_abc_40344_n603), .B(_abc_40344_n611_1), .C(DATAI_17_), .Y(_abc_40344_n1177) );
  OAI21X1 OAI21X1_990 ( .A(_abc_40344_n1183), .B(_abc_40344_n4237), .C(_abc_40344_n4286_1), .Y(n743) );
  OAI21X1 OAI21X1_991 ( .A(_abc_40344_n3464), .B(_abc_40344_n4152), .C(_abc_40344_n4237), .Y(_abc_40344_n4288) );
  OAI21X1 OAI21X1_992 ( .A(_abc_40344_n1132_1), .B(_abc_40344_n4237), .C(_abc_40344_n4289_1), .Y(n748) );
  OAI21X1 OAI21X1_993 ( .A(_abc_40344_n4160), .B(_abc_40344_n4156), .C(_abc_40344_n4237), .Y(_abc_40344_n4291) );
  OAI21X1 OAI21X1_994 ( .A(_abc_40344_n1412), .B(_abc_40344_n4237), .C(_abc_40344_n4292_1), .Y(n753) );
  OAI21X1 OAI21X1_995 ( .A(_abc_40344_n4166), .B(_abc_40344_n3436), .C(_abc_40344_n4237), .Y(_abc_40344_n4294) );
  OAI21X1 OAI21X1_996 ( .A(_abc_40344_n4172), .B(_abc_40344_n3415), .C(_abc_40344_n4237), .Y(_abc_40344_n4297) );
  OAI21X1 OAI21X1_997 ( .A(_abc_40344_n4238_1), .B(_abc_40344_n4179_1), .C(_abc_40344_n4300), .Y(n768) );
  OAI21X1 OAI21X1_998 ( .A(_abc_40344_n4185_1), .B(_abc_40344_n3369), .C(_abc_40344_n4237), .Y(_abc_40344_n4302_1) );
  OAI21X1 OAI21X1_999 ( .A(_abc_40344_n4191_1), .B(_abc_40344_n3339), .C(_abc_40344_n4237), .Y(_abc_40344_n4305_1) );
  OAI22X1 OAI22X1_1 ( .A(_abc_40344_n667), .B(_abc_40344_n753), .C(_abc_40344_n651_1), .D(_abc_40344_n752), .Y(_abc_40344_n754_1) );
  OAI22X1 OAI22X1_10 ( .A(_abc_40344_n633_1), .B(_abc_40344_n565_1), .C(D_REG_0_), .D(_abc_40344_n950), .Y(_abc_40344_n979) );
  OAI22X1 OAI22X1_100 ( .A(_abc_40344_n2403), .B(_abc_40344_n2405), .C(_abc_40344_n2409), .D(_abc_40344_n2408_1), .Y(_abc_40344_n2410) );
  OAI22X1 OAI22X1_101 ( .A(_abc_40344_n2216), .B(_abc_40344_n2215), .C(_abc_40344_n2433), .D(_abc_40344_n2434), .Y(_abc_40344_n2437) );
  OAI22X1 OAI22X1_102 ( .A(_abc_40344_n2252), .B(_abc_40344_n2251), .C(_abc_40344_n2236), .D(_abc_40344_n2235), .Y(_abc_40344_n2440) );
  OAI22X1 OAI22X1_103 ( .A(_abc_40344_n538_1), .B(_abc_40344_n603), .C(_abc_40344_n2681), .D(_abc_40344_n2682), .Y(_abc_40344_n2683) );
  OAI22X1 OAI22X1_104 ( .A(_abc_40344_n2679), .B(_abc_40344_n2683), .C(_abc_40344_n2677), .D(_abc_40344_n2684), .Y(_abc_40344_n2685) );
  OAI22X1 OAI22X1_105 ( .A(_abc_40344_n603), .B(_abc_40344_n774), .C(_abc_40344_n2667), .D(_abc_40344_n2756), .Y(_abc_40344_n2757) );
  OAI22X1 OAI22X1_106 ( .A(_abc_40344_n603), .B(_abc_40344_n917), .C(_abc_40344_n2806), .D(_abc_40344_n2808), .Y(_abc_40344_n2809) );
  OAI22X1 OAI22X1_107 ( .A(_abc_40344_n603), .B(_abc_40344_n1967), .C(_abc_40344_n2667), .D(_abc_40344_n2859), .Y(_abc_40344_n2860) );
  OAI22X1 OAI22X1_108 ( .A(_abc_40344_n603), .B(_abc_40344_n1196), .C(_abc_40344_n2667), .D(_abc_40344_n2966), .Y(_abc_40344_n2967) );
  OAI22X1 OAI22X1_109 ( .A(_abc_40344_n3052), .B(_abc_40344_n3058), .C(_abc_40344_n3056), .D(_abc_40344_n3051), .Y(_abc_40344_n3059) );
  OAI22X1 OAI22X1_11 ( .A(_abc_40344_n1008), .B(_abc_40344_n754_1), .C(_abc_40344_n1007), .D(_abc_40344_n761_1), .Y(_abc_40344_n1009) );
  OAI22X1 OAI22X1_110 ( .A(_abc_40344_n1440), .B(_abc_40344_n3379), .C(_abc_40344_n3261), .D(_abc_40344_n3380), .Y(_abc_40344_n3381) );
  OAI22X1 OAI22X1_111 ( .A(_abc_40344_n1031), .B(_abc_40344_n1104), .C(_abc_40344_n1090_1), .D(_abc_40344_n3244), .Y(_abc_40344_n3389) );
  OAI22X1 OAI22X1_112 ( .A(_abc_40344_n1031), .B(_abc_40344_n1693), .C(_abc_40344_n1110), .D(_abc_40344_n3244), .Y(_abc_40344_n3416) );
  OAI22X1 OAI22X1_113 ( .A(_abc_40344_n3109), .B(_abc_40344_n1421_1), .C(_abc_40344_n3232), .D(_abc_40344_n1440), .Y(_abc_40344_n3437) );
  OAI22X1 OAI22X1_114 ( .A(_abc_40344_n1031), .B(_abc_40344_n1408), .C(_abc_40344_n1429), .D(_abc_40344_n3244), .Y(_abc_40344_n3447) );
  OAI22X1 OAI22X1_115 ( .A(_abc_40344_n1138), .B(_abc_40344_n3379), .C(_abc_40344_n3261), .D(_abc_40344_n3455), .Y(_abc_40344_n3456) );
  OAI22X1 OAI22X1_116 ( .A(_abc_40344_n3109), .B(_abc_40344_n1137), .C(_abc_40344_n3232), .D(_abc_40344_n1414), .Y(_abc_40344_n3470) );
  OAI22X1 OAI22X1_117 ( .A(_abc_40344_n3067), .B(_abc_40344_n3585), .C(_abc_40344_n1259), .D(_abc_40344_n3244), .Y(_abc_40344_n3586) );
  OAI22X1 OAI22X1_118 ( .A(_abc_40344_n648), .B(_abc_40344_n3728), .C(_abc_40344_n3217), .D(_abc_40344_n3724), .Y(_abc_40344_n3729) );
  OAI22X1 OAI22X1_119 ( .A(_abc_40344_n763), .B(_abc_40344_n3232), .C(_abc_40344_n809), .D(_abc_40344_n3379), .Y(_abc_40344_n3732) );
  OAI22X1 OAI22X1_12 ( .A(_abc_40344_n1016), .B(_abc_40344_n921), .C(_abc_40344_n1010), .D(_abc_40344_n759), .Y(_abc_40344_n1017) );
  OAI22X1 OAI22X1_120 ( .A(_abc_40344_n648), .B(_abc_40344_n3749_1), .C(_abc_40344_n3217), .D(_abc_40344_n3744), .Y(_abc_40344_n3750) );
  OAI22X1 OAI22X1_121 ( .A(_abc_40344_n2095), .B(_abc_40344_n3104), .C(_abc_40344_n3379), .D(_abc_40344_n1550), .Y(_abc_40344_n3997) );
  OAI22X1 OAI22X1_122 ( .A(_abc_40344_n985), .B(_abc_40344_n627), .C(_abc_40344_n2657), .D(_abc_40344_n987), .Y(_abc_40344_n4044) );
  OAI22X1 OAI22X1_123 ( .A(_abc_40344_n1994), .B(_abc_40344_n3109), .C(_abc_40344_n4049), .D(_abc_40344_n3688), .Y(_abc_40344_n4075) );
  OAI22X1 OAI22X1_124 ( .A(_abc_40344_n3109), .B(_abc_40344_n1375), .C(_abc_40344_n1361), .D(_abc_40344_n3232), .Y(_abc_40344_n4086) );
  OAI22X1 OAI22X1_125 ( .A(_abc_40344_n3109), .B(_abc_40344_n1906), .C(_abc_40344_n1787), .D(_abc_40344_n3232), .Y(_abc_40344_n4092) );
  OAI22X1 OAI22X1_126 ( .A(_abc_40344_n3109), .B(_abc_40344_n1973), .C(_abc_40344_n1305), .D(_abc_40344_n3232), .Y(_abc_40344_n4104) );
  OAI22X1 OAI22X1_127 ( .A(_abc_40344_n3109), .B(_abc_40344_n1418), .C(_abc_40344_n3232), .D(_abc_40344_n1429), .Y(_abc_40344_n4158_1) );
  OAI22X1 OAI22X1_128 ( .A(_abc_40344_n3109), .B(_abc_40344_n1433), .C(_abc_40344_n3232), .D(_abc_40344_n1110), .Y(_abc_40344_n4170) );
  OAI22X1 OAI22X1_129 ( .A(_abc_40344_n3109), .B(_abc_40344_n1477), .C(_abc_40344_n3232), .D(_abc_40344_n1506), .Y(_abc_40344_n4195_1) );
  OAI22X1 OAI22X1_13 ( .A(_abc_40344_n922_1), .B(_abc_40344_n982), .C(_abc_40344_n1021), .D(_abc_40344_n1023_1), .Y(_abc_40344_n1024) );
  OAI22X1 OAI22X1_130 ( .A(_abc_40344_n3109), .B(_abc_40344_n1494), .C(_abc_40344_n3232), .D(_abc_40344_n1074), .Y(_abc_40344_n4201_1) );
  OAI22X1 OAI22X1_131 ( .A(_abc_40344_n3109), .B(_abc_40344_n1040), .C(_abc_40344_n3232), .D(_abc_40344_n1550), .Y(_abc_40344_n4207_1) );
  OAI22X1 OAI22X1_132 ( .A(_abc_40344_n3109), .B(_abc_40344_n1630), .C(_abc_40344_n3232), .D(_abc_40344_n1646), .Y(_abc_40344_n4213_1) );
  OAI22X1 OAI22X1_14 ( .A(_abc_40344_n745), .B(_abc_40344_n1040), .C(_abc_40344_n1039), .D(_abc_40344_n1074), .Y(_abc_40344_n1075) );
  OAI22X1 OAI22X1_15 ( .A(_abc_40344_n747), .B(_abc_40344_n1083), .C(_abc_40344_n745), .D(_abc_40344_n1090_1), .Y(_abc_40344_n1093) );
  OAI22X1 OAI22X1_16 ( .A(_abc_40344_n747), .B(_abc_40344_n1099), .C(_abc_40344_n745), .D(_abc_40344_n1110), .Y(_abc_40344_n1114) );
  OAI22X1 OAI22X1_17 ( .A(_abc_40344_n1132_1), .B(_abc_40344_n761_1), .C(_abc_40344_n1131), .D(_abc_40344_n759), .Y(_abc_40344_n1133) );
  OAI22X1 OAI22X1_18 ( .A(_abc_40344_n747), .B(_abc_40344_n1137), .C(_abc_40344_n745), .D(_abc_40344_n1138), .Y(_abc_40344_n1139) );
  OAI22X1 OAI22X1_19 ( .A(_abc_40344_n1165), .B(_abc_40344_n761_1), .C(_abc_40344_n1164), .D(_abc_40344_n759), .Y(_abc_40344_n1166_1) );
  OAI22X1 OAI22X1_2 ( .A(_abc_40344_n757), .B(_abc_40344_n761_1), .C(_abc_40344_n756), .D(_abc_40344_n759), .Y(_abc_40344_n762) );
  OAI22X1 OAI22X1_20 ( .A(_abc_40344_n747), .B(_abc_40344_n1152_1), .C(_abc_40344_n745), .D(_abc_40344_n1167), .Y(_abc_40344_n1170) );
  OAI22X1 OAI22X1_21 ( .A(_abc_40344_n1183), .B(_abc_40344_n761_1), .C(_abc_40344_n1182), .D(_abc_40344_n759), .Y(_abc_40344_n1184) );
  OAI22X1 OAI22X1_22 ( .A(_abc_40344_n1206), .B(_abc_40344_n761_1), .C(_abc_40344_n1207), .D(_abc_40344_n759), .Y(_abc_40344_n1208) );
  OAI22X1 OAI22X1_23 ( .A(_abc_40344_n745), .B(_abc_40344_n1209_1), .C(_abc_40344_n747), .D(_abc_40344_n1200), .Y(_abc_40344_n1212) );
  OAI22X1 OAI22X1_24 ( .A(_abc_40344_n1232), .B(_abc_40344_n761_1), .C(_abc_40344_n1231), .D(_abc_40344_n759), .Y(_abc_40344_n1233) );
  OAI22X1 OAI22X1_25 ( .A(_abc_40344_n1253), .B(_abc_40344_n754_1), .C(_abc_40344_n1252), .D(_abc_40344_n761_1), .Y(_abc_40344_n1254_1) );
  OAI22X1 OAI22X1_26 ( .A(_abc_40344_n1257), .B(_abc_40344_n921), .C(_abc_40344_n1255), .D(_abc_40344_n759), .Y(_abc_40344_n1258) );
  OAI22X1 OAI22X1_27 ( .A(_abc_40344_n745), .B(_abc_40344_n1259), .C(_abc_40344_n747), .D(_abc_40344_n1264), .Y(_abc_40344_n1265_1) );
  OAI22X1 OAI22X1_28 ( .A(_abc_40344_n1279), .B(_abc_40344_n921), .C(_abc_40344_n1274), .D(_abc_40344_n759), .Y(_abc_40344_n1280) );
  OAI22X1 OAI22X1_29 ( .A(_abc_40344_n1282_1), .B(_abc_40344_n754_1), .C(_abc_40344_n1281), .D(_abc_40344_n761_1), .Y(_abc_40344_n1283) );
  OAI22X1 OAI22X1_3 ( .A(_abc_40344_n745), .B(_abc_40344_n763), .C(_abc_40344_n747), .D(_abc_40344_n750), .Y(_abc_40344_n764) );
  OAI22X1 OAI22X1_30 ( .A(_abc_40344_n1297), .B(_abc_40344_n754_1), .C(_abc_40344_n1296), .D(_abc_40344_n761_1), .Y(_abc_40344_n1298) );
  OAI22X1 OAI22X1_31 ( .A(_abc_40344_n1039), .B(_abc_40344_n1305), .C(_abc_40344_n745), .D(_abc_40344_n1295), .Y(_abc_40344_n1306) );
  OAI22X1 OAI22X1_32 ( .A(_abc_40344_n1328), .B(_abc_40344_n754_1), .C(_abc_40344_n1330), .D(_abc_40344_n921), .Y(_abc_40344_n1331_1) );
  OAI22X1 OAI22X1_33 ( .A(_abc_40344_n1352), .B(_abc_40344_n754_1), .C(_abc_40344_n1351), .D(_abc_40344_n761_1), .Y(_abc_40344_n1353) );
  OAI22X1 OAI22X1_34 ( .A(_abc_40344_n1359_1), .B(_abc_40344_n921), .C(_abc_40344_n1354), .D(_abc_40344_n759), .Y(_abc_40344_n1360) );
  OAI22X1 OAI22X1_35 ( .A(_abc_40344_n745), .B(_abc_40344_n1375), .C(_abc_40344_n1018), .D(_abc_40344_n1039), .Y(_abc_40344_n1376) );
  OAI22X1 OAI22X1_36 ( .A(_abc_40344_n745), .B(_abc_40344_n1018), .C(_abc_40344_n747), .D(_abc_40344_n1375), .Y(_abc_40344_n1377) );
  OAI22X1 OAI22X1_37 ( .A(_abc_40344_n1412), .B(_abc_40344_n761_1), .C(_abc_40344_n1411), .D(_abc_40344_n759), .Y(_abc_40344_n1413) );
  OAI22X1 OAI22X1_38 ( .A(_abc_40344_n747), .B(_abc_40344_n1418), .C(_abc_40344_n745), .D(_abc_40344_n1414), .Y(_abc_40344_n1419) );
  OAI22X1 OAI22X1_39 ( .A(_abc_40344_n745), .B(_abc_40344_n1421_1), .C(_abc_40344_n1039), .D(_abc_40344_n1429), .Y(_abc_40344_n1430) );
  OAI22X1 OAI22X1_4 ( .A(_abc_40344_n745), .B(_abc_40344_n787_1), .C(_abc_40344_n776), .D(_abc_40344_n747), .Y(_abc_40344_n788) );
  OAI22X1 OAI22X1_40 ( .A(_abc_40344_n747), .B(_abc_40344_n1421_1), .C(_abc_40344_n745), .D(_abc_40344_n1429), .Y(_abc_40344_n1431) );
  OAI22X1 OAI22X1_41 ( .A(_abc_40344_n747), .B(_abc_40344_n1433), .C(_abc_40344_n745), .D(_abc_40344_n1440), .Y(_abc_40344_n1443) );
  OAI22X1 OAI22X1_42 ( .A(_abc_40344_n745), .B(_abc_40344_n1477), .C(_abc_40344_n1039), .D(_abc_40344_n1489), .Y(_abc_40344_n1490) );
  OAI22X1 OAI22X1_43 ( .A(_abc_40344_n747), .B(_abc_40344_n1494), .C(_abc_40344_n745), .D(_abc_40344_n1506), .Y(_abc_40344_n1509) );
  OAI22X1 OAI22X1_44 ( .A(_abc_40344_n1023_1), .B(_abc_40344_n1506), .C(_abc_40344_n1537), .D(_abc_40344_n1550), .Y(_abc_40344_n1551) );
  OAI22X1 OAI22X1_45 ( .A(_abc_40344_n1209_1), .B(_abc_40344_n1537), .C(_abc_40344_n1023_1), .D(_abc_40344_n1259), .Y(_abc_40344_n1565) );
  OAI22X1 OAI22X1_46 ( .A(_abc_40344_n1284), .B(_abc_40344_n1537), .C(_abc_40344_n1023_1), .D(_abc_40344_n1361), .Y(_abc_40344_n1593) );
  OAI22X1 OAI22X1_47 ( .A(_abc_40344_n787_1), .B(_abc_40344_n1537), .C(_abc_40344_n841), .D(_abc_40344_n1023_1), .Y(_abc_40344_n1605) );
  OAI22X1 OAI22X1_48 ( .A(_abc_40344_n1138), .B(_abc_40344_n1023_1), .C(_abc_40344_n1537), .D(_abc_40344_n1429), .Y(_abc_40344_n1622) );
  OAI22X1 OAI22X1_49 ( .A(_abc_40344_n747), .B(_abc_40344_n1630), .C(_abc_40344_n745), .D(_abc_40344_n1550), .Y(_abc_40344_n1631) );
  OAI22X1 OAI22X1_5 ( .A(_abc_40344_n837), .B(_abc_40344_n754_1), .C(_abc_40344_n836), .D(_abc_40344_n761_1), .Y(_abc_40344_n838) );
  OAI22X1 OAI22X1_50 ( .A(_abc_40344_n745), .B(_abc_40344_n1630), .C(_abc_40344_n1039), .D(_abc_40344_n1550), .Y(_abc_40344_n1632) );
  OAI22X1 OAI22X1_51 ( .A(_abc_40344_n1537), .B(_abc_40344_n1646), .C(_abc_40344_n1023_1), .D(_abc_40344_n1074), .Y(_abc_40344_n1647) );
  OAI22X1 OAI22X1_52 ( .A(_abc_40344_n927_1), .B(_abc_40344_n1023_1), .C(_abc_40344_n1537), .D(_abc_40344_n1361), .Y(_abc_40344_n1662) );
  OAI22X1 OAI22X1_53 ( .A(_abc_40344_n982), .B(_abc_40344_n1693), .C(_abc_40344_n1429), .D(_abc_40344_n1023_1), .Y(_abc_40344_n1694) );
  OAI22X1 OAI22X1_54 ( .A(_abc_40344_n1259), .B(_abc_40344_n1537), .C(_abc_40344_n1023_1), .D(_abc_40344_n1284), .Y(_abc_40344_n1709) );
  OAI22X1 OAI22X1_55 ( .A(_abc_40344_n1185), .B(_abc_40344_n1537), .C(_abc_40344_n1023_1), .D(_abc_40344_n1209_1), .Y(_abc_40344_n1736) );
  OAI22X1 OAI22X1_56 ( .A(_abc_40344_n1021), .B(_abc_40344_n1537), .C(_abc_40344_n787_1), .D(_abc_40344_n1023_1), .Y(_abc_40344_n1744) );
  OAI22X1 OAI22X1_57 ( .A(_abc_40344_n1138), .B(_abc_40344_n1537), .C(_abc_40344_n1023_1), .D(_abc_40344_n1167), .Y(_abc_40344_n1756) );
  OAI22X1 OAI22X1_58 ( .A(_abc_40344_n1023_1), .B(_abc_40344_n1090_1), .C(_abc_40344_n1537), .D(_abc_40344_n1489), .Y(_abc_40344_n1767) );
  OAI22X1 OAI22X1_59 ( .A(_abc_40344_n1018), .B(_abc_40344_n1023_1), .C(_abc_40344_n1537), .D(_abc_40344_n1787), .Y(_abc_40344_n1788) );
  OAI22X1 OAI22X1_6 ( .A(_abc_40344_n884), .B(_abc_40344_n754_1), .C(_abc_40344_n885), .D(_abc_40344_n761_1), .Y(_abc_40344_n886) );
  OAI22X1 OAI22X1_60 ( .A(_abc_40344_n1414), .B(_abc_40344_n1023_1), .C(_abc_40344_n1537), .D(_abc_40344_n1440), .Y(_abc_40344_n1811) );
  OAI22X1 OAI22X1_61 ( .A(_abc_40344_n1818), .B(_abc_40344_n1537), .C(_abc_40344_n1023_1), .D(_abc_40344_n1305), .Y(_abc_40344_n1819) );
  OAI22X1 OAI22X1_62 ( .A(_abc_40344_n1090_1), .B(_abc_40344_n1537), .C(_abc_40344_n1023_1), .D(_abc_40344_n1440), .Y(_abc_40344_n1834) );
  OAI22X1 OAI22X1_63 ( .A(_abc_40344_n809), .B(_abc_40344_n1537), .C(_abc_40344_n863), .D(_abc_40344_n1023_1), .Y(_abc_40344_n1853) );
  OAI22X1 OAI22X1_64 ( .A(_abc_40344_n1185), .B(_abc_40344_n1023_1), .C(_abc_40344_n1537), .D(_abc_40344_n1414), .Y(_abc_40344_n1863) );
  OAI22X1 OAI22X1_65 ( .A(_abc_40344_n763), .B(_abc_40344_n1023_1), .C(_abc_40344_n927_1), .D(_abc_40344_n1537), .Y(_abc_40344_n1871) );
  OAI22X1 OAI22X1_66 ( .A(_abc_40344_n1023_1), .B(_abc_40344_n1489), .C(_abc_40344_n1537), .D(_abc_40344_n1074), .Y(_abc_40344_n1886) );
  OAI22X1 OAI22X1_67 ( .A(_abc_40344_n1167), .B(_abc_40344_n1537), .C(_abc_40344_n1023_1), .D(_abc_40344_n1818), .Y(_abc_40344_n1898) );
  OAI22X1 OAI22X1_68 ( .A(_abc_40344_n1987), .B(_abc_40344_n754_1), .C(_abc_40344_n1872), .D(_abc_40344_n921), .Y(_abc_40344_n1988) );
  OAI22X1 OAI22X1_69 ( .A(_abc_40344_n1930), .B(_abc_40344_n1979), .C(_abc_40344_n1981), .D(_abc_40344_n2006), .Y(_abc_40344_n2007) );
  OAI22X1 OAI22X1_7 ( .A(_abc_40344_n922_1), .B(_abc_40344_n921), .C(_abc_40344_n920), .D(_abc_40344_n759), .Y(_abc_40344_n923_1) );
  OAI22X1 OAI22X1_70 ( .A(_abc_40344_n2015), .B(_abc_40344_n754_1), .C(_abc_40344_n2014), .D(_abc_40344_n761_1), .Y(_abc_40344_n2016) );
  OAI22X1 OAI22X1_71 ( .A(_abc_40344_n808), .B(_abc_40344_n2172), .C(_abc_40344_n2179), .D(_abc_40344_n813), .Y(_abc_40344_n2180) );
  OAI22X1 OAI22X1_72 ( .A(_abc_40344_n698), .B(_abc_40344_n2172), .C(_abc_40344_n2179), .D(_abc_40344_n714), .Y(_abc_40344_n2184) );
  OAI22X1 OAI22X1_73 ( .A(_abc_40344_n2184), .B(_abc_40344_n2183), .C(_abc_40344_n2186), .D(_abc_40344_n2189), .Y(_abc_40344_n2190) );
  OAI22X1 OAI22X1_74 ( .A(_abc_40344_n915_1), .B(_abc_40344_n2172), .C(_abc_40344_n2179), .D(_abc_40344_n908), .Y(_abc_40344_n2195) );
  OAI22X1 OAI22X1_75 ( .A(_abc_40344_n2191), .B(_abc_40344_n2192), .C(_abc_40344_n2195), .D(_abc_40344_n2194), .Y(_abc_40344_n2196) );
  OAI22X1 OAI22X1_76 ( .A(_abc_40344_n2207), .B(_abc_40344_n2208), .C(_abc_40344_n2199), .D(_abc_40344_n2206), .Y(_abc_40344_n2209) );
  OAI22X1 OAI22X1_77 ( .A(_abc_40344_n2172), .B(_abc_40344_n864), .C(_abc_40344_n2179), .D(_abc_40344_n856), .Y(_abc_40344_n2221) );
  OAI22X1 OAI22X1_78 ( .A(_abc_40344_n829_1), .B(_abc_40344_n2172), .C(_abc_40344_n2179), .D(_abc_40344_n825), .Y(_abc_40344_n2229) );
  OAI22X1 OAI22X1_79 ( .A(_abc_40344_n2242), .B(_abc_40344_n2241), .C(_abc_40344_n2246), .D(_abc_40344_n2247), .Y(_abc_40344_n2248) );
  OAI22X1 OAI22X1_8 ( .A(_abc_40344_n925), .B(_abc_40344_n754_1), .C(_abc_40344_n924), .D(_abc_40344_n761_1), .Y(_abc_40344_n926) );
  OAI22X1 OAI22X1_80 ( .A(_abc_40344_n2265), .B(_abc_40344_n2240), .C(_abc_40344_n2268), .D(_abc_40344_n2266), .Y(_abc_40344_n2269) );
  OAI22X1 OAI22X1_81 ( .A(_abc_40344_n2179), .B(_abc_40344_n1259), .C(_abc_40344_n585), .D(_abc_40344_n1305), .Y(_abc_40344_n2274) );
  OAI22X1 OAI22X1_82 ( .A(_abc_40344_n585), .B(_abc_40344_n1284), .C(_abc_40344_n2179), .D(_abc_40344_n1305), .Y(_abc_40344_n2278) );
  OAI22X1 OAI22X1_83 ( .A(_abc_40344_n2179), .B(_abc_40344_n1284), .C(_abc_40344_n585), .D(_abc_40344_n1787), .Y(_abc_40344_n2282) );
  OAI22X1 OAI22X1_84 ( .A(_abc_40344_n1234), .B(_abc_40344_n2172), .C(_abc_40344_n2179), .D(_abc_40344_n1224), .Y(_abc_40344_n2296) );
  OAI22X1 OAI22X1_85 ( .A(_abc_40344_n1209_1), .B(_abc_40344_n2179), .C(_abc_40344_n585), .D(_abc_40344_n1818), .Y(_abc_40344_n2301) );
  OAI22X1 OAI22X1_86 ( .A(_abc_40344_n2295), .B(_abc_40344_n2296), .C(_abc_40344_n2305), .D(_abc_40344_n2303), .Y(_abc_40344_n2306) );
  OAI22X1 OAI22X1_87 ( .A(_abc_40344_n585), .B(_abc_40344_n1209_1), .C(_abc_40344_n2179), .D(_abc_40344_n1167), .Y(_abc_40344_n2310) );
  OAI22X1 OAI22X1_88 ( .A(_abc_40344_n1185), .B(_abc_40344_n2179), .C(_abc_40344_n585), .D(_abc_40344_n1167), .Y(_abc_40344_n2317) );
  OAI22X1 OAI22X1_89 ( .A(_abc_40344_n585), .B(_abc_40344_n1185), .C(_abc_40344_n2179), .D(_abc_40344_n1138), .Y(_abc_40344_n2324) );
  OAI22X1 OAI22X1_9 ( .A(_abc_40344_n745), .B(_abc_40344_n927_1), .C(_abc_40344_n747), .D(_abc_40344_n919), .Y(_abc_40344_n928) );
  OAI22X1 OAI22X1_90 ( .A(_abc_40344_n2318), .B(_abc_40344_n2319), .C(_abc_40344_n2326), .D(_abc_40344_n2325), .Y(_abc_40344_n2327) );
  OAI22X1 OAI22X1_91 ( .A(_abc_40344_n585), .B(_abc_40344_n1138), .C(_abc_40344_n2179), .D(_abc_40344_n1414), .Y(_abc_40344_n2329) );
  OAI22X1 OAI22X1_92 ( .A(_abc_40344_n2161), .B(_abc_40344_n1421_1), .C(_abc_40344_n585), .D(_abc_40344_n1414), .Y(_abc_40344_n2336) );
  OAI22X1 OAI22X1_93 ( .A(_abc_40344_n2338), .B(_abc_40344_n2337), .C(_abc_40344_n2331_1), .D(_abc_40344_n2330), .Y(_abc_40344_n2339) );
  OAI22X1 OAI22X1_94 ( .A(_abc_40344_n2161), .B(_abc_40344_n1083), .C(_abc_40344_n585), .D(_abc_40344_n1110), .Y(_abc_40344_n2357) );
  OAI22X1 OAI22X1_95 ( .A(_abc_40344_n2358), .B(_abc_40344_n2359), .C(_abc_40344_n2367), .D(_abc_40344_n2366), .Y(_abc_40344_n2368) );
  OAI22X1 OAI22X1_96 ( .A(_abc_40344_n1491), .B(_abc_40344_n2179), .C(_abc_40344_n2172), .D(_abc_40344_n1488), .Y(_abc_40344_n2372) );
  OAI22X1 OAI22X1_97 ( .A(_abc_40344_n2377), .B(_abc_40344_n2379), .C(_abc_40344_n2385), .D(_abc_40344_n2383), .Y(_abc_40344_n2386) );
  OAI22X1 OAI22X1_98 ( .A(_abc_40344_n1649), .B(_abc_40344_n2179), .C(_abc_40344_n2172), .D(_abc_40344_n2391), .Y(_abc_40344_n2392) );
  OAI22X1 OAI22X1_99 ( .A(_abc_40344_n2396), .B(_abc_40344_n2398), .C(_abc_40344_n2390), .D(_abc_40344_n2392), .Y(_abc_40344_n2399) );
  OR2X2 OR2X2_1 ( .A(_abc_40344_n706), .B(IR_REG_4_), .Y(_abc_40344_n707_1) );
  OR2X2 OR2X2_10 ( .A(_abc_40344_n1060), .B(_abc_40344_n1046), .Y(_abc_40344_n1061) );
  OR2X2 OR2X2_11 ( .A(_abc_40344_n1058), .B(_abc_40344_n1047), .Y(_abc_40344_n1125) );
  OR2X2 OR2X2_12 ( .A(_abc_40344_n1130), .B(_abc_40344_n1133), .Y(_abc_40344_n1134) );
  OR2X2 OR2X2_13 ( .A(_abc_40344_n1230), .B(_abc_40344_n1233), .Y(_abc_40344_n1234) );
  OR2X2 OR2X2_14 ( .A(_abc_40344_n1266), .B(_abc_40344_n1262), .Y(_abc_40344_n1267) );
  OR2X2 OR2X2_15 ( .A(_abc_40344_n1288), .B(_abc_40344_n1286), .Y(_abc_40344_n1289) );
  OR2X2 OR2X2_16 ( .A(_abc_40344_n1311), .B(_abc_40344_n1306), .Y(_abc_40344_n1317_1) );
  OR2X2 OR2X2_17 ( .A(_abc_40344_n1334), .B(_abc_40344_n1331_1), .Y(_abc_40344_n1335) );
  OR2X2 OR2X2_18 ( .A(_abc_40344_n1444), .B(_abc_40344_n1442), .Y(_abc_40344_n1453) );
  OR2X2 OR2X2_19 ( .A(_abc_40344_n1063), .B(_abc_40344_n1043), .Y(_abc_40344_n1464) );
  OR2X2 OR2X2_2 ( .A(_abc_40344_n723), .B(_abc_40344_n720), .Y(_abc_40344_n725) );
  OR2X2 OR2X2_20 ( .A(_abc_40344_n1067), .B(_abc_40344_n1538), .Y(_abc_40344_n1640) );
  OR2X2 OR2X2_21 ( .A(_abc_40344_n1383_1), .B(_abc_40344_n1379), .Y(_abc_40344_n1655) );
  OR2X2 OR2X2_22 ( .A(_abc_40344_n1424), .B(_abc_40344_n1428), .Y(_abc_40344_n2037) );
  OR2X2 OR2X2_23 ( .A(_abc_40344_n2043), .B(_abc_40344_n1957), .Y(_abc_40344_n2044) );
  OR2X2 OR2X2_24 ( .A(_abc_40344_n1986), .B(_abc_40344_n2060), .Y(_abc_40344_n2061) );
  OR2X2 OR2X2_25 ( .A(_abc_40344_n2110), .B(_abc_40344_n2111), .Y(_abc_40344_n2112) );
  OR2X2 OR2X2_26 ( .A(_abc_40344_n2248), .B(_abc_40344_n2253_1), .Y(_abc_40344_n2254) );
  OR2X2 OR2X2_27 ( .A(_abc_40344_n2246), .B(_abc_40344_n2247), .Y(_abc_40344_n2270) );
  OR2X2 OR2X2_28 ( .A(_abc_40344_n2298), .B(_abc_40344_n2289), .Y(_abc_40344_n2299) );
  OR2X2 OR2X2_29 ( .A(IR_REG_31_), .B(IR_REG_19_), .Y(_abc_40344_n2416_1) );
  OR2X2 OR2X2_3 ( .A(_abc_40344_n764), .B(_abc_40344_n719), .Y(_abc_40344_n765) );
  OR2X2 OR2X2_30 ( .A(_abc_40344_n2506), .B(_abc_40344_n2499), .Y(_abc_40344_n2507) );
  OR2X2 OR2X2_31 ( .A(_abc_40344_n2038), .B(_abc_40344_n1954), .Y(_abc_40344_n2527) );
  OR2X2 OR2X2_32 ( .A(_abc_40344_n2546), .B(_abc_40344_n2545), .Y(_abc_40344_n2547) );
  OR2X2 OR2X2_33 ( .A(_abc_40344_n2557), .B(_abc_40344_n2098), .Y(_abc_40344_n2558) );
  OR2X2 OR2X2_34 ( .A(_abc_40344_n2125), .B(_abc_40344_n2151), .Y(_abc_40344_n2613) );
  OR2X2 OR2X2_35 ( .A(_abc_40344_n2608), .B(_abc_40344_n2621), .Y(_abc_40344_n2622) );
  OR2X2 OR2X2_36 ( .A(_abc_40344_n2643), .B(_abc_40344_n2644_1), .Y(_abc_40344_n2645) );
  OR2X2 OR2X2_37 ( .A(_abc_40344_n2826), .B(_abc_40344_n2820), .Y(n1022) );
  OR2X2 OR2X2_38 ( .A(_abc_40344_n2845), .B(REG1_REG_10_), .Y(_abc_40344_n2846) );
  OR2X2 OR2X2_39 ( .A(_abc_40344_n3099), .B(_abc_40344_n1916), .Y(_abc_40344_n3101) );
  OR2X2 OR2X2_4 ( .A(_abc_40344_n789), .B(_abc_40344_n786), .Y(_abc_40344_n791) );
  OR2X2 OR2X2_40 ( .A(_abc_40344_n3102), .B(_abc_40344_n3112), .Y(n973) );
  OR2X2 OR2X2_41 ( .A(_abc_40344_n3116), .B(_abc_40344_n3118), .Y(n968) );
  OR2X2 OR2X2_42 ( .A(_abc_40344_n3154), .B(_abc_40344_n3144), .Y(_abc_40344_n3155) );
  OR2X2 OR2X2_43 ( .A(_abc_40344_n3212), .B(_abc_40344_n3120), .Y(_abc_40344_n3214) );
  OR2X2 OR2X2_44 ( .A(_abc_40344_n3255), .B(_abc_40344_n3253), .Y(_abc_40344_n3256) );
  OR2X2 OR2X2_45 ( .A(_abc_40344_n3277), .B(_abc_40344_n3275), .Y(_abc_40344_n3278) );
  OR2X2 OR2X2_46 ( .A(_abc_40344_n3410), .B(_abc_40344_n3398), .Y(_abc_40344_n3412) );
  OR2X2 OR2X2_47 ( .A(_abc_40344_n3401), .B(_abc_40344_n3414), .Y(_abc_40344_n3415) );
  OR2X2 OR2X2_48 ( .A(_abc_40344_n3430), .B(_abc_40344_n2527), .Y(_abc_40344_n3431_1) );
  OR2X2 OR2X2_49 ( .A(_abc_40344_n3487), .B(_abc_40344_n3481), .Y(_abc_40344_n3488) );
  OR2X2 OR2X2_5 ( .A(_abc_40344_n883), .B(_abc_40344_n886), .Y(_abc_40344_n887) );
  OR2X2 OR2X2_50 ( .A(_abc_40344_n3734), .B(_abc_40344_n3731), .Y(_abc_40344_n3735) );
  OR2X2 OR2X2_51 ( .A(_abc_40344_n3219), .B(_abc_40344_n3770_1), .Y(_abc_40344_n3780_1) );
  OR2X2 OR2X2_52 ( .A(_abc_40344_n3198), .B(_abc_40344_n3202), .Y(_abc_40344_n4003) );
  OR2X2 OR2X2_53 ( .A(_abc_40344_n4075), .B(_abc_40344_n4074), .Y(_abc_40344_n4076) );
  OR2X2 OR2X2_54 ( .A(_abc_40344_n4118), .B(_abc_40344_n4116), .Y(_abc_40344_n4119_1) );
  OR2X2 OR2X2_55 ( .A(_abc_40344_n3456), .B(_abc_40344_n3454), .Y(_abc_40344_n4156) );
  OR2X2 OR2X2_56 ( .A(_abc_40344_n4189_1), .B(_abc_40344_n4190), .Y(_abc_40344_n4191_1) );
  OR2X2 OR2X2_6 ( .A(_abc_40344_n935_1), .B(_abc_40344_n932), .Y(_abc_40344_n936) );
  OR2X2 OR2X2_7 ( .A(_abc_40344_n991), .B(_abc_40344_n988), .Y(_abc_40344_n992) );
  OR2X2 OR2X2_8 ( .A(_abc_40344_n909), .B(_abc_40344_n1011), .Y(_abc_40344_n1014) );
  OR2X2 OR2X2_9 ( .A(_abc_40344_n1057), .B(_abc_40344_n1048), .Y(_abc_40344_n1058) );
  XNOR2X1 XNOR2X1_1 ( .A(_abc_40344_n709), .B(IR_REG_6_), .Y(_abc_40344_n710_1) );
  XNOR2X1 XNOR2X1_10 ( .A(_abc_40344_n1145), .B(_abc_40344_n1144), .Y(_abc_40344_n1146) );
  XNOR2X1 XNOR2X1_11 ( .A(_abc_40344_n1170), .B(_abc_40344_n720), .Y(_abc_40344_n1171) );
  XNOR2X1 XNOR2X1_12 ( .A(_abc_40344_n1189), .B(_abc_40344_n720), .Y(_abc_40344_n1190) );
  XNOR2X1 XNOR2X1_13 ( .A(_abc_40344_n1156), .B(REG3_REG_15_), .Y(_abc_40344_n1202) );
  XNOR2X1 XNOR2X1_14 ( .A(_abc_40344_n1212), .B(_abc_40344_n719), .Y(_abc_40344_n1213) );
  XNOR2X1 XNOR2X1_15 ( .A(_abc_40344_n574), .B(IR_REG_14_), .Y(_abc_40344_n1218) );
  XNOR2X1 XNOR2X1_16 ( .A(_abc_40344_n1236), .B(_abc_40344_n720), .Y(_abc_40344_n1237) );
  XNOR2X1 XNOR2X1_17 ( .A(_abc_40344_n1055), .B(REG3_REG_13_), .Y(_abc_40344_n1256) );
  XNOR2X1 XNOR2X1_18 ( .A(_abc_40344_n1265_1), .B(_abc_40344_n719), .Y(_abc_40344_n1266) );
  XNOR2X1 XNOR2X1_19 ( .A(_abc_40344_n1268), .B(IR_REG_11_), .Y(_abc_40344_n1269) );
  XNOR2X1 XNOR2X1_2 ( .A(_abc_40344_n788), .B(_abc_40344_n720), .Y(_abc_40344_n789) );
  XNOR2X1 XNOR2X1_20 ( .A(_abc_40344_n1287), .B(_abc_40344_n719), .Y(_abc_40344_n1288) );
  XNOR2X1 XNOR2X1_21 ( .A(_abc_40344_n1310), .B(_abc_40344_n720), .Y(_abc_40344_n1311) );
  XNOR2X1 XNOR2X1_22 ( .A(_abc_40344_n1051_1), .B(_abc_40344_n1052_1), .Y(_abc_40344_n1329) );
  XNOR2X1 XNOR2X1_23 ( .A(_abc_40344_n1337), .B(_abc_40344_n719), .Y(_abc_40344_n1338) );
  XNOR2X1 XNOR2X1_24 ( .A(_abc_40344_n1365), .B(_abc_40344_n720), .Y(_abc_40344_n1366) );
  XNOR2X1 XNOR2X1_25 ( .A(_abc_40344_n1377), .B(_abc_40344_n719), .Y(_abc_40344_n1378) );
  XNOR2X1 XNOR2X1_26 ( .A(_abc_40344_n1419), .B(_abc_40344_n719), .Y(_abc_40344_n1420) );
  XNOR2X1 XNOR2X1_27 ( .A(_abc_40344_n1431), .B(_abc_40344_n719), .Y(_abc_40344_n1432) );
  XNOR2X1 XNOR2X1_28 ( .A(_abc_40344_n1443), .B(_abc_40344_n720), .Y(_abc_40344_n1444) );
  XNOR2X1 XNOR2X1_29 ( .A(_abc_40344_n1474), .B(_abc_40344_n720), .Y(_abc_40344_n1475) );
  XNOR2X1 XNOR2X1_3 ( .A(_abc_40344_n1077), .B(_abc_40344_n720), .Y(_abc_40344_n1078_1) );
  XNOR2X1 XNOR2X1_30 ( .A(_abc_40344_n1492), .B(_abc_40344_n720), .Y(_abc_40344_n1493) );
  XNOR2X1 XNOR2X1_31 ( .A(_abc_40344_n1509), .B(_abc_40344_n720), .Y(_abc_40344_n1510) );
  XNOR2X1 XNOR2X1_32 ( .A(_abc_40344_n1632), .B(_abc_40344_n720), .Y(_abc_40344_n1633) );
  XNOR2X1 XNOR2X1_33 ( .A(_abc_40344_n1633), .B(_abc_40344_n1631), .Y(_abc_40344_n1634) );
  XNOR2X1 XNOR2X1_34 ( .A(_abc_40344_n1656), .B(_abc_40344_n1742), .Y(_abc_40344_n1743) );
  XNOR2X1 XNOR2X1_35 ( .A(_abc_40344_n889), .B(_abc_40344_n720), .Y(_abc_40344_n1795) );
  XNOR2X1 XNOR2X1_36 ( .A(_abc_40344_n1798), .B(_abc_40344_n720), .Y(_abc_40344_n1799) );
  XNOR2X1 XNOR2X1_37 ( .A(_abc_40344_n1795), .B(_abc_40344_n1799), .Y(_abc_40344_n1800) );
  XNOR2X1 XNOR2X1_38 ( .A(_abc_40344_n900), .B(_abc_40344_n1869), .Y(_abc_40344_n1870) );
  XNOR2X1 XNOR2X1_39 ( .A(_abc_40344_n823), .B(REG1_REG_2_), .Y(_abc_40344_n2720) );
  XNOR2X1 XNOR2X1_4 ( .A(_abc_40344_n1085), .B(REG3_REG_23_), .Y(_abc_40344_n1086) );
  XNOR2X1 XNOR2X1_40 ( .A(_abc_40344_n2720), .B(_abc_40344_n2721), .Y(_abc_40344_n2722_1) );
  XNOR2X1 XNOR2X1_41 ( .A(_abc_40344_n773), .B(_abc_40344_n2748), .Y(_abc_40344_n2749) );
  XNOR2X1 XNOR2X1_42 ( .A(_abc_40344_n2762), .B(REG1_REG_5_), .Y(_abc_40344_n2763) );
  XNOR2X1 XNOR2X1_43 ( .A(_abc_40344_n732_1), .B(REG2_REG_5_), .Y(_abc_40344_n2766) );
  XNOR2X1 XNOR2X1_44 ( .A(_abc_40344_n1372), .B(_abc_40344_n1010), .Y(_abc_40344_n2822) );
  XNOR2X1 XNOR2X1_45 ( .A(_abc_40344_n2823_1), .B(_abc_40344_n2822), .Y(_abc_40344_n2824) );
  XNOR2X1 XNOR2X1_46 ( .A(_abc_40344_n1347), .B(_abc_40344_n1354), .Y(_abc_40344_n2829) );
  XNOR2X1 XNOR2X1_47 ( .A(_abc_40344_n2838), .B(_abc_40344_n2837), .Y(_abc_40344_n2839) );
  XNOR2X1 XNOR2X1_48 ( .A(_abc_40344_n2858), .B(_abc_40344_n2856), .Y(_abc_40344_n2859) );
  XNOR2X1 XNOR2X1_49 ( .A(_abc_40344_n2868), .B(_abc_40344_n2867), .Y(_abc_40344_n2869) );
  XNOR2X1 XNOR2X1_5 ( .A(_abc_40344_n1093), .B(_abc_40344_n719), .Y(_abc_40344_n1094) );
  XNOR2X1 XNOR2X1_50 ( .A(_abc_40344_n2888), .B(_abc_40344_n2885), .Y(_abc_40344_n2889) );
  XNOR2X1 XNOR2X1_51 ( .A(_abc_40344_n2895), .B(_abc_40344_n2893), .Y(_abc_40344_n2896) );
  XNOR2X1 XNOR2X1_52 ( .A(_abc_40344_n2908), .B(_abc_40344_n1249), .Y(_abc_40344_n2909) );
  XNOR2X1 XNOR2X1_53 ( .A(_abc_40344_n2916), .B(_abc_40344_n2913), .Y(_abc_40344_n2917) );
  XNOR2X1 XNOR2X1_54 ( .A(_abc_40344_n2965), .B(_abc_40344_n2963), .Y(_abc_40344_n2966) );
  XNOR2X1 XNOR2X1_55 ( .A(_abc_40344_n3211), .B(_abc_40344_n2512), .Y(_abc_40344_n3245) );
  XNOR2X1 XNOR2X1_56 ( .A(_abc_40344_n2512), .B(_abc_40344_n2001), .Y(_abc_40344_n3248) );
  XNOR2X1 XNOR2X1_57 ( .A(_abc_40344_n3095), .B(_abc_40344_n1076), .Y(_abc_40344_n3252) );
  XNOR2X1 XNOR2X1_58 ( .A(_abc_40344_n3265), .B(_abc_40344_n2469), .Y(_abc_40344_n3266) );
  XNOR2X1 XNOR2X1_59 ( .A(_abc_40344_n3272), .B(_abc_40344_n1477), .Y(_abc_40344_n3291) );
  XNOR2X1 XNOR2X1_6 ( .A(_abc_40344_n1103_1), .B(_abc_40344_n1101), .Y(_abc_40344_n1104) );
  XNOR2X1 XNOR2X1_60 ( .A(_abc_40344_n3198), .B(_abc_40344_n2521), .Y(_abc_40344_n3296) );
  XNOR2X1 XNOR2X1_61 ( .A(_abc_40344_n3197), .B(_abc_40344_n2524), .Y(_abc_40344_n3351) );
  XNOR2X1 XNOR2X1_62 ( .A(_abc_40344_n3091), .B(_abc_40344_n1083), .Y(_abc_40344_n3372) );
  XNOR2X1 XNOR2X1_63 ( .A(_abc_40344_n3195), .B(_abc_40344_n2516), .Y(_abc_40344_n3380) );
  XNOR2X1 XNOR2X1_64 ( .A(_abc_40344_n3386), .B(_abc_40344_n1433), .Y(_abc_40344_n3396) );
  XNOR2X1 XNOR2X1_65 ( .A(_abc_40344_n3408), .B(_abc_40344_n2472), .Y(_abc_40344_n3445) );
  XNOR2X1 XNOR2X1_66 ( .A(_abc_40344_n3086), .B(_abc_40344_n1418), .Y(_abc_40344_n3446) );
  XNOR2X1 XNOR2X1_67 ( .A(_abc_40344_n3406), .B(_abc_40344_n2526), .Y(_abc_40344_n3459) );
  XNOR2X1 XNOR2X1_68 ( .A(_abc_40344_n3461), .B(_abc_40344_n2526), .Y(_abc_40344_n3462) );
  XNOR2X1 XNOR2X1_69 ( .A(_abc_40344_n3479), .B(_abc_40344_n3478_1), .Y(_abc_40344_n3480) );
  XNOR2X1 XNOR2X1_7 ( .A(_abc_40344_n1114), .B(_abc_40344_n719), .Y(_abc_40344_n1115) );
  XNOR2X1 XNOR2X1_70 ( .A(_abc_40344_n3465), .B(_abc_40344_n1178), .Y(_abc_40344_n3490) );
  XNOR2X1 XNOR2X1_71 ( .A(_abc_40344_n3176), .B(_abc_40344_n2503), .Y(_abc_40344_n3500) );
  XNOR2X1 XNOR2X1_72 ( .A(_abc_40344_n3503), .B(_abc_40344_n2503), .Y(_abc_40344_n3504) );
  XNOR2X1 XNOR2X1_73 ( .A(_abc_40344_n3483), .B(_abc_40344_n2480), .Y(_abc_40344_n3539) );
  XNOR2X1 XNOR2X1_74 ( .A(_abc_40344_n3563), .B(_abc_40344_n2545), .Y(_abc_40344_n3564) );
  XNOR2X1 XNOR2X1_75 ( .A(_abc_40344_n3159), .B(_abc_40344_n2484_1), .Y(_abc_40344_n3593) );
  XNOR2X1 XNOR2X1_76 ( .A(_abc_40344_n3313), .B(_abc_40344_n2536), .Y(_abc_40344_n3638) );
  XNOR2X1 XNOR2X1_77 ( .A(_abc_40344_n3616), .B(_abc_40344_n2536), .Y(_abc_40344_n3639) );
  XNOR2X1 XNOR2X1_78 ( .A(_abc_40344_n3652), .B(_abc_40344_n2532), .Y(_abc_40344_n3653) );
  XNOR2X1 XNOR2X1_79 ( .A(_abc_40344_n3614), .B(_abc_40344_n2532), .Y(_abc_40344_n3654) );
  XNOR2X1 XNOR2X1_8 ( .A(_abc_40344_n544), .B(_abc_40344_n1119), .Y(_abc_40344_n1120) );
  XNOR2X1 XNOR2X1_80 ( .A(_abc_40344_n3155), .B(_abc_40344_n2477), .Y(_abc_40344_n3688) );
  XNOR2X1 XNOR2X1_81 ( .A(_abc_40344_n3692), .B(_abc_40344_n2477), .Y(_abc_40344_n3693) );
  XNOR2X1 XNOR2X1_82 ( .A(_abc_40344_n3706_1), .B(_abc_40344_n2483), .Y(_abc_40344_n3707) );
  XNOR2X1 XNOR2X1_83 ( .A(_abc_40344_n3705), .B(_abc_40344_n2499), .Y(_abc_40344_n3724) );
  XNOR2X1 XNOR2X1_84 ( .A(_abc_40344_n3308), .B(_abc_40344_n2499), .Y(_abc_40344_n3730) );
  XNOR2X1 XNOR2X1_85 ( .A(_abc_40344_n3070), .B(_abc_40344_n825), .Y(_abc_40344_n3763) );
  XNOR2X1 XNOR2X1_86 ( .A(_abc_40344_n2488), .B(_abc_40344_n3136), .Y(_abc_40344_n3770_1) );
  XNOR2X1 XNOR2X1_9 ( .A(_abc_40344_n1139), .B(_abc_40344_n719), .Y(_abc_40344_n1140) );
  XOR2X1 XOR2X1_1 ( .A(_abc_40344_n816), .B(_abc_40344_n818_1), .Y(_abc_40344_n1599) );
  XOR2X1 XOR2X1_10 ( .A(_abc_40344_n2875), .B(_abc_40344_n2874), .Y(_abc_40344_n2876) );
  XOR2X1 XOR2X1_11 ( .A(_abc_40344_n2976), .B(_abc_40344_n2974), .Y(_abc_40344_n2977) );
  XOR2X1 XOR2X1_12 ( .A(_abc_40344_n3023), .B(_abc_40344_n3019), .Y(_abc_40344_n3024) );
  XOR2X1 XOR2X1_13 ( .A(_abc_40344_n3267), .B(_abc_40344_n2469), .Y(_abc_40344_n3268) );
  XOR2X1 XOR2X1_14 ( .A(_abc_40344_n3263), .B(_abc_40344_n2514), .Y(_abc_40344_n3283) );
  XOR2X1 XOR2X1_15 ( .A(_abc_40344_n3519), .B(_abc_40344_n2538), .Y(_abc_40344_n3520) );
  XOR2X1 XOR2X1_16 ( .A(_abc_40344_n3502), .B(_abc_40344_n2538), .Y(_abc_40344_n3522) );
  XOR2X1 XOR2X1_17 ( .A(_abc_40344_n3540), .B(_abc_40344_n2480), .Y(_abc_40344_n3541) );
  XOR2X1 XOR2X1_18 ( .A(_abc_40344_n3562), .B(_abc_40344_n3580), .Y(_abc_40344_n3581_1) );
  XOR2X1 XOR2X1_19 ( .A(_abc_40344_n3598), .B(_abc_40344_n2484_1), .Y(_abc_40344_n3599) );
  XOR2X1 XOR2X1_2 ( .A(_abc_40344_n1603), .B(_abc_40344_n1599), .Y(_abc_40344_n1604) );
  XOR2X1 XOR2X1_20 ( .A(_abc_40344_n3596), .B(_abc_40344_n2494), .Y(_abc_40344_n3610) );
  XOR2X1 XOR2X1_21 ( .A(_abc_40344_n3618), .B(_abc_40344_n2494), .Y(_abc_40344_n3619) );
  XOR2X1 XOR2X1_22 ( .A(_abc_40344_n3310), .B(_abc_40344_n2487), .Y(_abc_40344_n3673) );
  XOR2X1 XOR2X1_23 ( .A(_abc_40344_n3613), .B(_abc_40344_n2487), .Y(_abc_40344_n3674) );
  XOR2X1 XOR2X1_24 ( .A(_abc_40344_n3743), .B(_abc_40344_n2491), .Y(_abc_40344_n3744) );
  XOR2X1 XOR2X1_25 ( .A(_abc_40344_n3138), .B(_abc_40344_n2546), .Y(_abc_40344_n3759) );
  XOR2X1 XOR2X1_3 ( .A(_abc_40344_n1773), .B(_abc_40344_n1774), .Y(_abc_40344_n1775) );
  XOR2X1 XOR2X1_4 ( .A(_abc_40344_n1600), .B(_abc_40344_n1851), .Y(_abc_40344_n1852) );
  XOR2X1 XOR2X1_5 ( .A(_abc_40344_n2732), .B(_abc_40344_n2731), .Y(_abc_40344_n2733) );
  XOR2X1 XOR2X1_6 ( .A(_abc_40344_n2755), .B(_abc_40344_n2754), .Y(_abc_40344_n2756) );
  XOR2X1 XOR2X1_7 ( .A(_abc_40344_n2778), .B(_abc_40344_n2781), .Y(_abc_40344_n2782) );
  XOR2X1 XOR2X1_8 ( .A(_abc_40344_n2788), .B(_abc_40344_n2786), .Y(_abc_40344_n2789) );
  XOR2X1 XOR2X1_9 ( .A(_abc_40344_n2797), .B(_abc_40344_n2800), .Y(_abc_40344_n2801) );
endmodule