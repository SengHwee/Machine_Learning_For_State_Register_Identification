module fpSqrt(rst, clk, ce, ld, \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] , \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] , \o[24] , \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] , \o[32] , \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] , \o[40] , \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] , \o[48] , \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] , \o[56] , \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63] , \o[64] , \o[65] , \o[66] , \o[67] , \o[68] , \o[69] , \o[70] , \o[71] , \o[72] , \o[73] , \o[74] , \o[75] , \o[76] , \o[77] , \o[78] , \o[79] , \o[80] , \o[81] , \o[82] , \o[83] , \o[84] , \o[85] , \o[86] , \o[87] , \o[88] , \o[89] , \o[90] , \o[91] , \o[92] , \o[93] , \o[94] , \o[95] , \o[96] , \o[97] , \o[98] , \o[99] , \o[100] , \o[101] , \o[102] , \o[103] , \o[104] , \o[105] , \o[106] , \o[107] , \o[108] , \o[109] , \o[110] , \o[111] , \o[112] , \o[113] , \o[114] , \o[115] , \o[116] , \o[117] , \o[118] , \o[119] , \o[120] , \o[121] , \o[122] , \o[123] , \o[124] , \o[125] , \o[126] , \o[127] , \o[128] , \o[129] , \o[130] , \o[131] , \o[132] , \o[133] , \o[134] , \o[135] , \o[136] , \o[137] , \o[138] , \o[139] , \o[140] , \o[141] , \o[142] , \o[143] , \o[144] , \o[145] , \o[146] , \o[147] , \o[148] , \o[149] , \o[150] , \o[151] , \o[152] , \o[153] , \o[154] , \o[155] , \o[156] , \o[157] , \o[158] , \o[159] , \o[160] , \o[161] , \o[162] , \o[163] , \o[164] , \o[165] , \o[166] , \o[167] , \o[168] , \o[169] , \o[170] , \o[171] , \o[172] , \o[173] , \o[174] , \o[175] , \o[176] , \o[177] , \o[178] , \o[179] , \o[180] , \o[181] , \o[182] , \o[183] , \o[184] , \o[185] , \o[186] , \o[187] , \o[188] , \o[189] , \o[190] , \o[191] , \o[192] , \o[193] , \o[194] , \o[195] , \o[196] , \o[197] , \o[198] , \o[199] , \o[200] , \o[201] , \o[202] , \o[203] , \o[204] , \o[205] , \o[206] , \o[207] , \o[208] , \o[209] , \o[210] , \o[211] , \o[212] , \o[213] , \o[214] , \o[215] , \o[216] , \o[217] , \o[218] , \o[219] , \o[220] , \o[221] , \o[222] , \o[223] , \o[224] , \o[225] , \o[226] , \o[227] , \o[228] , \o[229] , \o[230] , \o[231] , \o[232] , \o[233] , \o[234] , \o[235] , \o[236] , \o[237] , \o[238] , \o[239] , \o[240] , \o[241] , done);

wire _abc_65734_new_n1001_; 
wire _abc_65734_new_n1002_; 
wire _abc_65734_new_n1004_; 
wire _abc_65734_new_n1005_; 
wire _abc_65734_new_n1007_; 
wire _abc_65734_new_n1008_; 
wire _abc_65734_new_n1010_; 
wire _abc_65734_new_n1011_; 
wire _abc_65734_new_n1013_; 
wire _abc_65734_new_n1014_; 
wire _abc_65734_new_n1016_; 
wire _abc_65734_new_n1017_; 
wire _abc_65734_new_n1019_; 
wire _abc_65734_new_n1020_; 
wire _abc_65734_new_n1022_; 
wire _abc_65734_new_n1023_; 
wire _abc_65734_new_n1025_; 
wire _abc_65734_new_n1026_; 
wire _abc_65734_new_n1028_; 
wire _abc_65734_new_n1029_; 
wire _abc_65734_new_n1031_; 
wire _abc_65734_new_n1032_; 
wire _abc_65734_new_n1034_; 
wire _abc_65734_new_n1035_; 
wire _abc_65734_new_n1037_; 
wire _abc_65734_new_n1038_; 
wire _abc_65734_new_n1040_; 
wire _abc_65734_new_n1041_; 
wire _abc_65734_new_n1043_; 
wire _abc_65734_new_n1044_; 
wire _abc_65734_new_n1046_; 
wire _abc_65734_new_n1047_; 
wire _abc_65734_new_n1049_; 
wire _abc_65734_new_n1050_; 
wire _abc_65734_new_n1052_; 
wire _abc_65734_new_n1053_; 
wire _abc_65734_new_n1055_; 
wire _abc_65734_new_n1056_; 
wire _abc_65734_new_n1058_; 
wire _abc_65734_new_n1059_; 
wire _abc_65734_new_n1061_; 
wire _abc_65734_new_n1062_; 
wire _abc_65734_new_n1064_; 
wire _abc_65734_new_n1065_; 
wire _abc_65734_new_n1067_; 
wire _abc_65734_new_n1068_; 
wire _abc_65734_new_n1070_; 
wire _abc_65734_new_n1071_; 
wire _abc_65734_new_n1073_; 
wire _abc_65734_new_n1074_; 
wire _abc_65734_new_n1076_; 
wire _abc_65734_new_n1077_; 
wire _abc_65734_new_n1079_; 
wire _abc_65734_new_n1080_; 
wire _abc_65734_new_n1082_; 
wire _abc_65734_new_n1083_; 
wire _abc_65734_new_n1085_; 
wire _abc_65734_new_n1086_; 
wire _abc_65734_new_n1088_; 
wire _abc_65734_new_n1089_; 
wire _abc_65734_new_n1091_; 
wire _abc_65734_new_n1092_; 
wire _abc_65734_new_n1094_; 
wire _abc_65734_new_n1095_; 
wire _abc_65734_new_n1097_; 
wire _abc_65734_new_n1098_; 
wire _abc_65734_new_n1100_; 
wire _abc_65734_new_n1101_; 
wire _abc_65734_new_n1103_; 
wire _abc_65734_new_n1104_; 
wire _abc_65734_new_n1106_; 
wire _abc_65734_new_n1107_; 
wire _abc_65734_new_n1109_; 
wire _abc_65734_new_n1110_; 
wire _abc_65734_new_n1112_; 
wire _abc_65734_new_n1113_; 
wire _abc_65734_new_n1115_; 
wire _abc_65734_new_n1116_; 
wire _abc_65734_new_n1118_; 
wire _abc_65734_new_n1119_; 
wire _abc_65734_new_n1121_; 
wire _abc_65734_new_n1122_; 
wire _abc_65734_new_n1124_; 
wire _abc_65734_new_n1125_; 
wire _abc_65734_new_n1127_; 
wire _abc_65734_new_n1128_; 
wire _abc_65734_new_n1130_; 
wire _abc_65734_new_n1131_; 
wire _abc_65734_new_n1133_; 
wire _abc_65734_new_n1134_; 
wire _abc_65734_new_n1136_; 
wire _abc_65734_new_n1137_; 
wire _abc_65734_new_n1139_; 
wire _abc_65734_new_n1140_; 
wire _abc_65734_new_n1142_; 
wire _abc_65734_new_n1143_; 
wire _abc_65734_new_n1145_; 
wire _abc_65734_new_n1146_; 
wire _abc_65734_new_n1148_; 
wire _abc_65734_new_n1149_; 
wire _abc_65734_new_n1151_; 
wire _abc_65734_new_n1152_; 
wire _abc_65734_new_n1154_; 
wire _abc_65734_new_n1155_; 
wire _abc_65734_new_n1157_; 
wire _abc_65734_new_n1158_; 
wire _abc_65734_new_n1160_; 
wire _abc_65734_new_n1161_; 
wire _abc_65734_new_n1163_; 
wire _abc_65734_new_n1164_; 
wire _abc_65734_new_n1168_; 
wire _abc_65734_new_n1169_; 
wire _abc_65734_new_n1171_; 
wire _abc_65734_new_n1173_; 
wire _abc_65734_new_n1174_; 
wire _abc_65734_new_n1176_; 
wire _abc_65734_new_n1178_; 
wire _abc_65734_new_n1179_; 
wire _abc_65734_new_n1181_; 
wire _abc_65734_new_n1183_; 
wire _abc_65734_new_n1184_; 
wire _abc_65734_new_n1186_; 
wire _abc_65734_new_n1188_; 
wire _abc_65734_new_n1189_; 
wire _abc_65734_new_n1191_; 
wire _abc_65734_new_n1193_; 
wire _abc_65734_new_n1194_; 
wire _abc_65734_new_n1196_; 
wire _abc_65734_new_n1198_; 
wire _abc_65734_new_n1199_; 
wire _abc_65734_new_n1201_; 
wire _abc_65734_new_n1203_; 
wire _abc_65734_new_n1204_; 
wire _abc_65734_new_n1206_; 
wire _abc_65734_new_n1208_; 
wire _abc_65734_new_n1209_; 
wire _abc_65734_new_n1211_; 
wire _abc_65734_new_n1213_; 
wire _abc_65734_new_n1214_; 
wire _abc_65734_new_n1216_; 
wire _abc_65734_new_n1218_; 
wire _abc_65734_new_n1219_; 
wire _abc_65734_new_n1221_; 
wire _abc_65734_new_n1223_; 
wire _abc_65734_new_n1224_; 
wire _abc_65734_new_n1226_; 
wire _abc_65734_new_n1228_; 
wire _abc_65734_new_n1229_; 
wire _abc_65734_new_n1231_; 
wire _abc_65734_new_n1233_; 
wire _abc_65734_new_n1234_; 
wire _abc_65734_new_n1236_; 
wire _abc_65734_new_n1238_; 
wire _abc_65734_new_n1239_; 
wire _abc_65734_new_n1241_; 
wire _abc_65734_new_n1243_; 
wire _abc_65734_new_n1244_; 
wire _abc_65734_new_n1246_; 
wire _abc_65734_new_n1248_; 
wire _abc_65734_new_n1249_; 
wire _abc_65734_new_n1251_; 
wire _abc_65734_new_n1253_; 
wire _abc_65734_new_n1254_; 
wire _abc_65734_new_n1256_; 
wire _abc_65734_new_n1258_; 
wire _abc_65734_new_n1259_; 
wire _abc_65734_new_n1261_; 
wire _abc_65734_new_n1263_; 
wire _abc_65734_new_n1264_; 
wire _abc_65734_new_n1266_; 
wire _abc_65734_new_n1268_; 
wire _abc_65734_new_n1269_; 
wire _abc_65734_new_n1271_; 
wire _abc_65734_new_n1273_; 
wire _abc_65734_new_n1274_; 
wire _abc_65734_new_n1276_; 
wire _abc_65734_new_n1278_; 
wire _abc_65734_new_n1279_; 
wire _abc_65734_new_n1281_; 
wire _abc_65734_new_n1283_; 
wire _abc_65734_new_n1284_; 
wire _abc_65734_new_n1286_; 
wire _abc_65734_new_n1288_; 
wire _abc_65734_new_n1289_; 
wire _abc_65734_new_n1291_; 
wire _abc_65734_new_n1293_; 
wire _abc_65734_new_n1294_; 
wire _abc_65734_new_n1296_; 
wire _abc_65734_new_n1298_; 
wire _abc_65734_new_n1299_; 
wire _abc_65734_new_n1301_; 
wire _abc_65734_new_n1303_; 
wire _abc_65734_new_n1304_; 
wire _abc_65734_new_n1306_; 
wire _abc_65734_new_n1308_; 
wire _abc_65734_new_n1309_; 
wire _abc_65734_new_n1311_; 
wire _abc_65734_new_n1313_; 
wire _abc_65734_new_n1314_; 
wire _abc_65734_new_n1316_; 
wire _abc_65734_new_n1318_; 
wire _abc_65734_new_n1319_; 
wire _abc_65734_new_n1321_; 
wire _abc_65734_new_n1323_; 
wire _abc_65734_new_n1324_; 
wire _abc_65734_new_n1326_; 
wire _abc_65734_new_n1328_; 
wire _abc_65734_new_n1329_; 
wire _abc_65734_new_n1331_; 
wire _abc_65734_new_n1333_; 
wire _abc_65734_new_n1334_; 
wire _abc_65734_new_n1336_; 
wire _abc_65734_new_n1338_; 
wire _abc_65734_new_n1339_; 
wire _abc_65734_new_n1341_; 
wire _abc_65734_new_n1343_; 
wire _abc_65734_new_n1344_; 
wire _abc_65734_new_n1346_; 
wire _abc_65734_new_n1348_; 
wire _abc_65734_new_n1349_; 
wire _abc_65734_new_n1351_; 
wire _abc_65734_new_n1353_; 
wire _abc_65734_new_n1354_; 
wire _abc_65734_new_n1356_; 
wire _abc_65734_new_n1358_; 
wire _abc_65734_new_n1359_; 
wire _abc_65734_new_n1361_; 
wire _abc_65734_new_n1363_; 
wire _abc_65734_new_n1364_; 
wire _abc_65734_new_n1366_; 
wire _abc_65734_new_n1368_; 
wire _abc_65734_new_n1369_; 
wire _abc_65734_new_n1371_; 
wire _abc_65734_new_n1373_; 
wire _abc_65734_new_n1374_; 
wire _abc_65734_new_n1376_; 
wire _abc_65734_new_n1378_; 
wire _abc_65734_new_n1379_; 
wire _abc_65734_new_n1381_; 
wire _abc_65734_new_n1383_; 
wire _abc_65734_new_n1384_; 
wire _abc_65734_new_n1386_; 
wire _abc_65734_new_n1388_; 
wire _abc_65734_new_n1389_; 
wire _abc_65734_new_n1391_; 
wire _abc_65734_new_n1393_; 
wire _abc_65734_new_n1394_; 
wire _abc_65734_new_n1396_; 
wire _abc_65734_new_n1398_; 
wire _abc_65734_new_n1399_; 
wire _abc_65734_new_n1401_; 
wire _abc_65734_new_n1403_; 
wire _abc_65734_new_n1404_; 
wire _abc_65734_new_n1406_; 
wire _abc_65734_new_n1408_; 
wire _abc_65734_new_n1409_; 
wire _abc_65734_new_n1411_; 
wire _abc_65734_new_n1413_; 
wire _abc_65734_new_n1414_; 
wire _abc_65734_new_n1416_; 
wire _abc_65734_new_n1418_; 
wire _abc_65734_new_n1419_; 
wire _abc_65734_new_n1421_; 
wire _abc_65734_new_n1423_; 
wire _abc_65734_new_n1424_; 
wire _abc_65734_new_n1426_; 
wire _abc_65734_new_n1428_; 
wire _abc_65734_new_n1429_; 
wire _abc_65734_new_n1431_; 
wire _abc_65734_new_n1433_; 
wire _abc_65734_new_n1434_; 
wire _abc_65734_new_n1436_; 
wire _abc_65734_new_n1438_; 
wire _abc_65734_new_n1439_; 
wire _abc_65734_new_n1441_; 
wire _abc_65734_new_n1443_; 
wire _abc_65734_new_n1444_; 
wire _abc_65734_new_n1446_; 
wire _abc_65734_new_n1448_; 
wire _abc_65734_new_n1449_; 
wire _abc_65734_new_n1452_; 
wire _abc_65734_new_n1453_; 
wire _abc_65734_new_n1454_; 
wire _abc_65734_new_n1456_; 
wire _abc_65734_new_n1457_; 
wire _abc_65734_new_n1458_; 
wire _abc_65734_new_n1459_; 
wire _abc_65734_new_n1461_; 
wire _abc_65734_new_n1462_; 
wire _abc_65734_new_n1463_; 
wire _abc_65734_new_n1464_; 
wire _abc_65734_new_n1465_; 
wire _abc_65734_new_n1466_; 
wire _abc_65734_new_n1467_; 
wire _abc_65734_new_n1468_; 
wire _abc_65734_new_n1470_; 
wire _abc_65734_new_n1471_; 
wire _abc_65734_new_n1472_; 
wire _abc_65734_new_n1473_; 
wire _abc_65734_new_n1474_; 
wire _abc_65734_new_n1475_; 
wire _abc_65734_new_n1476_; 
wire _abc_65734_new_n1477_; 
wire _abc_65734_new_n1479_; 
wire _abc_65734_new_n1480_; 
wire _abc_65734_new_n1481_; 
wire _abc_65734_new_n1482_; 
wire _abc_65734_new_n1483_; 
wire _abc_65734_new_n1484_; 
wire _abc_65734_new_n1485_; 
wire _abc_65734_new_n1486_; 
wire _abc_65734_new_n1487_; 
wire _abc_65734_new_n1488_; 
wire _abc_65734_new_n1489_; 
wire _abc_65734_new_n1490_; 
wire _abc_65734_new_n1492_; 
wire _abc_65734_new_n1493_; 
wire _abc_65734_new_n1494_; 
wire _abc_65734_new_n1495_; 
wire _abc_65734_new_n1496_; 
wire _abc_65734_new_n1497_; 
wire _abc_65734_new_n1498_; 
wire _abc_65734_new_n1500_; 
wire _abc_65734_new_n1501_; 
wire _abc_65734_new_n1502_; 
wire _abc_65734_new_n1503_; 
wire _abc_65734_new_n1504_; 
wire _abc_65734_new_n1505_; 
wire _abc_65734_new_n1506_; 
wire _abc_65734_new_n1507_; 
wire _abc_65734_new_n1508_; 
wire _abc_65734_new_n1510_; 
wire _abc_65734_new_n1511_; 
wire _abc_65734_new_n1512_; 
wire _abc_65734_new_n1513_; 
wire _abc_65734_new_n1514_; 
wire _abc_65734_new_n1515_; 
wire _abc_65734_new_n1516_; 
wire _abc_65734_new_n1517_; 
wire _abc_65734_new_n1518_; 
wire _abc_65734_new_n1519_; 
wire _abc_65734_new_n1520_; 
wire _abc_65734_new_n1522_; 
wire _abc_65734_new_n1523_; 
wire _abc_65734_new_n1524_; 
wire _abc_65734_new_n1525_; 
wire _abc_65734_new_n1526_; 
wire _abc_65734_new_n1527_; 
wire _abc_65734_new_n1528_; 
wire _abc_65734_new_n1529_; 
wire _abc_65734_new_n1530_; 
wire _abc_65734_new_n1531_; 
wire _abc_65734_new_n1533_; 
wire _abc_65734_new_n1534_; 
wire _abc_65734_new_n1535_; 
wire _abc_65734_new_n1536_; 
wire _abc_65734_new_n1537_; 
wire _abc_65734_new_n1538_; 
wire _abc_65734_new_n1539_; 
wire _abc_65734_new_n1540_; 
wire _abc_65734_new_n1541_; 
wire _abc_65734_new_n1542_; 
wire _abc_65734_new_n1544_; 
wire _abc_65734_new_n1545_; 
wire _abc_65734_new_n1546_; 
wire _abc_65734_new_n1547_; 
wire _abc_65734_new_n1548_; 
wire _abc_65734_new_n1549_; 
wire _abc_65734_new_n1550_; 
wire _abc_65734_new_n1551_; 
wire _abc_65734_new_n1552_; 
wire _abc_65734_new_n1554_; 
wire _abc_65734_new_n1555_; 
wire _abc_65734_new_n1556_; 
wire _abc_65734_new_n1557_; 
wire _abc_65734_new_n1558_; 
wire _abc_65734_new_n1559_; 
wire _abc_65734_new_n1560_; 
wire _abc_65734_new_n1561_; 
wire _abc_65734_new_n1563_; 
wire _abc_65734_new_n1564_; 
wire _abc_65734_new_n1565_; 
wire _abc_65734_new_n1566_; 
wire _abc_65734_new_n1567_; 
wire _abc_65734_new_n1568_; 
wire _abc_65734_new_n1569_; 
wire _abc_65734_new_n1571_; 
wire _abc_65734_new_n1572_; 
wire _abc_65734_new_n1573_; 
wire _abc_65734_new_n1574_; 
wire _abc_65734_new_n1575_; 
wire _abc_65734_new_n1576_; 
wire _abc_65734_new_n1577_; 
wire _abc_65734_new_n1578_; 
wire _abc_65734_new_n1580_; 
wire _abc_65734_new_n1581_; 
wire _abc_65734_new_n1582_; 
wire _abc_65734_new_n1583_; 
wire _abc_65734_new_n1584_; 
wire _abc_65734_new_n753_; 
wire _abc_65734_new_n830_; 
wire _abc_65734_new_n831_; 
wire _abc_65734_new_n833_; 
wire _abc_65734_new_n834_; 
wire _abc_65734_new_n836_; 
wire _abc_65734_new_n837_; 
wire _abc_65734_new_n839_; 
wire _abc_65734_new_n840_; 
wire _abc_65734_new_n842_; 
wire _abc_65734_new_n843_; 
wire _abc_65734_new_n845_; 
wire _abc_65734_new_n846_; 
wire _abc_65734_new_n848_; 
wire _abc_65734_new_n849_; 
wire _abc_65734_new_n851_; 
wire _abc_65734_new_n852_; 
wire _abc_65734_new_n854_; 
wire _abc_65734_new_n855_; 
wire _abc_65734_new_n857_; 
wire _abc_65734_new_n858_; 
wire _abc_65734_new_n860_; 
wire _abc_65734_new_n861_; 
wire _abc_65734_new_n863_; 
wire _abc_65734_new_n864_; 
wire _abc_65734_new_n866_; 
wire _abc_65734_new_n867_; 
wire _abc_65734_new_n869_; 
wire _abc_65734_new_n870_; 
wire _abc_65734_new_n872_; 
wire _abc_65734_new_n873_; 
wire _abc_65734_new_n875_; 
wire _abc_65734_new_n876_; 
wire _abc_65734_new_n878_; 
wire _abc_65734_new_n879_; 
wire _abc_65734_new_n881_; 
wire _abc_65734_new_n882_; 
wire _abc_65734_new_n884_; 
wire _abc_65734_new_n885_; 
wire _abc_65734_new_n887_; 
wire _abc_65734_new_n888_; 
wire _abc_65734_new_n890_; 
wire _abc_65734_new_n891_; 
wire _abc_65734_new_n893_; 
wire _abc_65734_new_n894_; 
wire _abc_65734_new_n896_; 
wire _abc_65734_new_n897_; 
wire _abc_65734_new_n899_; 
wire _abc_65734_new_n900_; 
wire _abc_65734_new_n902_; 
wire _abc_65734_new_n903_; 
wire _abc_65734_new_n905_; 
wire _abc_65734_new_n906_; 
wire _abc_65734_new_n908_; 
wire _abc_65734_new_n909_; 
wire _abc_65734_new_n911_; 
wire _abc_65734_new_n912_; 
wire _abc_65734_new_n914_; 
wire _abc_65734_new_n915_; 
wire _abc_65734_new_n917_; 
wire _abc_65734_new_n918_; 
wire _abc_65734_new_n920_; 
wire _abc_65734_new_n921_; 
wire _abc_65734_new_n923_; 
wire _abc_65734_new_n924_; 
wire _abc_65734_new_n926_; 
wire _abc_65734_new_n927_; 
wire _abc_65734_new_n929_; 
wire _abc_65734_new_n930_; 
wire _abc_65734_new_n932_; 
wire _abc_65734_new_n933_; 
wire _abc_65734_new_n935_; 
wire _abc_65734_new_n936_; 
wire _abc_65734_new_n938_; 
wire _abc_65734_new_n939_; 
wire _abc_65734_new_n941_; 
wire _abc_65734_new_n942_; 
wire _abc_65734_new_n944_; 
wire _abc_65734_new_n945_; 
wire _abc_65734_new_n947_; 
wire _abc_65734_new_n948_; 
wire _abc_65734_new_n950_; 
wire _abc_65734_new_n951_; 
wire _abc_65734_new_n953_; 
wire _abc_65734_new_n954_; 
wire _abc_65734_new_n956_; 
wire _abc_65734_new_n957_; 
wire _abc_65734_new_n959_; 
wire _abc_65734_new_n960_; 
wire _abc_65734_new_n962_; 
wire _abc_65734_new_n963_; 
wire _abc_65734_new_n965_; 
wire _abc_65734_new_n966_; 
wire _abc_65734_new_n968_; 
wire _abc_65734_new_n969_; 
wire _abc_65734_new_n971_; 
wire _abc_65734_new_n972_; 
wire _abc_65734_new_n974_; 
wire _abc_65734_new_n975_; 
wire _abc_65734_new_n977_; 
wire _abc_65734_new_n978_; 
wire _abc_65734_new_n980_; 
wire _abc_65734_new_n981_; 
wire _abc_65734_new_n983_; 
wire _abc_65734_new_n984_; 
wire _abc_65734_new_n986_; 
wire _abc_65734_new_n987_; 
wire _abc_65734_new_n989_; 
wire _abc_65734_new_n990_; 
wire _abc_65734_new_n992_; 
wire _abc_65734_new_n993_; 
wire _abc_65734_new_n995_; 
wire _abc_65734_new_n996_; 
wire _abc_65734_new_n998_; 
wire _abc_65734_new_n999_; 
wire aNan; 
input \a[0] ;
input \a[100] ;
input \a[101] ;
input \a[102] ;
input \a[103] ;
input \a[104] ;
input \a[105] ;
input \a[106] ;
input \a[107] ;
input \a[108] ;
input \a[109] ;
input \a[10] ;
input \a[110] ;
input \a[111] ;
input \a[112] ;
input \a[113] ;
input \a[114] ;
input \a[115] ;
input \a[116] ;
input \a[117] ;
input \a[118] ;
input \a[119] ;
input \a[11] ;
input \a[120] ;
input \a[121] ;
input \a[122] ;
input \a[123] ;
input \a[124] ;
input \a[125] ;
input \a[126] ;
input \a[127] ;
input \a[12] ;
input \a[13] ;
input \a[14] ;
input \a[15] ;
input \a[16] ;
input \a[17] ;
input \a[18] ;
input \a[19] ;
input \a[1] ;
input \a[20] ;
input \a[21] ;
input \a[22] ;
input \a[23] ;
input \a[24] ;
input \a[25] ;
input \a[26] ;
input \a[27] ;
input \a[28] ;
input \a[29] ;
input \a[2] ;
input \a[30] ;
input \a[31] ;
input \a[32] ;
input \a[33] ;
input \a[34] ;
input \a[35] ;
input \a[36] ;
input \a[37] ;
input \a[38] ;
input \a[39] ;
input \a[3] ;
input \a[40] ;
input \a[41] ;
input \a[42] ;
input \a[43] ;
input \a[44] ;
input \a[45] ;
input \a[46] ;
input \a[47] ;
input \a[48] ;
input \a[49] ;
input \a[4] ;
input \a[50] ;
input \a[51] ;
input \a[52] ;
input \a[53] ;
input \a[54] ;
input \a[55] ;
input \a[56] ;
input \a[57] ;
input \a[58] ;
input \a[59] ;
input \a[5] ;
input \a[60] ;
input \a[61] ;
input \a[62] ;
input \a[63] ;
input \a[64] ;
input \a[65] ;
input \a[66] ;
input \a[67] ;
input \a[68] ;
input \a[69] ;
input \a[6] ;
input \a[70] ;
input \a[71] ;
input \a[72] ;
input \a[73] ;
input \a[74] ;
input \a[75] ;
input \a[76] ;
input \a[77] ;
input \a[78] ;
input \a[79] ;
input \a[7] ;
input \a[80] ;
input \a[81] ;
input \a[82] ;
input \a[83] ;
input \a[84] ;
input \a[85] ;
input \a[86] ;
input \a[87] ;
input \a[88] ;
input \a[89] ;
input \a[8] ;
input \a[90] ;
input \a[91] ;
input \a[92] ;
input \a[93] ;
input \a[94] ;
input \a[95] ;
input \a[96] ;
input \a[97] ;
input \a[98] ;
input \a[99] ;
input \a[9] ;
input ce;
input clk;
output done;
wire fracta1_0_; 
wire fracta1_100_; 
wire fracta1_101_; 
wire fracta1_102_; 
wire fracta1_103_; 
wire fracta1_104_; 
wire fracta1_105_; 
wire fracta1_106_; 
wire fracta1_107_; 
wire fracta1_108_; 
wire fracta1_109_; 
wire fracta1_10_; 
wire fracta1_110_; 
wire fracta1_111_; 
wire fracta1_112_; 
wire fracta1_113_; 
wire fracta1_11_; 
wire fracta1_12_; 
wire fracta1_13_; 
wire fracta1_14_; 
wire fracta1_15_; 
wire fracta1_16_; 
wire fracta1_17_; 
wire fracta1_18_; 
wire fracta1_19_; 
wire fracta1_1_; 
wire fracta1_20_; 
wire fracta1_21_; 
wire fracta1_22_; 
wire fracta1_23_; 
wire fracta1_24_; 
wire fracta1_25_; 
wire fracta1_26_; 
wire fracta1_27_; 
wire fracta1_28_; 
wire fracta1_29_; 
wire fracta1_2_; 
wire fracta1_30_; 
wire fracta1_31_; 
wire fracta1_32_; 
wire fracta1_33_; 
wire fracta1_34_; 
wire fracta1_35_; 
wire fracta1_36_; 
wire fracta1_37_; 
wire fracta1_38_; 
wire fracta1_39_; 
wire fracta1_3_; 
wire fracta1_40_; 
wire fracta1_41_; 
wire fracta1_42_; 
wire fracta1_43_; 
wire fracta1_44_; 
wire fracta1_45_; 
wire fracta1_46_; 
wire fracta1_47_; 
wire fracta1_48_; 
wire fracta1_49_; 
wire fracta1_4_; 
wire fracta1_50_; 
wire fracta1_51_; 
wire fracta1_52_; 
wire fracta1_53_; 
wire fracta1_54_; 
wire fracta1_55_; 
wire fracta1_56_; 
wire fracta1_57_; 
wire fracta1_58_; 
wire fracta1_59_; 
wire fracta1_5_; 
wire fracta1_60_; 
wire fracta1_61_; 
wire fracta1_62_; 
wire fracta1_63_; 
wire fracta1_64_; 
wire fracta1_65_; 
wire fracta1_66_; 
wire fracta1_67_; 
wire fracta1_68_; 
wire fracta1_69_; 
wire fracta1_6_; 
wire fracta1_70_; 
wire fracta1_71_; 
wire fracta1_72_; 
wire fracta1_73_; 
wire fracta1_74_; 
wire fracta1_75_; 
wire fracta1_76_; 
wire fracta1_77_; 
wire fracta1_78_; 
wire fracta1_79_; 
wire fracta1_7_; 
wire fracta1_80_; 
wire fracta1_81_; 
wire fracta1_82_; 
wire fracta1_83_; 
wire fracta1_84_; 
wire fracta1_85_; 
wire fracta1_86_; 
wire fracta1_87_; 
wire fracta1_88_; 
wire fracta1_89_; 
wire fracta1_8_; 
wire fracta1_90_; 
wire fracta1_91_; 
wire fracta1_92_; 
wire fracta1_93_; 
wire fracta1_94_; 
wire fracta1_95_; 
wire fracta1_96_; 
wire fracta1_97_; 
wire fracta1_98_; 
wire fracta1_99_; 
wire fracta1_9_; 
wire fracta_112_; 
input ld;
output \o[0] ;
output \o[100] ;
output \o[101] ;
output \o[102] ;
output \o[103] ;
output \o[104] ;
output \o[105] ;
output \o[106] ;
output \o[107] ;
output \o[108] ;
output \o[109] ;
output \o[10] ;
output \o[110] ;
output \o[111] ;
output \o[112] ;
output \o[113] ;
output \o[114] ;
output \o[115] ;
output \o[116] ;
output \o[117] ;
output \o[118] ;
output \o[119] ;
output \o[11] ;
output \o[120] ;
output \o[121] ;
output \o[122] ;
output \o[123] ;
output \o[124] ;
output \o[125] ;
output \o[126] ;
output \o[127] ;
output \o[128] ;
output \o[129] ;
output \o[12] ;
output \o[130] ;
output \o[131] ;
output \o[132] ;
output \o[133] ;
output \o[134] ;
output \o[135] ;
output \o[136] ;
output \o[137] ;
output \o[138] ;
output \o[139] ;
output \o[13] ;
output \o[140] ;
output \o[141] ;
output \o[142] ;
output \o[143] ;
output \o[144] ;
output \o[145] ;
output \o[146] ;
output \o[147] ;
output \o[148] ;
output \o[149] ;
output \o[14] ;
output \o[150] ;
output \o[151] ;
output \o[152] ;
output \o[153] ;
output \o[154] ;
output \o[155] ;
output \o[156] ;
output \o[157] ;
output \o[158] ;
output \o[159] ;
output \o[15] ;
output \o[160] ;
output \o[161] ;
output \o[162] ;
output \o[163] ;
output \o[164] ;
output \o[165] ;
output \o[166] ;
output \o[167] ;
output \o[168] ;
output \o[169] ;
output \o[16] ;
output \o[170] ;
output \o[171] ;
output \o[172] ;
output \o[173] ;
output \o[174] ;
output \o[175] ;
output \o[176] ;
output \o[177] ;
output \o[178] ;
output \o[179] ;
output \o[17] ;
output \o[180] ;
output \o[181] ;
output \o[182] ;
output \o[183] ;
output \o[184] ;
output \o[185] ;
output \o[186] ;
output \o[187] ;
output \o[188] ;
output \o[189] ;
output \o[18] ;
output \o[190] ;
output \o[191] ;
output \o[192] ;
output \o[193] ;
output \o[194] ;
output \o[195] ;
output \o[196] ;
output \o[197] ;
output \o[198] ;
output \o[199] ;
output \o[19] ;
output \o[1] ;
output \o[200] ;
output \o[201] ;
output \o[202] ;
output \o[203] ;
output \o[204] ;
output \o[205] ;
output \o[206] ;
output \o[207] ;
output \o[208] ;
output \o[209] ;
output \o[20] ;
output \o[210] ;
output \o[211] ;
output \o[212] ;
output \o[213] ;
output \o[214] ;
output \o[215] ;
output \o[216] ;
output \o[217] ;
output \o[218] ;
output \o[219] ;
output \o[21] ;
output \o[220] ;
output \o[221] ;
output \o[222] ;
output \o[223] ;
output \o[224] ;
output \o[225] ;
output \o[226] ;
output \o[227] ;
output \o[228] ;
output \o[229] ;
output \o[22] ;
output \o[230] ;
output \o[231] ;
output \o[232] ;
output \o[233] ;
output \o[234] ;
output \o[235] ;
output \o[236] ;
output \o[237] ;
output \o[238] ;
output \o[239] ;
output \o[23] ;
output \o[240] ;
output \o[241] ;
output \o[24] ;
output \o[25] ;
output \o[26] ;
output \o[27] ;
output \o[28] ;
output \o[29] ;
output \o[2] ;
output \o[30] ;
output \o[31] ;
output \o[32] ;
output \o[33] ;
output \o[34] ;
output \o[35] ;
output \o[36] ;
output \o[37] ;
output \o[38] ;
output \o[39] ;
output \o[3] ;
output \o[40] ;
output \o[41] ;
output \o[42] ;
output \o[43] ;
output \o[44] ;
output \o[45] ;
output \o[46] ;
output \o[47] ;
output \o[48] ;
output \o[49] ;
output \o[4] ;
output \o[50] ;
output \o[51] ;
output \o[52] ;
output \o[53] ;
output \o[54] ;
output \o[55] ;
output \o[56] ;
output \o[57] ;
output \o[58] ;
output \o[59] ;
output \o[5] ;
output \o[60] ;
output \o[61] ;
output \o[62] ;
output \o[63] ;
output \o[64] ;
output \o[65] ;
output \o[66] ;
output \o[67] ;
output \o[68] ;
output \o[69] ;
output \o[6] ;
output \o[70] ;
output \o[71] ;
output \o[72] ;
output \o[73] ;
output \o[74] ;
output \o[75] ;
output \o[76] ;
output \o[77] ;
output \o[78] ;
output \o[79] ;
output \o[7] ;
output \o[80] ;
output \o[81] ;
output \o[82] ;
output \o[83] ;
output \o[84] ;
output \o[85] ;
output \o[86] ;
output \o[87] ;
output \o[88] ;
output \o[89] ;
output \o[8] ;
output \o[90] ;
output \o[91] ;
output \o[92] ;
output \o[93] ;
output \o[94] ;
output \o[95] ;
output \o[96] ;
output \o[97] ;
output \o[98] ;
output \o[99] ;
output \o[9] ;
input rst;
wire sqrto_0_; 
wire sqrto_100_; 
wire sqrto_101_; 
wire sqrto_102_; 
wire sqrto_103_; 
wire sqrto_104_; 
wire sqrto_105_; 
wire sqrto_106_; 
wire sqrto_107_; 
wire sqrto_108_; 
wire sqrto_109_; 
wire sqrto_10_; 
wire sqrto_110_; 
wire sqrto_111_; 
wire sqrto_112_; 
wire sqrto_113_; 
wire sqrto_114_; 
wire sqrto_115_; 
wire sqrto_116_; 
wire sqrto_117_; 
wire sqrto_118_; 
wire sqrto_119_; 
wire sqrto_11_; 
wire sqrto_120_; 
wire sqrto_121_; 
wire sqrto_122_; 
wire sqrto_123_; 
wire sqrto_124_; 
wire sqrto_125_; 
wire sqrto_126_; 
wire sqrto_127_; 
wire sqrto_128_; 
wire sqrto_129_; 
wire sqrto_12_; 
wire sqrto_130_; 
wire sqrto_131_; 
wire sqrto_132_; 
wire sqrto_133_; 
wire sqrto_134_; 
wire sqrto_135_; 
wire sqrto_136_; 
wire sqrto_137_; 
wire sqrto_138_; 
wire sqrto_139_; 
wire sqrto_13_; 
wire sqrto_140_; 
wire sqrto_141_; 
wire sqrto_142_; 
wire sqrto_143_; 
wire sqrto_144_; 
wire sqrto_145_; 
wire sqrto_146_; 
wire sqrto_147_; 
wire sqrto_148_; 
wire sqrto_149_; 
wire sqrto_14_; 
wire sqrto_150_; 
wire sqrto_151_; 
wire sqrto_152_; 
wire sqrto_153_; 
wire sqrto_154_; 
wire sqrto_155_; 
wire sqrto_156_; 
wire sqrto_157_; 
wire sqrto_158_; 
wire sqrto_159_; 
wire sqrto_15_; 
wire sqrto_160_; 
wire sqrto_161_; 
wire sqrto_162_; 
wire sqrto_163_; 
wire sqrto_164_; 
wire sqrto_165_; 
wire sqrto_166_; 
wire sqrto_167_; 
wire sqrto_168_; 
wire sqrto_169_; 
wire sqrto_16_; 
wire sqrto_170_; 
wire sqrto_171_; 
wire sqrto_172_; 
wire sqrto_173_; 
wire sqrto_174_; 
wire sqrto_175_; 
wire sqrto_176_; 
wire sqrto_177_; 
wire sqrto_178_; 
wire sqrto_179_; 
wire sqrto_17_; 
wire sqrto_180_; 
wire sqrto_181_; 
wire sqrto_182_; 
wire sqrto_183_; 
wire sqrto_184_; 
wire sqrto_185_; 
wire sqrto_186_; 
wire sqrto_187_; 
wire sqrto_188_; 
wire sqrto_189_; 
wire sqrto_18_; 
wire sqrto_190_; 
wire sqrto_191_; 
wire sqrto_192_; 
wire sqrto_193_; 
wire sqrto_194_; 
wire sqrto_195_; 
wire sqrto_196_; 
wire sqrto_197_; 
wire sqrto_198_; 
wire sqrto_199_; 
wire sqrto_19_; 
wire sqrto_1_; 
wire sqrto_200_; 
wire sqrto_201_; 
wire sqrto_202_; 
wire sqrto_203_; 
wire sqrto_204_; 
wire sqrto_205_; 
wire sqrto_206_; 
wire sqrto_207_; 
wire sqrto_208_; 
wire sqrto_209_; 
wire sqrto_20_; 
wire sqrto_210_; 
wire sqrto_211_; 
wire sqrto_212_; 
wire sqrto_213_; 
wire sqrto_214_; 
wire sqrto_215_; 
wire sqrto_216_; 
wire sqrto_217_; 
wire sqrto_218_; 
wire sqrto_219_; 
wire sqrto_21_; 
wire sqrto_220_; 
wire sqrto_221_; 
wire sqrto_222_; 
wire sqrto_223_; 
wire sqrto_224_; 
wire sqrto_225_; 
wire sqrto_22_; 
wire sqrto_23_; 
wire sqrto_24_; 
wire sqrto_25_; 
wire sqrto_26_; 
wire sqrto_27_; 
wire sqrto_28_; 
wire sqrto_29_; 
wire sqrto_2_; 
wire sqrto_30_; 
wire sqrto_31_; 
wire sqrto_32_; 
wire sqrto_33_; 
wire sqrto_34_; 
wire sqrto_35_; 
wire sqrto_36_; 
wire sqrto_37_; 
wire sqrto_38_; 
wire sqrto_39_; 
wire sqrto_3_; 
wire sqrto_40_; 
wire sqrto_41_; 
wire sqrto_42_; 
wire sqrto_43_; 
wire sqrto_44_; 
wire sqrto_45_; 
wire sqrto_46_; 
wire sqrto_47_; 
wire sqrto_48_; 
wire sqrto_49_; 
wire sqrto_4_; 
wire sqrto_50_; 
wire sqrto_51_; 
wire sqrto_52_; 
wire sqrto_53_; 
wire sqrto_54_; 
wire sqrto_55_; 
wire sqrto_56_; 
wire sqrto_57_; 
wire sqrto_58_; 
wire sqrto_59_; 
wire sqrto_5_; 
wire sqrto_60_; 
wire sqrto_61_; 
wire sqrto_62_; 
wire sqrto_63_; 
wire sqrto_64_; 
wire sqrto_65_; 
wire sqrto_66_; 
wire sqrto_67_; 
wire sqrto_68_; 
wire sqrto_69_; 
wire sqrto_6_; 
wire sqrto_70_; 
wire sqrto_71_; 
wire sqrto_72_; 
wire sqrto_73_; 
wire sqrto_74_; 
wire sqrto_75_; 
wire sqrto_76_; 
wire sqrto_77_; 
wire sqrto_78_; 
wire sqrto_79_; 
wire sqrto_7_; 
wire sqrto_80_; 
wire sqrto_81_; 
wire sqrto_82_; 
wire sqrto_83_; 
wire sqrto_84_; 
wire sqrto_85_; 
wire sqrto_86_; 
wire sqrto_87_; 
wire sqrto_88_; 
wire sqrto_89_; 
wire sqrto_8_; 
wire sqrto_90_; 
wire sqrto_91_; 
wire sqrto_92_; 
wire sqrto_93_; 
wire sqrto_94_; 
wire sqrto_95_; 
wire sqrto_96_; 
wire sqrto_97_; 
wire sqrto_98_; 
wire sqrto_99_; 
wire sqrto_9_; 
wire u1__abc_51895_new_n137_; 
wire u1__abc_51895_new_n138_; 
wire u1__abc_51895_new_n139_; 
wire u1__abc_51895_new_n140_; 
wire u1__abc_51895_new_n141_; 
wire u1__abc_51895_new_n142_; 
wire u1__abc_51895_new_n143_; 
wire u1__abc_51895_new_n144_; 
wire u1__abc_51895_new_n145_; 
wire u1__abc_51895_new_n146_; 
wire u1__abc_51895_new_n147_; 
wire u1__abc_51895_new_n148_; 
wire u1__abc_51895_new_n149_; 
wire u1__abc_51895_new_n150_; 
wire u1__abc_51895_new_n153_; 
wire u1__abc_51895_new_n154_; 
wire u1__abc_51895_new_n155_; 
wire u1__abc_51895_new_n156_; 
wire u1__abc_51895_new_n157_; 
wire u1__abc_51895_new_n158_; 
wire u1__abc_51895_new_n159_; 
wire u1__abc_51895_new_n160_; 
wire u1__abc_51895_new_n161_; 
wire u1__abc_51895_new_n162_; 
wire u1__abc_51895_new_n163_; 
wire u1__abc_51895_new_n164_; 
wire u1__abc_51895_new_n166_; 
wire u1__abc_51895_new_n167_; 
wire u1__abc_51895_new_n168_; 
wire u1__abc_51895_new_n169_; 
wire u1__abc_51895_new_n170_; 
wire u1__abc_51895_new_n171_; 
wire u1__abc_51895_new_n172_; 
wire u1__abc_51895_new_n173_; 
wire u1__abc_51895_new_n174_; 
wire u1__abc_51895_new_n175_; 
wire u1__abc_51895_new_n176_; 
wire u1__abc_51895_new_n177_; 
wire u1__abc_51895_new_n178_; 
wire u1__abc_51895_new_n179_; 
wire u1__abc_51895_new_n180_; 
wire u1__abc_51895_new_n278_; 
wire u1__abc_51895_new_n282_; 
wire u1__abc_51895_new_n283_; 
wire u1__abc_51895_new_n284_; 
wire u1__abc_51895_new_n285_; 
wire u1__abc_51895_new_n286_; 
wire u1__abc_51895_new_n287_; 
wire u1__abc_51895_new_n288_; 
wire u1__abc_51895_new_n289_; 
wire u1__abc_51895_new_n290_; 
wire u1__abc_51895_new_n291_; 
wire u1__abc_51895_new_n292_; 
wire u1__abc_51895_new_n293_; 
wire u1__abc_51895_new_n294_; 
wire u1__abc_51895_new_n295_; 
wire u1__abc_51895_new_n296_; 
wire u1__abc_51895_new_n297_; 
wire u1__abc_51895_new_n298_; 
wire u1__abc_51895_new_n299_; 
wire u1__abc_51895_new_n300_; 
wire u1__abc_51895_new_n301_; 
wire u1__abc_51895_new_n302_; 
wire u1__abc_51895_new_n303_; 
wire u1__abc_51895_new_n304_; 
wire u1__abc_51895_new_n305_; 
wire u1__abc_51895_new_n306_; 
wire u1__abc_51895_new_n307_; 
wire u1__abc_51895_new_n308_; 
wire u1__abc_51895_new_n309_; 
wire u1__abc_51895_new_n310_; 
wire u1__abc_51895_new_n311_; 
wire u1__abc_51895_new_n312_; 
wire u1__abc_51895_new_n313_; 
wire u1__abc_51895_new_n314_; 
wire u1__abc_51895_new_n315_; 
wire u1__abc_51895_new_n316_; 
wire u1__abc_51895_new_n317_; 
wire u1__abc_51895_new_n318_; 
wire u1__abc_51895_new_n319_; 
wire u1__abc_51895_new_n320_; 
wire u1__abc_51895_new_n321_; 
wire u1__abc_51895_new_n322_; 
wire u1__abc_51895_new_n323_; 
wire u1__abc_51895_new_n324_; 
wire u1__abc_51895_new_n325_; 
wire u1__abc_51895_new_n326_; 
wire u1__abc_51895_new_n327_; 
wire u1__abc_51895_new_n328_; 
wire u1__abc_51895_new_n329_; 
wire u1__abc_51895_new_n330_; 
wire u1__abc_51895_new_n331_; 
wire u1__abc_51895_new_n332_; 
wire u1__abc_51895_new_n333_; 
wire u1__abc_51895_new_n334_; 
wire u1__abc_51895_new_n335_; 
wire u1__abc_51895_new_n336_; 
wire u1__abc_51895_new_n337_; 
wire u1__abc_51895_new_n338_; 
wire u1__abc_51895_new_n339_; 
wire u1__abc_51895_new_n340_; 
wire u1__abc_51895_new_n341_; 
wire u1__abc_51895_new_n342_; 
wire u1__abc_51895_new_n343_; 
wire u1__abc_51895_new_n344_; 
wire u1__abc_51895_new_n345_; 
wire u1__abc_51895_new_n346_; 
wire u1__abc_51895_new_n347_; 
wire u1__abc_51895_new_n348_; 
wire u1__abc_51895_new_n349_; 
wire u1__abc_51895_new_n350_; 
wire u1__abc_51895_new_n351_; 
wire u1__abc_51895_new_n352_; 
wire u1__abc_51895_new_n353_; 
wire u1__abc_51895_new_n354_; 
wire u1__abc_51895_new_n355_; 
wire u1__abc_51895_new_n356_; 
wire u1__abc_51895_new_n357_; 
wire u1__abc_51895_new_n358_; 
wire u1__abc_51895_new_n359_; 
wire u1__abc_51895_new_n360_; 
wire u1__abc_51895_new_n361_; 
wire u1__abc_51895_new_n362_; 
wire u1__abc_51895_new_n363_; 
wire u1__abc_51895_new_n364_; 
wire u1__abc_51895_new_n365_; 
wire u1__abc_51895_new_n366_; 
wire u1__abc_51895_new_n367_; 
wire u1__abc_51895_new_n368_; 
wire u1__abc_51895_new_n369_; 
wire u1__abc_51895_new_n370_; 
wire u1__abc_51895_new_n371_; 
wire u1__abc_51895_new_n372_; 
wire u1__abc_51895_new_n373_; 
wire u1__abc_51895_new_n374_; 
wire u1__abc_51895_new_n375_; 
wire u1_xinf; 
wire u2__0cnt_7_0__0_; 
wire u2__0cnt_7_0__1_; 
wire u2__0cnt_7_0__2_; 
wire u2__0cnt_7_0__3_; 
wire u2__0cnt_7_0__4_; 
wire u2__0cnt_7_0__5_; 
wire u2__0cnt_7_0__6_; 
wire u2__0cnt_7_0__7_; 
wire u2__0remHi_451_0__0_; 
wire u2__0remHi_451_0__100_; 
wire u2__0remHi_451_0__101_; 
wire u2__0remHi_451_0__102_; 
wire u2__0remHi_451_0__103_; 
wire u2__0remHi_451_0__104_; 
wire u2__0remHi_451_0__105_; 
wire u2__0remHi_451_0__106_; 
wire u2__0remHi_451_0__107_; 
wire u2__0remHi_451_0__108_; 
wire u2__0remHi_451_0__109_; 
wire u2__0remHi_451_0__10_; 
wire u2__0remHi_451_0__110_; 
wire u2__0remHi_451_0__111_; 
wire u2__0remHi_451_0__112_; 
wire u2__0remHi_451_0__113_; 
wire u2__0remHi_451_0__114_; 
wire u2__0remHi_451_0__115_; 
wire u2__0remHi_451_0__116_; 
wire u2__0remHi_451_0__117_; 
wire u2__0remHi_451_0__118_; 
wire u2__0remHi_451_0__119_; 
wire u2__0remHi_451_0__11_; 
wire u2__0remHi_451_0__120_; 
wire u2__0remHi_451_0__121_; 
wire u2__0remHi_451_0__122_; 
wire u2__0remHi_451_0__123_; 
wire u2__0remHi_451_0__124_; 
wire u2__0remHi_451_0__125_; 
wire u2__0remHi_451_0__126_; 
wire u2__0remHi_451_0__127_; 
wire u2__0remHi_451_0__128_; 
wire u2__0remHi_451_0__129_; 
wire u2__0remHi_451_0__12_; 
wire u2__0remHi_451_0__130_; 
wire u2__0remHi_451_0__131_; 
wire u2__0remHi_451_0__132_; 
wire u2__0remHi_451_0__133_; 
wire u2__0remHi_451_0__134_; 
wire u2__0remHi_451_0__135_; 
wire u2__0remHi_451_0__136_; 
wire u2__0remHi_451_0__137_; 
wire u2__0remHi_451_0__138_; 
wire u2__0remHi_451_0__139_; 
wire u2__0remHi_451_0__13_; 
wire u2__0remHi_451_0__140_; 
wire u2__0remHi_451_0__141_; 
wire u2__0remHi_451_0__142_; 
wire u2__0remHi_451_0__143_; 
wire u2__0remHi_451_0__144_; 
wire u2__0remHi_451_0__145_; 
wire u2__0remHi_451_0__146_; 
wire u2__0remHi_451_0__147_; 
wire u2__0remHi_451_0__148_; 
wire u2__0remHi_451_0__149_; 
wire u2__0remHi_451_0__14_; 
wire u2__0remHi_451_0__150_; 
wire u2__0remHi_451_0__151_; 
wire u2__0remHi_451_0__152_; 
wire u2__0remHi_451_0__153_; 
wire u2__0remHi_451_0__154_; 
wire u2__0remHi_451_0__155_; 
wire u2__0remHi_451_0__156_; 
wire u2__0remHi_451_0__157_; 
wire u2__0remHi_451_0__158_; 
wire u2__0remHi_451_0__159_; 
wire u2__0remHi_451_0__15_; 
wire u2__0remHi_451_0__160_; 
wire u2__0remHi_451_0__161_; 
wire u2__0remHi_451_0__162_; 
wire u2__0remHi_451_0__163_; 
wire u2__0remHi_451_0__164_; 
wire u2__0remHi_451_0__165_; 
wire u2__0remHi_451_0__166_; 
wire u2__0remHi_451_0__167_; 
wire u2__0remHi_451_0__168_; 
wire u2__0remHi_451_0__169_; 
wire u2__0remHi_451_0__16_; 
wire u2__0remHi_451_0__170_; 
wire u2__0remHi_451_0__171_; 
wire u2__0remHi_451_0__172_; 
wire u2__0remHi_451_0__173_; 
wire u2__0remHi_451_0__174_; 
wire u2__0remHi_451_0__175_; 
wire u2__0remHi_451_0__176_; 
wire u2__0remHi_451_0__177_; 
wire u2__0remHi_451_0__178_; 
wire u2__0remHi_451_0__179_; 
wire u2__0remHi_451_0__17_; 
wire u2__0remHi_451_0__180_; 
wire u2__0remHi_451_0__181_; 
wire u2__0remHi_451_0__182_; 
wire u2__0remHi_451_0__183_; 
wire u2__0remHi_451_0__184_; 
wire u2__0remHi_451_0__185_; 
wire u2__0remHi_451_0__186_; 
wire u2__0remHi_451_0__187_; 
wire u2__0remHi_451_0__188_; 
wire u2__0remHi_451_0__189_; 
wire u2__0remHi_451_0__18_; 
wire u2__0remHi_451_0__190_; 
wire u2__0remHi_451_0__191_; 
wire u2__0remHi_451_0__192_; 
wire u2__0remHi_451_0__193_; 
wire u2__0remHi_451_0__194_; 
wire u2__0remHi_451_0__195_; 
wire u2__0remHi_451_0__196_; 
wire u2__0remHi_451_0__197_; 
wire u2__0remHi_451_0__198_; 
wire u2__0remHi_451_0__199_; 
wire u2__0remHi_451_0__19_; 
wire u2__0remHi_451_0__1_; 
wire u2__0remHi_451_0__200_; 
wire u2__0remHi_451_0__201_; 
wire u2__0remHi_451_0__202_; 
wire u2__0remHi_451_0__203_; 
wire u2__0remHi_451_0__204_; 
wire u2__0remHi_451_0__205_; 
wire u2__0remHi_451_0__206_; 
wire u2__0remHi_451_0__207_; 
wire u2__0remHi_451_0__208_; 
wire u2__0remHi_451_0__209_; 
wire u2__0remHi_451_0__20_; 
wire u2__0remHi_451_0__210_; 
wire u2__0remHi_451_0__211_; 
wire u2__0remHi_451_0__212_; 
wire u2__0remHi_451_0__213_; 
wire u2__0remHi_451_0__214_; 
wire u2__0remHi_451_0__215_; 
wire u2__0remHi_451_0__216_; 
wire u2__0remHi_451_0__217_; 
wire u2__0remHi_451_0__218_; 
wire u2__0remHi_451_0__219_; 
wire u2__0remHi_451_0__21_; 
wire u2__0remHi_451_0__220_; 
wire u2__0remHi_451_0__221_; 
wire u2__0remHi_451_0__222_; 
wire u2__0remHi_451_0__223_; 
wire u2__0remHi_451_0__224_; 
wire u2__0remHi_451_0__225_; 
wire u2__0remHi_451_0__226_; 
wire u2__0remHi_451_0__227_; 
wire u2__0remHi_451_0__228_; 
wire u2__0remHi_451_0__229_; 
wire u2__0remHi_451_0__22_; 
wire u2__0remHi_451_0__230_; 
wire u2__0remHi_451_0__231_; 
wire u2__0remHi_451_0__232_; 
wire u2__0remHi_451_0__233_; 
wire u2__0remHi_451_0__234_; 
wire u2__0remHi_451_0__235_; 
wire u2__0remHi_451_0__236_; 
wire u2__0remHi_451_0__237_; 
wire u2__0remHi_451_0__238_; 
wire u2__0remHi_451_0__239_; 
wire u2__0remHi_451_0__23_; 
wire u2__0remHi_451_0__240_; 
wire u2__0remHi_451_0__241_; 
wire u2__0remHi_451_0__242_; 
wire u2__0remHi_451_0__243_; 
wire u2__0remHi_451_0__244_; 
wire u2__0remHi_451_0__245_; 
wire u2__0remHi_451_0__246_; 
wire u2__0remHi_451_0__247_; 
wire u2__0remHi_451_0__248_; 
wire u2__0remHi_451_0__249_; 
wire u2__0remHi_451_0__24_; 
wire u2__0remHi_451_0__250_; 
wire u2__0remHi_451_0__251_; 
wire u2__0remHi_451_0__252_; 
wire u2__0remHi_451_0__253_; 
wire u2__0remHi_451_0__254_; 
wire u2__0remHi_451_0__255_; 
wire u2__0remHi_451_0__256_; 
wire u2__0remHi_451_0__257_; 
wire u2__0remHi_451_0__258_; 
wire u2__0remHi_451_0__259_; 
wire u2__0remHi_451_0__25_; 
wire u2__0remHi_451_0__260_; 
wire u2__0remHi_451_0__261_; 
wire u2__0remHi_451_0__262_; 
wire u2__0remHi_451_0__263_; 
wire u2__0remHi_451_0__264_; 
wire u2__0remHi_451_0__265_; 
wire u2__0remHi_451_0__266_; 
wire u2__0remHi_451_0__267_; 
wire u2__0remHi_451_0__268_; 
wire u2__0remHi_451_0__269_; 
wire u2__0remHi_451_0__26_; 
wire u2__0remHi_451_0__270_; 
wire u2__0remHi_451_0__271_; 
wire u2__0remHi_451_0__272_; 
wire u2__0remHi_451_0__273_; 
wire u2__0remHi_451_0__274_; 
wire u2__0remHi_451_0__275_; 
wire u2__0remHi_451_0__276_; 
wire u2__0remHi_451_0__277_; 
wire u2__0remHi_451_0__278_; 
wire u2__0remHi_451_0__279_; 
wire u2__0remHi_451_0__27_; 
wire u2__0remHi_451_0__280_; 
wire u2__0remHi_451_0__281_; 
wire u2__0remHi_451_0__282_; 
wire u2__0remHi_451_0__283_; 
wire u2__0remHi_451_0__284_; 
wire u2__0remHi_451_0__285_; 
wire u2__0remHi_451_0__286_; 
wire u2__0remHi_451_0__287_; 
wire u2__0remHi_451_0__288_; 
wire u2__0remHi_451_0__289_; 
wire u2__0remHi_451_0__28_; 
wire u2__0remHi_451_0__290_; 
wire u2__0remHi_451_0__291_; 
wire u2__0remHi_451_0__292_; 
wire u2__0remHi_451_0__293_; 
wire u2__0remHi_451_0__294_; 
wire u2__0remHi_451_0__295_; 
wire u2__0remHi_451_0__296_; 
wire u2__0remHi_451_0__297_; 
wire u2__0remHi_451_0__298_; 
wire u2__0remHi_451_0__299_; 
wire u2__0remHi_451_0__29_; 
wire u2__0remHi_451_0__2_; 
wire u2__0remHi_451_0__300_; 
wire u2__0remHi_451_0__301_; 
wire u2__0remHi_451_0__302_; 
wire u2__0remHi_451_0__303_; 
wire u2__0remHi_451_0__304_; 
wire u2__0remHi_451_0__305_; 
wire u2__0remHi_451_0__306_; 
wire u2__0remHi_451_0__307_; 
wire u2__0remHi_451_0__308_; 
wire u2__0remHi_451_0__309_; 
wire u2__0remHi_451_0__30_; 
wire u2__0remHi_451_0__310_; 
wire u2__0remHi_451_0__311_; 
wire u2__0remHi_451_0__312_; 
wire u2__0remHi_451_0__313_; 
wire u2__0remHi_451_0__314_; 
wire u2__0remHi_451_0__315_; 
wire u2__0remHi_451_0__316_; 
wire u2__0remHi_451_0__317_; 
wire u2__0remHi_451_0__318_; 
wire u2__0remHi_451_0__319_; 
wire u2__0remHi_451_0__31_; 
wire u2__0remHi_451_0__320_; 
wire u2__0remHi_451_0__321_; 
wire u2__0remHi_451_0__322_; 
wire u2__0remHi_451_0__323_; 
wire u2__0remHi_451_0__324_; 
wire u2__0remHi_451_0__325_; 
wire u2__0remHi_451_0__326_; 
wire u2__0remHi_451_0__327_; 
wire u2__0remHi_451_0__328_; 
wire u2__0remHi_451_0__329_; 
wire u2__0remHi_451_0__32_; 
wire u2__0remHi_451_0__330_; 
wire u2__0remHi_451_0__331_; 
wire u2__0remHi_451_0__332_; 
wire u2__0remHi_451_0__333_; 
wire u2__0remHi_451_0__334_; 
wire u2__0remHi_451_0__335_; 
wire u2__0remHi_451_0__336_; 
wire u2__0remHi_451_0__337_; 
wire u2__0remHi_451_0__338_; 
wire u2__0remHi_451_0__339_; 
wire u2__0remHi_451_0__33_; 
wire u2__0remHi_451_0__340_; 
wire u2__0remHi_451_0__341_; 
wire u2__0remHi_451_0__342_; 
wire u2__0remHi_451_0__343_; 
wire u2__0remHi_451_0__344_; 
wire u2__0remHi_451_0__345_; 
wire u2__0remHi_451_0__346_; 
wire u2__0remHi_451_0__347_; 
wire u2__0remHi_451_0__348_; 
wire u2__0remHi_451_0__349_; 
wire u2__0remHi_451_0__34_; 
wire u2__0remHi_451_0__350_; 
wire u2__0remHi_451_0__351_; 
wire u2__0remHi_451_0__352_; 
wire u2__0remHi_451_0__353_; 
wire u2__0remHi_451_0__354_; 
wire u2__0remHi_451_0__355_; 
wire u2__0remHi_451_0__356_; 
wire u2__0remHi_451_0__357_; 
wire u2__0remHi_451_0__358_; 
wire u2__0remHi_451_0__359_; 
wire u2__0remHi_451_0__35_; 
wire u2__0remHi_451_0__360_; 
wire u2__0remHi_451_0__361_; 
wire u2__0remHi_451_0__362_; 
wire u2__0remHi_451_0__363_; 
wire u2__0remHi_451_0__364_; 
wire u2__0remHi_451_0__365_; 
wire u2__0remHi_451_0__366_; 
wire u2__0remHi_451_0__367_; 
wire u2__0remHi_451_0__368_; 
wire u2__0remHi_451_0__369_; 
wire u2__0remHi_451_0__36_; 
wire u2__0remHi_451_0__370_; 
wire u2__0remHi_451_0__371_; 
wire u2__0remHi_451_0__372_; 
wire u2__0remHi_451_0__373_; 
wire u2__0remHi_451_0__374_; 
wire u2__0remHi_451_0__375_; 
wire u2__0remHi_451_0__376_; 
wire u2__0remHi_451_0__377_; 
wire u2__0remHi_451_0__378_; 
wire u2__0remHi_451_0__379_; 
wire u2__0remHi_451_0__37_; 
wire u2__0remHi_451_0__380_; 
wire u2__0remHi_451_0__381_; 
wire u2__0remHi_451_0__382_; 
wire u2__0remHi_451_0__383_; 
wire u2__0remHi_451_0__384_; 
wire u2__0remHi_451_0__385_; 
wire u2__0remHi_451_0__386_; 
wire u2__0remHi_451_0__387_; 
wire u2__0remHi_451_0__388_; 
wire u2__0remHi_451_0__389_; 
wire u2__0remHi_451_0__38_; 
wire u2__0remHi_451_0__390_; 
wire u2__0remHi_451_0__391_; 
wire u2__0remHi_451_0__392_; 
wire u2__0remHi_451_0__393_; 
wire u2__0remHi_451_0__394_; 
wire u2__0remHi_451_0__395_; 
wire u2__0remHi_451_0__396_; 
wire u2__0remHi_451_0__397_; 
wire u2__0remHi_451_0__398_; 
wire u2__0remHi_451_0__399_; 
wire u2__0remHi_451_0__39_; 
wire u2__0remHi_451_0__3_; 
wire u2__0remHi_451_0__400_; 
wire u2__0remHi_451_0__401_; 
wire u2__0remHi_451_0__402_; 
wire u2__0remHi_451_0__403_; 
wire u2__0remHi_451_0__404_; 
wire u2__0remHi_451_0__405_; 
wire u2__0remHi_451_0__406_; 
wire u2__0remHi_451_0__407_; 
wire u2__0remHi_451_0__408_; 
wire u2__0remHi_451_0__409_; 
wire u2__0remHi_451_0__40_; 
wire u2__0remHi_451_0__410_; 
wire u2__0remHi_451_0__411_; 
wire u2__0remHi_451_0__412_; 
wire u2__0remHi_451_0__413_; 
wire u2__0remHi_451_0__414_; 
wire u2__0remHi_451_0__415_; 
wire u2__0remHi_451_0__416_; 
wire u2__0remHi_451_0__417_; 
wire u2__0remHi_451_0__418_; 
wire u2__0remHi_451_0__419_; 
wire u2__0remHi_451_0__41_; 
wire u2__0remHi_451_0__420_; 
wire u2__0remHi_451_0__421_; 
wire u2__0remHi_451_0__422_; 
wire u2__0remHi_451_0__423_; 
wire u2__0remHi_451_0__424_; 
wire u2__0remHi_451_0__425_; 
wire u2__0remHi_451_0__426_; 
wire u2__0remHi_451_0__427_; 
wire u2__0remHi_451_0__428_; 
wire u2__0remHi_451_0__429_; 
wire u2__0remHi_451_0__42_; 
wire u2__0remHi_451_0__430_; 
wire u2__0remHi_451_0__431_; 
wire u2__0remHi_451_0__432_; 
wire u2__0remHi_451_0__433_; 
wire u2__0remHi_451_0__434_; 
wire u2__0remHi_451_0__435_; 
wire u2__0remHi_451_0__436_; 
wire u2__0remHi_451_0__437_; 
wire u2__0remHi_451_0__438_; 
wire u2__0remHi_451_0__439_; 
wire u2__0remHi_451_0__43_; 
wire u2__0remHi_451_0__440_; 
wire u2__0remHi_451_0__441_; 
wire u2__0remHi_451_0__442_; 
wire u2__0remHi_451_0__443_; 
wire u2__0remHi_451_0__444_; 
wire u2__0remHi_451_0__445_; 
wire u2__0remHi_451_0__446_; 
wire u2__0remHi_451_0__447_; 
wire u2__0remHi_451_0__448_; 
wire u2__0remHi_451_0__449_; 
wire u2__0remHi_451_0__44_; 
wire u2__0remHi_451_0__45_; 
wire u2__0remHi_451_0__46_; 
wire u2__0remHi_451_0__47_; 
wire u2__0remHi_451_0__48_; 
wire u2__0remHi_451_0__49_; 
wire u2__0remHi_451_0__4_; 
wire u2__0remHi_451_0__50_; 
wire u2__0remHi_451_0__51_; 
wire u2__0remHi_451_0__52_; 
wire u2__0remHi_451_0__53_; 
wire u2__0remHi_451_0__54_; 
wire u2__0remHi_451_0__55_; 
wire u2__0remHi_451_0__56_; 
wire u2__0remHi_451_0__57_; 
wire u2__0remHi_451_0__58_; 
wire u2__0remHi_451_0__59_; 
wire u2__0remHi_451_0__5_; 
wire u2__0remHi_451_0__60_; 
wire u2__0remHi_451_0__61_; 
wire u2__0remHi_451_0__62_; 
wire u2__0remHi_451_0__63_; 
wire u2__0remHi_451_0__64_; 
wire u2__0remHi_451_0__65_; 
wire u2__0remHi_451_0__66_; 
wire u2__0remHi_451_0__67_; 
wire u2__0remHi_451_0__68_; 
wire u2__0remHi_451_0__69_; 
wire u2__0remHi_451_0__6_; 
wire u2__0remHi_451_0__70_; 
wire u2__0remHi_451_0__71_; 
wire u2__0remHi_451_0__72_; 
wire u2__0remHi_451_0__73_; 
wire u2__0remHi_451_0__74_; 
wire u2__0remHi_451_0__75_; 
wire u2__0remHi_451_0__76_; 
wire u2__0remHi_451_0__77_; 
wire u2__0remHi_451_0__78_; 
wire u2__0remHi_451_0__79_; 
wire u2__0remHi_451_0__7_; 
wire u2__0remHi_451_0__80_; 
wire u2__0remHi_451_0__81_; 
wire u2__0remHi_451_0__82_; 
wire u2__0remHi_451_0__83_; 
wire u2__0remHi_451_0__84_; 
wire u2__0remHi_451_0__85_; 
wire u2__0remHi_451_0__86_; 
wire u2__0remHi_451_0__87_; 
wire u2__0remHi_451_0__88_; 
wire u2__0remHi_451_0__89_; 
wire u2__0remHi_451_0__8_; 
wire u2__0remHi_451_0__90_; 
wire u2__0remHi_451_0__91_; 
wire u2__0remHi_451_0__92_; 
wire u2__0remHi_451_0__93_; 
wire u2__0remHi_451_0__94_; 
wire u2__0remHi_451_0__95_; 
wire u2__0remHi_451_0__96_; 
wire u2__0remHi_451_0__97_; 
wire u2__0remHi_451_0__98_; 
wire u2__0remHi_451_0__99_; 
wire u2__0remHi_451_0__9_; 
wire u2__0remLo_451_0__0_; 
wire u2__0remLo_451_0__100_; 
wire u2__0remLo_451_0__101_; 
wire u2__0remLo_451_0__102_; 
wire u2__0remLo_451_0__103_; 
wire u2__0remLo_451_0__104_; 
wire u2__0remLo_451_0__105_; 
wire u2__0remLo_451_0__106_; 
wire u2__0remLo_451_0__107_; 
wire u2__0remLo_451_0__108_; 
wire u2__0remLo_451_0__109_; 
wire u2__0remLo_451_0__10_; 
wire u2__0remLo_451_0__110_; 
wire u2__0remLo_451_0__111_; 
wire u2__0remLo_451_0__112_; 
wire u2__0remLo_451_0__113_; 
wire u2__0remLo_451_0__114_; 
wire u2__0remLo_451_0__115_; 
wire u2__0remLo_451_0__116_; 
wire u2__0remLo_451_0__117_; 
wire u2__0remLo_451_0__118_; 
wire u2__0remLo_451_0__119_; 
wire u2__0remLo_451_0__11_; 
wire u2__0remLo_451_0__120_; 
wire u2__0remLo_451_0__121_; 
wire u2__0remLo_451_0__122_; 
wire u2__0remLo_451_0__123_; 
wire u2__0remLo_451_0__124_; 
wire u2__0remLo_451_0__125_; 
wire u2__0remLo_451_0__126_; 
wire u2__0remLo_451_0__127_; 
wire u2__0remLo_451_0__128_; 
wire u2__0remLo_451_0__129_; 
wire u2__0remLo_451_0__12_; 
wire u2__0remLo_451_0__130_; 
wire u2__0remLo_451_0__131_; 
wire u2__0remLo_451_0__132_; 
wire u2__0remLo_451_0__133_; 
wire u2__0remLo_451_0__134_; 
wire u2__0remLo_451_0__135_; 
wire u2__0remLo_451_0__136_; 
wire u2__0remLo_451_0__137_; 
wire u2__0remLo_451_0__138_; 
wire u2__0remLo_451_0__139_; 
wire u2__0remLo_451_0__13_; 
wire u2__0remLo_451_0__140_; 
wire u2__0remLo_451_0__141_; 
wire u2__0remLo_451_0__142_; 
wire u2__0remLo_451_0__143_; 
wire u2__0remLo_451_0__144_; 
wire u2__0remLo_451_0__145_; 
wire u2__0remLo_451_0__146_; 
wire u2__0remLo_451_0__147_; 
wire u2__0remLo_451_0__148_; 
wire u2__0remLo_451_0__149_; 
wire u2__0remLo_451_0__14_; 
wire u2__0remLo_451_0__150_; 
wire u2__0remLo_451_0__151_; 
wire u2__0remLo_451_0__152_; 
wire u2__0remLo_451_0__153_; 
wire u2__0remLo_451_0__154_; 
wire u2__0remLo_451_0__155_; 
wire u2__0remLo_451_0__156_; 
wire u2__0remLo_451_0__157_; 
wire u2__0remLo_451_0__158_; 
wire u2__0remLo_451_0__159_; 
wire u2__0remLo_451_0__15_; 
wire u2__0remLo_451_0__160_; 
wire u2__0remLo_451_0__161_; 
wire u2__0remLo_451_0__162_; 
wire u2__0remLo_451_0__163_; 
wire u2__0remLo_451_0__164_; 
wire u2__0remLo_451_0__165_; 
wire u2__0remLo_451_0__166_; 
wire u2__0remLo_451_0__167_; 
wire u2__0remLo_451_0__168_; 
wire u2__0remLo_451_0__169_; 
wire u2__0remLo_451_0__16_; 
wire u2__0remLo_451_0__170_; 
wire u2__0remLo_451_0__171_; 
wire u2__0remLo_451_0__172_; 
wire u2__0remLo_451_0__173_; 
wire u2__0remLo_451_0__174_; 
wire u2__0remLo_451_0__175_; 
wire u2__0remLo_451_0__176_; 
wire u2__0remLo_451_0__177_; 
wire u2__0remLo_451_0__178_; 
wire u2__0remLo_451_0__179_; 
wire u2__0remLo_451_0__17_; 
wire u2__0remLo_451_0__180_; 
wire u2__0remLo_451_0__181_; 
wire u2__0remLo_451_0__182_; 
wire u2__0remLo_451_0__183_; 
wire u2__0remLo_451_0__184_; 
wire u2__0remLo_451_0__185_; 
wire u2__0remLo_451_0__186_; 
wire u2__0remLo_451_0__187_; 
wire u2__0remLo_451_0__188_; 
wire u2__0remLo_451_0__189_; 
wire u2__0remLo_451_0__18_; 
wire u2__0remLo_451_0__190_; 
wire u2__0remLo_451_0__191_; 
wire u2__0remLo_451_0__192_; 
wire u2__0remLo_451_0__193_; 
wire u2__0remLo_451_0__194_; 
wire u2__0remLo_451_0__195_; 
wire u2__0remLo_451_0__196_; 
wire u2__0remLo_451_0__197_; 
wire u2__0remLo_451_0__198_; 
wire u2__0remLo_451_0__199_; 
wire u2__0remLo_451_0__19_; 
wire u2__0remLo_451_0__1_; 
wire u2__0remLo_451_0__200_; 
wire u2__0remLo_451_0__201_; 
wire u2__0remLo_451_0__202_; 
wire u2__0remLo_451_0__203_; 
wire u2__0remLo_451_0__204_; 
wire u2__0remLo_451_0__205_; 
wire u2__0remLo_451_0__206_; 
wire u2__0remLo_451_0__207_; 
wire u2__0remLo_451_0__208_; 
wire u2__0remLo_451_0__209_; 
wire u2__0remLo_451_0__20_; 
wire u2__0remLo_451_0__210_; 
wire u2__0remLo_451_0__211_; 
wire u2__0remLo_451_0__212_; 
wire u2__0remLo_451_0__213_; 
wire u2__0remLo_451_0__214_; 
wire u2__0remLo_451_0__215_; 
wire u2__0remLo_451_0__216_; 
wire u2__0remLo_451_0__217_; 
wire u2__0remLo_451_0__218_; 
wire u2__0remLo_451_0__219_; 
wire u2__0remLo_451_0__21_; 
wire u2__0remLo_451_0__220_; 
wire u2__0remLo_451_0__221_; 
wire u2__0remLo_451_0__222_; 
wire u2__0remLo_451_0__223_; 
wire u2__0remLo_451_0__224_; 
wire u2__0remLo_451_0__225_; 
wire u2__0remLo_451_0__226_; 
wire u2__0remLo_451_0__227_; 
wire u2__0remLo_451_0__228_; 
wire u2__0remLo_451_0__229_; 
wire u2__0remLo_451_0__22_; 
wire u2__0remLo_451_0__230_; 
wire u2__0remLo_451_0__231_; 
wire u2__0remLo_451_0__232_; 
wire u2__0remLo_451_0__233_; 
wire u2__0remLo_451_0__234_; 
wire u2__0remLo_451_0__235_; 
wire u2__0remLo_451_0__236_; 
wire u2__0remLo_451_0__237_; 
wire u2__0remLo_451_0__238_; 
wire u2__0remLo_451_0__239_; 
wire u2__0remLo_451_0__23_; 
wire u2__0remLo_451_0__240_; 
wire u2__0remLo_451_0__241_; 
wire u2__0remLo_451_0__242_; 
wire u2__0remLo_451_0__243_; 
wire u2__0remLo_451_0__244_; 
wire u2__0remLo_451_0__245_; 
wire u2__0remLo_451_0__246_; 
wire u2__0remLo_451_0__247_; 
wire u2__0remLo_451_0__248_; 
wire u2__0remLo_451_0__249_; 
wire u2__0remLo_451_0__24_; 
wire u2__0remLo_451_0__250_; 
wire u2__0remLo_451_0__251_; 
wire u2__0remLo_451_0__252_; 
wire u2__0remLo_451_0__253_; 
wire u2__0remLo_451_0__254_; 
wire u2__0remLo_451_0__255_; 
wire u2__0remLo_451_0__256_; 
wire u2__0remLo_451_0__257_; 
wire u2__0remLo_451_0__258_; 
wire u2__0remLo_451_0__259_; 
wire u2__0remLo_451_0__25_; 
wire u2__0remLo_451_0__260_; 
wire u2__0remLo_451_0__261_; 
wire u2__0remLo_451_0__262_; 
wire u2__0remLo_451_0__263_; 
wire u2__0remLo_451_0__264_; 
wire u2__0remLo_451_0__265_; 
wire u2__0remLo_451_0__266_; 
wire u2__0remLo_451_0__267_; 
wire u2__0remLo_451_0__268_; 
wire u2__0remLo_451_0__269_; 
wire u2__0remLo_451_0__26_; 
wire u2__0remLo_451_0__270_; 
wire u2__0remLo_451_0__271_; 
wire u2__0remLo_451_0__272_; 
wire u2__0remLo_451_0__273_; 
wire u2__0remLo_451_0__274_; 
wire u2__0remLo_451_0__275_; 
wire u2__0remLo_451_0__276_; 
wire u2__0remLo_451_0__277_; 
wire u2__0remLo_451_0__278_; 
wire u2__0remLo_451_0__279_; 
wire u2__0remLo_451_0__27_; 
wire u2__0remLo_451_0__280_; 
wire u2__0remLo_451_0__281_; 
wire u2__0remLo_451_0__282_; 
wire u2__0remLo_451_0__283_; 
wire u2__0remLo_451_0__284_; 
wire u2__0remLo_451_0__285_; 
wire u2__0remLo_451_0__286_; 
wire u2__0remLo_451_0__287_; 
wire u2__0remLo_451_0__288_; 
wire u2__0remLo_451_0__289_; 
wire u2__0remLo_451_0__28_; 
wire u2__0remLo_451_0__290_; 
wire u2__0remLo_451_0__291_; 
wire u2__0remLo_451_0__292_; 
wire u2__0remLo_451_0__293_; 
wire u2__0remLo_451_0__294_; 
wire u2__0remLo_451_0__295_; 
wire u2__0remLo_451_0__296_; 
wire u2__0remLo_451_0__297_; 
wire u2__0remLo_451_0__298_; 
wire u2__0remLo_451_0__299_; 
wire u2__0remLo_451_0__29_; 
wire u2__0remLo_451_0__2_; 
wire u2__0remLo_451_0__300_; 
wire u2__0remLo_451_0__301_; 
wire u2__0remLo_451_0__302_; 
wire u2__0remLo_451_0__303_; 
wire u2__0remLo_451_0__304_; 
wire u2__0remLo_451_0__305_; 
wire u2__0remLo_451_0__306_; 
wire u2__0remLo_451_0__307_; 
wire u2__0remLo_451_0__308_; 
wire u2__0remLo_451_0__309_; 
wire u2__0remLo_451_0__30_; 
wire u2__0remLo_451_0__310_; 
wire u2__0remLo_451_0__311_; 
wire u2__0remLo_451_0__312_; 
wire u2__0remLo_451_0__313_; 
wire u2__0remLo_451_0__314_; 
wire u2__0remLo_451_0__315_; 
wire u2__0remLo_451_0__316_; 
wire u2__0remLo_451_0__317_; 
wire u2__0remLo_451_0__318_; 
wire u2__0remLo_451_0__319_; 
wire u2__0remLo_451_0__31_; 
wire u2__0remLo_451_0__320_; 
wire u2__0remLo_451_0__321_; 
wire u2__0remLo_451_0__322_; 
wire u2__0remLo_451_0__323_; 
wire u2__0remLo_451_0__324_; 
wire u2__0remLo_451_0__325_; 
wire u2__0remLo_451_0__326_; 
wire u2__0remLo_451_0__327_; 
wire u2__0remLo_451_0__328_; 
wire u2__0remLo_451_0__329_; 
wire u2__0remLo_451_0__32_; 
wire u2__0remLo_451_0__330_; 
wire u2__0remLo_451_0__331_; 
wire u2__0remLo_451_0__332_; 
wire u2__0remLo_451_0__333_; 
wire u2__0remLo_451_0__334_; 
wire u2__0remLo_451_0__335_; 
wire u2__0remLo_451_0__336_; 
wire u2__0remLo_451_0__337_; 
wire u2__0remLo_451_0__338_; 
wire u2__0remLo_451_0__339_; 
wire u2__0remLo_451_0__33_; 
wire u2__0remLo_451_0__340_; 
wire u2__0remLo_451_0__341_; 
wire u2__0remLo_451_0__342_; 
wire u2__0remLo_451_0__343_; 
wire u2__0remLo_451_0__344_; 
wire u2__0remLo_451_0__345_; 
wire u2__0remLo_451_0__346_; 
wire u2__0remLo_451_0__347_; 
wire u2__0remLo_451_0__348_; 
wire u2__0remLo_451_0__349_; 
wire u2__0remLo_451_0__34_; 
wire u2__0remLo_451_0__350_; 
wire u2__0remLo_451_0__351_; 
wire u2__0remLo_451_0__352_; 
wire u2__0remLo_451_0__353_; 
wire u2__0remLo_451_0__354_; 
wire u2__0remLo_451_0__355_; 
wire u2__0remLo_451_0__356_; 
wire u2__0remLo_451_0__357_; 
wire u2__0remLo_451_0__358_; 
wire u2__0remLo_451_0__359_; 
wire u2__0remLo_451_0__35_; 
wire u2__0remLo_451_0__360_; 
wire u2__0remLo_451_0__361_; 
wire u2__0remLo_451_0__362_; 
wire u2__0remLo_451_0__363_; 
wire u2__0remLo_451_0__364_; 
wire u2__0remLo_451_0__365_; 
wire u2__0remLo_451_0__366_; 
wire u2__0remLo_451_0__367_; 
wire u2__0remLo_451_0__368_; 
wire u2__0remLo_451_0__369_; 
wire u2__0remLo_451_0__36_; 
wire u2__0remLo_451_0__370_; 
wire u2__0remLo_451_0__371_; 
wire u2__0remLo_451_0__372_; 
wire u2__0remLo_451_0__373_; 
wire u2__0remLo_451_0__374_; 
wire u2__0remLo_451_0__375_; 
wire u2__0remLo_451_0__376_; 
wire u2__0remLo_451_0__377_; 
wire u2__0remLo_451_0__378_; 
wire u2__0remLo_451_0__379_; 
wire u2__0remLo_451_0__37_; 
wire u2__0remLo_451_0__380_; 
wire u2__0remLo_451_0__381_; 
wire u2__0remLo_451_0__382_; 
wire u2__0remLo_451_0__383_; 
wire u2__0remLo_451_0__384_; 
wire u2__0remLo_451_0__385_; 
wire u2__0remLo_451_0__386_; 
wire u2__0remLo_451_0__387_; 
wire u2__0remLo_451_0__388_; 
wire u2__0remLo_451_0__389_; 
wire u2__0remLo_451_0__38_; 
wire u2__0remLo_451_0__390_; 
wire u2__0remLo_451_0__391_; 
wire u2__0remLo_451_0__392_; 
wire u2__0remLo_451_0__393_; 
wire u2__0remLo_451_0__394_; 
wire u2__0remLo_451_0__395_; 
wire u2__0remLo_451_0__396_; 
wire u2__0remLo_451_0__397_; 
wire u2__0remLo_451_0__398_; 
wire u2__0remLo_451_0__399_; 
wire u2__0remLo_451_0__39_; 
wire u2__0remLo_451_0__3_; 
wire u2__0remLo_451_0__400_; 
wire u2__0remLo_451_0__401_; 
wire u2__0remLo_451_0__402_; 
wire u2__0remLo_451_0__403_; 
wire u2__0remLo_451_0__404_; 
wire u2__0remLo_451_0__405_; 
wire u2__0remLo_451_0__406_; 
wire u2__0remLo_451_0__407_; 
wire u2__0remLo_451_0__408_; 
wire u2__0remLo_451_0__409_; 
wire u2__0remLo_451_0__40_; 
wire u2__0remLo_451_0__410_; 
wire u2__0remLo_451_0__411_; 
wire u2__0remLo_451_0__412_; 
wire u2__0remLo_451_0__413_; 
wire u2__0remLo_451_0__414_; 
wire u2__0remLo_451_0__415_; 
wire u2__0remLo_451_0__416_; 
wire u2__0remLo_451_0__417_; 
wire u2__0remLo_451_0__418_; 
wire u2__0remLo_451_0__419_; 
wire u2__0remLo_451_0__41_; 
wire u2__0remLo_451_0__420_; 
wire u2__0remLo_451_0__421_; 
wire u2__0remLo_451_0__422_; 
wire u2__0remLo_451_0__423_; 
wire u2__0remLo_451_0__424_; 
wire u2__0remLo_451_0__425_; 
wire u2__0remLo_451_0__426_; 
wire u2__0remLo_451_0__427_; 
wire u2__0remLo_451_0__428_; 
wire u2__0remLo_451_0__429_; 
wire u2__0remLo_451_0__42_; 
wire u2__0remLo_451_0__430_; 
wire u2__0remLo_451_0__431_; 
wire u2__0remLo_451_0__432_; 
wire u2__0remLo_451_0__433_; 
wire u2__0remLo_451_0__434_; 
wire u2__0remLo_451_0__435_; 
wire u2__0remLo_451_0__436_; 
wire u2__0remLo_451_0__437_; 
wire u2__0remLo_451_0__438_; 
wire u2__0remLo_451_0__439_; 
wire u2__0remLo_451_0__43_; 
wire u2__0remLo_451_0__440_; 
wire u2__0remLo_451_0__441_; 
wire u2__0remLo_451_0__442_; 
wire u2__0remLo_451_0__443_; 
wire u2__0remLo_451_0__444_; 
wire u2__0remLo_451_0__445_; 
wire u2__0remLo_451_0__446_; 
wire u2__0remLo_451_0__447_; 
wire u2__0remLo_451_0__448_; 
wire u2__0remLo_451_0__449_; 
wire u2__0remLo_451_0__44_; 
wire u2__0remLo_451_0__450_; 
wire u2__0remLo_451_0__451_; 
wire u2__0remLo_451_0__45_; 
wire u2__0remLo_451_0__46_; 
wire u2__0remLo_451_0__47_; 
wire u2__0remLo_451_0__48_; 
wire u2__0remLo_451_0__49_; 
wire u2__0remLo_451_0__4_; 
wire u2__0remLo_451_0__50_; 
wire u2__0remLo_451_0__51_; 
wire u2__0remLo_451_0__52_; 
wire u2__0remLo_451_0__53_; 
wire u2__0remLo_451_0__54_; 
wire u2__0remLo_451_0__55_; 
wire u2__0remLo_451_0__56_; 
wire u2__0remLo_451_0__57_; 
wire u2__0remLo_451_0__58_; 
wire u2__0remLo_451_0__59_; 
wire u2__0remLo_451_0__5_; 
wire u2__0remLo_451_0__60_; 
wire u2__0remLo_451_0__61_; 
wire u2__0remLo_451_0__62_; 
wire u2__0remLo_451_0__63_; 
wire u2__0remLo_451_0__64_; 
wire u2__0remLo_451_0__65_; 
wire u2__0remLo_451_0__66_; 
wire u2__0remLo_451_0__67_; 
wire u2__0remLo_451_0__68_; 
wire u2__0remLo_451_0__69_; 
wire u2__0remLo_451_0__6_; 
wire u2__0remLo_451_0__70_; 
wire u2__0remLo_451_0__71_; 
wire u2__0remLo_451_0__72_; 
wire u2__0remLo_451_0__73_; 
wire u2__0remLo_451_0__74_; 
wire u2__0remLo_451_0__75_; 
wire u2__0remLo_451_0__76_; 
wire u2__0remLo_451_0__77_; 
wire u2__0remLo_451_0__78_; 
wire u2__0remLo_451_0__79_; 
wire u2__0remLo_451_0__7_; 
wire u2__0remLo_451_0__80_; 
wire u2__0remLo_451_0__81_; 
wire u2__0remLo_451_0__82_; 
wire u2__0remLo_451_0__83_; 
wire u2__0remLo_451_0__84_; 
wire u2__0remLo_451_0__85_; 
wire u2__0remLo_451_0__86_; 
wire u2__0remLo_451_0__87_; 
wire u2__0remLo_451_0__88_; 
wire u2__0remLo_451_0__89_; 
wire u2__0remLo_451_0__8_; 
wire u2__0remLo_451_0__90_; 
wire u2__0remLo_451_0__91_; 
wire u2__0remLo_451_0__92_; 
wire u2__0remLo_451_0__93_; 
wire u2__0remLo_451_0__94_; 
wire u2__0remLo_451_0__95_; 
wire u2__0remLo_451_0__96_; 
wire u2__0remLo_451_0__97_; 
wire u2__0remLo_451_0__98_; 
wire u2__0remLo_451_0__99_; 
wire u2__0remLo_451_0__9_; 
wire u2__0root_452_0__0_; 
wire u2__0root_452_0__100_; 
wire u2__0root_452_0__101_; 
wire u2__0root_452_0__102_; 
wire u2__0root_452_0__103_; 
wire u2__0root_452_0__104_; 
wire u2__0root_452_0__105_; 
wire u2__0root_452_0__106_; 
wire u2__0root_452_0__107_; 
wire u2__0root_452_0__108_; 
wire u2__0root_452_0__109_; 
wire u2__0root_452_0__10_; 
wire u2__0root_452_0__110_; 
wire u2__0root_452_0__111_; 
wire u2__0root_452_0__112_; 
wire u2__0root_452_0__113_; 
wire u2__0root_452_0__114_; 
wire u2__0root_452_0__115_; 
wire u2__0root_452_0__116_; 
wire u2__0root_452_0__117_; 
wire u2__0root_452_0__118_; 
wire u2__0root_452_0__119_; 
wire u2__0root_452_0__11_; 
wire u2__0root_452_0__120_; 
wire u2__0root_452_0__121_; 
wire u2__0root_452_0__122_; 
wire u2__0root_452_0__123_; 
wire u2__0root_452_0__124_; 
wire u2__0root_452_0__125_; 
wire u2__0root_452_0__126_; 
wire u2__0root_452_0__127_; 
wire u2__0root_452_0__128_; 
wire u2__0root_452_0__129_; 
wire u2__0root_452_0__12_; 
wire u2__0root_452_0__130_; 
wire u2__0root_452_0__131_; 
wire u2__0root_452_0__132_; 
wire u2__0root_452_0__133_; 
wire u2__0root_452_0__134_; 
wire u2__0root_452_0__135_; 
wire u2__0root_452_0__136_; 
wire u2__0root_452_0__137_; 
wire u2__0root_452_0__138_; 
wire u2__0root_452_0__139_; 
wire u2__0root_452_0__13_; 
wire u2__0root_452_0__140_; 
wire u2__0root_452_0__141_; 
wire u2__0root_452_0__142_; 
wire u2__0root_452_0__143_; 
wire u2__0root_452_0__144_; 
wire u2__0root_452_0__145_; 
wire u2__0root_452_0__146_; 
wire u2__0root_452_0__147_; 
wire u2__0root_452_0__148_; 
wire u2__0root_452_0__149_; 
wire u2__0root_452_0__14_; 
wire u2__0root_452_0__150_; 
wire u2__0root_452_0__151_; 
wire u2__0root_452_0__152_; 
wire u2__0root_452_0__153_; 
wire u2__0root_452_0__154_; 
wire u2__0root_452_0__155_; 
wire u2__0root_452_0__156_; 
wire u2__0root_452_0__157_; 
wire u2__0root_452_0__158_; 
wire u2__0root_452_0__159_; 
wire u2__0root_452_0__15_; 
wire u2__0root_452_0__160_; 
wire u2__0root_452_0__161_; 
wire u2__0root_452_0__162_; 
wire u2__0root_452_0__163_; 
wire u2__0root_452_0__164_; 
wire u2__0root_452_0__165_; 
wire u2__0root_452_0__166_; 
wire u2__0root_452_0__167_; 
wire u2__0root_452_0__168_; 
wire u2__0root_452_0__169_; 
wire u2__0root_452_0__16_; 
wire u2__0root_452_0__170_; 
wire u2__0root_452_0__171_; 
wire u2__0root_452_0__172_; 
wire u2__0root_452_0__173_; 
wire u2__0root_452_0__174_; 
wire u2__0root_452_0__175_; 
wire u2__0root_452_0__176_; 
wire u2__0root_452_0__177_; 
wire u2__0root_452_0__178_; 
wire u2__0root_452_0__179_; 
wire u2__0root_452_0__17_; 
wire u2__0root_452_0__180_; 
wire u2__0root_452_0__181_; 
wire u2__0root_452_0__182_; 
wire u2__0root_452_0__183_; 
wire u2__0root_452_0__184_; 
wire u2__0root_452_0__185_; 
wire u2__0root_452_0__186_; 
wire u2__0root_452_0__187_; 
wire u2__0root_452_0__188_; 
wire u2__0root_452_0__189_; 
wire u2__0root_452_0__18_; 
wire u2__0root_452_0__190_; 
wire u2__0root_452_0__191_; 
wire u2__0root_452_0__192_; 
wire u2__0root_452_0__193_; 
wire u2__0root_452_0__194_; 
wire u2__0root_452_0__195_; 
wire u2__0root_452_0__196_; 
wire u2__0root_452_0__197_; 
wire u2__0root_452_0__198_; 
wire u2__0root_452_0__199_; 
wire u2__0root_452_0__19_; 
wire u2__0root_452_0__1_; 
wire u2__0root_452_0__200_; 
wire u2__0root_452_0__201_; 
wire u2__0root_452_0__202_; 
wire u2__0root_452_0__203_; 
wire u2__0root_452_0__204_; 
wire u2__0root_452_0__205_; 
wire u2__0root_452_0__206_; 
wire u2__0root_452_0__207_; 
wire u2__0root_452_0__208_; 
wire u2__0root_452_0__209_; 
wire u2__0root_452_0__20_; 
wire u2__0root_452_0__210_; 
wire u2__0root_452_0__211_; 
wire u2__0root_452_0__212_; 
wire u2__0root_452_0__213_; 
wire u2__0root_452_0__214_; 
wire u2__0root_452_0__215_; 
wire u2__0root_452_0__216_; 
wire u2__0root_452_0__217_; 
wire u2__0root_452_0__218_; 
wire u2__0root_452_0__219_; 
wire u2__0root_452_0__21_; 
wire u2__0root_452_0__220_; 
wire u2__0root_452_0__221_; 
wire u2__0root_452_0__222_; 
wire u2__0root_452_0__223_; 
wire u2__0root_452_0__224_; 
wire u2__0root_452_0__225_; 
wire u2__0root_452_0__226_; 
wire u2__0root_452_0__227_; 
wire u2__0root_452_0__228_; 
wire u2__0root_452_0__229_; 
wire u2__0root_452_0__22_; 
wire u2__0root_452_0__230_; 
wire u2__0root_452_0__231_; 
wire u2__0root_452_0__232_; 
wire u2__0root_452_0__233_; 
wire u2__0root_452_0__234_; 
wire u2__0root_452_0__235_; 
wire u2__0root_452_0__236_; 
wire u2__0root_452_0__237_; 
wire u2__0root_452_0__238_; 
wire u2__0root_452_0__239_; 
wire u2__0root_452_0__23_; 
wire u2__0root_452_0__240_; 
wire u2__0root_452_0__241_; 
wire u2__0root_452_0__242_; 
wire u2__0root_452_0__243_; 
wire u2__0root_452_0__244_; 
wire u2__0root_452_0__245_; 
wire u2__0root_452_0__246_; 
wire u2__0root_452_0__247_; 
wire u2__0root_452_0__248_; 
wire u2__0root_452_0__249_; 
wire u2__0root_452_0__24_; 
wire u2__0root_452_0__250_; 
wire u2__0root_452_0__251_; 
wire u2__0root_452_0__252_; 
wire u2__0root_452_0__253_; 
wire u2__0root_452_0__254_; 
wire u2__0root_452_0__255_; 
wire u2__0root_452_0__256_; 
wire u2__0root_452_0__257_; 
wire u2__0root_452_0__258_; 
wire u2__0root_452_0__259_; 
wire u2__0root_452_0__25_; 
wire u2__0root_452_0__260_; 
wire u2__0root_452_0__261_; 
wire u2__0root_452_0__262_; 
wire u2__0root_452_0__263_; 
wire u2__0root_452_0__264_; 
wire u2__0root_452_0__265_; 
wire u2__0root_452_0__266_; 
wire u2__0root_452_0__267_; 
wire u2__0root_452_0__268_; 
wire u2__0root_452_0__269_; 
wire u2__0root_452_0__26_; 
wire u2__0root_452_0__270_; 
wire u2__0root_452_0__271_; 
wire u2__0root_452_0__272_; 
wire u2__0root_452_0__273_; 
wire u2__0root_452_0__274_; 
wire u2__0root_452_0__275_; 
wire u2__0root_452_0__276_; 
wire u2__0root_452_0__277_; 
wire u2__0root_452_0__278_; 
wire u2__0root_452_0__279_; 
wire u2__0root_452_0__27_; 
wire u2__0root_452_0__280_; 
wire u2__0root_452_0__281_; 
wire u2__0root_452_0__282_; 
wire u2__0root_452_0__283_; 
wire u2__0root_452_0__284_; 
wire u2__0root_452_0__285_; 
wire u2__0root_452_0__286_; 
wire u2__0root_452_0__287_; 
wire u2__0root_452_0__288_; 
wire u2__0root_452_0__289_; 
wire u2__0root_452_0__28_; 
wire u2__0root_452_0__290_; 
wire u2__0root_452_0__291_; 
wire u2__0root_452_0__292_; 
wire u2__0root_452_0__293_; 
wire u2__0root_452_0__294_; 
wire u2__0root_452_0__295_; 
wire u2__0root_452_0__296_; 
wire u2__0root_452_0__297_; 
wire u2__0root_452_0__298_; 
wire u2__0root_452_0__299_; 
wire u2__0root_452_0__29_; 
wire u2__0root_452_0__2_; 
wire u2__0root_452_0__300_; 
wire u2__0root_452_0__301_; 
wire u2__0root_452_0__302_; 
wire u2__0root_452_0__303_; 
wire u2__0root_452_0__304_; 
wire u2__0root_452_0__305_; 
wire u2__0root_452_0__306_; 
wire u2__0root_452_0__307_; 
wire u2__0root_452_0__308_; 
wire u2__0root_452_0__309_; 
wire u2__0root_452_0__30_; 
wire u2__0root_452_0__310_; 
wire u2__0root_452_0__311_; 
wire u2__0root_452_0__312_; 
wire u2__0root_452_0__313_; 
wire u2__0root_452_0__314_; 
wire u2__0root_452_0__315_; 
wire u2__0root_452_0__316_; 
wire u2__0root_452_0__317_; 
wire u2__0root_452_0__318_; 
wire u2__0root_452_0__319_; 
wire u2__0root_452_0__31_; 
wire u2__0root_452_0__320_; 
wire u2__0root_452_0__321_; 
wire u2__0root_452_0__322_; 
wire u2__0root_452_0__323_; 
wire u2__0root_452_0__324_; 
wire u2__0root_452_0__325_; 
wire u2__0root_452_0__326_; 
wire u2__0root_452_0__327_; 
wire u2__0root_452_0__328_; 
wire u2__0root_452_0__329_; 
wire u2__0root_452_0__32_; 
wire u2__0root_452_0__330_; 
wire u2__0root_452_0__331_; 
wire u2__0root_452_0__332_; 
wire u2__0root_452_0__333_; 
wire u2__0root_452_0__334_; 
wire u2__0root_452_0__335_; 
wire u2__0root_452_0__336_; 
wire u2__0root_452_0__337_; 
wire u2__0root_452_0__338_; 
wire u2__0root_452_0__339_; 
wire u2__0root_452_0__33_; 
wire u2__0root_452_0__340_; 
wire u2__0root_452_0__341_; 
wire u2__0root_452_0__342_; 
wire u2__0root_452_0__343_; 
wire u2__0root_452_0__344_; 
wire u2__0root_452_0__345_; 
wire u2__0root_452_0__346_; 
wire u2__0root_452_0__347_; 
wire u2__0root_452_0__348_; 
wire u2__0root_452_0__349_; 
wire u2__0root_452_0__34_; 
wire u2__0root_452_0__350_; 
wire u2__0root_452_0__351_; 
wire u2__0root_452_0__352_; 
wire u2__0root_452_0__353_; 
wire u2__0root_452_0__354_; 
wire u2__0root_452_0__355_; 
wire u2__0root_452_0__356_; 
wire u2__0root_452_0__357_; 
wire u2__0root_452_0__358_; 
wire u2__0root_452_0__359_; 
wire u2__0root_452_0__35_; 
wire u2__0root_452_0__360_; 
wire u2__0root_452_0__361_; 
wire u2__0root_452_0__362_; 
wire u2__0root_452_0__363_; 
wire u2__0root_452_0__364_; 
wire u2__0root_452_0__365_; 
wire u2__0root_452_0__366_; 
wire u2__0root_452_0__367_; 
wire u2__0root_452_0__368_; 
wire u2__0root_452_0__369_; 
wire u2__0root_452_0__36_; 
wire u2__0root_452_0__370_; 
wire u2__0root_452_0__371_; 
wire u2__0root_452_0__372_; 
wire u2__0root_452_0__373_; 
wire u2__0root_452_0__374_; 
wire u2__0root_452_0__375_; 
wire u2__0root_452_0__376_; 
wire u2__0root_452_0__377_; 
wire u2__0root_452_0__378_; 
wire u2__0root_452_0__379_; 
wire u2__0root_452_0__37_; 
wire u2__0root_452_0__380_; 
wire u2__0root_452_0__381_; 
wire u2__0root_452_0__382_; 
wire u2__0root_452_0__383_; 
wire u2__0root_452_0__384_; 
wire u2__0root_452_0__385_; 
wire u2__0root_452_0__386_; 
wire u2__0root_452_0__387_; 
wire u2__0root_452_0__388_; 
wire u2__0root_452_0__389_; 
wire u2__0root_452_0__38_; 
wire u2__0root_452_0__390_; 
wire u2__0root_452_0__391_; 
wire u2__0root_452_0__392_; 
wire u2__0root_452_0__393_; 
wire u2__0root_452_0__394_; 
wire u2__0root_452_0__395_; 
wire u2__0root_452_0__396_; 
wire u2__0root_452_0__397_; 
wire u2__0root_452_0__398_; 
wire u2__0root_452_0__399_; 
wire u2__0root_452_0__39_; 
wire u2__0root_452_0__3_; 
wire u2__0root_452_0__400_; 
wire u2__0root_452_0__401_; 
wire u2__0root_452_0__402_; 
wire u2__0root_452_0__403_; 
wire u2__0root_452_0__404_; 
wire u2__0root_452_0__405_; 
wire u2__0root_452_0__406_; 
wire u2__0root_452_0__407_; 
wire u2__0root_452_0__408_; 
wire u2__0root_452_0__409_; 
wire u2__0root_452_0__40_; 
wire u2__0root_452_0__410_; 
wire u2__0root_452_0__411_; 
wire u2__0root_452_0__412_; 
wire u2__0root_452_0__413_; 
wire u2__0root_452_0__414_; 
wire u2__0root_452_0__415_; 
wire u2__0root_452_0__416_; 
wire u2__0root_452_0__417_; 
wire u2__0root_452_0__418_; 
wire u2__0root_452_0__419_; 
wire u2__0root_452_0__41_; 
wire u2__0root_452_0__420_; 
wire u2__0root_452_0__421_; 
wire u2__0root_452_0__422_; 
wire u2__0root_452_0__423_; 
wire u2__0root_452_0__424_; 
wire u2__0root_452_0__425_; 
wire u2__0root_452_0__426_; 
wire u2__0root_452_0__427_; 
wire u2__0root_452_0__428_; 
wire u2__0root_452_0__429_; 
wire u2__0root_452_0__42_; 
wire u2__0root_452_0__430_; 
wire u2__0root_452_0__431_; 
wire u2__0root_452_0__432_; 
wire u2__0root_452_0__433_; 
wire u2__0root_452_0__434_; 
wire u2__0root_452_0__435_; 
wire u2__0root_452_0__436_; 
wire u2__0root_452_0__437_; 
wire u2__0root_452_0__438_; 
wire u2__0root_452_0__439_; 
wire u2__0root_452_0__43_; 
wire u2__0root_452_0__440_; 
wire u2__0root_452_0__441_; 
wire u2__0root_452_0__442_; 
wire u2__0root_452_0__443_; 
wire u2__0root_452_0__444_; 
wire u2__0root_452_0__445_; 
wire u2__0root_452_0__446_; 
wire u2__0root_452_0__447_; 
wire u2__0root_452_0__448_; 
wire u2__0root_452_0__449_; 
wire u2__0root_452_0__44_; 
wire u2__0root_452_0__450_; 
wire u2__0root_452_0__45_; 
wire u2__0root_452_0__46_; 
wire u2__0root_452_0__47_; 
wire u2__0root_452_0__48_; 
wire u2__0root_452_0__49_; 
wire u2__0root_452_0__4_; 
wire u2__0root_452_0__50_; 
wire u2__0root_452_0__51_; 
wire u2__0root_452_0__52_; 
wire u2__0root_452_0__53_; 
wire u2__0root_452_0__54_; 
wire u2__0root_452_0__55_; 
wire u2__0root_452_0__56_; 
wire u2__0root_452_0__57_; 
wire u2__0root_452_0__58_; 
wire u2__0root_452_0__59_; 
wire u2__0root_452_0__5_; 
wire u2__0root_452_0__60_; 
wire u2__0root_452_0__61_; 
wire u2__0root_452_0__62_; 
wire u2__0root_452_0__63_; 
wire u2__0root_452_0__64_; 
wire u2__0root_452_0__65_; 
wire u2__0root_452_0__66_; 
wire u2__0root_452_0__67_; 
wire u2__0root_452_0__68_; 
wire u2__0root_452_0__69_; 
wire u2__0root_452_0__6_; 
wire u2__0root_452_0__70_; 
wire u2__0root_452_0__71_; 
wire u2__0root_452_0__72_; 
wire u2__0root_452_0__73_; 
wire u2__0root_452_0__74_; 
wire u2__0root_452_0__75_; 
wire u2__0root_452_0__76_; 
wire u2__0root_452_0__77_; 
wire u2__0root_452_0__78_; 
wire u2__0root_452_0__79_; 
wire u2__0root_452_0__7_; 
wire u2__0root_452_0__80_; 
wire u2__0root_452_0__81_; 
wire u2__0root_452_0__82_; 
wire u2__0root_452_0__83_; 
wire u2__0root_452_0__84_; 
wire u2__0root_452_0__85_; 
wire u2__0root_452_0__86_; 
wire u2__0root_452_0__87_; 
wire u2__0root_452_0__88_; 
wire u2__0root_452_0__89_; 
wire u2__0root_452_0__8_; 
wire u2__0root_452_0__90_; 
wire u2__0root_452_0__91_; 
wire u2__0root_452_0__92_; 
wire u2__0root_452_0__93_; 
wire u2__0root_452_0__94_; 
wire u2__0root_452_0__95_; 
wire u2__0root_452_0__96_; 
wire u2__0root_452_0__97_; 
wire u2__0root_452_0__98_; 
wire u2__0root_452_0__99_; 
wire u2__0root_452_0__9_; 
wire u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_0_; 
wire u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_1_; 
wire u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_2_; 
wire u2__abc_52138_new_n10000_; 
wire u2__abc_52138_new_n10001_; 
wire u2__abc_52138_new_n10002_; 
wire u2__abc_52138_new_n10003_; 
wire u2__abc_52138_new_n10005_; 
wire u2__abc_52138_new_n10006_; 
wire u2__abc_52138_new_n10007_; 
wire u2__abc_52138_new_n10008_; 
wire u2__abc_52138_new_n10009_; 
wire u2__abc_52138_new_n10010_; 
wire u2__abc_52138_new_n10011_; 
wire u2__abc_52138_new_n10012_; 
wire u2__abc_52138_new_n10013_; 
wire u2__abc_52138_new_n10014_; 
wire u2__abc_52138_new_n10015_; 
wire u2__abc_52138_new_n10016_; 
wire u2__abc_52138_new_n10018_; 
wire u2__abc_52138_new_n10019_; 
wire u2__abc_52138_new_n10020_; 
wire u2__abc_52138_new_n10021_; 
wire u2__abc_52138_new_n10022_; 
wire u2__abc_52138_new_n10023_; 
wire u2__abc_52138_new_n10024_; 
wire u2__abc_52138_new_n10026_; 
wire u2__abc_52138_new_n10027_; 
wire u2__abc_52138_new_n10028_; 
wire u2__abc_52138_new_n10029_; 
wire u2__abc_52138_new_n10030_; 
wire u2__abc_52138_new_n10031_; 
wire u2__abc_52138_new_n10032_; 
wire u2__abc_52138_new_n10033_; 
wire u2__abc_52138_new_n10034_; 
wire u2__abc_52138_new_n10036_; 
wire u2__abc_52138_new_n10037_; 
wire u2__abc_52138_new_n10038_; 
wire u2__abc_52138_new_n10039_; 
wire u2__abc_52138_new_n10040_; 
wire u2__abc_52138_new_n10041_; 
wire u2__abc_52138_new_n10042_; 
wire u2__abc_52138_new_n10043_; 
wire u2__abc_52138_new_n10045_; 
wire u2__abc_52138_new_n10046_; 
wire u2__abc_52138_new_n10047_; 
wire u2__abc_52138_new_n10048_; 
wire u2__abc_52138_new_n10049_; 
wire u2__abc_52138_new_n10050_; 
wire u2__abc_52138_new_n10051_; 
wire u2__abc_52138_new_n10052_; 
wire u2__abc_52138_new_n10053_; 
wire u2__abc_52138_new_n10054_; 
wire u2__abc_52138_new_n10055_; 
wire u2__abc_52138_new_n10056_; 
wire u2__abc_52138_new_n10057_; 
wire u2__abc_52138_new_n10059_; 
wire u2__abc_52138_new_n10060_; 
wire u2__abc_52138_new_n10061_; 
wire u2__abc_52138_new_n10062_; 
wire u2__abc_52138_new_n10063_; 
wire u2__abc_52138_new_n10064_; 
wire u2__abc_52138_new_n10065_; 
wire u2__abc_52138_new_n10066_; 
wire u2__abc_52138_new_n10067_; 
wire u2__abc_52138_new_n10069_; 
wire u2__abc_52138_new_n10070_; 
wire u2__abc_52138_new_n10071_; 
wire u2__abc_52138_new_n10072_; 
wire u2__abc_52138_new_n10073_; 
wire u2__abc_52138_new_n10074_; 
wire u2__abc_52138_new_n10075_; 
wire u2__abc_52138_new_n10076_; 
wire u2__abc_52138_new_n10077_; 
wire u2__abc_52138_new_n10079_; 
wire u2__abc_52138_new_n10080_; 
wire u2__abc_52138_new_n10081_; 
wire u2__abc_52138_new_n10082_; 
wire u2__abc_52138_new_n10083_; 
wire u2__abc_52138_new_n10084_; 
wire u2__abc_52138_new_n10085_; 
wire u2__abc_52138_new_n10086_; 
wire u2__abc_52138_new_n10088_; 
wire u2__abc_52138_new_n10089_; 
wire u2__abc_52138_new_n10090_; 
wire u2__abc_52138_new_n10091_; 
wire u2__abc_52138_new_n10092_; 
wire u2__abc_52138_new_n10093_; 
wire u2__abc_52138_new_n10094_; 
wire u2__abc_52138_new_n10095_; 
wire u2__abc_52138_new_n10096_; 
wire u2__abc_52138_new_n10097_; 
wire u2__abc_52138_new_n10098_; 
wire u2__abc_52138_new_n10099_; 
wire u2__abc_52138_new_n10101_; 
wire u2__abc_52138_new_n10102_; 
wire u2__abc_52138_new_n10103_; 
wire u2__abc_52138_new_n10104_; 
wire u2__abc_52138_new_n10105_; 
wire u2__abc_52138_new_n10106_; 
wire u2__abc_52138_new_n10107_; 
wire u2__abc_52138_new_n10108_; 
wire u2__abc_52138_new_n10110_; 
wire u2__abc_52138_new_n10111_; 
wire u2__abc_52138_new_n10112_; 
wire u2__abc_52138_new_n10113_; 
wire u2__abc_52138_new_n10114_; 
wire u2__abc_52138_new_n10115_; 
wire u2__abc_52138_new_n10116_; 
wire u2__abc_52138_new_n10117_; 
wire u2__abc_52138_new_n10118_; 
wire u2__abc_52138_new_n10119_; 
wire u2__abc_52138_new_n10121_; 
wire u2__abc_52138_new_n10122_; 
wire u2__abc_52138_new_n10123_; 
wire u2__abc_52138_new_n10124_; 
wire u2__abc_52138_new_n10125_; 
wire u2__abc_52138_new_n10126_; 
wire u2__abc_52138_new_n10127_; 
wire u2__abc_52138_new_n10128_; 
wire u2__abc_52138_new_n10130_; 
wire u2__abc_52138_new_n10131_; 
wire u2__abc_52138_new_n10132_; 
wire u2__abc_52138_new_n10133_; 
wire u2__abc_52138_new_n10134_; 
wire u2__abc_52138_new_n10135_; 
wire u2__abc_52138_new_n10136_; 
wire u2__abc_52138_new_n10137_; 
wire u2__abc_52138_new_n10138_; 
wire u2__abc_52138_new_n10139_; 
wire u2__abc_52138_new_n10140_; 
wire u2__abc_52138_new_n10141_; 
wire u2__abc_52138_new_n10142_; 
wire u2__abc_52138_new_n10143_; 
wire u2__abc_52138_new_n10144_; 
wire u2__abc_52138_new_n10146_; 
wire u2__abc_52138_new_n10147_; 
wire u2__abc_52138_new_n10148_; 
wire u2__abc_52138_new_n10149_; 
wire u2__abc_52138_new_n10150_; 
wire u2__abc_52138_new_n10151_; 
wire u2__abc_52138_new_n10152_; 
wire u2__abc_52138_new_n10154_; 
wire u2__abc_52138_new_n10155_; 
wire u2__abc_52138_new_n10156_; 
wire u2__abc_52138_new_n10157_; 
wire u2__abc_52138_new_n10158_; 
wire u2__abc_52138_new_n10159_; 
wire u2__abc_52138_new_n10160_; 
wire u2__abc_52138_new_n10161_; 
wire u2__abc_52138_new_n10162_; 
wire u2__abc_52138_new_n10164_; 
wire u2__abc_52138_new_n10165_; 
wire u2__abc_52138_new_n10166_; 
wire u2__abc_52138_new_n10167_; 
wire u2__abc_52138_new_n10168_; 
wire u2__abc_52138_new_n10169_; 
wire u2__abc_52138_new_n10170_; 
wire u2__abc_52138_new_n10171_; 
wire u2__abc_52138_new_n10173_; 
wire u2__abc_52138_new_n10174_; 
wire u2__abc_52138_new_n10175_; 
wire u2__abc_52138_new_n10176_; 
wire u2__abc_52138_new_n10177_; 
wire u2__abc_52138_new_n10178_; 
wire u2__abc_52138_new_n10179_; 
wire u2__abc_52138_new_n10180_; 
wire u2__abc_52138_new_n10181_; 
wire u2__abc_52138_new_n10182_; 
wire u2__abc_52138_new_n10183_; 
wire u2__abc_52138_new_n10184_; 
wire u2__abc_52138_new_n10185_; 
wire u2__abc_52138_new_n10186_; 
wire u2__abc_52138_new_n10187_; 
wire u2__abc_52138_new_n10189_; 
wire u2__abc_52138_new_n10190_; 
wire u2__abc_52138_new_n10191_; 
wire u2__abc_52138_new_n10192_; 
wire u2__abc_52138_new_n10193_; 
wire u2__abc_52138_new_n10194_; 
wire u2__abc_52138_new_n10195_; 
wire u2__abc_52138_new_n10197_; 
wire u2__abc_52138_new_n10198_; 
wire u2__abc_52138_new_n10199_; 
wire u2__abc_52138_new_n10200_; 
wire u2__abc_52138_new_n10201_; 
wire u2__abc_52138_new_n10202_; 
wire u2__abc_52138_new_n10203_; 
wire u2__abc_52138_new_n10204_; 
wire u2__abc_52138_new_n10205_; 
wire u2__abc_52138_new_n10207_; 
wire u2__abc_52138_new_n10208_; 
wire u2__abc_52138_new_n10209_; 
wire u2__abc_52138_new_n10210_; 
wire u2__abc_52138_new_n10211_; 
wire u2__abc_52138_new_n10212_; 
wire u2__abc_52138_new_n10213_; 
wire u2__abc_52138_new_n10214_; 
wire u2__abc_52138_new_n10216_; 
wire u2__abc_52138_new_n10217_; 
wire u2__abc_52138_new_n10218_; 
wire u2__abc_52138_new_n10219_; 
wire u2__abc_52138_new_n10220_; 
wire u2__abc_52138_new_n10221_; 
wire u2__abc_52138_new_n10222_; 
wire u2__abc_52138_new_n10223_; 
wire u2__abc_52138_new_n10224_; 
wire u2__abc_52138_new_n10225_; 
wire u2__abc_52138_new_n10226_; 
wire u2__abc_52138_new_n10227_; 
wire u2__abc_52138_new_n10228_; 
wire u2__abc_52138_new_n10229_; 
wire u2__abc_52138_new_n10230_; 
wire u2__abc_52138_new_n10232_; 
wire u2__abc_52138_new_n10233_; 
wire u2__abc_52138_new_n10234_; 
wire u2__abc_52138_new_n10235_; 
wire u2__abc_52138_new_n10236_; 
wire u2__abc_52138_new_n10237_; 
wire u2__abc_52138_new_n10238_; 
wire u2__abc_52138_new_n10239_; 
wire u2__abc_52138_new_n10241_; 
wire u2__abc_52138_new_n10242_; 
wire u2__abc_52138_new_n10243_; 
wire u2__abc_52138_new_n10244_; 
wire u2__abc_52138_new_n10245_; 
wire u2__abc_52138_new_n10246_; 
wire u2__abc_52138_new_n10247_; 
wire u2__abc_52138_new_n10248_; 
wire u2__abc_52138_new_n10249_; 
wire u2__abc_52138_new_n10250_; 
wire u2__abc_52138_new_n10252_; 
wire u2__abc_52138_new_n10253_; 
wire u2__abc_52138_new_n10254_; 
wire u2__abc_52138_new_n10255_; 
wire u2__abc_52138_new_n10256_; 
wire u2__abc_52138_new_n10257_; 
wire u2__abc_52138_new_n10258_; 
wire u2__abc_52138_new_n10259_; 
wire u2__abc_52138_new_n10261_; 
wire u2__abc_52138_new_n10262_; 
wire u2__abc_52138_new_n10263_; 
wire u2__abc_52138_new_n10264_; 
wire u2__abc_52138_new_n10265_; 
wire u2__abc_52138_new_n10266_; 
wire u2__abc_52138_new_n10267_; 
wire u2__abc_52138_new_n10268_; 
wire u2__abc_52138_new_n10269_; 
wire u2__abc_52138_new_n10270_; 
wire u2__abc_52138_new_n10271_; 
wire u2__abc_52138_new_n10272_; 
wire u2__abc_52138_new_n10273_; 
wire u2__abc_52138_new_n10274_; 
wire u2__abc_52138_new_n10276_; 
wire u2__abc_52138_new_n10277_; 
wire u2__abc_52138_new_n10278_; 
wire u2__abc_52138_new_n10279_; 
wire u2__abc_52138_new_n10280_; 
wire u2__abc_52138_new_n10281_; 
wire u2__abc_52138_new_n10282_; 
wire u2__abc_52138_new_n10284_; 
wire u2__abc_52138_new_n10285_; 
wire u2__abc_52138_new_n10286_; 
wire u2__abc_52138_new_n10287_; 
wire u2__abc_52138_new_n10288_; 
wire u2__abc_52138_new_n10289_; 
wire u2__abc_52138_new_n10290_; 
wire u2__abc_52138_new_n10291_; 
wire u2__abc_52138_new_n10292_; 
wire u2__abc_52138_new_n10293_; 
wire u2__abc_52138_new_n10294_; 
wire u2__abc_52138_new_n10296_; 
wire u2__abc_52138_new_n10297_; 
wire u2__abc_52138_new_n10298_; 
wire u2__abc_52138_new_n10299_; 
wire u2__abc_52138_new_n10300_; 
wire u2__abc_52138_new_n10301_; 
wire u2__abc_52138_new_n10302_; 
wire u2__abc_52138_new_n10304_; 
wire u2__abc_52138_new_n10305_; 
wire u2__abc_52138_new_n10306_; 
wire u2__abc_52138_new_n10307_; 
wire u2__abc_52138_new_n10308_; 
wire u2__abc_52138_new_n10309_; 
wire u2__abc_52138_new_n10310_; 
wire u2__abc_52138_new_n10311_; 
wire u2__abc_52138_new_n10312_; 
wire u2__abc_52138_new_n10313_; 
wire u2__abc_52138_new_n10314_; 
wire u2__abc_52138_new_n10315_; 
wire u2__abc_52138_new_n10316_; 
wire u2__abc_52138_new_n10317_; 
wire u2__abc_52138_new_n10318_; 
wire u2__abc_52138_new_n10319_; 
wire u2__abc_52138_new_n10320_; 
wire u2__abc_52138_new_n10322_; 
wire u2__abc_52138_new_n10323_; 
wire u2__abc_52138_new_n10324_; 
wire u2__abc_52138_new_n10325_; 
wire u2__abc_52138_new_n10326_; 
wire u2__abc_52138_new_n10327_; 
wire u2__abc_52138_new_n10328_; 
wire u2__abc_52138_new_n10330_; 
wire u2__abc_52138_new_n10331_; 
wire u2__abc_52138_new_n10332_; 
wire u2__abc_52138_new_n10333_; 
wire u2__abc_52138_new_n10334_; 
wire u2__abc_52138_new_n10335_; 
wire u2__abc_52138_new_n10336_; 
wire u2__abc_52138_new_n10337_; 
wire u2__abc_52138_new_n10338_; 
wire u2__abc_52138_new_n10340_; 
wire u2__abc_52138_new_n10341_; 
wire u2__abc_52138_new_n10342_; 
wire u2__abc_52138_new_n10343_; 
wire u2__abc_52138_new_n10344_; 
wire u2__abc_52138_new_n10345_; 
wire u2__abc_52138_new_n10346_; 
wire u2__abc_52138_new_n10347_; 
wire u2__abc_52138_new_n10349_; 
wire u2__abc_52138_new_n10350_; 
wire u2__abc_52138_new_n10351_; 
wire u2__abc_52138_new_n10352_; 
wire u2__abc_52138_new_n10353_; 
wire u2__abc_52138_new_n10354_; 
wire u2__abc_52138_new_n10355_; 
wire u2__abc_52138_new_n10356_; 
wire u2__abc_52138_new_n10357_; 
wire u2__abc_52138_new_n10358_; 
wire u2__abc_52138_new_n10359_; 
wire u2__abc_52138_new_n10360_; 
wire u2__abc_52138_new_n10361_; 
wire u2__abc_52138_new_n10362_; 
wire u2__abc_52138_new_n10364_; 
wire u2__abc_52138_new_n10365_; 
wire u2__abc_52138_new_n10366_; 
wire u2__abc_52138_new_n10367_; 
wire u2__abc_52138_new_n10368_; 
wire u2__abc_52138_new_n10369_; 
wire u2__abc_52138_new_n10370_; 
wire u2__abc_52138_new_n10371_; 
wire u2__abc_52138_new_n10373_; 
wire u2__abc_52138_new_n10374_; 
wire u2__abc_52138_new_n10375_; 
wire u2__abc_52138_new_n10376_; 
wire u2__abc_52138_new_n10377_; 
wire u2__abc_52138_new_n10378_; 
wire u2__abc_52138_new_n10379_; 
wire u2__abc_52138_new_n10380_; 
wire u2__abc_52138_new_n10381_; 
wire u2__abc_52138_new_n10382_; 
wire u2__abc_52138_new_n10384_; 
wire u2__abc_52138_new_n10385_; 
wire u2__abc_52138_new_n10386_; 
wire u2__abc_52138_new_n10387_; 
wire u2__abc_52138_new_n10388_; 
wire u2__abc_52138_new_n10389_; 
wire u2__abc_52138_new_n10390_; 
wire u2__abc_52138_new_n10391_; 
wire u2__abc_52138_new_n10393_; 
wire u2__abc_52138_new_n10394_; 
wire u2__abc_52138_new_n10395_; 
wire u2__abc_52138_new_n10396_; 
wire u2__abc_52138_new_n10397_; 
wire u2__abc_52138_new_n10398_; 
wire u2__abc_52138_new_n10399_; 
wire u2__abc_52138_new_n10400_; 
wire u2__abc_52138_new_n10401_; 
wire u2__abc_52138_new_n10402_; 
wire u2__abc_52138_new_n10403_; 
wire u2__abc_52138_new_n10404_; 
wire u2__abc_52138_new_n10405_; 
wire u2__abc_52138_new_n10406_; 
wire u2__abc_52138_new_n10408_; 
wire u2__abc_52138_new_n10409_; 
wire u2__abc_52138_new_n10410_; 
wire u2__abc_52138_new_n10411_; 
wire u2__abc_52138_new_n10412_; 
wire u2__abc_52138_new_n10413_; 
wire u2__abc_52138_new_n10414_; 
wire u2__abc_52138_new_n10415_; 
wire u2__abc_52138_new_n10417_; 
wire u2__abc_52138_new_n10418_; 
wire u2__abc_52138_new_n10419_; 
wire u2__abc_52138_new_n10420_; 
wire u2__abc_52138_new_n10421_; 
wire u2__abc_52138_new_n10422_; 
wire u2__abc_52138_new_n10423_; 
wire u2__abc_52138_new_n10424_; 
wire u2__abc_52138_new_n10425_; 
wire u2__abc_52138_new_n10426_; 
wire u2__abc_52138_new_n10427_; 
wire u2__abc_52138_new_n10429_; 
wire u2__abc_52138_new_n10430_; 
wire u2__abc_52138_new_n10431_; 
wire u2__abc_52138_new_n10432_; 
wire u2__abc_52138_new_n10433_; 
wire u2__abc_52138_new_n10434_; 
wire u2__abc_52138_new_n10435_; 
wire u2__abc_52138_new_n10436_; 
wire u2__abc_52138_new_n10438_; 
wire u2__abc_52138_new_n10439_; 
wire u2__abc_52138_new_n10440_; 
wire u2__abc_52138_new_n10441_; 
wire u2__abc_52138_new_n10442_; 
wire u2__abc_52138_new_n10443_; 
wire u2__abc_52138_new_n10444_; 
wire u2__abc_52138_new_n10445_; 
wire u2__abc_52138_new_n10446_; 
wire u2__abc_52138_new_n10447_; 
wire u2__abc_52138_new_n10448_; 
wire u2__abc_52138_new_n10449_; 
wire u2__abc_52138_new_n10450_; 
wire u2__abc_52138_new_n10452_; 
wire u2__abc_52138_new_n10453_; 
wire u2__abc_52138_new_n10454_; 
wire u2__abc_52138_new_n10455_; 
wire u2__abc_52138_new_n10456_; 
wire u2__abc_52138_new_n10457_; 
wire u2__abc_52138_new_n10458_; 
wire u2__abc_52138_new_n10460_; 
wire u2__abc_52138_new_n10461_; 
wire u2__abc_52138_new_n10462_; 
wire u2__abc_52138_new_n10463_; 
wire u2__abc_52138_new_n10464_; 
wire u2__abc_52138_new_n10465_; 
wire u2__abc_52138_new_n10466_; 
wire u2__abc_52138_new_n10467_; 
wire u2__abc_52138_new_n10468_; 
wire u2__abc_52138_new_n10470_; 
wire u2__abc_52138_new_n10471_; 
wire u2__abc_52138_new_n10472_; 
wire u2__abc_52138_new_n10473_; 
wire u2__abc_52138_new_n10474_; 
wire u2__abc_52138_new_n10475_; 
wire u2__abc_52138_new_n10476_; 
wire u2__abc_52138_new_n10477_; 
wire u2__abc_52138_new_n10479_; 
wire u2__abc_52138_new_n10480_; 
wire u2__abc_52138_new_n10481_; 
wire u2__abc_52138_new_n10482_; 
wire u2__abc_52138_new_n10483_; 
wire u2__abc_52138_new_n10484_; 
wire u2__abc_52138_new_n10485_; 
wire u2__abc_52138_new_n10486_; 
wire u2__abc_52138_new_n10487_; 
wire u2__abc_52138_new_n10488_; 
wire u2__abc_52138_new_n10489_; 
wire u2__abc_52138_new_n10490_; 
wire u2__abc_52138_new_n10491_; 
wire u2__abc_52138_new_n10492_; 
wire u2__abc_52138_new_n10493_; 
wire u2__abc_52138_new_n10494_; 
wire u2__abc_52138_new_n10496_; 
wire u2__abc_52138_new_n10497_; 
wire u2__abc_52138_new_n10498_; 
wire u2__abc_52138_new_n10499_; 
wire u2__abc_52138_new_n10500_; 
wire u2__abc_52138_new_n10501_; 
wire u2__abc_52138_new_n10502_; 
wire u2__abc_52138_new_n10504_; 
wire u2__abc_52138_new_n10505_; 
wire u2__abc_52138_new_n10506_; 
wire u2__abc_52138_new_n10507_; 
wire u2__abc_52138_new_n10508_; 
wire u2__abc_52138_new_n10509_; 
wire u2__abc_52138_new_n10510_; 
wire u2__abc_52138_new_n10511_; 
wire u2__abc_52138_new_n10512_; 
wire u2__abc_52138_new_n10514_; 
wire u2__abc_52138_new_n10515_; 
wire u2__abc_52138_new_n10516_; 
wire u2__abc_52138_new_n10517_; 
wire u2__abc_52138_new_n10518_; 
wire u2__abc_52138_new_n10519_; 
wire u2__abc_52138_new_n10520_; 
wire u2__abc_52138_new_n10521_; 
wire u2__abc_52138_new_n10523_; 
wire u2__abc_52138_new_n10524_; 
wire u2__abc_52138_new_n10525_; 
wire u2__abc_52138_new_n10526_; 
wire u2__abc_52138_new_n10527_; 
wire u2__abc_52138_new_n10528_; 
wire u2__abc_52138_new_n10529_; 
wire u2__abc_52138_new_n10530_; 
wire u2__abc_52138_new_n10531_; 
wire u2__abc_52138_new_n10532_; 
wire u2__abc_52138_new_n10533_; 
wire u2__abc_52138_new_n10535_; 
wire u2__abc_52138_new_n10536_; 
wire u2__abc_52138_new_n10537_; 
wire u2__abc_52138_new_n10538_; 
wire u2__abc_52138_new_n10539_; 
wire u2__abc_52138_new_n10540_; 
wire u2__abc_52138_new_n10541_; 
wire u2__abc_52138_new_n10542_; 
wire u2__abc_52138_new_n10544_; 
wire u2__abc_52138_new_n10545_; 
wire u2__abc_52138_new_n10546_; 
wire u2__abc_52138_new_n10547_; 
wire u2__abc_52138_new_n10548_; 
wire u2__abc_52138_new_n10549_; 
wire u2__abc_52138_new_n10550_; 
wire u2__abc_52138_new_n10551_; 
wire u2__abc_52138_new_n10553_; 
wire u2__abc_52138_new_n10554_; 
wire u2__abc_52138_new_n10555_; 
wire u2__abc_52138_new_n10556_; 
wire u2__abc_52138_new_n10557_; 
wire u2__abc_52138_new_n10558_; 
wire u2__abc_52138_new_n10559_; 
wire u2__abc_52138_new_n10560_; 
wire u2__abc_52138_new_n10562_; 
wire u2__abc_52138_new_n10563_; 
wire u2__abc_52138_new_n10564_; 
wire u2__abc_52138_new_n10565_; 
wire u2__abc_52138_new_n10566_; 
wire u2__abc_52138_new_n10567_; 
wire u2__abc_52138_new_n10568_; 
wire u2__abc_52138_new_n10569_; 
wire u2__abc_52138_new_n10570_; 
wire u2__abc_52138_new_n10571_; 
wire u2__abc_52138_new_n10572_; 
wire u2__abc_52138_new_n10573_; 
wire u2__abc_52138_new_n10575_; 
wire u2__abc_52138_new_n10576_; 
wire u2__abc_52138_new_n10577_; 
wire u2__abc_52138_new_n10578_; 
wire u2__abc_52138_new_n10579_; 
wire u2__abc_52138_new_n10580_; 
wire u2__abc_52138_new_n10581_; 
wire u2__abc_52138_new_n10582_; 
wire u2__abc_52138_new_n10584_; 
wire u2__abc_52138_new_n10585_; 
wire u2__abc_52138_new_n10586_; 
wire u2__abc_52138_new_n10587_; 
wire u2__abc_52138_new_n10588_; 
wire u2__abc_52138_new_n10589_; 
wire u2__abc_52138_new_n10590_; 
wire u2__abc_52138_new_n10591_; 
wire u2__abc_52138_new_n10592_; 
wire u2__abc_52138_new_n10593_; 
wire u2__abc_52138_new_n10594_; 
wire u2__abc_52138_new_n10595_; 
wire u2__abc_52138_new_n10597_; 
wire u2__abc_52138_new_n10598_; 
wire u2__abc_52138_new_n10599_; 
wire u2__abc_52138_new_n10600_; 
wire u2__abc_52138_new_n10601_; 
wire u2__abc_52138_new_n10602_; 
wire u2__abc_52138_new_n10603_; 
wire u2__abc_52138_new_n10604_; 
wire u2__abc_52138_new_n10606_; 
wire u2__abc_52138_new_n10607_; 
wire u2__abc_52138_new_n10608_; 
wire u2__abc_52138_new_n10609_; 
wire u2__abc_52138_new_n10610_; 
wire u2__abc_52138_new_n10611_; 
wire u2__abc_52138_new_n10612_; 
wire u2__abc_52138_new_n10613_; 
wire u2__abc_52138_new_n10614_; 
wire u2__abc_52138_new_n10615_; 
wire u2__abc_52138_new_n10617_; 
wire u2__abc_52138_new_n10618_; 
wire u2__abc_52138_new_n10619_; 
wire u2__abc_52138_new_n10620_; 
wire u2__abc_52138_new_n10621_; 
wire u2__abc_52138_new_n10622_; 
wire u2__abc_52138_new_n10623_; 
wire u2__abc_52138_new_n10625_; 
wire u2__abc_52138_new_n10626_; 
wire u2__abc_52138_new_n10627_; 
wire u2__abc_52138_new_n10628_; 
wire u2__abc_52138_new_n10629_; 
wire u2__abc_52138_new_n10630_; 
wire u2__abc_52138_new_n10631_; 
wire u2__abc_52138_new_n10632_; 
wire u2__abc_52138_new_n10633_; 
wire u2__abc_52138_new_n10634_; 
wire u2__abc_52138_new_n10636_; 
wire u2__abc_52138_new_n10637_; 
wire u2__abc_52138_new_n10638_; 
wire u2__abc_52138_new_n10639_; 
wire u2__abc_52138_new_n10640_; 
wire u2__abc_52138_new_n10641_; 
wire u2__abc_52138_new_n10642_; 
wire u2__abc_52138_new_n10643_; 
wire u2__abc_52138_new_n10645_; 
wire u2__abc_52138_new_n10646_; 
wire u2__abc_52138_new_n10647_; 
wire u2__abc_52138_new_n10648_; 
wire u2__abc_52138_new_n10649_; 
wire u2__abc_52138_new_n10650_; 
wire u2__abc_52138_new_n10651_; 
wire u2__abc_52138_new_n10652_; 
wire u2__abc_52138_new_n10653_; 
wire u2__abc_52138_new_n10654_; 
wire u2__abc_52138_new_n10655_; 
wire u2__abc_52138_new_n10656_; 
wire u2__abc_52138_new_n10657_; 
wire u2__abc_52138_new_n10658_; 
wire u2__abc_52138_new_n10659_; 
wire u2__abc_52138_new_n10660_; 
wire u2__abc_52138_new_n10661_; 
wire u2__abc_52138_new_n10662_; 
wire u2__abc_52138_new_n10663_; 
wire u2__abc_52138_new_n10664_; 
wire u2__abc_52138_new_n10665_; 
wire u2__abc_52138_new_n10666_; 
wire u2__abc_52138_new_n10667_; 
wire u2__abc_52138_new_n10668_; 
wire u2__abc_52138_new_n10670_; 
wire u2__abc_52138_new_n10671_; 
wire u2__abc_52138_new_n10672_; 
wire u2__abc_52138_new_n10673_; 
wire u2__abc_52138_new_n10674_; 
wire u2__abc_52138_new_n10675_; 
wire u2__abc_52138_new_n10676_; 
wire u2__abc_52138_new_n10678_; 
wire u2__abc_52138_new_n10679_; 
wire u2__abc_52138_new_n10680_; 
wire u2__abc_52138_new_n10681_; 
wire u2__abc_52138_new_n10682_; 
wire u2__abc_52138_new_n10683_; 
wire u2__abc_52138_new_n10684_; 
wire u2__abc_52138_new_n10685_; 
wire u2__abc_52138_new_n10686_; 
wire u2__abc_52138_new_n10687_; 
wire u2__abc_52138_new_n10689_; 
wire u2__abc_52138_new_n10690_; 
wire u2__abc_52138_new_n10691_; 
wire u2__abc_52138_new_n10692_; 
wire u2__abc_52138_new_n10693_; 
wire u2__abc_52138_new_n10694_; 
wire u2__abc_52138_new_n10695_; 
wire u2__abc_52138_new_n10696_; 
wire u2__abc_52138_new_n10698_; 
wire u2__abc_52138_new_n10699_; 
wire u2__abc_52138_new_n10700_; 
wire u2__abc_52138_new_n10701_; 
wire u2__abc_52138_new_n10702_; 
wire u2__abc_52138_new_n10703_; 
wire u2__abc_52138_new_n10704_; 
wire u2__abc_52138_new_n10705_; 
wire u2__abc_52138_new_n10706_; 
wire u2__abc_52138_new_n10707_; 
wire u2__abc_52138_new_n10708_; 
wire u2__abc_52138_new_n10709_; 
wire u2__abc_52138_new_n10710_; 
wire u2__abc_52138_new_n10711_; 
wire u2__abc_52138_new_n10713_; 
wire u2__abc_52138_new_n10714_; 
wire u2__abc_52138_new_n10715_; 
wire u2__abc_52138_new_n10716_; 
wire u2__abc_52138_new_n10717_; 
wire u2__abc_52138_new_n10718_; 
wire u2__abc_52138_new_n10719_; 
wire u2__abc_52138_new_n10721_; 
wire u2__abc_52138_new_n10722_; 
wire u2__abc_52138_new_n10723_; 
wire u2__abc_52138_new_n10724_; 
wire u2__abc_52138_new_n10725_; 
wire u2__abc_52138_new_n10726_; 
wire u2__abc_52138_new_n10727_; 
wire u2__abc_52138_new_n10728_; 
wire u2__abc_52138_new_n10729_; 
wire u2__abc_52138_new_n10730_; 
wire u2__abc_52138_new_n10731_; 
wire u2__abc_52138_new_n10732_; 
wire u2__abc_52138_new_n10734_; 
wire u2__abc_52138_new_n10735_; 
wire u2__abc_52138_new_n10736_; 
wire u2__abc_52138_new_n10737_; 
wire u2__abc_52138_new_n10738_; 
wire u2__abc_52138_new_n10739_; 
wire u2__abc_52138_new_n10740_; 
wire u2__abc_52138_new_n10741_; 
wire u2__abc_52138_new_n10743_; 
wire u2__abc_52138_new_n10744_; 
wire u2__abc_52138_new_n10745_; 
wire u2__abc_52138_new_n10746_; 
wire u2__abc_52138_new_n10747_; 
wire u2__abc_52138_new_n10748_; 
wire u2__abc_52138_new_n10749_; 
wire u2__abc_52138_new_n10750_; 
wire u2__abc_52138_new_n10751_; 
wire u2__abc_52138_new_n10752_; 
wire u2__abc_52138_new_n10753_; 
wire u2__abc_52138_new_n10754_; 
wire u2__abc_52138_new_n10755_; 
wire u2__abc_52138_new_n10756_; 
wire u2__abc_52138_new_n10758_; 
wire u2__abc_52138_new_n10759_; 
wire u2__abc_52138_new_n10760_; 
wire u2__abc_52138_new_n10761_; 
wire u2__abc_52138_new_n10762_; 
wire u2__abc_52138_new_n10763_; 
wire u2__abc_52138_new_n10764_; 
wire u2__abc_52138_new_n10765_; 
wire u2__abc_52138_new_n10766_; 
wire u2__abc_52138_new_n10767_; 
wire u2__abc_52138_new_n10769_; 
wire u2__abc_52138_new_n10770_; 
wire u2__abc_52138_new_n10771_; 
wire u2__abc_52138_new_n10772_; 
wire u2__abc_52138_new_n10773_; 
wire u2__abc_52138_new_n10774_; 
wire u2__abc_52138_new_n10775_; 
wire u2__abc_52138_new_n10777_; 
wire u2__abc_52138_new_n10778_; 
wire u2__abc_52138_new_n10779_; 
wire u2__abc_52138_new_n10780_; 
wire u2__abc_52138_new_n10781_; 
wire u2__abc_52138_new_n10782_; 
wire u2__abc_52138_new_n10783_; 
wire u2__abc_52138_new_n10784_; 
wire u2__abc_52138_new_n10786_; 
wire u2__abc_52138_new_n10787_; 
wire u2__abc_52138_new_n10788_; 
wire u2__abc_52138_new_n10789_; 
wire u2__abc_52138_new_n10790_; 
wire u2__abc_52138_new_n10791_; 
wire u2__abc_52138_new_n10792_; 
wire u2__abc_52138_new_n10793_; 
wire u2__abc_52138_new_n10794_; 
wire u2__abc_52138_new_n10795_; 
wire u2__abc_52138_new_n10796_; 
wire u2__abc_52138_new_n10797_; 
wire u2__abc_52138_new_n10798_; 
wire u2__abc_52138_new_n10799_; 
wire u2__abc_52138_new_n10800_; 
wire u2__abc_52138_new_n10802_; 
wire u2__abc_52138_new_n10803_; 
wire u2__abc_52138_new_n10804_; 
wire u2__abc_52138_new_n10805_; 
wire u2__abc_52138_new_n10806_; 
wire u2__abc_52138_new_n10807_; 
wire u2__abc_52138_new_n10808_; 
wire u2__abc_52138_new_n10810_; 
wire u2__abc_52138_new_n10811_; 
wire u2__abc_52138_new_n10812_; 
wire u2__abc_52138_new_n10813_; 
wire u2__abc_52138_new_n10814_; 
wire u2__abc_52138_new_n10815_; 
wire u2__abc_52138_new_n10816_; 
wire u2__abc_52138_new_n10817_; 
wire u2__abc_52138_new_n10818_; 
wire u2__abc_52138_new_n10820_; 
wire u2__abc_52138_new_n10821_; 
wire u2__abc_52138_new_n10822_; 
wire u2__abc_52138_new_n10823_; 
wire u2__abc_52138_new_n10824_; 
wire u2__abc_52138_new_n10825_; 
wire u2__abc_52138_new_n10826_; 
wire u2__abc_52138_new_n10827_; 
wire u2__abc_52138_new_n10829_; 
wire u2__abc_52138_new_n10830_; 
wire u2__abc_52138_new_n10831_; 
wire u2__abc_52138_new_n10832_; 
wire u2__abc_52138_new_n10833_; 
wire u2__abc_52138_new_n10834_; 
wire u2__abc_52138_new_n10835_; 
wire u2__abc_52138_new_n10836_; 
wire u2__abc_52138_new_n10837_; 
wire u2__abc_52138_new_n10838_; 
wire u2__abc_52138_new_n10839_; 
wire u2__abc_52138_new_n10840_; 
wire u2__abc_52138_new_n10841_; 
wire u2__abc_52138_new_n10843_; 
wire u2__abc_52138_new_n10844_; 
wire u2__abc_52138_new_n10845_; 
wire u2__abc_52138_new_n10846_; 
wire u2__abc_52138_new_n10847_; 
wire u2__abc_52138_new_n10848_; 
wire u2__abc_52138_new_n10849_; 
wire u2__abc_52138_new_n10850_; 
wire u2__abc_52138_new_n10852_; 
wire u2__abc_52138_new_n10853_; 
wire u2__abc_52138_new_n10854_; 
wire u2__abc_52138_new_n10855_; 
wire u2__abc_52138_new_n10856_; 
wire u2__abc_52138_new_n10857_; 
wire u2__abc_52138_new_n10858_; 
wire u2__abc_52138_new_n10859_; 
wire u2__abc_52138_new_n10860_; 
wire u2__abc_52138_new_n10862_; 
wire u2__abc_52138_new_n10863_; 
wire u2__abc_52138_new_n10864_; 
wire u2__abc_52138_new_n10865_; 
wire u2__abc_52138_new_n10866_; 
wire u2__abc_52138_new_n10867_; 
wire u2__abc_52138_new_n10868_; 
wire u2__abc_52138_new_n10869_; 
wire u2__abc_52138_new_n10871_; 
wire u2__abc_52138_new_n10872_; 
wire u2__abc_52138_new_n10873_; 
wire u2__abc_52138_new_n10874_; 
wire u2__abc_52138_new_n10875_; 
wire u2__abc_52138_new_n10876_; 
wire u2__abc_52138_new_n10877_; 
wire u2__abc_52138_new_n10878_; 
wire u2__abc_52138_new_n10879_; 
wire u2__abc_52138_new_n10880_; 
wire u2__abc_52138_new_n10881_; 
wire u2__abc_52138_new_n10882_; 
wire u2__abc_52138_new_n10883_; 
wire u2__abc_52138_new_n10884_; 
wire u2__abc_52138_new_n10886_; 
wire u2__abc_52138_new_n10887_; 
wire u2__abc_52138_new_n10888_; 
wire u2__abc_52138_new_n10889_; 
wire u2__abc_52138_new_n10890_; 
wire u2__abc_52138_new_n10891_; 
wire u2__abc_52138_new_n10892_; 
wire u2__abc_52138_new_n10894_; 
wire u2__abc_52138_new_n10895_; 
wire u2__abc_52138_new_n10896_; 
wire u2__abc_52138_new_n10897_; 
wire u2__abc_52138_new_n10898_; 
wire u2__abc_52138_new_n10899_; 
wire u2__abc_52138_new_n10900_; 
wire u2__abc_52138_new_n10901_; 
wire u2__abc_52138_new_n10902_; 
wire u2__abc_52138_new_n10903_; 
wire u2__abc_52138_new_n10905_; 
wire u2__abc_52138_new_n10906_; 
wire u2__abc_52138_new_n10907_; 
wire u2__abc_52138_new_n10908_; 
wire u2__abc_52138_new_n10909_; 
wire u2__abc_52138_new_n10910_; 
wire u2__abc_52138_new_n10911_; 
wire u2__abc_52138_new_n10912_; 
wire u2__abc_52138_new_n10914_; 
wire u2__abc_52138_new_n10915_; 
wire u2__abc_52138_new_n10916_; 
wire u2__abc_52138_new_n10917_; 
wire u2__abc_52138_new_n10918_; 
wire u2__abc_52138_new_n10919_; 
wire u2__abc_52138_new_n10920_; 
wire u2__abc_52138_new_n10921_; 
wire u2__abc_52138_new_n10922_; 
wire u2__abc_52138_new_n10923_; 
wire u2__abc_52138_new_n10924_; 
wire u2__abc_52138_new_n10925_; 
wire u2__abc_52138_new_n10926_; 
wire u2__abc_52138_new_n10927_; 
wire u2__abc_52138_new_n10928_; 
wire u2__abc_52138_new_n10930_; 
wire u2__abc_52138_new_n10931_; 
wire u2__abc_52138_new_n10932_; 
wire u2__abc_52138_new_n10933_; 
wire u2__abc_52138_new_n10934_; 
wire u2__abc_52138_new_n10935_; 
wire u2__abc_52138_new_n10936_; 
wire u2__abc_52138_new_n10938_; 
wire u2__abc_52138_new_n10939_; 
wire u2__abc_52138_new_n10940_; 
wire u2__abc_52138_new_n10941_; 
wire u2__abc_52138_new_n10942_; 
wire u2__abc_52138_new_n10943_; 
wire u2__abc_52138_new_n10944_; 
wire u2__abc_52138_new_n10945_; 
wire u2__abc_52138_new_n10946_; 
wire u2__abc_52138_new_n10947_; 
wire u2__abc_52138_new_n10949_; 
wire u2__abc_52138_new_n10950_; 
wire u2__abc_52138_new_n10951_; 
wire u2__abc_52138_new_n10952_; 
wire u2__abc_52138_new_n10953_; 
wire u2__abc_52138_new_n10954_; 
wire u2__abc_52138_new_n10955_; 
wire u2__abc_52138_new_n10956_; 
wire u2__abc_52138_new_n10958_; 
wire u2__abc_52138_new_n10959_; 
wire u2__abc_52138_new_n10960_; 
wire u2__abc_52138_new_n10961_; 
wire u2__abc_52138_new_n10962_; 
wire u2__abc_52138_new_n10963_; 
wire u2__abc_52138_new_n10964_; 
wire u2__abc_52138_new_n10965_; 
wire u2__abc_52138_new_n10966_; 
wire u2__abc_52138_new_n10967_; 
wire u2__abc_52138_new_n10968_; 
wire u2__abc_52138_new_n10969_; 
wire u2__abc_52138_new_n10970_; 
wire u2__abc_52138_new_n10971_; 
wire u2__abc_52138_new_n10973_; 
wire u2__abc_52138_new_n10974_; 
wire u2__abc_52138_new_n10975_; 
wire u2__abc_52138_new_n10976_; 
wire u2__abc_52138_new_n10977_; 
wire u2__abc_52138_new_n10978_; 
wire u2__abc_52138_new_n10979_; 
wire u2__abc_52138_new_n10980_; 
wire u2__abc_52138_new_n10982_; 
wire u2__abc_52138_new_n10983_; 
wire u2__abc_52138_new_n10984_; 
wire u2__abc_52138_new_n10985_; 
wire u2__abc_52138_new_n10986_; 
wire u2__abc_52138_new_n10987_; 
wire u2__abc_52138_new_n10988_; 
wire u2__abc_52138_new_n10989_; 
wire u2__abc_52138_new_n10990_; 
wire u2__abc_52138_new_n10992_; 
wire u2__abc_52138_new_n10993_; 
wire u2__abc_52138_new_n10994_; 
wire u2__abc_52138_new_n10995_; 
wire u2__abc_52138_new_n10996_; 
wire u2__abc_52138_new_n10997_; 
wire u2__abc_52138_new_n10998_; 
wire u2__abc_52138_new_n10999_; 
wire u2__abc_52138_new_n11001_; 
wire u2__abc_52138_new_n11002_; 
wire u2__abc_52138_new_n11003_; 
wire u2__abc_52138_new_n11004_; 
wire u2__abc_52138_new_n11005_; 
wire u2__abc_52138_new_n11006_; 
wire u2__abc_52138_new_n11007_; 
wire u2__abc_52138_new_n11008_; 
wire u2__abc_52138_new_n11009_; 
wire u2__abc_52138_new_n11010_; 
wire u2__abc_52138_new_n11011_; 
wire u2__abc_52138_new_n11012_; 
wire u2__abc_52138_new_n11013_; 
wire u2__abc_52138_new_n11014_; 
wire u2__abc_52138_new_n11015_; 
wire u2__abc_52138_new_n11016_; 
wire u2__abc_52138_new_n11017_; 
wire u2__abc_52138_new_n11018_; 
wire u2__abc_52138_new_n11020_; 
wire u2__abc_52138_new_n11021_; 
wire u2__abc_52138_new_n11022_; 
wire u2__abc_52138_new_n11023_; 
wire u2__abc_52138_new_n11024_; 
wire u2__abc_52138_new_n11025_; 
wire u2__abc_52138_new_n11026_; 
wire u2__abc_52138_new_n11028_; 
wire u2__abc_52138_new_n11029_; 
wire u2__abc_52138_new_n11030_; 
wire u2__abc_52138_new_n11031_; 
wire u2__abc_52138_new_n11032_; 
wire u2__abc_52138_new_n11033_; 
wire u2__abc_52138_new_n11034_; 
wire u2__abc_52138_new_n11035_; 
wire u2__abc_52138_new_n11036_; 
wire u2__abc_52138_new_n11037_; 
wire u2__abc_52138_new_n11038_; 
wire u2__abc_52138_new_n11040_; 
wire u2__abc_52138_new_n11041_; 
wire u2__abc_52138_new_n11042_; 
wire u2__abc_52138_new_n11043_; 
wire u2__abc_52138_new_n11044_; 
wire u2__abc_52138_new_n11045_; 
wire u2__abc_52138_new_n11046_; 
wire u2__abc_52138_new_n11047_; 
wire u2__abc_52138_new_n11049_; 
wire u2__abc_52138_new_n11050_; 
wire u2__abc_52138_new_n11051_; 
wire u2__abc_52138_new_n11052_; 
wire u2__abc_52138_new_n11053_; 
wire u2__abc_52138_new_n11054_; 
wire u2__abc_52138_new_n11055_; 
wire u2__abc_52138_new_n11056_; 
wire u2__abc_52138_new_n11057_; 
wire u2__abc_52138_new_n11058_; 
wire u2__abc_52138_new_n11059_; 
wire u2__abc_52138_new_n11060_; 
wire u2__abc_52138_new_n11061_; 
wire u2__abc_52138_new_n11062_; 
wire u2__abc_52138_new_n11064_; 
wire u2__abc_52138_new_n11065_; 
wire u2__abc_52138_new_n11066_; 
wire u2__abc_52138_new_n11067_; 
wire u2__abc_52138_new_n11068_; 
wire u2__abc_52138_new_n11069_; 
wire u2__abc_52138_new_n11070_; 
wire u2__abc_52138_new_n11071_; 
wire u2__abc_52138_new_n11073_; 
wire u2__abc_52138_new_n11074_; 
wire u2__abc_52138_new_n11075_; 
wire u2__abc_52138_new_n11076_; 
wire u2__abc_52138_new_n11077_; 
wire u2__abc_52138_new_n11078_; 
wire u2__abc_52138_new_n11079_; 
wire u2__abc_52138_new_n11080_; 
wire u2__abc_52138_new_n11081_; 
wire u2__abc_52138_new_n11082_; 
wire u2__abc_52138_new_n11084_; 
wire u2__abc_52138_new_n11085_; 
wire u2__abc_52138_new_n11086_; 
wire u2__abc_52138_new_n11087_; 
wire u2__abc_52138_new_n11088_; 
wire u2__abc_52138_new_n11089_; 
wire u2__abc_52138_new_n11090_; 
wire u2__abc_52138_new_n11091_; 
wire u2__abc_52138_new_n11093_; 
wire u2__abc_52138_new_n11094_; 
wire u2__abc_52138_new_n11095_; 
wire u2__abc_52138_new_n11096_; 
wire u2__abc_52138_new_n11097_; 
wire u2__abc_52138_new_n11098_; 
wire u2__abc_52138_new_n11099_; 
wire u2__abc_52138_new_n11100_; 
wire u2__abc_52138_new_n11101_; 
wire u2__abc_52138_new_n11102_; 
wire u2__abc_52138_new_n11103_; 
wire u2__abc_52138_new_n11104_; 
wire u2__abc_52138_new_n11105_; 
wire u2__abc_52138_new_n11107_; 
wire u2__abc_52138_new_n11108_; 
wire u2__abc_52138_new_n11109_; 
wire u2__abc_52138_new_n11110_; 
wire u2__abc_52138_new_n11111_; 
wire u2__abc_52138_new_n11112_; 
wire u2__abc_52138_new_n11113_; 
wire u2__abc_52138_new_n11114_; 
wire u2__abc_52138_new_n11116_; 
wire u2__abc_52138_new_n11117_; 
wire u2__abc_52138_new_n11118_; 
wire u2__abc_52138_new_n11119_; 
wire u2__abc_52138_new_n11120_; 
wire u2__abc_52138_new_n11121_; 
wire u2__abc_52138_new_n11122_; 
wire u2__abc_52138_new_n11123_; 
wire u2__abc_52138_new_n11124_; 
wire u2__abc_52138_new_n11125_; 
wire u2__abc_52138_new_n11127_; 
wire u2__abc_52138_new_n11128_; 
wire u2__abc_52138_new_n11129_; 
wire u2__abc_52138_new_n11130_; 
wire u2__abc_52138_new_n11131_; 
wire u2__abc_52138_new_n11132_; 
wire u2__abc_52138_new_n11133_; 
wire u2__abc_52138_new_n11134_; 
wire u2__abc_52138_new_n11136_; 
wire u2__abc_52138_new_n11137_; 
wire u2__abc_52138_new_n11138_; 
wire u2__abc_52138_new_n11139_; 
wire u2__abc_52138_new_n11140_; 
wire u2__abc_52138_new_n11141_; 
wire u2__abc_52138_new_n11142_; 
wire u2__abc_52138_new_n11143_; 
wire u2__abc_52138_new_n11144_; 
wire u2__abc_52138_new_n11145_; 
wire u2__abc_52138_new_n11146_; 
wire u2__abc_52138_new_n11147_; 
wire u2__abc_52138_new_n11149_; 
wire u2__abc_52138_new_n11150_; 
wire u2__abc_52138_new_n11151_; 
wire u2__abc_52138_new_n11152_; 
wire u2__abc_52138_new_n11153_; 
wire u2__abc_52138_new_n11154_; 
wire u2__abc_52138_new_n11155_; 
wire u2__abc_52138_new_n11157_; 
wire u2__abc_52138_new_n11158_; 
wire u2__abc_52138_new_n11159_; 
wire u2__abc_52138_new_n11160_; 
wire u2__abc_52138_new_n11161_; 
wire u2__abc_52138_new_n11162_; 
wire u2__abc_52138_new_n11163_; 
wire u2__abc_52138_new_n11164_; 
wire u2__abc_52138_new_n11165_; 
wire u2__abc_52138_new_n11166_; 
wire u2__abc_52138_new_n11167_; 
wire u2__abc_52138_new_n11169_; 
wire u2__abc_52138_new_n11170_; 
wire u2__abc_52138_new_n11171_; 
wire u2__abc_52138_new_n11172_; 
wire u2__abc_52138_new_n11173_; 
wire u2__abc_52138_new_n11174_; 
wire u2__abc_52138_new_n11175_; 
wire u2__abc_52138_new_n11176_; 
wire u2__abc_52138_new_n11178_; 
wire u2__abc_52138_new_n11179_; 
wire u2__abc_52138_new_n11180_; 
wire u2__abc_52138_new_n11181_; 
wire u2__abc_52138_new_n11182_; 
wire u2__abc_52138_new_n11183_; 
wire u2__abc_52138_new_n11184_; 
wire u2__abc_52138_new_n11185_; 
wire u2__abc_52138_new_n11186_; 
wire u2__abc_52138_new_n11187_; 
wire u2__abc_52138_new_n11188_; 
wire u2__abc_52138_new_n11189_; 
wire u2__abc_52138_new_n11190_; 
wire u2__abc_52138_new_n11192_; 
wire u2__abc_52138_new_n11193_; 
wire u2__abc_52138_new_n11194_; 
wire u2__abc_52138_new_n11195_; 
wire u2__abc_52138_new_n11196_; 
wire u2__abc_52138_new_n11197_; 
wire u2__abc_52138_new_n11198_; 
wire u2__abc_52138_new_n11199_; 
wire u2__abc_52138_new_n11200_; 
wire u2__abc_52138_new_n11202_; 
wire u2__abc_52138_new_n11203_; 
wire u2__abc_52138_new_n11204_; 
wire u2__abc_52138_new_n11205_; 
wire u2__abc_52138_new_n11206_; 
wire u2__abc_52138_new_n11207_; 
wire u2__abc_52138_new_n11208_; 
wire u2__abc_52138_new_n11209_; 
wire u2__abc_52138_new_n11210_; 
wire u2__abc_52138_new_n11211_; 
wire u2__abc_52138_new_n11212_; 
wire u2__abc_52138_new_n11214_; 
wire u2__abc_52138_new_n11215_; 
wire u2__abc_52138_new_n11216_; 
wire u2__abc_52138_new_n11217_; 
wire u2__abc_52138_new_n11218_; 
wire u2__abc_52138_new_n11219_; 
wire u2__abc_52138_new_n11220_; 
wire u2__abc_52138_new_n11222_; 
wire u2__abc_52138_new_n11223_; 
wire u2__abc_52138_new_n11224_; 
wire u2__abc_52138_new_n11225_; 
wire u2__abc_52138_new_n11226_; 
wire u2__abc_52138_new_n11227_; 
wire u2__abc_52138_new_n11228_; 
wire u2__abc_52138_new_n11229_; 
wire u2__abc_52138_new_n11230_; 
wire u2__abc_52138_new_n11231_; 
wire u2__abc_52138_new_n11233_; 
wire u2__abc_52138_new_n11234_; 
wire u2__abc_52138_new_n11235_; 
wire u2__abc_52138_new_n11236_; 
wire u2__abc_52138_new_n11237_; 
wire u2__abc_52138_new_n11238_; 
wire u2__abc_52138_new_n11239_; 
wire u2__abc_52138_new_n11240_; 
wire u2__abc_52138_new_n11241_; 
wire u2__abc_52138_new_n11242_; 
wire u2__abc_52138_new_n11244_; 
wire u2__abc_52138_new_n11245_; 
wire u2__abc_52138_new_n11246_; 
wire u2__abc_52138_new_n11247_; 
wire u2__abc_52138_new_n11248_; 
wire u2__abc_52138_new_n11249_; 
wire u2__abc_52138_new_n11250_; 
wire u2__abc_52138_new_n11251_; 
wire u2__abc_52138_new_n11252_; 
wire u2__abc_52138_new_n11254_; 
wire u2__abc_52138_new_n11255_; 
wire u2__abc_52138_new_n11256_; 
wire u2__abc_52138_new_n11257_; 
wire u2__abc_52138_new_n11258_; 
wire u2__abc_52138_new_n11259_; 
wire u2__abc_52138_new_n11260_; 
wire u2__abc_52138_new_n11262_; 
wire u2__abc_52138_new_n11263_; 
wire u2__abc_52138_new_n11264_; 
wire u2__abc_52138_new_n11265_; 
wire u2__abc_52138_new_n11266_; 
wire u2__abc_52138_new_n11267_; 
wire u2__abc_52138_new_n11268_; 
wire u2__abc_52138_new_n11269_; 
wire u2__abc_52138_new_n11270_; 
wire u2__abc_52138_new_n11271_; 
wire u2__abc_52138_new_n11272_; 
wire u2__abc_52138_new_n11273_; 
wire u2__abc_52138_new_n11274_; 
wire u2__abc_52138_new_n11276_; 
wire u2__abc_52138_new_n11277_; 
wire u2__abc_52138_new_n11278_; 
wire u2__abc_52138_new_n11279_; 
wire u2__abc_52138_new_n11280_; 
wire u2__abc_52138_new_n11281_; 
wire u2__abc_52138_new_n11282_; 
wire u2__abc_52138_new_n11283_; 
wire u2__abc_52138_new_n11285_; 
wire u2__abc_52138_new_n11286_; 
wire u2__abc_52138_new_n11287_; 
wire u2__abc_52138_new_n11288_; 
wire u2__abc_52138_new_n11289_; 
wire u2__abc_52138_new_n11290_; 
wire u2__abc_52138_new_n11291_; 
wire u2__abc_52138_new_n11292_; 
wire u2__abc_52138_new_n11293_; 
wire u2__abc_52138_new_n11294_; 
wire u2__abc_52138_new_n11295_; 
wire u2__abc_52138_new_n11296_; 
wire u2__abc_52138_new_n11297_; 
wire u2__abc_52138_new_n11299_; 
wire u2__abc_52138_new_n11300_; 
wire u2__abc_52138_new_n11301_; 
wire u2__abc_52138_new_n11302_; 
wire u2__abc_52138_new_n11303_; 
wire u2__abc_52138_new_n11304_; 
wire u2__abc_52138_new_n11305_; 
wire u2__abc_52138_new_n11306_; 
wire u2__abc_52138_new_n11308_; 
wire u2__abc_52138_new_n11309_; 
wire u2__abc_52138_new_n11310_; 
wire u2__abc_52138_new_n11311_; 
wire u2__abc_52138_new_n11312_; 
wire u2__abc_52138_new_n11313_; 
wire u2__abc_52138_new_n11314_; 
wire u2__abc_52138_new_n11315_; 
wire u2__abc_52138_new_n11316_; 
wire u2__abc_52138_new_n11317_; 
wire u2__abc_52138_new_n11318_; 
wire u2__abc_52138_new_n11319_; 
wire u2__abc_52138_new_n11320_; 
wire u2__abc_52138_new_n11322_; 
wire u2__abc_52138_new_n11323_; 
wire u2__abc_52138_new_n11324_; 
wire u2__abc_52138_new_n11325_; 
wire u2__abc_52138_new_n11326_; 
wire u2__abc_52138_new_n11327_; 
wire u2__abc_52138_new_n11328_; 
wire u2__abc_52138_new_n11330_; 
wire u2__abc_52138_new_n11331_; 
wire u2__abc_52138_new_n11332_; 
wire u2__abc_52138_new_n11333_; 
wire u2__abc_52138_new_n11334_; 
wire u2__abc_52138_new_n11335_; 
wire u2__abc_52138_new_n11336_; 
wire u2__abc_52138_new_n11337_; 
wire u2__abc_52138_new_n11338_; 
wire u2__abc_52138_new_n11339_; 
wire u2__abc_52138_new_n11340_; 
wire u2__abc_52138_new_n11342_; 
wire u2__abc_52138_new_n11343_; 
wire u2__abc_52138_new_n11344_; 
wire u2__abc_52138_new_n11345_; 
wire u2__abc_52138_new_n11346_; 
wire u2__abc_52138_new_n11347_; 
wire u2__abc_52138_new_n11348_; 
wire u2__abc_52138_new_n11349_; 
wire u2__abc_52138_new_n11351_; 
wire u2__abc_52138_new_n11352_; 
wire u2__abc_52138_new_n11353_; 
wire u2__abc_52138_new_n11354_; 
wire u2__abc_52138_new_n11355_; 
wire u2__abc_52138_new_n11356_; 
wire u2__abc_52138_new_n11357_; 
wire u2__abc_52138_new_n11358_; 
wire u2__abc_52138_new_n11359_; 
wire u2__abc_52138_new_n11360_; 
wire u2__abc_52138_new_n11361_; 
wire u2__abc_52138_new_n11362_; 
wire u2__abc_52138_new_n11363_; 
wire u2__abc_52138_new_n11364_; 
wire u2__abc_52138_new_n11365_; 
wire u2__abc_52138_new_n11366_; 
wire u2__abc_52138_new_n11368_; 
wire u2__abc_52138_new_n11369_; 
wire u2__abc_52138_new_n11370_; 
wire u2__abc_52138_new_n11371_; 
wire u2__abc_52138_new_n11372_; 
wire u2__abc_52138_new_n11373_; 
wire u2__abc_52138_new_n11374_; 
wire u2__abc_52138_new_n11375_; 
wire u2__abc_52138_new_n11377_; 
wire u2__abc_52138_new_n11378_; 
wire u2__abc_52138_new_n11379_; 
wire u2__abc_52138_new_n11380_; 
wire u2__abc_52138_new_n11382_; 
wire u2__abc_52138_new_n11383_; 
wire u2__abc_52138_new_n11384_; 
wire u2__abc_52138_new_n11386_; 
wire u2__abc_52138_new_n11387_; 
wire u2__abc_52138_new_n11388_; 
wire u2__abc_52138_new_n11389_; 
wire u2__abc_52138_new_n11391_; 
wire u2__abc_52138_new_n11392_; 
wire u2__abc_52138_new_n11393_; 
wire u2__abc_52138_new_n11394_; 
wire u2__abc_52138_new_n11395_; 
wire u2__abc_52138_new_n11396_; 
wire u2__abc_52138_new_n11398_; 
wire u2__abc_52138_new_n11399_; 
wire u2__abc_52138_new_n11401_; 
wire u2__abc_52138_new_n11402_; 
wire u2__abc_52138_new_n11403_; 
wire u2__abc_52138_new_n11405_; 
wire u2__abc_52138_new_n11406_; 
wire u2__abc_52138_new_n11407_; 
wire u2__abc_52138_new_n11409_; 
wire u2__abc_52138_new_n11410_; 
wire u2__abc_52138_new_n11412_; 
wire u2__abc_52138_new_n11413_; 
wire u2__abc_52138_new_n11415_; 
wire u2__abc_52138_new_n11417_; 
wire u2__abc_52138_new_n11418_; 
wire u2__abc_52138_new_n11420_; 
wire u2__abc_52138_new_n11421_; 
wire u2__abc_52138_new_n11423_; 
wire u2__abc_52138_new_n11424_; 
wire u2__abc_52138_new_n11426_; 
wire u2__abc_52138_new_n11427_; 
wire u2__abc_52138_new_n11429_; 
wire u2__abc_52138_new_n11430_; 
wire u2__abc_52138_new_n11432_; 
wire u2__abc_52138_new_n11433_; 
wire u2__abc_52138_new_n11435_; 
wire u2__abc_52138_new_n11436_; 
wire u2__abc_52138_new_n11438_; 
wire u2__abc_52138_new_n11439_; 
wire u2__abc_52138_new_n11441_; 
wire u2__abc_52138_new_n11442_; 
wire u2__abc_52138_new_n11444_; 
wire u2__abc_52138_new_n11445_; 
wire u2__abc_52138_new_n11447_; 
wire u2__abc_52138_new_n11448_; 
wire u2__abc_52138_new_n11450_; 
wire u2__abc_52138_new_n11451_; 
wire u2__abc_52138_new_n11453_; 
wire u2__abc_52138_new_n11454_; 
wire u2__abc_52138_new_n11456_; 
wire u2__abc_52138_new_n11457_; 
wire u2__abc_52138_new_n11459_; 
wire u2__abc_52138_new_n11460_; 
wire u2__abc_52138_new_n11462_; 
wire u2__abc_52138_new_n11463_; 
wire u2__abc_52138_new_n11465_; 
wire u2__abc_52138_new_n11466_; 
wire u2__abc_52138_new_n11468_; 
wire u2__abc_52138_new_n11469_; 
wire u2__abc_52138_new_n11471_; 
wire u2__abc_52138_new_n11472_; 
wire u2__abc_52138_new_n11474_; 
wire u2__abc_52138_new_n11475_; 
wire u2__abc_52138_new_n11477_; 
wire u2__abc_52138_new_n11478_; 
wire u2__abc_52138_new_n11480_; 
wire u2__abc_52138_new_n11481_; 
wire u2__abc_52138_new_n11483_; 
wire u2__abc_52138_new_n11484_; 
wire u2__abc_52138_new_n11486_; 
wire u2__abc_52138_new_n11487_; 
wire u2__abc_52138_new_n11489_; 
wire u2__abc_52138_new_n11490_; 
wire u2__abc_52138_new_n11492_; 
wire u2__abc_52138_new_n11493_; 
wire u2__abc_52138_new_n11495_; 
wire u2__abc_52138_new_n11496_; 
wire u2__abc_52138_new_n11498_; 
wire u2__abc_52138_new_n11499_; 
wire u2__abc_52138_new_n11501_; 
wire u2__abc_52138_new_n11502_; 
wire u2__abc_52138_new_n11504_; 
wire u2__abc_52138_new_n11505_; 
wire u2__abc_52138_new_n11507_; 
wire u2__abc_52138_new_n11508_; 
wire u2__abc_52138_new_n11509_; 
wire u2__abc_52138_new_n11510_; 
wire u2__abc_52138_new_n11512_; 
wire u2__abc_52138_new_n11513_; 
wire u2__abc_52138_new_n11514_; 
wire u2__abc_52138_new_n11515_; 
wire u2__abc_52138_new_n11516_; 
wire u2__abc_52138_new_n11518_; 
wire u2__abc_52138_new_n11519_; 
wire u2__abc_52138_new_n11521_; 
wire u2__abc_52138_new_n11522_; 
wire u2__abc_52138_new_n11524_; 
wire u2__abc_52138_new_n11525_; 
wire u2__abc_52138_new_n11526_; 
wire u2__abc_52138_new_n11527_; 
wire u2__abc_52138_new_n11528_; 
wire u2__abc_52138_new_n11530_; 
wire u2__abc_52138_new_n11531_; 
wire u2__abc_52138_new_n11533_; 
wire u2__abc_52138_new_n11534_; 
wire u2__abc_52138_new_n11536_; 
wire u2__abc_52138_new_n11537_; 
wire u2__abc_52138_new_n11539_; 
wire u2__abc_52138_new_n11540_; 
wire u2__abc_52138_new_n11542_; 
wire u2__abc_52138_new_n11543_; 
wire u2__abc_52138_new_n11545_; 
wire u2__abc_52138_new_n11546_; 
wire u2__abc_52138_new_n11548_; 
wire u2__abc_52138_new_n11549_; 
wire u2__abc_52138_new_n11551_; 
wire u2__abc_52138_new_n11552_; 
wire u2__abc_52138_new_n11554_; 
wire u2__abc_52138_new_n11555_; 
wire u2__abc_52138_new_n11557_; 
wire u2__abc_52138_new_n11558_; 
wire u2__abc_52138_new_n11560_; 
wire u2__abc_52138_new_n11561_; 
wire u2__abc_52138_new_n11563_; 
wire u2__abc_52138_new_n11564_; 
wire u2__abc_52138_new_n11565_; 
wire u2__abc_52138_new_n11566_; 
wire u2__abc_52138_new_n11567_; 
wire u2__abc_52138_new_n11569_; 
wire u2__abc_52138_new_n11570_; 
wire u2__abc_52138_new_n11572_; 
wire u2__abc_52138_new_n11573_; 
wire u2__abc_52138_new_n11575_; 
wire u2__abc_52138_new_n11576_; 
wire u2__abc_52138_new_n11578_; 
wire u2__abc_52138_new_n11579_; 
wire u2__abc_52138_new_n11581_; 
wire u2__abc_52138_new_n11582_; 
wire u2__abc_52138_new_n11584_; 
wire u2__abc_52138_new_n11585_; 
wire u2__abc_52138_new_n11587_; 
wire u2__abc_52138_new_n11588_; 
wire u2__abc_52138_new_n11590_; 
wire u2__abc_52138_new_n11591_; 
wire u2__abc_52138_new_n11593_; 
wire u2__abc_52138_new_n11594_; 
wire u2__abc_52138_new_n11596_; 
wire u2__abc_52138_new_n11597_; 
wire u2__abc_52138_new_n11599_; 
wire u2__abc_52138_new_n11600_; 
wire u2__abc_52138_new_n11602_; 
wire u2__abc_52138_new_n11603_; 
wire u2__abc_52138_new_n11605_; 
wire u2__abc_52138_new_n11606_; 
wire u2__abc_52138_new_n11608_; 
wire u2__abc_52138_new_n11609_; 
wire u2__abc_52138_new_n11611_; 
wire u2__abc_52138_new_n11612_; 
wire u2__abc_52138_new_n11614_; 
wire u2__abc_52138_new_n11615_; 
wire u2__abc_52138_new_n11617_; 
wire u2__abc_52138_new_n11618_; 
wire u2__abc_52138_new_n11620_; 
wire u2__abc_52138_new_n11621_; 
wire u2__abc_52138_new_n11623_; 
wire u2__abc_52138_new_n11624_; 
wire u2__abc_52138_new_n11625_; 
wire u2__abc_52138_new_n11626_; 
wire u2__abc_52138_new_n11627_; 
wire u2__abc_52138_new_n11629_; 
wire u2__abc_52138_new_n11630_; 
wire u2__abc_52138_new_n11632_; 
wire u2__abc_52138_new_n11633_; 
wire u2__abc_52138_new_n11635_; 
wire u2__abc_52138_new_n11636_; 
wire u2__abc_52138_new_n11638_; 
wire u2__abc_52138_new_n11639_; 
wire u2__abc_52138_new_n11641_; 
wire u2__abc_52138_new_n11642_; 
wire u2__abc_52138_new_n11644_; 
wire u2__abc_52138_new_n11645_; 
wire u2__abc_52138_new_n11647_; 
wire u2__abc_52138_new_n11648_; 
wire u2__abc_52138_new_n11650_; 
wire u2__abc_52138_new_n11651_; 
wire u2__abc_52138_new_n11653_; 
wire u2__abc_52138_new_n11654_; 
wire u2__abc_52138_new_n11655_; 
wire u2__abc_52138_new_n11656_; 
wire u2__abc_52138_new_n11657_; 
wire u2__abc_52138_new_n11659_; 
wire u2__abc_52138_new_n11660_; 
wire u2__abc_52138_new_n11662_; 
wire u2__abc_52138_new_n11663_; 
wire u2__abc_52138_new_n11665_; 
wire u2__abc_52138_new_n11666_; 
wire u2__abc_52138_new_n11668_; 
wire u2__abc_52138_new_n11669_; 
wire u2__abc_52138_new_n11671_; 
wire u2__abc_52138_new_n11672_; 
wire u2__abc_52138_new_n11674_; 
wire u2__abc_52138_new_n11675_; 
wire u2__abc_52138_new_n11677_; 
wire u2__abc_52138_new_n11678_; 
wire u2__abc_52138_new_n11680_; 
wire u2__abc_52138_new_n11681_; 
wire u2__abc_52138_new_n11683_; 
wire u2__abc_52138_new_n11684_; 
wire u2__abc_52138_new_n11686_; 
wire u2__abc_52138_new_n11687_; 
wire u2__abc_52138_new_n11689_; 
wire u2__abc_52138_new_n11690_; 
wire u2__abc_52138_new_n11692_; 
wire u2__abc_52138_new_n11693_; 
wire u2__abc_52138_new_n11695_; 
wire u2__abc_52138_new_n11696_; 
wire u2__abc_52138_new_n11698_; 
wire u2__abc_52138_new_n11699_; 
wire u2__abc_52138_new_n11701_; 
wire u2__abc_52138_new_n11702_; 
wire u2__abc_52138_new_n11704_; 
wire u2__abc_52138_new_n11705_; 
wire u2__abc_52138_new_n11707_; 
wire u2__abc_52138_new_n11708_; 
wire u2__abc_52138_new_n11710_; 
wire u2__abc_52138_new_n11711_; 
wire u2__abc_52138_new_n11713_; 
wire u2__abc_52138_new_n11714_; 
wire u2__abc_52138_new_n11716_; 
wire u2__abc_52138_new_n11717_; 
wire u2__abc_52138_new_n11718_; 
wire u2__abc_52138_new_n11719_; 
wire u2__abc_52138_new_n11721_; 
wire u2__abc_52138_new_n11722_; 
wire u2__abc_52138_new_n11724_; 
wire u2__abc_52138_new_n11725_; 
wire u2__abc_52138_new_n11726_; 
wire u2__abc_52138_new_n11728_; 
wire u2__abc_52138_new_n11729_; 
wire u2__abc_52138_new_n11730_; 
wire u2__abc_52138_new_n11731_; 
wire u2__abc_52138_new_n11732_; 
wire u2__abc_52138_new_n11734_; 
wire u2__abc_52138_new_n11735_; 
wire u2__abc_52138_new_n11737_; 
wire u2__abc_52138_new_n11738_; 
wire u2__abc_52138_new_n11740_; 
wire u2__abc_52138_new_n11741_; 
wire u2__abc_52138_new_n11743_; 
wire u2__abc_52138_new_n11744_; 
wire u2__abc_52138_new_n11746_; 
wire u2__abc_52138_new_n11747_; 
wire u2__abc_52138_new_n11749_; 
wire u2__abc_52138_new_n11750_; 
wire u2__abc_52138_new_n11752_; 
wire u2__abc_52138_new_n11753_; 
wire u2__abc_52138_new_n11755_; 
wire u2__abc_52138_new_n11756_; 
wire u2__abc_52138_new_n11758_; 
wire u2__abc_52138_new_n11759_; 
wire u2__abc_52138_new_n11761_; 
wire u2__abc_52138_new_n11762_; 
wire u2__abc_52138_new_n11764_; 
wire u2__abc_52138_new_n11765_; 
wire u2__abc_52138_new_n11767_; 
wire u2__abc_52138_new_n11768_; 
wire u2__abc_52138_new_n11770_; 
wire u2__abc_52138_new_n11771_; 
wire u2__abc_52138_new_n11773_; 
wire u2__abc_52138_new_n11774_; 
wire u2__abc_52138_new_n11776_; 
wire u2__abc_52138_new_n11777_; 
wire u2__abc_52138_new_n11779_; 
wire u2__abc_52138_new_n11780_; 
wire u2__abc_52138_new_n11782_; 
wire u2__abc_52138_new_n11783_; 
wire u2__abc_52138_new_n11784_; 
wire u2__abc_52138_new_n11785_; 
wire u2__abc_52138_new_n11786_; 
wire u2__abc_52138_new_n11788_; 
wire u2__abc_52138_new_n11789_; 
wire u2__abc_52138_new_n11791_; 
wire u2__abc_52138_new_n11792_; 
wire u2__abc_52138_new_n11794_; 
wire u2__abc_52138_new_n11795_; 
wire u2__abc_52138_new_n11797_; 
wire u2__abc_52138_new_n11798_; 
wire u2__abc_52138_new_n11800_; 
wire u2__abc_52138_new_n11801_; 
wire u2__abc_52138_new_n11803_; 
wire u2__abc_52138_new_n11804_; 
wire u2__abc_52138_new_n11806_; 
wire u2__abc_52138_new_n11807_; 
wire u2__abc_52138_new_n11809_; 
wire u2__abc_52138_new_n11810_; 
wire u2__abc_52138_new_n11812_; 
wire u2__abc_52138_new_n11813_; 
wire u2__abc_52138_new_n11815_; 
wire u2__abc_52138_new_n11816_; 
wire u2__abc_52138_new_n11818_; 
wire u2__abc_52138_new_n11819_; 
wire u2__abc_52138_new_n11821_; 
wire u2__abc_52138_new_n11822_; 
wire u2__abc_52138_new_n11824_; 
wire u2__abc_52138_new_n11825_; 
wire u2__abc_52138_new_n11827_; 
wire u2__abc_52138_new_n11828_; 
wire u2__abc_52138_new_n11830_; 
wire u2__abc_52138_new_n11831_; 
wire u2__abc_52138_new_n11832_; 
wire u2__abc_52138_new_n11833_; 
wire u2__abc_52138_new_n11834_; 
wire u2__abc_52138_new_n11836_; 
wire u2__abc_52138_new_n11837_; 
wire u2__abc_52138_new_n11839_; 
wire u2__abc_52138_new_n11840_; 
wire u2__abc_52138_new_n11841_; 
wire u2__abc_52138_new_n11843_; 
wire u2__abc_52138_new_n11844_; 
wire u2__abc_52138_new_n11846_; 
wire u2__abc_52138_new_n11847_; 
wire u2__abc_52138_new_n11849_; 
wire u2__abc_52138_new_n11850_; 
wire u2__abc_52138_new_n11852_; 
wire u2__abc_52138_new_n11853_; 
wire u2__abc_52138_new_n11855_; 
wire u2__abc_52138_new_n11856_; 
wire u2__abc_52138_new_n11858_; 
wire u2__abc_52138_new_n11859_; 
wire u2__abc_52138_new_n11861_; 
wire u2__abc_52138_new_n11862_; 
wire u2__abc_52138_new_n11864_; 
wire u2__abc_52138_new_n11865_; 
wire u2__abc_52138_new_n11867_; 
wire u2__abc_52138_new_n11868_; 
wire u2__abc_52138_new_n11870_; 
wire u2__abc_52138_new_n11871_; 
wire u2__abc_52138_new_n11873_; 
wire u2__abc_52138_new_n11874_; 
wire u2__abc_52138_new_n11876_; 
wire u2__abc_52138_new_n11877_; 
wire u2__abc_52138_new_n11879_; 
wire u2__abc_52138_new_n11880_; 
wire u2__abc_52138_new_n11882_; 
wire u2__abc_52138_new_n11883_; 
wire u2__abc_52138_new_n11885_; 
wire u2__abc_52138_new_n11886_; 
wire u2__abc_52138_new_n11888_; 
wire u2__abc_52138_new_n11889_; 
wire u2__abc_52138_new_n11891_; 
wire u2__abc_52138_new_n11892_; 
wire u2__abc_52138_new_n11894_; 
wire u2__abc_52138_new_n11895_; 
wire u2__abc_52138_new_n11897_; 
wire u2__abc_52138_new_n11898_; 
wire u2__abc_52138_new_n11900_; 
wire u2__abc_52138_new_n11901_; 
wire u2__abc_52138_new_n11903_; 
wire u2__abc_52138_new_n11904_; 
wire u2__abc_52138_new_n11906_; 
wire u2__abc_52138_new_n11907_; 
wire u2__abc_52138_new_n11909_; 
wire u2__abc_52138_new_n11910_; 
wire u2__abc_52138_new_n11912_; 
wire u2__abc_52138_new_n11913_; 
wire u2__abc_52138_new_n11915_; 
wire u2__abc_52138_new_n11916_; 
wire u2__abc_52138_new_n11918_; 
wire u2__abc_52138_new_n11919_; 
wire u2__abc_52138_new_n11921_; 
wire u2__abc_52138_new_n11922_; 
wire u2__abc_52138_new_n11924_; 
wire u2__abc_52138_new_n11925_; 
wire u2__abc_52138_new_n11927_; 
wire u2__abc_52138_new_n11928_; 
wire u2__abc_52138_new_n11930_; 
wire u2__abc_52138_new_n11931_; 
wire u2__abc_52138_new_n11932_; 
wire u2__abc_52138_new_n11933_; 
wire u2__abc_52138_new_n11934_; 
wire u2__abc_52138_new_n11936_; 
wire u2__abc_52138_new_n11937_; 
wire u2__abc_52138_new_n11939_; 
wire u2__abc_52138_new_n11940_; 
wire u2__abc_52138_new_n11942_; 
wire u2__abc_52138_new_n11943_; 
wire u2__abc_52138_new_n11945_; 
wire u2__abc_52138_new_n11946_; 
wire u2__abc_52138_new_n11948_; 
wire u2__abc_52138_new_n11949_; 
wire u2__abc_52138_new_n11951_; 
wire u2__abc_52138_new_n11952_; 
wire u2__abc_52138_new_n11954_; 
wire u2__abc_52138_new_n11955_; 
wire u2__abc_52138_new_n11957_; 
wire u2__abc_52138_new_n11958_; 
wire u2__abc_52138_new_n11960_; 
wire u2__abc_52138_new_n11961_; 
wire u2__abc_52138_new_n11963_; 
wire u2__abc_52138_new_n11964_; 
wire u2__abc_52138_new_n11966_; 
wire u2__abc_52138_new_n11967_; 
wire u2__abc_52138_new_n11968_; 
wire u2__abc_52138_new_n11970_; 
wire u2__abc_52138_new_n11971_; 
wire u2__abc_52138_new_n11973_; 
wire u2__abc_52138_new_n11974_; 
wire u2__abc_52138_new_n11976_; 
wire u2__abc_52138_new_n11977_; 
wire u2__abc_52138_new_n11979_; 
wire u2__abc_52138_new_n11980_; 
wire u2__abc_52138_new_n11982_; 
wire u2__abc_52138_new_n11983_; 
wire u2__abc_52138_new_n11985_; 
wire u2__abc_52138_new_n11986_; 
wire u2__abc_52138_new_n11988_; 
wire u2__abc_52138_new_n11989_; 
wire u2__abc_52138_new_n11991_; 
wire u2__abc_52138_new_n11992_; 
wire u2__abc_52138_new_n11994_; 
wire u2__abc_52138_new_n11995_; 
wire u2__abc_52138_new_n11997_; 
wire u2__abc_52138_new_n11998_; 
wire u2__abc_52138_new_n12000_; 
wire u2__abc_52138_new_n12001_; 
wire u2__abc_52138_new_n12003_; 
wire u2__abc_52138_new_n12004_; 
wire u2__abc_52138_new_n12006_; 
wire u2__abc_52138_new_n12007_; 
wire u2__abc_52138_new_n12009_; 
wire u2__abc_52138_new_n12010_; 
wire u2__abc_52138_new_n12012_; 
wire u2__abc_52138_new_n12013_; 
wire u2__abc_52138_new_n12015_; 
wire u2__abc_52138_new_n12016_; 
wire u2__abc_52138_new_n12018_; 
wire u2__abc_52138_new_n12019_; 
wire u2__abc_52138_new_n12021_; 
wire u2__abc_52138_new_n12022_; 
wire u2__abc_52138_new_n12024_; 
wire u2__abc_52138_new_n12025_; 
wire u2__abc_52138_new_n12027_; 
wire u2__abc_52138_new_n12028_; 
wire u2__abc_52138_new_n12030_; 
wire u2__abc_52138_new_n12031_; 
wire u2__abc_52138_new_n12032_; 
wire u2__abc_52138_new_n12033_; 
wire u2__abc_52138_new_n12034_; 
wire u2__abc_52138_new_n12036_; 
wire u2__abc_52138_new_n12037_; 
wire u2__abc_52138_new_n12039_; 
wire u2__abc_52138_new_n12040_; 
wire u2__abc_52138_new_n12042_; 
wire u2__abc_52138_new_n12043_; 
wire u2__abc_52138_new_n12045_; 
wire u2__abc_52138_new_n12046_; 
wire u2__abc_52138_new_n12048_; 
wire u2__abc_52138_new_n12049_; 
wire u2__abc_52138_new_n12051_; 
wire u2__abc_52138_new_n12052_; 
wire u2__abc_52138_new_n12054_; 
wire u2__abc_52138_new_n12055_; 
wire u2__abc_52138_new_n12057_; 
wire u2__abc_52138_new_n12058_; 
wire u2__abc_52138_new_n12060_; 
wire u2__abc_52138_new_n12061_; 
wire u2__abc_52138_new_n12062_; 
wire u2__abc_52138_new_n12063_; 
wire u2__abc_52138_new_n12064_; 
wire u2__abc_52138_new_n12066_; 
wire u2__abc_52138_new_n12067_; 
wire u2__abc_52138_new_n12069_; 
wire u2__abc_52138_new_n12070_; 
wire u2__abc_52138_new_n12071_; 
wire u2__abc_52138_new_n12073_; 
wire u2__abc_52138_new_n12074_; 
wire u2__abc_52138_new_n12076_; 
wire u2__abc_52138_new_n12077_; 
wire u2__abc_52138_new_n12079_; 
wire u2__abc_52138_new_n12080_; 
wire u2__abc_52138_new_n12082_; 
wire u2__abc_52138_new_n12083_; 
wire u2__abc_52138_new_n12085_; 
wire u2__abc_52138_new_n12086_; 
wire u2__abc_52138_new_n12088_; 
wire u2__abc_52138_new_n12089_; 
wire u2__abc_52138_new_n12091_; 
wire u2__abc_52138_new_n12092_; 
wire u2__abc_52138_new_n12094_; 
wire u2__abc_52138_new_n12095_; 
wire u2__abc_52138_new_n12097_; 
wire u2__abc_52138_new_n12098_; 
wire u2__abc_52138_new_n12100_; 
wire u2__abc_52138_new_n12101_; 
wire u2__abc_52138_new_n12103_; 
wire u2__abc_52138_new_n12104_; 
wire u2__abc_52138_new_n12106_; 
wire u2__abc_52138_new_n12107_; 
wire u2__abc_52138_new_n12109_; 
wire u2__abc_52138_new_n12110_; 
wire u2__abc_52138_new_n12112_; 
wire u2__abc_52138_new_n12113_; 
wire u2__abc_52138_new_n12115_; 
wire u2__abc_52138_new_n12116_; 
wire u2__abc_52138_new_n12118_; 
wire u2__abc_52138_new_n12119_; 
wire u2__abc_52138_new_n12121_; 
wire u2__abc_52138_new_n12122_; 
wire u2__abc_52138_new_n12124_; 
wire u2__abc_52138_new_n12125_; 
wire u2__abc_52138_new_n12127_; 
wire u2__abc_52138_new_n12128_; 
wire u2__abc_52138_new_n12130_; 
wire u2__abc_52138_new_n12131_; 
wire u2__abc_52138_new_n12133_; 
wire u2__abc_52138_new_n12134_; 
wire u2__abc_52138_new_n12135_; 
wire u2__abc_52138_new_n12136_; 
wire u2__abc_52138_new_n12137_; 
wire u2__abc_52138_new_n12139_; 
wire u2__abc_52138_new_n12140_; 
wire u2__abc_52138_new_n12141_; 
wire u2__abc_52138_new_n12142_; 
wire u2__abc_52138_new_n12143_; 
wire u2__abc_52138_new_n12145_; 
wire u2__abc_52138_new_n12146_; 
wire u2__abc_52138_new_n12148_; 
wire u2__abc_52138_new_n12149_; 
wire u2__abc_52138_new_n12151_; 
wire u2__abc_52138_new_n12152_; 
wire u2__abc_52138_new_n12154_; 
wire u2__abc_52138_new_n12155_; 
wire u2__abc_52138_new_n12157_; 
wire u2__abc_52138_new_n12158_; 
wire u2__abc_52138_new_n12160_; 
wire u2__abc_52138_new_n12161_; 
wire u2__abc_52138_new_n12162_; 
wire u2__abc_52138_new_n12164_; 
wire u2__abc_52138_new_n12165_; 
wire u2__abc_52138_new_n12167_; 
wire u2__abc_52138_new_n12168_; 
wire u2__abc_52138_new_n12170_; 
wire u2__abc_52138_new_n12171_; 
wire u2__abc_52138_new_n12173_; 
wire u2__abc_52138_new_n12174_; 
wire u2__abc_52138_new_n12176_; 
wire u2__abc_52138_new_n12177_; 
wire u2__abc_52138_new_n12179_; 
wire u2__abc_52138_new_n12180_; 
wire u2__abc_52138_new_n12182_; 
wire u2__abc_52138_new_n12183_; 
wire u2__abc_52138_new_n12185_; 
wire u2__abc_52138_new_n12186_; 
wire u2__abc_52138_new_n12188_; 
wire u2__abc_52138_new_n12189_; 
wire u2__abc_52138_new_n12191_; 
wire u2__abc_52138_new_n12192_; 
wire u2__abc_52138_new_n12194_; 
wire u2__abc_52138_new_n12195_; 
wire u2__abc_52138_new_n12197_; 
wire u2__abc_52138_new_n12198_; 
wire u2__abc_52138_new_n12200_; 
wire u2__abc_52138_new_n12201_; 
wire u2__abc_52138_new_n12203_; 
wire u2__abc_52138_new_n12204_; 
wire u2__abc_52138_new_n12206_; 
wire u2__abc_52138_new_n12207_; 
wire u2__abc_52138_new_n12209_; 
wire u2__abc_52138_new_n12210_; 
wire u2__abc_52138_new_n12212_; 
wire u2__abc_52138_new_n12213_; 
wire u2__abc_52138_new_n12215_; 
wire u2__abc_52138_new_n12216_; 
wire u2__abc_52138_new_n12218_; 
wire u2__abc_52138_new_n12219_; 
wire u2__abc_52138_new_n12221_; 
wire u2__abc_52138_new_n12222_; 
wire u2__abc_52138_new_n12224_; 
wire u2__abc_52138_new_n12225_; 
wire u2__abc_52138_new_n12227_; 
wire u2__abc_52138_new_n12228_; 
wire u2__abc_52138_new_n12229_; 
wire u2__abc_52138_new_n12231_; 
wire u2__abc_52138_new_n12232_; 
wire u2__abc_52138_new_n12234_; 
wire u2__abc_52138_new_n12235_; 
wire u2__abc_52138_new_n12237_; 
wire u2__abc_52138_new_n12238_; 
wire u2__abc_52138_new_n12240_; 
wire u2__abc_52138_new_n12241_; 
wire u2__abc_52138_new_n12243_; 
wire u2__abc_52138_new_n12244_; 
wire u2__abc_52138_new_n12246_; 
wire u2__abc_52138_new_n12247_; 
wire u2__abc_52138_new_n12249_; 
wire u2__abc_52138_new_n12250_; 
wire u2__abc_52138_new_n12252_; 
wire u2__abc_52138_new_n12253_; 
wire u2__abc_52138_new_n12255_; 
wire u2__abc_52138_new_n12256_; 
wire u2__abc_52138_new_n12258_; 
wire u2__abc_52138_new_n12259_; 
wire u2__abc_52138_new_n12261_; 
wire u2__abc_52138_new_n12262_; 
wire u2__abc_52138_new_n12264_; 
wire u2__abc_52138_new_n12265_; 
wire u2__abc_52138_new_n12267_; 
wire u2__abc_52138_new_n12268_; 
wire u2__abc_52138_new_n12270_; 
wire u2__abc_52138_new_n12271_; 
wire u2__abc_52138_new_n12273_; 
wire u2__abc_52138_new_n12274_; 
wire u2__abc_52138_new_n12276_; 
wire u2__abc_52138_new_n12277_; 
wire u2__abc_52138_new_n12279_; 
wire u2__abc_52138_new_n12280_; 
wire u2__abc_52138_new_n12282_; 
wire u2__abc_52138_new_n12283_; 
wire u2__abc_52138_new_n12285_; 
wire u2__abc_52138_new_n12286_; 
wire u2__abc_52138_new_n12288_; 
wire u2__abc_52138_new_n12289_; 
wire u2__abc_52138_new_n12291_; 
wire u2__abc_52138_new_n12292_; 
wire u2__abc_52138_new_n12294_; 
wire u2__abc_52138_new_n12295_; 
wire u2__abc_52138_new_n12297_; 
wire u2__abc_52138_new_n12298_; 
wire u2__abc_52138_new_n12300_; 
wire u2__abc_52138_new_n12301_; 
wire u2__abc_52138_new_n12303_; 
wire u2__abc_52138_new_n12304_; 
wire u2__abc_52138_new_n12306_; 
wire u2__abc_52138_new_n12307_; 
wire u2__abc_52138_new_n12309_; 
wire u2__abc_52138_new_n12310_; 
wire u2__abc_52138_new_n12312_; 
wire u2__abc_52138_new_n12313_; 
wire u2__abc_52138_new_n12315_; 
wire u2__abc_52138_new_n12316_; 
wire u2__abc_52138_new_n12318_; 
wire u2__abc_52138_new_n12319_; 
wire u2__abc_52138_new_n12321_; 
wire u2__abc_52138_new_n12322_; 
wire u2__abc_52138_new_n12324_; 
wire u2__abc_52138_new_n12325_; 
wire u2__abc_52138_new_n12327_; 
wire u2__abc_52138_new_n12328_; 
wire u2__abc_52138_new_n12330_; 
wire u2__abc_52138_new_n12331_; 
wire u2__abc_52138_new_n12333_; 
wire u2__abc_52138_new_n12334_; 
wire u2__abc_52138_new_n12336_; 
wire u2__abc_52138_new_n12337_; 
wire u2__abc_52138_new_n12339_; 
wire u2__abc_52138_new_n12340_; 
wire u2__abc_52138_new_n12342_; 
wire u2__abc_52138_new_n12343_; 
wire u2__abc_52138_new_n12345_; 
wire u2__abc_52138_new_n12346_; 
wire u2__abc_52138_new_n12348_; 
wire u2__abc_52138_new_n12349_; 
wire u2__abc_52138_new_n12351_; 
wire u2__abc_52138_new_n12352_; 
wire u2__abc_52138_new_n12354_; 
wire u2__abc_52138_new_n12355_; 
wire u2__abc_52138_new_n12357_; 
wire u2__abc_52138_new_n12358_; 
wire u2__abc_52138_new_n12360_; 
wire u2__abc_52138_new_n12361_; 
wire u2__abc_52138_new_n12363_; 
wire u2__abc_52138_new_n12364_; 
wire u2__abc_52138_new_n12366_; 
wire u2__abc_52138_new_n12367_; 
wire u2__abc_52138_new_n12369_; 
wire u2__abc_52138_new_n12370_; 
wire u2__abc_52138_new_n12372_; 
wire u2__abc_52138_new_n12373_; 
wire u2__abc_52138_new_n12375_; 
wire u2__abc_52138_new_n12376_; 
wire u2__abc_52138_new_n12378_; 
wire u2__abc_52138_new_n12379_; 
wire u2__abc_52138_new_n12381_; 
wire u2__abc_52138_new_n12382_; 
wire u2__abc_52138_new_n12384_; 
wire u2__abc_52138_new_n12385_; 
wire u2__abc_52138_new_n12387_; 
wire u2__abc_52138_new_n12388_; 
wire u2__abc_52138_new_n12390_; 
wire u2__abc_52138_new_n12391_; 
wire u2__abc_52138_new_n12393_; 
wire u2__abc_52138_new_n12394_; 
wire u2__abc_52138_new_n12396_; 
wire u2__abc_52138_new_n12397_; 
wire u2__abc_52138_new_n12399_; 
wire u2__abc_52138_new_n12400_; 
wire u2__abc_52138_new_n12402_; 
wire u2__abc_52138_new_n12403_; 
wire u2__abc_52138_new_n12405_; 
wire u2__abc_52138_new_n12406_; 
wire u2__abc_52138_new_n12408_; 
wire u2__abc_52138_new_n12409_; 
wire u2__abc_52138_new_n12411_; 
wire u2__abc_52138_new_n12412_; 
wire u2__abc_52138_new_n12414_; 
wire u2__abc_52138_new_n12415_; 
wire u2__abc_52138_new_n12417_; 
wire u2__abc_52138_new_n12418_; 
wire u2__abc_52138_new_n12420_; 
wire u2__abc_52138_new_n12421_; 
wire u2__abc_52138_new_n12423_; 
wire u2__abc_52138_new_n12424_; 
wire u2__abc_52138_new_n12426_; 
wire u2__abc_52138_new_n12427_; 
wire u2__abc_52138_new_n12429_; 
wire u2__abc_52138_new_n12430_; 
wire u2__abc_52138_new_n12432_; 
wire u2__abc_52138_new_n12433_; 
wire u2__abc_52138_new_n12435_; 
wire u2__abc_52138_new_n12436_; 
wire u2__abc_52138_new_n12438_; 
wire u2__abc_52138_new_n12439_; 
wire u2__abc_52138_new_n12441_; 
wire u2__abc_52138_new_n12442_; 
wire u2__abc_52138_new_n12444_; 
wire u2__abc_52138_new_n12445_; 
wire u2__abc_52138_new_n12447_; 
wire u2__abc_52138_new_n12448_; 
wire u2__abc_52138_new_n12450_; 
wire u2__abc_52138_new_n12451_; 
wire u2__abc_52138_new_n12453_; 
wire u2__abc_52138_new_n12454_; 
wire u2__abc_52138_new_n12456_; 
wire u2__abc_52138_new_n12457_; 
wire u2__abc_52138_new_n12459_; 
wire u2__abc_52138_new_n12460_; 
wire u2__abc_52138_new_n12462_; 
wire u2__abc_52138_new_n12463_; 
wire u2__abc_52138_new_n12465_; 
wire u2__abc_52138_new_n12466_; 
wire u2__abc_52138_new_n12468_; 
wire u2__abc_52138_new_n12469_; 
wire u2__abc_52138_new_n12471_; 
wire u2__abc_52138_new_n12472_; 
wire u2__abc_52138_new_n12474_; 
wire u2__abc_52138_new_n12475_; 
wire u2__abc_52138_new_n12477_; 
wire u2__abc_52138_new_n12478_; 
wire u2__abc_52138_new_n12480_; 
wire u2__abc_52138_new_n12481_; 
wire u2__abc_52138_new_n12483_; 
wire u2__abc_52138_new_n12484_; 
wire u2__abc_52138_new_n12486_; 
wire u2__abc_52138_new_n12487_; 
wire u2__abc_52138_new_n12489_; 
wire u2__abc_52138_new_n12490_; 
wire u2__abc_52138_new_n12492_; 
wire u2__abc_52138_new_n12493_; 
wire u2__abc_52138_new_n12495_; 
wire u2__abc_52138_new_n12496_; 
wire u2__abc_52138_new_n12498_; 
wire u2__abc_52138_new_n12499_; 
wire u2__abc_52138_new_n12501_; 
wire u2__abc_52138_new_n12502_; 
wire u2__abc_52138_new_n12504_; 
wire u2__abc_52138_new_n12505_; 
wire u2__abc_52138_new_n12507_; 
wire u2__abc_52138_new_n12508_; 
wire u2__abc_52138_new_n12510_; 
wire u2__abc_52138_new_n12511_; 
wire u2__abc_52138_new_n12513_; 
wire u2__abc_52138_new_n12514_; 
wire u2__abc_52138_new_n12516_; 
wire u2__abc_52138_new_n12517_; 
wire u2__abc_52138_new_n12519_; 
wire u2__abc_52138_new_n12520_; 
wire u2__abc_52138_new_n12522_; 
wire u2__abc_52138_new_n12523_; 
wire u2__abc_52138_new_n12525_; 
wire u2__abc_52138_new_n12526_; 
wire u2__abc_52138_new_n12528_; 
wire u2__abc_52138_new_n12529_; 
wire u2__abc_52138_new_n12531_; 
wire u2__abc_52138_new_n12532_; 
wire u2__abc_52138_new_n12534_; 
wire u2__abc_52138_new_n12535_; 
wire u2__abc_52138_new_n12537_; 
wire u2__abc_52138_new_n12538_; 
wire u2__abc_52138_new_n12540_; 
wire u2__abc_52138_new_n12541_; 
wire u2__abc_52138_new_n12543_; 
wire u2__abc_52138_new_n12544_; 
wire u2__abc_52138_new_n12546_; 
wire u2__abc_52138_new_n12547_; 
wire u2__abc_52138_new_n12549_; 
wire u2__abc_52138_new_n12550_; 
wire u2__abc_52138_new_n12552_; 
wire u2__abc_52138_new_n12553_; 
wire u2__abc_52138_new_n12555_; 
wire u2__abc_52138_new_n12556_; 
wire u2__abc_52138_new_n12558_; 
wire u2__abc_52138_new_n12559_; 
wire u2__abc_52138_new_n12561_; 
wire u2__abc_52138_new_n12562_; 
wire u2__abc_52138_new_n12564_; 
wire u2__abc_52138_new_n12565_; 
wire u2__abc_52138_new_n12567_; 
wire u2__abc_52138_new_n12568_; 
wire u2__abc_52138_new_n12570_; 
wire u2__abc_52138_new_n12571_; 
wire u2__abc_52138_new_n12573_; 
wire u2__abc_52138_new_n12574_; 
wire u2__abc_52138_new_n12576_; 
wire u2__abc_52138_new_n12577_; 
wire u2__abc_52138_new_n12579_; 
wire u2__abc_52138_new_n12580_; 
wire u2__abc_52138_new_n12582_; 
wire u2__abc_52138_new_n12583_; 
wire u2__abc_52138_new_n12585_; 
wire u2__abc_52138_new_n12586_; 
wire u2__abc_52138_new_n12588_; 
wire u2__abc_52138_new_n12589_; 
wire u2__abc_52138_new_n12591_; 
wire u2__abc_52138_new_n12592_; 
wire u2__abc_52138_new_n12594_; 
wire u2__abc_52138_new_n12595_; 
wire u2__abc_52138_new_n12597_; 
wire u2__abc_52138_new_n12598_; 
wire u2__abc_52138_new_n12600_; 
wire u2__abc_52138_new_n12601_; 
wire u2__abc_52138_new_n12603_; 
wire u2__abc_52138_new_n12604_; 
wire u2__abc_52138_new_n12606_; 
wire u2__abc_52138_new_n12607_; 
wire u2__abc_52138_new_n12609_; 
wire u2__abc_52138_new_n12610_; 
wire u2__abc_52138_new_n12612_; 
wire u2__abc_52138_new_n12613_; 
wire u2__abc_52138_new_n12615_; 
wire u2__abc_52138_new_n12616_; 
wire u2__abc_52138_new_n12618_; 
wire u2__abc_52138_new_n12619_; 
wire u2__abc_52138_new_n12621_; 
wire u2__abc_52138_new_n12622_; 
wire u2__abc_52138_new_n12624_; 
wire u2__abc_52138_new_n12625_; 
wire u2__abc_52138_new_n12627_; 
wire u2__abc_52138_new_n12628_; 
wire u2__abc_52138_new_n12630_; 
wire u2__abc_52138_new_n12631_; 
wire u2__abc_52138_new_n12633_; 
wire u2__abc_52138_new_n12634_; 
wire u2__abc_52138_new_n12636_; 
wire u2__abc_52138_new_n12637_; 
wire u2__abc_52138_new_n12639_; 
wire u2__abc_52138_new_n12640_; 
wire u2__abc_52138_new_n12642_; 
wire u2__abc_52138_new_n12643_; 
wire u2__abc_52138_new_n12645_; 
wire u2__abc_52138_new_n12646_; 
wire u2__abc_52138_new_n12648_; 
wire u2__abc_52138_new_n12649_; 
wire u2__abc_52138_new_n12651_; 
wire u2__abc_52138_new_n12652_; 
wire u2__abc_52138_new_n12654_; 
wire u2__abc_52138_new_n12655_; 
wire u2__abc_52138_new_n12657_; 
wire u2__abc_52138_new_n12658_; 
wire u2__abc_52138_new_n12660_; 
wire u2__abc_52138_new_n12661_; 
wire u2__abc_52138_new_n12663_; 
wire u2__abc_52138_new_n12664_; 
wire u2__abc_52138_new_n12666_; 
wire u2__abc_52138_new_n12667_; 
wire u2__abc_52138_new_n12669_; 
wire u2__abc_52138_new_n12670_; 
wire u2__abc_52138_new_n12672_; 
wire u2__abc_52138_new_n12673_; 
wire u2__abc_52138_new_n12675_; 
wire u2__abc_52138_new_n12676_; 
wire u2__abc_52138_new_n12678_; 
wire u2__abc_52138_new_n12679_; 
wire u2__abc_52138_new_n12681_; 
wire u2__abc_52138_new_n12682_; 
wire u2__abc_52138_new_n12684_; 
wire u2__abc_52138_new_n12685_; 
wire u2__abc_52138_new_n12687_; 
wire u2__abc_52138_new_n12688_; 
wire u2__abc_52138_new_n12690_; 
wire u2__abc_52138_new_n12691_; 
wire u2__abc_52138_new_n12693_; 
wire u2__abc_52138_new_n12694_; 
wire u2__abc_52138_new_n12696_; 
wire u2__abc_52138_new_n12697_; 
wire u2__abc_52138_new_n12699_; 
wire u2__abc_52138_new_n12700_; 
wire u2__abc_52138_new_n12702_; 
wire u2__abc_52138_new_n12703_; 
wire u2__abc_52138_new_n12705_; 
wire u2__abc_52138_new_n12706_; 
wire u2__abc_52138_new_n12708_; 
wire u2__abc_52138_new_n12709_; 
wire u2__abc_52138_new_n12711_; 
wire u2__abc_52138_new_n12712_; 
wire u2__abc_52138_new_n12714_; 
wire u2__abc_52138_new_n12715_; 
wire u2__abc_52138_new_n12717_; 
wire u2__abc_52138_new_n12718_; 
wire u2__abc_52138_new_n12720_; 
wire u2__abc_52138_new_n12721_; 
wire u2__abc_52138_new_n12723_; 
wire u2__abc_52138_new_n12724_; 
wire u2__abc_52138_new_n12726_; 
wire u2__abc_52138_new_n12727_; 
wire u2__abc_52138_new_n12729_; 
wire u2__abc_52138_new_n12730_; 
wire u2__abc_52138_new_n12732_; 
wire u2__abc_52138_new_n12733_; 
wire u2__abc_52138_new_n12735_; 
wire u2__abc_52138_new_n12736_; 
wire u2__abc_52138_new_n12738_; 
wire u2__abc_52138_new_n12739_; 
wire u2__abc_52138_new_n12741_; 
wire u2__abc_52138_new_n12742_; 
wire u2__abc_52138_new_n12744_; 
wire u2__abc_52138_new_n12745_; 
wire u2__abc_52138_new_n12747_; 
wire u2__abc_52138_new_n12748_; 
wire u2__abc_52138_new_n12750_; 
wire u2__abc_52138_new_n12751_; 
wire u2__abc_52138_new_n12753_; 
wire u2__abc_52138_new_n12754_; 
wire u2__abc_52138_new_n12756_; 
wire u2__abc_52138_new_n12757_; 
wire u2__abc_52138_new_n12759_; 
wire u2__abc_52138_new_n12760_; 
wire u2__abc_52138_new_n12762_; 
wire u2__abc_52138_new_n12763_; 
wire u2__abc_52138_new_n12765_; 
wire u2__abc_52138_new_n12766_; 
wire u2__abc_52138_new_n12768_; 
wire u2__abc_52138_new_n12769_; 
wire u2__abc_52138_new_n12771_; 
wire u2__abc_52138_new_n12772_; 
wire u2__abc_52138_new_n12774_; 
wire u2__abc_52138_new_n12775_; 
wire u2__abc_52138_new_n12777_; 
wire u2__abc_52138_new_n12778_; 
wire u2__abc_52138_new_n12780_; 
wire u2__abc_52138_new_n12781_; 
wire u2__abc_52138_new_n12783_; 
wire u2__abc_52138_new_n12784_; 
wire u2__abc_52138_new_n12786_; 
wire u2__abc_52138_new_n12787_; 
wire u2__abc_52138_new_n12789_; 
wire u2__abc_52138_new_n12790_; 
wire u2__abc_52138_new_n12792_; 
wire u2__abc_52138_new_n12793_; 
wire u2__abc_52138_new_n12795_; 
wire u2__abc_52138_new_n12796_; 
wire u2__abc_52138_new_n12798_; 
wire u2__abc_52138_new_n12799_; 
wire u2__abc_52138_new_n12801_; 
wire u2__abc_52138_new_n12802_; 
wire u2__abc_52138_new_n12804_; 
wire u2__abc_52138_new_n12805_; 
wire u2__abc_52138_new_n12807_; 
wire u2__abc_52138_new_n12808_; 
wire u2__abc_52138_new_n12810_; 
wire u2__abc_52138_new_n12811_; 
wire u2__abc_52138_new_n12813_; 
wire u2__abc_52138_new_n12814_; 
wire u2__abc_52138_new_n12816_; 
wire u2__abc_52138_new_n12818_; 
wire u2__abc_52138_new_n12819_; 
wire u2__abc_52138_new_n12820_; 
wire u2__abc_52138_new_n12821_; 
wire u2__abc_52138_new_n12822_; 
wire u2__abc_52138_new_n12823_; 
wire u2__abc_52138_new_n12824_; 
wire u2__abc_52138_new_n12825_; 
wire u2__abc_52138_new_n12826_; 
wire u2__abc_52138_new_n12827_; 
wire u2__abc_52138_new_n12828_; 
wire u2__abc_52138_new_n12829_; 
wire u2__abc_52138_new_n12830_; 
wire u2__abc_52138_new_n12831_; 
wire u2__abc_52138_new_n12832_; 
wire u2__abc_52138_new_n12833_; 
wire u2__abc_52138_new_n12834_; 
wire u2__abc_52138_new_n12835_; 
wire u2__abc_52138_new_n12836_; 
wire u2__abc_52138_new_n12837_; 
wire u2__abc_52138_new_n12838_; 
wire u2__abc_52138_new_n12839_; 
wire u2__abc_52138_new_n12840_; 
wire u2__abc_52138_new_n12841_; 
wire u2__abc_52138_new_n12842_; 
wire u2__abc_52138_new_n12843_; 
wire u2__abc_52138_new_n12844_; 
wire u2__abc_52138_new_n12845_; 
wire u2__abc_52138_new_n12846_; 
wire u2__abc_52138_new_n12847_; 
wire u2__abc_52138_new_n12848_; 
wire u2__abc_52138_new_n12849_; 
wire u2__abc_52138_new_n12850_; 
wire u2__abc_52138_new_n12851_; 
wire u2__abc_52138_new_n12852_; 
wire u2__abc_52138_new_n12853_; 
wire u2__abc_52138_new_n12854_; 
wire u2__abc_52138_new_n12855_; 
wire u2__abc_52138_new_n12856_; 
wire u2__abc_52138_new_n12857_; 
wire u2__abc_52138_new_n12858_; 
wire u2__abc_52138_new_n12859_; 
wire u2__abc_52138_new_n12860_; 
wire u2__abc_52138_new_n12861_; 
wire u2__abc_52138_new_n12862_; 
wire u2__abc_52138_new_n12863_; 
wire u2__abc_52138_new_n12864_; 
wire u2__abc_52138_new_n12865_; 
wire u2__abc_52138_new_n12866_; 
wire u2__abc_52138_new_n12867_; 
wire u2__abc_52138_new_n12868_; 
wire u2__abc_52138_new_n12869_; 
wire u2__abc_52138_new_n12870_; 
wire u2__abc_52138_new_n12871_; 
wire u2__abc_52138_new_n12872_; 
wire u2__abc_52138_new_n12873_; 
wire u2__abc_52138_new_n12874_; 
wire u2__abc_52138_new_n12875_; 
wire u2__abc_52138_new_n12876_; 
wire u2__abc_52138_new_n12877_; 
wire u2__abc_52138_new_n12878_; 
wire u2__abc_52138_new_n12879_; 
wire u2__abc_52138_new_n12880_; 
wire u2__abc_52138_new_n12881_; 
wire u2__abc_52138_new_n12882_; 
wire u2__abc_52138_new_n12883_; 
wire u2__abc_52138_new_n12884_; 
wire u2__abc_52138_new_n12885_; 
wire u2__abc_52138_new_n12886_; 
wire u2__abc_52138_new_n12887_; 
wire u2__abc_52138_new_n12888_; 
wire u2__abc_52138_new_n12889_; 
wire u2__abc_52138_new_n12890_; 
wire u2__abc_52138_new_n12891_; 
wire u2__abc_52138_new_n12892_; 
wire u2__abc_52138_new_n12893_; 
wire u2__abc_52138_new_n12894_; 
wire u2__abc_52138_new_n12895_; 
wire u2__abc_52138_new_n12896_; 
wire u2__abc_52138_new_n12897_; 
wire u2__abc_52138_new_n12898_; 
wire u2__abc_52138_new_n12899_; 
wire u2__abc_52138_new_n12900_; 
wire u2__abc_52138_new_n12901_; 
wire u2__abc_52138_new_n12902_; 
wire u2__abc_52138_new_n12903_; 
wire u2__abc_52138_new_n12904_; 
wire u2__abc_52138_new_n12905_; 
wire u2__abc_52138_new_n12906_; 
wire u2__abc_52138_new_n12907_; 
wire u2__abc_52138_new_n12908_; 
wire u2__abc_52138_new_n12909_; 
wire u2__abc_52138_new_n12910_; 
wire u2__abc_52138_new_n12911_; 
wire u2__abc_52138_new_n12912_; 
wire u2__abc_52138_new_n12913_; 
wire u2__abc_52138_new_n12914_; 
wire u2__abc_52138_new_n12915_; 
wire u2__abc_52138_new_n12916_; 
wire u2__abc_52138_new_n12917_; 
wire u2__abc_52138_new_n12918_; 
wire u2__abc_52138_new_n12919_; 
wire u2__abc_52138_new_n12920_; 
wire u2__abc_52138_new_n12921_; 
wire u2__abc_52138_new_n12922_; 
wire u2__abc_52138_new_n12923_; 
wire u2__abc_52138_new_n12924_; 
wire u2__abc_52138_new_n12925_; 
wire u2__abc_52138_new_n12926_; 
wire u2__abc_52138_new_n12927_; 
wire u2__abc_52138_new_n12928_; 
wire u2__abc_52138_new_n12929_; 
wire u2__abc_52138_new_n12930_; 
wire u2__abc_52138_new_n12931_; 
wire u2__abc_52138_new_n12932_; 
wire u2__abc_52138_new_n12933_; 
wire u2__abc_52138_new_n12934_; 
wire u2__abc_52138_new_n12935_; 
wire u2__abc_52138_new_n12936_; 
wire u2__abc_52138_new_n12937_; 
wire u2__abc_52138_new_n12938_; 
wire u2__abc_52138_new_n12939_; 
wire u2__abc_52138_new_n12940_; 
wire u2__abc_52138_new_n12941_; 
wire u2__abc_52138_new_n12942_; 
wire u2__abc_52138_new_n12943_; 
wire u2__abc_52138_new_n12944_; 
wire u2__abc_52138_new_n12945_; 
wire u2__abc_52138_new_n12946_; 
wire u2__abc_52138_new_n12947_; 
wire u2__abc_52138_new_n12948_; 
wire u2__abc_52138_new_n12949_; 
wire u2__abc_52138_new_n12950_; 
wire u2__abc_52138_new_n12951_; 
wire u2__abc_52138_new_n12952_; 
wire u2__abc_52138_new_n12953_; 
wire u2__abc_52138_new_n12954_; 
wire u2__abc_52138_new_n12955_; 
wire u2__abc_52138_new_n12956_; 
wire u2__abc_52138_new_n12957_; 
wire u2__abc_52138_new_n12958_; 
wire u2__abc_52138_new_n12959_; 
wire u2__abc_52138_new_n12960_; 
wire u2__abc_52138_new_n12961_; 
wire u2__abc_52138_new_n12962_; 
wire u2__abc_52138_new_n12963_; 
wire u2__abc_52138_new_n12964_; 
wire u2__abc_52138_new_n12965_; 
wire u2__abc_52138_new_n12966_; 
wire u2__abc_52138_new_n12967_; 
wire u2__abc_52138_new_n12968_; 
wire u2__abc_52138_new_n12969_; 
wire u2__abc_52138_new_n12970_; 
wire u2__abc_52138_new_n12971_; 
wire u2__abc_52138_new_n12972_; 
wire u2__abc_52138_new_n12973_; 
wire u2__abc_52138_new_n12974_; 
wire u2__abc_52138_new_n12975_; 
wire u2__abc_52138_new_n12976_; 
wire u2__abc_52138_new_n12977_; 
wire u2__abc_52138_new_n12978_; 
wire u2__abc_52138_new_n12979_; 
wire u2__abc_52138_new_n12980_; 
wire u2__abc_52138_new_n12981_; 
wire u2__abc_52138_new_n12982_; 
wire u2__abc_52138_new_n12983_; 
wire u2__abc_52138_new_n12984_; 
wire u2__abc_52138_new_n12985_; 
wire u2__abc_52138_new_n12986_; 
wire u2__abc_52138_new_n12987_; 
wire u2__abc_52138_new_n12988_; 
wire u2__abc_52138_new_n12989_; 
wire u2__abc_52138_new_n12990_; 
wire u2__abc_52138_new_n12991_; 
wire u2__abc_52138_new_n12992_; 
wire u2__abc_52138_new_n12993_; 
wire u2__abc_52138_new_n12994_; 
wire u2__abc_52138_new_n12995_; 
wire u2__abc_52138_new_n12996_; 
wire u2__abc_52138_new_n12997_; 
wire u2__abc_52138_new_n12998_; 
wire u2__abc_52138_new_n12999_; 
wire u2__abc_52138_new_n13000_; 
wire u2__abc_52138_new_n13001_; 
wire u2__abc_52138_new_n13002_; 
wire u2__abc_52138_new_n13003_; 
wire u2__abc_52138_new_n13004_; 
wire u2__abc_52138_new_n13005_; 
wire u2__abc_52138_new_n13006_; 
wire u2__abc_52138_new_n13007_; 
wire u2__abc_52138_new_n13008_; 
wire u2__abc_52138_new_n13009_; 
wire u2__abc_52138_new_n13010_; 
wire u2__abc_52138_new_n13011_; 
wire u2__abc_52138_new_n13012_; 
wire u2__abc_52138_new_n13013_; 
wire u2__abc_52138_new_n13014_; 
wire u2__abc_52138_new_n13015_; 
wire u2__abc_52138_new_n13016_; 
wire u2__abc_52138_new_n13017_; 
wire u2__abc_52138_new_n13018_; 
wire u2__abc_52138_new_n13019_; 
wire u2__abc_52138_new_n13020_; 
wire u2__abc_52138_new_n13021_; 
wire u2__abc_52138_new_n13022_; 
wire u2__abc_52138_new_n13023_; 
wire u2__abc_52138_new_n13024_; 
wire u2__abc_52138_new_n13025_; 
wire u2__abc_52138_new_n13026_; 
wire u2__abc_52138_new_n13027_; 
wire u2__abc_52138_new_n13028_; 
wire u2__abc_52138_new_n13029_; 
wire u2__abc_52138_new_n13030_; 
wire u2__abc_52138_new_n13031_; 
wire u2__abc_52138_new_n13032_; 
wire u2__abc_52138_new_n13033_; 
wire u2__abc_52138_new_n13034_; 
wire u2__abc_52138_new_n13035_; 
wire u2__abc_52138_new_n13036_; 
wire u2__abc_52138_new_n13037_; 
wire u2__abc_52138_new_n13038_; 
wire u2__abc_52138_new_n13039_; 
wire u2__abc_52138_new_n13040_; 
wire u2__abc_52138_new_n13041_; 
wire u2__abc_52138_new_n13042_; 
wire u2__abc_52138_new_n13043_; 
wire u2__abc_52138_new_n13044_; 
wire u2__abc_52138_new_n13045_; 
wire u2__abc_52138_new_n13046_; 
wire u2__abc_52138_new_n13047_; 
wire u2__abc_52138_new_n13048_; 
wire u2__abc_52138_new_n13050_; 
wire u2__abc_52138_new_n13051_; 
wire u2__abc_52138_new_n13052_; 
wire u2__abc_52138_new_n13053_; 
wire u2__abc_52138_new_n13054_; 
wire u2__abc_52138_new_n13055_; 
wire u2__abc_52138_new_n13057_; 
wire u2__abc_52138_new_n13058_; 
wire u2__abc_52138_new_n13059_; 
wire u2__abc_52138_new_n13060_; 
wire u2__abc_52138_new_n13061_; 
wire u2__abc_52138_new_n13062_; 
wire u2__abc_52138_new_n13063_; 
wire u2__abc_52138_new_n13065_; 
wire u2__abc_52138_new_n13066_; 
wire u2__abc_52138_new_n13067_; 
wire u2__abc_52138_new_n13068_; 
wire u2__abc_52138_new_n13069_; 
wire u2__abc_52138_new_n13070_; 
wire u2__abc_52138_new_n13071_; 
wire u2__abc_52138_new_n13073_; 
wire u2__abc_52138_new_n13074_; 
wire u2__abc_52138_new_n13075_; 
wire u2__abc_52138_new_n13076_; 
wire u2__abc_52138_new_n13077_; 
wire u2__abc_52138_new_n13078_; 
wire u2__abc_52138_new_n13079_; 
wire u2__abc_52138_new_n13081_; 
wire u2__abc_52138_new_n13082_; 
wire u2__abc_52138_new_n13083_; 
wire u2__abc_52138_new_n13084_; 
wire u2__abc_52138_new_n13085_; 
wire u2__abc_52138_new_n13086_; 
wire u2__abc_52138_new_n13088_; 
wire u2__abc_52138_new_n13089_; 
wire u2__abc_52138_new_n13090_; 
wire u2__abc_52138_new_n13091_; 
wire u2__abc_52138_new_n13092_; 
wire u2__abc_52138_new_n13093_; 
wire u2__abc_52138_new_n13094_; 
wire u2__abc_52138_new_n13096_; 
wire u2__abc_52138_new_n13097_; 
wire u2__abc_52138_new_n13098_; 
wire u2__abc_52138_new_n13099_; 
wire u2__abc_52138_new_n13100_; 
wire u2__abc_52138_new_n13101_; 
wire u2__abc_52138_new_n13102_; 
wire u2__abc_52138_new_n13104_; 
wire u2__abc_52138_new_n13105_; 
wire u2__abc_52138_new_n13106_; 
wire u2__abc_52138_new_n13107_; 
wire u2__abc_52138_new_n13108_; 
wire u2__abc_52138_new_n13109_; 
wire u2__abc_52138_new_n13110_; 
wire u2__abc_52138_new_n13112_; 
wire u2__abc_52138_new_n13113_; 
wire u2__abc_52138_new_n13114_; 
wire u2__abc_52138_new_n13115_; 
wire u2__abc_52138_new_n13116_; 
wire u2__abc_52138_new_n13117_; 
wire u2__abc_52138_new_n13119_; 
wire u2__abc_52138_new_n13120_; 
wire u2__abc_52138_new_n13121_; 
wire u2__abc_52138_new_n13122_; 
wire u2__abc_52138_new_n13123_; 
wire u2__abc_52138_new_n13124_; 
wire u2__abc_52138_new_n13125_; 
wire u2__abc_52138_new_n13127_; 
wire u2__abc_52138_new_n13128_; 
wire u2__abc_52138_new_n13129_; 
wire u2__abc_52138_new_n13130_; 
wire u2__abc_52138_new_n13131_; 
wire u2__abc_52138_new_n13132_; 
wire u2__abc_52138_new_n13133_; 
wire u2__abc_52138_new_n13135_; 
wire u2__abc_52138_new_n13136_; 
wire u2__abc_52138_new_n13137_; 
wire u2__abc_52138_new_n13138_; 
wire u2__abc_52138_new_n13139_; 
wire u2__abc_52138_new_n13140_; 
wire u2__abc_52138_new_n13141_; 
wire u2__abc_52138_new_n13143_; 
wire u2__abc_52138_new_n13144_; 
wire u2__abc_52138_new_n13145_; 
wire u2__abc_52138_new_n13146_; 
wire u2__abc_52138_new_n13147_; 
wire u2__abc_52138_new_n13148_; 
wire u2__abc_52138_new_n13150_; 
wire u2__abc_52138_new_n13151_; 
wire u2__abc_52138_new_n13152_; 
wire u2__abc_52138_new_n13153_; 
wire u2__abc_52138_new_n13154_; 
wire u2__abc_52138_new_n13155_; 
wire u2__abc_52138_new_n13156_; 
wire u2__abc_52138_new_n13158_; 
wire u2__abc_52138_new_n13159_; 
wire u2__abc_52138_new_n13160_; 
wire u2__abc_52138_new_n13161_; 
wire u2__abc_52138_new_n13162_; 
wire u2__abc_52138_new_n13163_; 
wire u2__abc_52138_new_n13164_; 
wire u2__abc_52138_new_n13166_; 
wire u2__abc_52138_new_n13167_; 
wire u2__abc_52138_new_n13168_; 
wire u2__abc_52138_new_n13169_; 
wire u2__abc_52138_new_n13170_; 
wire u2__abc_52138_new_n13171_; 
wire u2__abc_52138_new_n13172_; 
wire u2__abc_52138_new_n13174_; 
wire u2__abc_52138_new_n13175_; 
wire u2__abc_52138_new_n13176_; 
wire u2__abc_52138_new_n13177_; 
wire u2__abc_52138_new_n13178_; 
wire u2__abc_52138_new_n13179_; 
wire u2__abc_52138_new_n13181_; 
wire u2__abc_52138_new_n13182_; 
wire u2__abc_52138_new_n13183_; 
wire u2__abc_52138_new_n13184_; 
wire u2__abc_52138_new_n13185_; 
wire u2__abc_52138_new_n13186_; 
wire u2__abc_52138_new_n13187_; 
wire u2__abc_52138_new_n13189_; 
wire u2__abc_52138_new_n13190_; 
wire u2__abc_52138_new_n13191_; 
wire u2__abc_52138_new_n13192_; 
wire u2__abc_52138_new_n13193_; 
wire u2__abc_52138_new_n13194_; 
wire u2__abc_52138_new_n13195_; 
wire u2__abc_52138_new_n13197_; 
wire u2__abc_52138_new_n13198_; 
wire u2__abc_52138_new_n13199_; 
wire u2__abc_52138_new_n13200_; 
wire u2__abc_52138_new_n13201_; 
wire u2__abc_52138_new_n13202_; 
wire u2__abc_52138_new_n13203_; 
wire u2__abc_52138_new_n13205_; 
wire u2__abc_52138_new_n13206_; 
wire u2__abc_52138_new_n13207_; 
wire u2__abc_52138_new_n13208_; 
wire u2__abc_52138_new_n13209_; 
wire u2__abc_52138_new_n13210_; 
wire u2__abc_52138_new_n13212_; 
wire u2__abc_52138_new_n13213_; 
wire u2__abc_52138_new_n13214_; 
wire u2__abc_52138_new_n13215_; 
wire u2__abc_52138_new_n13216_; 
wire u2__abc_52138_new_n13217_; 
wire u2__abc_52138_new_n13218_; 
wire u2__abc_52138_new_n13220_; 
wire u2__abc_52138_new_n13221_; 
wire u2__abc_52138_new_n13222_; 
wire u2__abc_52138_new_n13223_; 
wire u2__abc_52138_new_n13224_; 
wire u2__abc_52138_new_n13225_; 
wire u2__abc_52138_new_n13226_; 
wire u2__abc_52138_new_n13228_; 
wire u2__abc_52138_new_n13229_; 
wire u2__abc_52138_new_n13230_; 
wire u2__abc_52138_new_n13231_; 
wire u2__abc_52138_new_n13232_; 
wire u2__abc_52138_new_n13233_; 
wire u2__abc_52138_new_n13234_; 
wire u2__abc_52138_new_n13236_; 
wire u2__abc_52138_new_n13237_; 
wire u2__abc_52138_new_n13238_; 
wire u2__abc_52138_new_n13239_; 
wire u2__abc_52138_new_n13240_; 
wire u2__abc_52138_new_n13241_; 
wire u2__abc_52138_new_n13243_; 
wire u2__abc_52138_new_n13244_; 
wire u2__abc_52138_new_n13245_; 
wire u2__abc_52138_new_n13246_; 
wire u2__abc_52138_new_n13247_; 
wire u2__abc_52138_new_n13248_; 
wire u2__abc_52138_new_n13249_; 
wire u2__abc_52138_new_n13251_; 
wire u2__abc_52138_new_n13252_; 
wire u2__abc_52138_new_n13253_; 
wire u2__abc_52138_new_n13254_; 
wire u2__abc_52138_new_n13255_; 
wire u2__abc_52138_new_n13256_; 
wire u2__abc_52138_new_n13257_; 
wire u2__abc_52138_new_n13259_; 
wire u2__abc_52138_new_n13260_; 
wire u2__abc_52138_new_n13261_; 
wire u2__abc_52138_new_n13262_; 
wire u2__abc_52138_new_n13263_; 
wire u2__abc_52138_new_n13264_; 
wire u2__abc_52138_new_n13265_; 
wire u2__abc_52138_new_n13267_; 
wire u2__abc_52138_new_n13268_; 
wire u2__abc_52138_new_n13269_; 
wire u2__abc_52138_new_n13270_; 
wire u2__abc_52138_new_n13271_; 
wire u2__abc_52138_new_n13272_; 
wire u2__abc_52138_new_n13274_; 
wire u2__abc_52138_new_n13275_; 
wire u2__abc_52138_new_n13276_; 
wire u2__abc_52138_new_n13277_; 
wire u2__abc_52138_new_n13278_; 
wire u2__abc_52138_new_n13279_; 
wire u2__abc_52138_new_n13280_; 
wire u2__abc_52138_new_n13282_; 
wire u2__abc_52138_new_n13283_; 
wire u2__abc_52138_new_n13284_; 
wire u2__abc_52138_new_n13285_; 
wire u2__abc_52138_new_n13286_; 
wire u2__abc_52138_new_n13287_; 
wire u2__abc_52138_new_n13288_; 
wire u2__abc_52138_new_n13290_; 
wire u2__abc_52138_new_n13291_; 
wire u2__abc_52138_new_n13292_; 
wire u2__abc_52138_new_n13293_; 
wire u2__abc_52138_new_n13294_; 
wire u2__abc_52138_new_n13295_; 
wire u2__abc_52138_new_n13296_; 
wire u2__abc_52138_new_n13298_; 
wire u2__abc_52138_new_n13299_; 
wire u2__abc_52138_new_n13300_; 
wire u2__abc_52138_new_n13301_; 
wire u2__abc_52138_new_n13302_; 
wire u2__abc_52138_new_n13303_; 
wire u2__abc_52138_new_n13305_; 
wire u2__abc_52138_new_n13306_; 
wire u2__abc_52138_new_n13307_; 
wire u2__abc_52138_new_n13308_; 
wire u2__abc_52138_new_n13309_; 
wire u2__abc_52138_new_n13310_; 
wire u2__abc_52138_new_n13311_; 
wire u2__abc_52138_new_n13312_; 
wire u2__abc_52138_new_n13314_; 
wire u2__abc_52138_new_n13315_; 
wire u2__abc_52138_new_n13316_; 
wire u2__abc_52138_new_n13317_; 
wire u2__abc_52138_new_n13318_; 
wire u2__abc_52138_new_n13319_; 
wire u2__abc_52138_new_n13320_; 
wire u2__abc_52138_new_n13322_; 
wire u2__abc_52138_new_n13323_; 
wire u2__abc_52138_new_n13324_; 
wire u2__abc_52138_new_n13325_; 
wire u2__abc_52138_new_n13326_; 
wire u2__abc_52138_new_n13327_; 
wire u2__abc_52138_new_n13328_; 
wire u2__abc_52138_new_n13330_; 
wire u2__abc_52138_new_n13331_; 
wire u2__abc_52138_new_n13332_; 
wire u2__abc_52138_new_n13333_; 
wire u2__abc_52138_new_n13334_; 
wire u2__abc_52138_new_n13335_; 
wire u2__abc_52138_new_n13337_; 
wire u2__abc_52138_new_n13338_; 
wire u2__abc_52138_new_n13339_; 
wire u2__abc_52138_new_n13340_; 
wire u2__abc_52138_new_n13341_; 
wire u2__abc_52138_new_n13342_; 
wire u2__abc_52138_new_n13343_; 
wire u2__abc_52138_new_n13345_; 
wire u2__abc_52138_new_n13346_; 
wire u2__abc_52138_new_n13347_; 
wire u2__abc_52138_new_n13348_; 
wire u2__abc_52138_new_n13349_; 
wire u2__abc_52138_new_n13350_; 
wire u2__abc_52138_new_n13351_; 
wire u2__abc_52138_new_n13353_; 
wire u2__abc_52138_new_n13354_; 
wire u2__abc_52138_new_n13355_; 
wire u2__abc_52138_new_n13356_; 
wire u2__abc_52138_new_n13357_; 
wire u2__abc_52138_new_n13358_; 
wire u2__abc_52138_new_n13359_; 
wire u2__abc_52138_new_n13361_; 
wire u2__abc_52138_new_n13362_; 
wire u2__abc_52138_new_n13363_; 
wire u2__abc_52138_new_n13364_; 
wire u2__abc_52138_new_n13365_; 
wire u2__abc_52138_new_n13366_; 
wire u2__abc_52138_new_n13368_; 
wire u2__abc_52138_new_n13369_; 
wire u2__abc_52138_new_n13370_; 
wire u2__abc_52138_new_n13371_; 
wire u2__abc_52138_new_n13372_; 
wire u2__abc_52138_new_n13373_; 
wire u2__abc_52138_new_n13374_; 
wire u2__abc_52138_new_n13376_; 
wire u2__abc_52138_new_n13377_; 
wire u2__abc_52138_new_n13378_; 
wire u2__abc_52138_new_n13379_; 
wire u2__abc_52138_new_n13380_; 
wire u2__abc_52138_new_n13381_; 
wire u2__abc_52138_new_n13382_; 
wire u2__abc_52138_new_n13384_; 
wire u2__abc_52138_new_n13385_; 
wire u2__abc_52138_new_n13386_; 
wire u2__abc_52138_new_n13387_; 
wire u2__abc_52138_new_n13388_; 
wire u2__abc_52138_new_n13389_; 
wire u2__abc_52138_new_n13390_; 
wire u2__abc_52138_new_n13392_; 
wire u2__abc_52138_new_n13393_; 
wire u2__abc_52138_new_n13394_; 
wire u2__abc_52138_new_n13395_; 
wire u2__abc_52138_new_n13396_; 
wire u2__abc_52138_new_n13397_; 
wire u2__abc_52138_new_n13399_; 
wire u2__abc_52138_new_n13400_; 
wire u2__abc_52138_new_n13401_; 
wire u2__abc_52138_new_n13402_; 
wire u2__abc_52138_new_n13403_; 
wire u2__abc_52138_new_n13404_; 
wire u2__abc_52138_new_n13405_; 
wire u2__abc_52138_new_n13407_; 
wire u2__abc_52138_new_n13408_; 
wire u2__abc_52138_new_n13409_; 
wire u2__abc_52138_new_n13410_; 
wire u2__abc_52138_new_n13411_; 
wire u2__abc_52138_new_n13412_; 
wire u2__abc_52138_new_n13413_; 
wire u2__abc_52138_new_n13415_; 
wire u2__abc_52138_new_n13416_; 
wire u2__abc_52138_new_n13417_; 
wire u2__abc_52138_new_n13418_; 
wire u2__abc_52138_new_n13419_; 
wire u2__abc_52138_new_n13420_; 
wire u2__abc_52138_new_n13421_; 
wire u2__abc_52138_new_n13423_; 
wire u2__abc_52138_new_n13424_; 
wire u2__abc_52138_new_n13425_; 
wire u2__abc_52138_new_n13426_; 
wire u2__abc_52138_new_n13427_; 
wire u2__abc_52138_new_n13428_; 
wire u2__abc_52138_new_n13430_; 
wire u2__abc_52138_new_n13431_; 
wire u2__abc_52138_new_n13432_; 
wire u2__abc_52138_new_n13433_; 
wire u2__abc_52138_new_n13434_; 
wire u2__abc_52138_new_n13435_; 
wire u2__abc_52138_new_n13436_; 
wire u2__abc_52138_new_n13438_; 
wire u2__abc_52138_new_n13439_; 
wire u2__abc_52138_new_n13440_; 
wire u2__abc_52138_new_n13441_; 
wire u2__abc_52138_new_n13442_; 
wire u2__abc_52138_new_n13443_; 
wire u2__abc_52138_new_n13444_; 
wire u2__abc_52138_new_n13446_; 
wire u2__abc_52138_new_n13447_; 
wire u2__abc_52138_new_n13448_; 
wire u2__abc_52138_new_n13449_; 
wire u2__abc_52138_new_n13450_; 
wire u2__abc_52138_new_n13451_; 
wire u2__abc_52138_new_n13452_; 
wire u2__abc_52138_new_n13454_; 
wire u2__abc_52138_new_n13455_; 
wire u2__abc_52138_new_n13456_; 
wire u2__abc_52138_new_n13457_; 
wire u2__abc_52138_new_n13458_; 
wire u2__abc_52138_new_n13459_; 
wire u2__abc_52138_new_n13461_; 
wire u2__abc_52138_new_n13462_; 
wire u2__abc_52138_new_n13463_; 
wire u2__abc_52138_new_n13464_; 
wire u2__abc_52138_new_n13465_; 
wire u2__abc_52138_new_n13466_; 
wire u2__abc_52138_new_n13467_; 
wire u2__abc_52138_new_n13469_; 
wire u2__abc_52138_new_n13470_; 
wire u2__abc_52138_new_n13471_; 
wire u2__abc_52138_new_n13472_; 
wire u2__abc_52138_new_n13473_; 
wire u2__abc_52138_new_n13474_; 
wire u2__abc_52138_new_n13475_; 
wire u2__abc_52138_new_n13477_; 
wire u2__abc_52138_new_n13478_; 
wire u2__abc_52138_new_n13479_; 
wire u2__abc_52138_new_n13480_; 
wire u2__abc_52138_new_n13481_; 
wire u2__abc_52138_new_n13482_; 
wire u2__abc_52138_new_n13483_; 
wire u2__abc_52138_new_n13485_; 
wire u2__abc_52138_new_n13486_; 
wire u2__abc_52138_new_n13487_; 
wire u2__abc_52138_new_n13488_; 
wire u2__abc_52138_new_n13489_; 
wire u2__abc_52138_new_n13490_; 
wire u2__abc_52138_new_n13492_; 
wire u2__abc_52138_new_n13493_; 
wire u2__abc_52138_new_n13494_; 
wire u2__abc_52138_new_n13495_; 
wire u2__abc_52138_new_n13496_; 
wire u2__abc_52138_new_n13497_; 
wire u2__abc_52138_new_n13498_; 
wire u2__abc_52138_new_n13500_; 
wire u2__abc_52138_new_n13501_; 
wire u2__abc_52138_new_n13502_; 
wire u2__abc_52138_new_n13503_; 
wire u2__abc_52138_new_n13504_; 
wire u2__abc_52138_new_n13505_; 
wire u2__abc_52138_new_n13506_; 
wire u2__abc_52138_new_n13508_; 
wire u2__abc_52138_new_n13509_; 
wire u2__abc_52138_new_n13510_; 
wire u2__abc_52138_new_n13511_; 
wire u2__abc_52138_new_n13512_; 
wire u2__abc_52138_new_n13513_; 
wire u2__abc_52138_new_n13514_; 
wire u2__abc_52138_new_n13516_; 
wire u2__abc_52138_new_n13517_; 
wire u2__abc_52138_new_n13518_; 
wire u2__abc_52138_new_n13519_; 
wire u2__abc_52138_new_n13520_; 
wire u2__abc_52138_new_n13521_; 
wire u2__abc_52138_new_n13523_; 
wire u2__abc_52138_new_n13524_; 
wire u2__abc_52138_new_n13525_; 
wire u2__abc_52138_new_n13526_; 
wire u2__abc_52138_new_n13527_; 
wire u2__abc_52138_new_n13528_; 
wire u2__abc_52138_new_n13529_; 
wire u2__abc_52138_new_n13531_; 
wire u2__abc_52138_new_n13532_; 
wire u2__abc_52138_new_n13533_; 
wire u2__abc_52138_new_n13534_; 
wire u2__abc_52138_new_n13535_; 
wire u2__abc_52138_new_n13536_; 
wire u2__abc_52138_new_n13537_; 
wire u2__abc_52138_new_n13539_; 
wire u2__abc_52138_new_n13540_; 
wire u2__abc_52138_new_n13541_; 
wire u2__abc_52138_new_n13542_; 
wire u2__abc_52138_new_n13543_; 
wire u2__abc_52138_new_n13544_; 
wire u2__abc_52138_new_n13545_; 
wire u2__abc_52138_new_n13547_; 
wire u2__abc_52138_new_n13548_; 
wire u2__abc_52138_new_n13549_; 
wire u2__abc_52138_new_n13550_; 
wire u2__abc_52138_new_n13551_; 
wire u2__abc_52138_new_n13552_; 
wire u2__abc_52138_new_n13554_; 
wire u2__abc_52138_new_n13555_; 
wire u2__abc_52138_new_n13556_; 
wire u2__abc_52138_new_n13557_; 
wire u2__abc_52138_new_n13558_; 
wire u2__abc_52138_new_n13559_; 
wire u2__abc_52138_new_n13560_; 
wire u2__abc_52138_new_n13562_; 
wire u2__abc_52138_new_n13563_; 
wire u2__abc_52138_new_n13564_; 
wire u2__abc_52138_new_n13565_; 
wire u2__abc_52138_new_n13566_; 
wire u2__abc_52138_new_n13567_; 
wire u2__abc_52138_new_n13568_; 
wire u2__abc_52138_new_n13570_; 
wire u2__abc_52138_new_n13571_; 
wire u2__abc_52138_new_n13572_; 
wire u2__abc_52138_new_n13573_; 
wire u2__abc_52138_new_n13574_; 
wire u2__abc_52138_new_n13575_; 
wire u2__abc_52138_new_n13576_; 
wire u2__abc_52138_new_n13578_; 
wire u2__abc_52138_new_n13579_; 
wire u2__abc_52138_new_n13580_; 
wire u2__abc_52138_new_n13581_; 
wire u2__abc_52138_new_n13582_; 
wire u2__abc_52138_new_n13583_; 
wire u2__abc_52138_new_n13585_; 
wire u2__abc_52138_new_n13586_; 
wire u2__abc_52138_new_n13587_; 
wire u2__abc_52138_new_n13588_; 
wire u2__abc_52138_new_n13589_; 
wire u2__abc_52138_new_n13590_; 
wire u2__abc_52138_new_n13591_; 
wire u2__abc_52138_new_n13593_; 
wire u2__abc_52138_new_n13594_; 
wire u2__abc_52138_new_n13595_; 
wire u2__abc_52138_new_n13596_; 
wire u2__abc_52138_new_n13597_; 
wire u2__abc_52138_new_n13598_; 
wire u2__abc_52138_new_n13599_; 
wire u2__abc_52138_new_n13601_; 
wire u2__abc_52138_new_n13602_; 
wire u2__abc_52138_new_n13603_; 
wire u2__abc_52138_new_n13604_; 
wire u2__abc_52138_new_n13605_; 
wire u2__abc_52138_new_n13606_; 
wire u2__abc_52138_new_n13607_; 
wire u2__abc_52138_new_n13609_; 
wire u2__abc_52138_new_n13610_; 
wire u2__abc_52138_new_n13611_; 
wire u2__abc_52138_new_n13612_; 
wire u2__abc_52138_new_n13613_; 
wire u2__abc_52138_new_n13614_; 
wire u2__abc_52138_new_n13616_; 
wire u2__abc_52138_new_n13617_; 
wire u2__abc_52138_new_n13618_; 
wire u2__abc_52138_new_n13619_; 
wire u2__abc_52138_new_n13620_; 
wire u2__abc_52138_new_n13621_; 
wire u2__abc_52138_new_n13622_; 
wire u2__abc_52138_new_n13624_; 
wire u2__abc_52138_new_n13625_; 
wire u2__abc_52138_new_n13626_; 
wire u2__abc_52138_new_n13627_; 
wire u2__abc_52138_new_n13628_; 
wire u2__abc_52138_new_n13629_; 
wire u2__abc_52138_new_n13630_; 
wire u2__abc_52138_new_n13632_; 
wire u2__abc_52138_new_n13633_; 
wire u2__abc_52138_new_n13634_; 
wire u2__abc_52138_new_n13635_; 
wire u2__abc_52138_new_n13636_; 
wire u2__abc_52138_new_n13637_; 
wire u2__abc_52138_new_n13638_; 
wire u2__abc_52138_new_n13640_; 
wire u2__abc_52138_new_n13641_; 
wire u2__abc_52138_new_n13642_; 
wire u2__abc_52138_new_n13643_; 
wire u2__abc_52138_new_n13644_; 
wire u2__abc_52138_new_n13645_; 
wire u2__abc_52138_new_n13647_; 
wire u2__abc_52138_new_n13648_; 
wire u2__abc_52138_new_n13649_; 
wire u2__abc_52138_new_n13650_; 
wire u2__abc_52138_new_n13651_; 
wire u2__abc_52138_new_n13652_; 
wire u2__abc_52138_new_n13653_; 
wire u2__abc_52138_new_n13655_; 
wire u2__abc_52138_new_n13656_; 
wire u2__abc_52138_new_n13657_; 
wire u2__abc_52138_new_n13658_; 
wire u2__abc_52138_new_n13659_; 
wire u2__abc_52138_new_n13660_; 
wire u2__abc_52138_new_n13661_; 
wire u2__abc_52138_new_n13663_; 
wire u2__abc_52138_new_n13664_; 
wire u2__abc_52138_new_n13665_; 
wire u2__abc_52138_new_n13666_; 
wire u2__abc_52138_new_n13667_; 
wire u2__abc_52138_new_n13668_; 
wire u2__abc_52138_new_n13669_; 
wire u2__abc_52138_new_n13671_; 
wire u2__abc_52138_new_n13672_; 
wire u2__abc_52138_new_n13673_; 
wire u2__abc_52138_new_n13674_; 
wire u2__abc_52138_new_n13675_; 
wire u2__abc_52138_new_n13676_; 
wire u2__abc_52138_new_n13678_; 
wire u2__abc_52138_new_n13679_; 
wire u2__abc_52138_new_n13680_; 
wire u2__abc_52138_new_n13681_; 
wire u2__abc_52138_new_n13682_; 
wire u2__abc_52138_new_n13683_; 
wire u2__abc_52138_new_n13684_; 
wire u2__abc_52138_new_n13686_; 
wire u2__abc_52138_new_n13687_; 
wire u2__abc_52138_new_n13688_; 
wire u2__abc_52138_new_n13689_; 
wire u2__abc_52138_new_n13690_; 
wire u2__abc_52138_new_n13691_; 
wire u2__abc_52138_new_n13692_; 
wire u2__abc_52138_new_n13694_; 
wire u2__abc_52138_new_n13695_; 
wire u2__abc_52138_new_n13696_; 
wire u2__abc_52138_new_n13697_; 
wire u2__abc_52138_new_n13698_; 
wire u2__abc_52138_new_n13699_; 
wire u2__abc_52138_new_n13700_; 
wire u2__abc_52138_new_n13702_; 
wire u2__abc_52138_new_n13703_; 
wire u2__abc_52138_new_n13704_; 
wire u2__abc_52138_new_n13705_; 
wire u2__abc_52138_new_n13706_; 
wire u2__abc_52138_new_n13707_; 
wire u2__abc_52138_new_n13709_; 
wire u2__abc_52138_new_n13710_; 
wire u2__abc_52138_new_n13711_; 
wire u2__abc_52138_new_n13712_; 
wire u2__abc_52138_new_n13713_; 
wire u2__abc_52138_new_n13714_; 
wire u2__abc_52138_new_n13715_; 
wire u2__abc_52138_new_n13717_; 
wire u2__abc_52138_new_n13718_; 
wire u2__abc_52138_new_n13719_; 
wire u2__abc_52138_new_n13720_; 
wire u2__abc_52138_new_n13721_; 
wire u2__abc_52138_new_n13722_; 
wire u2__abc_52138_new_n13723_; 
wire u2__abc_52138_new_n13725_; 
wire u2__abc_52138_new_n13726_; 
wire u2__abc_52138_new_n13727_; 
wire u2__abc_52138_new_n13728_; 
wire u2__abc_52138_new_n13729_; 
wire u2__abc_52138_new_n13730_; 
wire u2__abc_52138_new_n13731_; 
wire u2__abc_52138_new_n13733_; 
wire u2__abc_52138_new_n13734_; 
wire u2__abc_52138_new_n13735_; 
wire u2__abc_52138_new_n13736_; 
wire u2__abc_52138_new_n13737_; 
wire u2__abc_52138_new_n13738_; 
wire u2__abc_52138_new_n13740_; 
wire u2__abc_52138_new_n13741_; 
wire u2__abc_52138_new_n13742_; 
wire u2__abc_52138_new_n13743_; 
wire u2__abc_52138_new_n13744_; 
wire u2__abc_52138_new_n13745_; 
wire u2__abc_52138_new_n13746_; 
wire u2__abc_52138_new_n13748_; 
wire u2__abc_52138_new_n13749_; 
wire u2__abc_52138_new_n13750_; 
wire u2__abc_52138_new_n13751_; 
wire u2__abc_52138_new_n13752_; 
wire u2__abc_52138_new_n13753_; 
wire u2__abc_52138_new_n13754_; 
wire u2__abc_52138_new_n13756_; 
wire u2__abc_52138_new_n13757_; 
wire u2__abc_52138_new_n13758_; 
wire u2__abc_52138_new_n13759_; 
wire u2__abc_52138_new_n13760_; 
wire u2__abc_52138_new_n13761_; 
wire u2__abc_52138_new_n13762_; 
wire u2__abc_52138_new_n13764_; 
wire u2__abc_52138_new_n13765_; 
wire u2__abc_52138_new_n13766_; 
wire u2__abc_52138_new_n13767_; 
wire u2__abc_52138_new_n13768_; 
wire u2__abc_52138_new_n13769_; 
wire u2__abc_52138_new_n13771_; 
wire u2__abc_52138_new_n13772_; 
wire u2__abc_52138_new_n13773_; 
wire u2__abc_52138_new_n13774_; 
wire u2__abc_52138_new_n13775_; 
wire u2__abc_52138_new_n13776_; 
wire u2__abc_52138_new_n13777_; 
wire u2__abc_52138_new_n13779_; 
wire u2__abc_52138_new_n13780_; 
wire u2__abc_52138_new_n13781_; 
wire u2__abc_52138_new_n13782_; 
wire u2__abc_52138_new_n13783_; 
wire u2__abc_52138_new_n13784_; 
wire u2__abc_52138_new_n13785_; 
wire u2__abc_52138_new_n13787_; 
wire u2__abc_52138_new_n13788_; 
wire u2__abc_52138_new_n13789_; 
wire u2__abc_52138_new_n13790_; 
wire u2__abc_52138_new_n13791_; 
wire u2__abc_52138_new_n13792_; 
wire u2__abc_52138_new_n13793_; 
wire u2__abc_52138_new_n13795_; 
wire u2__abc_52138_new_n13796_; 
wire u2__abc_52138_new_n13797_; 
wire u2__abc_52138_new_n13798_; 
wire u2__abc_52138_new_n13799_; 
wire u2__abc_52138_new_n13800_; 
wire u2__abc_52138_new_n13802_; 
wire u2__abc_52138_new_n13803_; 
wire u2__abc_52138_new_n13804_; 
wire u2__abc_52138_new_n13805_; 
wire u2__abc_52138_new_n13806_; 
wire u2__abc_52138_new_n13807_; 
wire u2__abc_52138_new_n13808_; 
wire u2__abc_52138_new_n13810_; 
wire u2__abc_52138_new_n13811_; 
wire u2__abc_52138_new_n13812_; 
wire u2__abc_52138_new_n13813_; 
wire u2__abc_52138_new_n13814_; 
wire u2__abc_52138_new_n13815_; 
wire u2__abc_52138_new_n13816_; 
wire u2__abc_52138_new_n13818_; 
wire u2__abc_52138_new_n13819_; 
wire u2__abc_52138_new_n13820_; 
wire u2__abc_52138_new_n13821_; 
wire u2__abc_52138_new_n13822_; 
wire u2__abc_52138_new_n13823_; 
wire u2__abc_52138_new_n13824_; 
wire u2__abc_52138_new_n13826_; 
wire u2__abc_52138_new_n13827_; 
wire u2__abc_52138_new_n13828_; 
wire u2__abc_52138_new_n13829_; 
wire u2__abc_52138_new_n13830_; 
wire u2__abc_52138_new_n13831_; 
wire u2__abc_52138_new_n13833_; 
wire u2__abc_52138_new_n13834_; 
wire u2__abc_52138_new_n13835_; 
wire u2__abc_52138_new_n13836_; 
wire u2__abc_52138_new_n13837_; 
wire u2__abc_52138_new_n13838_; 
wire u2__abc_52138_new_n13839_; 
wire u2__abc_52138_new_n13841_; 
wire u2__abc_52138_new_n13842_; 
wire u2__abc_52138_new_n13843_; 
wire u2__abc_52138_new_n13844_; 
wire u2__abc_52138_new_n13845_; 
wire u2__abc_52138_new_n13846_; 
wire u2__abc_52138_new_n13847_; 
wire u2__abc_52138_new_n13849_; 
wire u2__abc_52138_new_n13850_; 
wire u2__abc_52138_new_n13851_; 
wire u2__abc_52138_new_n13852_; 
wire u2__abc_52138_new_n13853_; 
wire u2__abc_52138_new_n13854_; 
wire u2__abc_52138_new_n13855_; 
wire u2__abc_52138_new_n13857_; 
wire u2__abc_52138_new_n13858_; 
wire u2__abc_52138_new_n13859_; 
wire u2__abc_52138_new_n13860_; 
wire u2__abc_52138_new_n13861_; 
wire u2__abc_52138_new_n13862_; 
wire u2__abc_52138_new_n13864_; 
wire u2__abc_52138_new_n13865_; 
wire u2__abc_52138_new_n13866_; 
wire u2__abc_52138_new_n13867_; 
wire u2__abc_52138_new_n13868_; 
wire u2__abc_52138_new_n13869_; 
wire u2__abc_52138_new_n13870_; 
wire u2__abc_52138_new_n13872_; 
wire u2__abc_52138_new_n13873_; 
wire u2__abc_52138_new_n13874_; 
wire u2__abc_52138_new_n13875_; 
wire u2__abc_52138_new_n13876_; 
wire u2__abc_52138_new_n13877_; 
wire u2__abc_52138_new_n13878_; 
wire u2__abc_52138_new_n13880_; 
wire u2__abc_52138_new_n13881_; 
wire u2__abc_52138_new_n13882_; 
wire u2__abc_52138_new_n13883_; 
wire u2__abc_52138_new_n13884_; 
wire u2__abc_52138_new_n13885_; 
wire u2__abc_52138_new_n13886_; 
wire u2__abc_52138_new_n13888_; 
wire u2__abc_52138_new_n13889_; 
wire u2__abc_52138_new_n13890_; 
wire u2__abc_52138_new_n13891_; 
wire u2__abc_52138_new_n13892_; 
wire u2__abc_52138_new_n13893_; 
wire u2__abc_52138_new_n13895_; 
wire u2__abc_52138_new_n13896_; 
wire u2__abc_52138_new_n13897_; 
wire u2__abc_52138_new_n13898_; 
wire u2__abc_52138_new_n13899_; 
wire u2__abc_52138_new_n13900_; 
wire u2__abc_52138_new_n13901_; 
wire u2__abc_52138_new_n13903_; 
wire u2__abc_52138_new_n13904_; 
wire u2__abc_52138_new_n13905_; 
wire u2__abc_52138_new_n13906_; 
wire u2__abc_52138_new_n13907_; 
wire u2__abc_52138_new_n13908_; 
wire u2__abc_52138_new_n13909_; 
wire u2__abc_52138_new_n13911_; 
wire u2__abc_52138_new_n13912_; 
wire u2__abc_52138_new_n13913_; 
wire u2__abc_52138_new_n13914_; 
wire u2__abc_52138_new_n13915_; 
wire u2__abc_52138_new_n13916_; 
wire u2__abc_52138_new_n13917_; 
wire u2__abc_52138_new_n13919_; 
wire u2__abc_52138_new_n13920_; 
wire u2__abc_52138_new_n13921_; 
wire u2__abc_52138_new_n13922_; 
wire u2__abc_52138_new_n13923_; 
wire u2__abc_52138_new_n13924_; 
wire u2__abc_52138_new_n13926_; 
wire u2__abc_52138_new_n13927_; 
wire u2__abc_52138_new_n13928_; 
wire u2__abc_52138_new_n13929_; 
wire u2__abc_52138_new_n13930_; 
wire u2__abc_52138_new_n13931_; 
wire u2__abc_52138_new_n13932_; 
wire u2__abc_52138_new_n13934_; 
wire u2__abc_52138_new_n13935_; 
wire u2__abc_52138_new_n13936_; 
wire u2__abc_52138_new_n13937_; 
wire u2__abc_52138_new_n13938_; 
wire u2__abc_52138_new_n13939_; 
wire u2__abc_52138_new_n13940_; 
wire u2__abc_52138_new_n13942_; 
wire u2__abc_52138_new_n13943_; 
wire u2__abc_52138_new_n13944_; 
wire u2__abc_52138_new_n13945_; 
wire u2__abc_52138_new_n13946_; 
wire u2__abc_52138_new_n13947_; 
wire u2__abc_52138_new_n13948_; 
wire u2__abc_52138_new_n13950_; 
wire u2__abc_52138_new_n13951_; 
wire u2__abc_52138_new_n13952_; 
wire u2__abc_52138_new_n13953_; 
wire u2__abc_52138_new_n13954_; 
wire u2__abc_52138_new_n13955_; 
wire u2__abc_52138_new_n13957_; 
wire u2__abc_52138_new_n13958_; 
wire u2__abc_52138_new_n13959_; 
wire u2__abc_52138_new_n13960_; 
wire u2__abc_52138_new_n13961_; 
wire u2__abc_52138_new_n13962_; 
wire u2__abc_52138_new_n13963_; 
wire u2__abc_52138_new_n13964_; 
wire u2__abc_52138_new_n13966_; 
wire u2__abc_52138_new_n13967_; 
wire u2__abc_52138_new_n13968_; 
wire u2__abc_52138_new_n13969_; 
wire u2__abc_52138_new_n13970_; 
wire u2__abc_52138_new_n13971_; 
wire u2__abc_52138_new_n13972_; 
wire u2__abc_52138_new_n13974_; 
wire u2__abc_52138_new_n13975_; 
wire u2__abc_52138_new_n13976_; 
wire u2__abc_52138_new_n13977_; 
wire u2__abc_52138_new_n13978_; 
wire u2__abc_52138_new_n13979_; 
wire u2__abc_52138_new_n13980_; 
wire u2__abc_52138_new_n13982_; 
wire u2__abc_52138_new_n13983_; 
wire u2__abc_52138_new_n13984_; 
wire u2__abc_52138_new_n13985_; 
wire u2__abc_52138_new_n13986_; 
wire u2__abc_52138_new_n13987_; 
wire u2__abc_52138_new_n13989_; 
wire u2__abc_52138_new_n13990_; 
wire u2__abc_52138_new_n13991_; 
wire u2__abc_52138_new_n13992_; 
wire u2__abc_52138_new_n13993_; 
wire u2__abc_52138_new_n13994_; 
wire u2__abc_52138_new_n13995_; 
wire u2__abc_52138_new_n13997_; 
wire u2__abc_52138_new_n13998_; 
wire u2__abc_52138_new_n13999_; 
wire u2__abc_52138_new_n14000_; 
wire u2__abc_52138_new_n14001_; 
wire u2__abc_52138_new_n14002_; 
wire u2__abc_52138_new_n14003_; 
wire u2__abc_52138_new_n14005_; 
wire u2__abc_52138_new_n14006_; 
wire u2__abc_52138_new_n14007_; 
wire u2__abc_52138_new_n14008_; 
wire u2__abc_52138_new_n14009_; 
wire u2__abc_52138_new_n14010_; 
wire u2__abc_52138_new_n14011_; 
wire u2__abc_52138_new_n14013_; 
wire u2__abc_52138_new_n14014_; 
wire u2__abc_52138_new_n14015_; 
wire u2__abc_52138_new_n14016_; 
wire u2__abc_52138_new_n14017_; 
wire u2__abc_52138_new_n14018_; 
wire u2__abc_52138_new_n14020_; 
wire u2__abc_52138_new_n14021_; 
wire u2__abc_52138_new_n14022_; 
wire u2__abc_52138_new_n14023_; 
wire u2__abc_52138_new_n14024_; 
wire u2__abc_52138_new_n14025_; 
wire u2__abc_52138_new_n14026_; 
wire u2__abc_52138_new_n14028_; 
wire u2__abc_52138_new_n14029_; 
wire u2__abc_52138_new_n14030_; 
wire u2__abc_52138_new_n14031_; 
wire u2__abc_52138_new_n14032_; 
wire u2__abc_52138_new_n14033_; 
wire u2__abc_52138_new_n14034_; 
wire u2__abc_52138_new_n14036_; 
wire u2__abc_52138_new_n14037_; 
wire u2__abc_52138_new_n14038_; 
wire u2__abc_52138_new_n14039_; 
wire u2__abc_52138_new_n14040_; 
wire u2__abc_52138_new_n14041_; 
wire u2__abc_52138_new_n14042_; 
wire u2__abc_52138_new_n14044_; 
wire u2__abc_52138_new_n14045_; 
wire u2__abc_52138_new_n14046_; 
wire u2__abc_52138_new_n14047_; 
wire u2__abc_52138_new_n14048_; 
wire u2__abc_52138_new_n14049_; 
wire u2__abc_52138_new_n14051_; 
wire u2__abc_52138_new_n14052_; 
wire u2__abc_52138_new_n14053_; 
wire u2__abc_52138_new_n14054_; 
wire u2__abc_52138_new_n14055_; 
wire u2__abc_52138_new_n14056_; 
wire u2__abc_52138_new_n14057_; 
wire u2__abc_52138_new_n14058_; 
wire u2__abc_52138_new_n14060_; 
wire u2__abc_52138_new_n14061_; 
wire u2__abc_52138_new_n14062_; 
wire u2__abc_52138_new_n14063_; 
wire u2__abc_52138_new_n14064_; 
wire u2__abc_52138_new_n14065_; 
wire u2__abc_52138_new_n14066_; 
wire u2__abc_52138_new_n14068_; 
wire u2__abc_52138_new_n14069_; 
wire u2__abc_52138_new_n14070_; 
wire u2__abc_52138_new_n14071_; 
wire u2__abc_52138_new_n14072_; 
wire u2__abc_52138_new_n14073_; 
wire u2__abc_52138_new_n14074_; 
wire u2__abc_52138_new_n14076_; 
wire u2__abc_52138_new_n14077_; 
wire u2__abc_52138_new_n14078_; 
wire u2__abc_52138_new_n14079_; 
wire u2__abc_52138_new_n14080_; 
wire u2__abc_52138_new_n14081_; 
wire u2__abc_52138_new_n14083_; 
wire u2__abc_52138_new_n14084_; 
wire u2__abc_52138_new_n14085_; 
wire u2__abc_52138_new_n14086_; 
wire u2__abc_52138_new_n14087_; 
wire u2__abc_52138_new_n14088_; 
wire u2__abc_52138_new_n14089_; 
wire u2__abc_52138_new_n14091_; 
wire u2__abc_52138_new_n14092_; 
wire u2__abc_52138_new_n14093_; 
wire u2__abc_52138_new_n14094_; 
wire u2__abc_52138_new_n14095_; 
wire u2__abc_52138_new_n14096_; 
wire u2__abc_52138_new_n14097_; 
wire u2__abc_52138_new_n14099_; 
wire u2__abc_52138_new_n14100_; 
wire u2__abc_52138_new_n14101_; 
wire u2__abc_52138_new_n14102_; 
wire u2__abc_52138_new_n14103_; 
wire u2__abc_52138_new_n14104_; 
wire u2__abc_52138_new_n14105_; 
wire u2__abc_52138_new_n14107_; 
wire u2__abc_52138_new_n14108_; 
wire u2__abc_52138_new_n14109_; 
wire u2__abc_52138_new_n14110_; 
wire u2__abc_52138_new_n14111_; 
wire u2__abc_52138_new_n14112_; 
wire u2__abc_52138_new_n14114_; 
wire u2__abc_52138_new_n14115_; 
wire u2__abc_52138_new_n14116_; 
wire u2__abc_52138_new_n14117_; 
wire u2__abc_52138_new_n14118_; 
wire u2__abc_52138_new_n14119_; 
wire u2__abc_52138_new_n14120_; 
wire u2__abc_52138_new_n14122_; 
wire u2__abc_52138_new_n14123_; 
wire u2__abc_52138_new_n14124_; 
wire u2__abc_52138_new_n14125_; 
wire u2__abc_52138_new_n14126_; 
wire u2__abc_52138_new_n14127_; 
wire u2__abc_52138_new_n14128_; 
wire u2__abc_52138_new_n14130_; 
wire u2__abc_52138_new_n14131_; 
wire u2__abc_52138_new_n14132_; 
wire u2__abc_52138_new_n14133_; 
wire u2__abc_52138_new_n14134_; 
wire u2__abc_52138_new_n14135_; 
wire u2__abc_52138_new_n14136_; 
wire u2__abc_52138_new_n14138_; 
wire u2__abc_52138_new_n14139_; 
wire u2__abc_52138_new_n14140_; 
wire u2__abc_52138_new_n14141_; 
wire u2__abc_52138_new_n14142_; 
wire u2__abc_52138_new_n14143_; 
wire u2__abc_52138_new_n14145_; 
wire u2__abc_52138_new_n14146_; 
wire u2__abc_52138_new_n14147_; 
wire u2__abc_52138_new_n14148_; 
wire u2__abc_52138_new_n14149_; 
wire u2__abc_52138_new_n14150_; 
wire u2__abc_52138_new_n14151_; 
wire u2__abc_52138_new_n14153_; 
wire u2__abc_52138_new_n14154_; 
wire u2__abc_52138_new_n14155_; 
wire u2__abc_52138_new_n14156_; 
wire u2__abc_52138_new_n14157_; 
wire u2__abc_52138_new_n14158_; 
wire u2__abc_52138_new_n14159_; 
wire u2__abc_52138_new_n14161_; 
wire u2__abc_52138_new_n14162_; 
wire u2__abc_52138_new_n14163_; 
wire u2__abc_52138_new_n14164_; 
wire u2__abc_52138_new_n14165_; 
wire u2__abc_52138_new_n14166_; 
wire u2__abc_52138_new_n14167_; 
wire u2__abc_52138_new_n14169_; 
wire u2__abc_52138_new_n14170_; 
wire u2__abc_52138_new_n14171_; 
wire u2__abc_52138_new_n14172_; 
wire u2__abc_52138_new_n14173_; 
wire u2__abc_52138_new_n14174_; 
wire u2__abc_52138_new_n14176_; 
wire u2__abc_52138_new_n14177_; 
wire u2__abc_52138_new_n14178_; 
wire u2__abc_52138_new_n14179_; 
wire u2__abc_52138_new_n14180_; 
wire u2__abc_52138_new_n14181_; 
wire u2__abc_52138_new_n14182_; 
wire u2__abc_52138_new_n14184_; 
wire u2__abc_52138_new_n14185_; 
wire u2__abc_52138_new_n14186_; 
wire u2__abc_52138_new_n14187_; 
wire u2__abc_52138_new_n14188_; 
wire u2__abc_52138_new_n14189_; 
wire u2__abc_52138_new_n14190_; 
wire u2__abc_52138_new_n14192_; 
wire u2__abc_52138_new_n14193_; 
wire u2__abc_52138_new_n14194_; 
wire u2__abc_52138_new_n14195_; 
wire u2__abc_52138_new_n14196_; 
wire u2__abc_52138_new_n14197_; 
wire u2__abc_52138_new_n14198_; 
wire u2__abc_52138_new_n14200_; 
wire u2__abc_52138_new_n14201_; 
wire u2__abc_52138_new_n14202_; 
wire u2__abc_52138_new_n14203_; 
wire u2__abc_52138_new_n14204_; 
wire u2__abc_52138_new_n14205_; 
wire u2__abc_52138_new_n14207_; 
wire u2__abc_52138_new_n14208_; 
wire u2__abc_52138_new_n14209_; 
wire u2__abc_52138_new_n14210_; 
wire u2__abc_52138_new_n14211_; 
wire u2__abc_52138_new_n14212_; 
wire u2__abc_52138_new_n14213_; 
wire u2__abc_52138_new_n14215_; 
wire u2__abc_52138_new_n14216_; 
wire u2__abc_52138_new_n14217_; 
wire u2__abc_52138_new_n14218_; 
wire u2__abc_52138_new_n14219_; 
wire u2__abc_52138_new_n14220_; 
wire u2__abc_52138_new_n14221_; 
wire u2__abc_52138_new_n14223_; 
wire u2__abc_52138_new_n14224_; 
wire u2__abc_52138_new_n14225_; 
wire u2__abc_52138_new_n14226_; 
wire u2__abc_52138_new_n14227_; 
wire u2__abc_52138_new_n14228_; 
wire u2__abc_52138_new_n14229_; 
wire u2__abc_52138_new_n14231_; 
wire u2__abc_52138_new_n14232_; 
wire u2__abc_52138_new_n14233_; 
wire u2__abc_52138_new_n14234_; 
wire u2__abc_52138_new_n14235_; 
wire u2__abc_52138_new_n14236_; 
wire u2__abc_52138_new_n14238_; 
wire u2__abc_52138_new_n14239_; 
wire u2__abc_52138_new_n14240_; 
wire u2__abc_52138_new_n14241_; 
wire u2__abc_52138_new_n14242_; 
wire u2__abc_52138_new_n14243_; 
wire u2__abc_52138_new_n14244_; 
wire u2__abc_52138_new_n14246_; 
wire u2__abc_52138_new_n14247_; 
wire u2__abc_52138_new_n14248_; 
wire u2__abc_52138_new_n14249_; 
wire u2__abc_52138_new_n14250_; 
wire u2__abc_52138_new_n14251_; 
wire u2__abc_52138_new_n14252_; 
wire u2__abc_52138_new_n14254_; 
wire u2__abc_52138_new_n14255_; 
wire u2__abc_52138_new_n14256_; 
wire u2__abc_52138_new_n14257_; 
wire u2__abc_52138_new_n14258_; 
wire u2__abc_52138_new_n14259_; 
wire u2__abc_52138_new_n14260_; 
wire u2__abc_52138_new_n14262_; 
wire u2__abc_52138_new_n14263_; 
wire u2__abc_52138_new_n14264_; 
wire u2__abc_52138_new_n14265_; 
wire u2__abc_52138_new_n14266_; 
wire u2__abc_52138_new_n14267_; 
wire u2__abc_52138_new_n14269_; 
wire u2__abc_52138_new_n14270_; 
wire u2__abc_52138_new_n14271_; 
wire u2__abc_52138_new_n14272_; 
wire u2__abc_52138_new_n14273_; 
wire u2__abc_52138_new_n14274_; 
wire u2__abc_52138_new_n14275_; 
wire u2__abc_52138_new_n14277_; 
wire u2__abc_52138_new_n14278_; 
wire u2__abc_52138_new_n14279_; 
wire u2__abc_52138_new_n14280_; 
wire u2__abc_52138_new_n14281_; 
wire u2__abc_52138_new_n14282_; 
wire u2__abc_52138_new_n14283_; 
wire u2__abc_52138_new_n14285_; 
wire u2__abc_52138_new_n14286_; 
wire u2__abc_52138_new_n14287_; 
wire u2__abc_52138_new_n14288_; 
wire u2__abc_52138_new_n14289_; 
wire u2__abc_52138_new_n14290_; 
wire u2__abc_52138_new_n14291_; 
wire u2__abc_52138_new_n14293_; 
wire u2__abc_52138_new_n14294_; 
wire u2__abc_52138_new_n14295_; 
wire u2__abc_52138_new_n14296_; 
wire u2__abc_52138_new_n14297_; 
wire u2__abc_52138_new_n14298_; 
wire u2__abc_52138_new_n14300_; 
wire u2__abc_52138_new_n14301_; 
wire u2__abc_52138_new_n14302_; 
wire u2__abc_52138_new_n14303_; 
wire u2__abc_52138_new_n14304_; 
wire u2__abc_52138_new_n14305_; 
wire u2__abc_52138_new_n14306_; 
wire u2__abc_52138_new_n14308_; 
wire u2__abc_52138_new_n14309_; 
wire u2__abc_52138_new_n14310_; 
wire u2__abc_52138_new_n14311_; 
wire u2__abc_52138_new_n14312_; 
wire u2__abc_52138_new_n14313_; 
wire u2__abc_52138_new_n14314_; 
wire u2__abc_52138_new_n14316_; 
wire u2__abc_52138_new_n14317_; 
wire u2__abc_52138_new_n14318_; 
wire u2__abc_52138_new_n14319_; 
wire u2__abc_52138_new_n14320_; 
wire u2__abc_52138_new_n14321_; 
wire u2__abc_52138_new_n14322_; 
wire u2__abc_52138_new_n14324_; 
wire u2__abc_52138_new_n14325_; 
wire u2__abc_52138_new_n14326_; 
wire u2__abc_52138_new_n14327_; 
wire u2__abc_52138_new_n14328_; 
wire u2__abc_52138_new_n14329_; 
wire u2__abc_52138_new_n14331_; 
wire u2__abc_52138_new_n14332_; 
wire u2__abc_52138_new_n14333_; 
wire u2__abc_52138_new_n14334_; 
wire u2__abc_52138_new_n14335_; 
wire u2__abc_52138_new_n14336_; 
wire u2__abc_52138_new_n14337_; 
wire u2__abc_52138_new_n14339_; 
wire u2__abc_52138_new_n14340_; 
wire u2__abc_52138_new_n14341_; 
wire u2__abc_52138_new_n14342_; 
wire u2__abc_52138_new_n14343_; 
wire u2__abc_52138_new_n14344_; 
wire u2__abc_52138_new_n14345_; 
wire u2__abc_52138_new_n14347_; 
wire u2__abc_52138_new_n14348_; 
wire u2__abc_52138_new_n14349_; 
wire u2__abc_52138_new_n14350_; 
wire u2__abc_52138_new_n14351_; 
wire u2__abc_52138_new_n14352_; 
wire u2__abc_52138_new_n14353_; 
wire u2__abc_52138_new_n14355_; 
wire u2__abc_52138_new_n14356_; 
wire u2__abc_52138_new_n14357_; 
wire u2__abc_52138_new_n14358_; 
wire u2__abc_52138_new_n14359_; 
wire u2__abc_52138_new_n14360_; 
wire u2__abc_52138_new_n14362_; 
wire u2__abc_52138_new_n14363_; 
wire u2__abc_52138_new_n14364_; 
wire u2__abc_52138_new_n14365_; 
wire u2__abc_52138_new_n14366_; 
wire u2__abc_52138_new_n14367_; 
wire u2__abc_52138_new_n14368_; 
wire u2__abc_52138_new_n14370_; 
wire u2__abc_52138_new_n14371_; 
wire u2__abc_52138_new_n14372_; 
wire u2__abc_52138_new_n14373_; 
wire u2__abc_52138_new_n14374_; 
wire u2__abc_52138_new_n14375_; 
wire u2__abc_52138_new_n14376_; 
wire u2__abc_52138_new_n14378_; 
wire u2__abc_52138_new_n14379_; 
wire u2__abc_52138_new_n14380_; 
wire u2__abc_52138_new_n14381_; 
wire u2__abc_52138_new_n14382_; 
wire u2__abc_52138_new_n14383_; 
wire u2__abc_52138_new_n14384_; 
wire u2__abc_52138_new_n14386_; 
wire u2__abc_52138_new_n14387_; 
wire u2__abc_52138_new_n14388_; 
wire u2__abc_52138_new_n14389_; 
wire u2__abc_52138_new_n14390_; 
wire u2__abc_52138_new_n14391_; 
wire u2__abc_52138_new_n14393_; 
wire u2__abc_52138_new_n14394_; 
wire u2__abc_52138_new_n14395_; 
wire u2__abc_52138_new_n14396_; 
wire u2__abc_52138_new_n14397_; 
wire u2__abc_52138_new_n14398_; 
wire u2__abc_52138_new_n14399_; 
wire u2__abc_52138_new_n14401_; 
wire u2__abc_52138_new_n14402_; 
wire u2__abc_52138_new_n14403_; 
wire u2__abc_52138_new_n14404_; 
wire u2__abc_52138_new_n14405_; 
wire u2__abc_52138_new_n14406_; 
wire u2__abc_52138_new_n14407_; 
wire u2__abc_52138_new_n14409_; 
wire u2__abc_52138_new_n14410_; 
wire u2__abc_52138_new_n14411_; 
wire u2__abc_52138_new_n14412_; 
wire u2__abc_52138_new_n14413_; 
wire u2__abc_52138_new_n14414_; 
wire u2__abc_52138_new_n14415_; 
wire u2__abc_52138_new_n14417_; 
wire u2__abc_52138_new_n14418_; 
wire u2__abc_52138_new_n14419_; 
wire u2__abc_52138_new_n14420_; 
wire u2__abc_52138_new_n14421_; 
wire u2__abc_52138_new_n14422_; 
wire u2__abc_52138_new_n14424_; 
wire u2__abc_52138_new_n14425_; 
wire u2__abc_52138_new_n14426_; 
wire u2__abc_52138_new_n14427_; 
wire u2__abc_52138_new_n14428_; 
wire u2__abc_52138_new_n14429_; 
wire u2__abc_52138_new_n14430_; 
wire u2__abc_52138_new_n14432_; 
wire u2__abc_52138_new_n14433_; 
wire u2__abc_52138_new_n14434_; 
wire u2__abc_52138_new_n14435_; 
wire u2__abc_52138_new_n14436_; 
wire u2__abc_52138_new_n14437_; 
wire u2__abc_52138_new_n14438_; 
wire u2__abc_52138_new_n14440_; 
wire u2__abc_52138_new_n14441_; 
wire u2__abc_52138_new_n14442_; 
wire u2__abc_52138_new_n14443_; 
wire u2__abc_52138_new_n14444_; 
wire u2__abc_52138_new_n14445_; 
wire u2__abc_52138_new_n14446_; 
wire u2__abc_52138_new_n14448_; 
wire u2__abc_52138_new_n14449_; 
wire u2__abc_52138_new_n14450_; 
wire u2__abc_52138_new_n14451_; 
wire u2__abc_52138_new_n14452_; 
wire u2__abc_52138_new_n14453_; 
wire u2__abc_52138_new_n14455_; 
wire u2__abc_52138_new_n14456_; 
wire u2__abc_52138_new_n14457_; 
wire u2__abc_52138_new_n14458_; 
wire u2__abc_52138_new_n14459_; 
wire u2__abc_52138_new_n14460_; 
wire u2__abc_52138_new_n14461_; 
wire u2__abc_52138_new_n14463_; 
wire u2__abc_52138_new_n14464_; 
wire u2__abc_52138_new_n14465_; 
wire u2__abc_52138_new_n14466_; 
wire u2__abc_52138_new_n14467_; 
wire u2__abc_52138_new_n14468_; 
wire u2__abc_52138_new_n14469_; 
wire u2__abc_52138_new_n14471_; 
wire u2__abc_52138_new_n14472_; 
wire u2__abc_52138_new_n14473_; 
wire u2__abc_52138_new_n14474_; 
wire u2__abc_52138_new_n14475_; 
wire u2__abc_52138_new_n14476_; 
wire u2__abc_52138_new_n14477_; 
wire u2__abc_52138_new_n14479_; 
wire u2__abc_52138_new_n14480_; 
wire u2__abc_52138_new_n14481_; 
wire u2__abc_52138_new_n14482_; 
wire u2__abc_52138_new_n14483_; 
wire u2__abc_52138_new_n14484_; 
wire u2__abc_52138_new_n14486_; 
wire u2__abc_52138_new_n14487_; 
wire u2__abc_52138_new_n14488_; 
wire u2__abc_52138_new_n14489_; 
wire u2__abc_52138_new_n14490_; 
wire u2__abc_52138_new_n14491_; 
wire u2__abc_52138_new_n14492_; 
wire u2__abc_52138_new_n14494_; 
wire u2__abc_52138_new_n14495_; 
wire u2__abc_52138_new_n14496_; 
wire u2__abc_52138_new_n14497_; 
wire u2__abc_52138_new_n14498_; 
wire u2__abc_52138_new_n14499_; 
wire u2__abc_52138_new_n14500_; 
wire u2__abc_52138_new_n14502_; 
wire u2__abc_52138_new_n14503_; 
wire u2__abc_52138_new_n14504_; 
wire u2__abc_52138_new_n14505_; 
wire u2__abc_52138_new_n14506_; 
wire u2__abc_52138_new_n14507_; 
wire u2__abc_52138_new_n14508_; 
wire u2__abc_52138_new_n14510_; 
wire u2__abc_52138_new_n14511_; 
wire u2__abc_52138_new_n14512_; 
wire u2__abc_52138_new_n14513_; 
wire u2__abc_52138_new_n14514_; 
wire u2__abc_52138_new_n14515_; 
wire u2__abc_52138_new_n14517_; 
wire u2__abc_52138_new_n14518_; 
wire u2__abc_52138_new_n14519_; 
wire u2__abc_52138_new_n14520_; 
wire u2__abc_52138_new_n14521_; 
wire u2__abc_52138_new_n14522_; 
wire u2__abc_52138_new_n14523_; 
wire u2__abc_52138_new_n14525_; 
wire u2__abc_52138_new_n14526_; 
wire u2__abc_52138_new_n14527_; 
wire u2__abc_52138_new_n14528_; 
wire u2__abc_52138_new_n14529_; 
wire u2__abc_52138_new_n14530_; 
wire u2__abc_52138_new_n14531_; 
wire u2__abc_52138_new_n14533_; 
wire u2__abc_52138_new_n14534_; 
wire u2__abc_52138_new_n14535_; 
wire u2__abc_52138_new_n14536_; 
wire u2__abc_52138_new_n14537_; 
wire u2__abc_52138_new_n14538_; 
wire u2__abc_52138_new_n14539_; 
wire u2__abc_52138_new_n14541_; 
wire u2__abc_52138_new_n14542_; 
wire u2__abc_52138_new_n14543_; 
wire u2__abc_52138_new_n14544_; 
wire u2__abc_52138_new_n14545_; 
wire u2__abc_52138_new_n14546_; 
wire u2__abc_52138_new_n14548_; 
wire u2__abc_52138_new_n14549_; 
wire u2__abc_52138_new_n14550_; 
wire u2__abc_52138_new_n14551_; 
wire u2__abc_52138_new_n14552_; 
wire u2__abc_52138_new_n14553_; 
wire u2__abc_52138_new_n14554_; 
wire u2__abc_52138_new_n14556_; 
wire u2__abc_52138_new_n14557_; 
wire u2__abc_52138_new_n14558_; 
wire u2__abc_52138_new_n14559_; 
wire u2__abc_52138_new_n14560_; 
wire u2__abc_52138_new_n14561_; 
wire u2__abc_52138_new_n14562_; 
wire u2__abc_52138_new_n14564_; 
wire u2__abc_52138_new_n14565_; 
wire u2__abc_52138_new_n14566_; 
wire u2__abc_52138_new_n14567_; 
wire u2__abc_52138_new_n14568_; 
wire u2__abc_52138_new_n14569_; 
wire u2__abc_52138_new_n14570_; 
wire u2__abc_52138_new_n14572_; 
wire u2__abc_52138_new_n14573_; 
wire u2__abc_52138_new_n14574_; 
wire u2__abc_52138_new_n14575_; 
wire u2__abc_52138_new_n14576_; 
wire u2__abc_52138_new_n14577_; 
wire u2__abc_52138_new_n14579_; 
wire u2__abc_52138_new_n14580_; 
wire u2__abc_52138_new_n14581_; 
wire u2__abc_52138_new_n14582_; 
wire u2__abc_52138_new_n14583_; 
wire u2__abc_52138_new_n14584_; 
wire u2__abc_52138_new_n14585_; 
wire u2__abc_52138_new_n14587_; 
wire u2__abc_52138_new_n14588_; 
wire u2__abc_52138_new_n14589_; 
wire u2__abc_52138_new_n14590_; 
wire u2__abc_52138_new_n14591_; 
wire u2__abc_52138_new_n14592_; 
wire u2__abc_52138_new_n14593_; 
wire u2__abc_52138_new_n14595_; 
wire u2__abc_52138_new_n14596_; 
wire u2__abc_52138_new_n14597_; 
wire u2__abc_52138_new_n14598_; 
wire u2__abc_52138_new_n14599_; 
wire u2__abc_52138_new_n14600_; 
wire u2__abc_52138_new_n14601_; 
wire u2__abc_52138_new_n14603_; 
wire u2__abc_52138_new_n14604_; 
wire u2__abc_52138_new_n14605_; 
wire u2__abc_52138_new_n14606_; 
wire u2__abc_52138_new_n14607_; 
wire u2__abc_52138_new_n14608_; 
wire u2__abc_52138_new_n14610_; 
wire u2__abc_52138_new_n14611_; 
wire u2__abc_52138_new_n14612_; 
wire u2__abc_52138_new_n14613_; 
wire u2__abc_52138_new_n14614_; 
wire u2__abc_52138_new_n14615_; 
wire u2__abc_52138_new_n14616_; 
wire u2__abc_52138_new_n14617_; 
wire u2__abc_52138_new_n14619_; 
wire u2__abc_52138_new_n14620_; 
wire u2__abc_52138_new_n14621_; 
wire u2__abc_52138_new_n14622_; 
wire u2__abc_52138_new_n14623_; 
wire u2__abc_52138_new_n14624_; 
wire u2__abc_52138_new_n14625_; 
wire u2__abc_52138_new_n14627_; 
wire u2__abc_52138_new_n14628_; 
wire u2__abc_52138_new_n14629_; 
wire u2__abc_52138_new_n14630_; 
wire u2__abc_52138_new_n14631_; 
wire u2__abc_52138_new_n14632_; 
wire u2__abc_52138_new_n14633_; 
wire u2__abc_52138_new_n14635_; 
wire u2__abc_52138_new_n14636_; 
wire u2__abc_52138_new_n14637_; 
wire u2__abc_52138_new_n14638_; 
wire u2__abc_52138_new_n14639_; 
wire u2__abc_52138_new_n14640_; 
wire u2__abc_52138_new_n14642_; 
wire u2__abc_52138_new_n14643_; 
wire u2__abc_52138_new_n14644_; 
wire u2__abc_52138_new_n14645_; 
wire u2__abc_52138_new_n14646_; 
wire u2__abc_52138_new_n14647_; 
wire u2__abc_52138_new_n14648_; 
wire u2__abc_52138_new_n14650_; 
wire u2__abc_52138_new_n14651_; 
wire u2__abc_52138_new_n14652_; 
wire u2__abc_52138_new_n14653_; 
wire u2__abc_52138_new_n14654_; 
wire u2__abc_52138_new_n14655_; 
wire u2__abc_52138_new_n14656_; 
wire u2__abc_52138_new_n14658_; 
wire u2__abc_52138_new_n14659_; 
wire u2__abc_52138_new_n14660_; 
wire u2__abc_52138_new_n14661_; 
wire u2__abc_52138_new_n14662_; 
wire u2__abc_52138_new_n14663_; 
wire u2__abc_52138_new_n14664_; 
wire u2__abc_52138_new_n14666_; 
wire u2__abc_52138_new_n14667_; 
wire u2__abc_52138_new_n14668_; 
wire u2__abc_52138_new_n14669_; 
wire u2__abc_52138_new_n14670_; 
wire u2__abc_52138_new_n14671_; 
wire u2__abc_52138_new_n14673_; 
wire u2__abc_52138_new_n14674_; 
wire u2__abc_52138_new_n14675_; 
wire u2__abc_52138_new_n14676_; 
wire u2__abc_52138_new_n14677_; 
wire u2__abc_52138_new_n14678_; 
wire u2__abc_52138_new_n14679_; 
wire u2__abc_52138_new_n14681_; 
wire u2__abc_52138_new_n14682_; 
wire u2__abc_52138_new_n14683_; 
wire u2__abc_52138_new_n14684_; 
wire u2__abc_52138_new_n14685_; 
wire u2__abc_52138_new_n14686_; 
wire u2__abc_52138_new_n14687_; 
wire u2__abc_52138_new_n14689_; 
wire u2__abc_52138_new_n14690_; 
wire u2__abc_52138_new_n14691_; 
wire u2__abc_52138_new_n14692_; 
wire u2__abc_52138_new_n14693_; 
wire u2__abc_52138_new_n14694_; 
wire u2__abc_52138_new_n14695_; 
wire u2__abc_52138_new_n14697_; 
wire u2__abc_52138_new_n14698_; 
wire u2__abc_52138_new_n14699_; 
wire u2__abc_52138_new_n14700_; 
wire u2__abc_52138_new_n14701_; 
wire u2__abc_52138_new_n14702_; 
wire u2__abc_52138_new_n14704_; 
wire u2__abc_52138_new_n14705_; 
wire u2__abc_52138_new_n14706_; 
wire u2__abc_52138_new_n14707_; 
wire u2__abc_52138_new_n14708_; 
wire u2__abc_52138_new_n14709_; 
wire u2__abc_52138_new_n14710_; 
wire u2__abc_52138_new_n14712_; 
wire u2__abc_52138_new_n14713_; 
wire u2__abc_52138_new_n14714_; 
wire u2__abc_52138_new_n14715_; 
wire u2__abc_52138_new_n14716_; 
wire u2__abc_52138_new_n14717_; 
wire u2__abc_52138_new_n14718_; 
wire u2__abc_52138_new_n14720_; 
wire u2__abc_52138_new_n14721_; 
wire u2__abc_52138_new_n14722_; 
wire u2__abc_52138_new_n14723_; 
wire u2__abc_52138_new_n14724_; 
wire u2__abc_52138_new_n14725_; 
wire u2__abc_52138_new_n14726_; 
wire u2__abc_52138_new_n14728_; 
wire u2__abc_52138_new_n14729_; 
wire u2__abc_52138_new_n14730_; 
wire u2__abc_52138_new_n14731_; 
wire u2__abc_52138_new_n14732_; 
wire u2__abc_52138_new_n14733_; 
wire u2__abc_52138_new_n14735_; 
wire u2__abc_52138_new_n14736_; 
wire u2__abc_52138_new_n14737_; 
wire u2__abc_52138_new_n14738_; 
wire u2__abc_52138_new_n14739_; 
wire u2__abc_52138_new_n14740_; 
wire u2__abc_52138_new_n14741_; 
wire u2__abc_52138_new_n14743_; 
wire u2__abc_52138_new_n14744_; 
wire u2__abc_52138_new_n14745_; 
wire u2__abc_52138_new_n14746_; 
wire u2__abc_52138_new_n14747_; 
wire u2__abc_52138_new_n14748_; 
wire u2__abc_52138_new_n14749_; 
wire u2__abc_52138_new_n14751_; 
wire u2__abc_52138_new_n14752_; 
wire u2__abc_52138_new_n14753_; 
wire u2__abc_52138_new_n14754_; 
wire u2__abc_52138_new_n14755_; 
wire u2__abc_52138_new_n14756_; 
wire u2__abc_52138_new_n14757_; 
wire u2__abc_52138_new_n14759_; 
wire u2__abc_52138_new_n14760_; 
wire u2__abc_52138_new_n14761_; 
wire u2__abc_52138_new_n14762_; 
wire u2__abc_52138_new_n14763_; 
wire u2__abc_52138_new_n14764_; 
wire u2__abc_52138_new_n14766_; 
wire u2__abc_52138_new_n14767_; 
wire u2__abc_52138_new_n14768_; 
wire u2__abc_52138_new_n14769_; 
wire u2__abc_52138_new_n14770_; 
wire u2__abc_52138_new_n14771_; 
wire u2__abc_52138_new_n14772_; 
wire u2__abc_52138_new_n14774_; 
wire u2__abc_52138_new_n14775_; 
wire u2__abc_52138_new_n14776_; 
wire u2__abc_52138_new_n14777_; 
wire u2__abc_52138_new_n14778_; 
wire u2__abc_52138_new_n14779_; 
wire u2__abc_52138_new_n14780_; 
wire u2__abc_52138_new_n14782_; 
wire u2__abc_52138_new_n14783_; 
wire u2__abc_52138_new_n14784_; 
wire u2__abc_52138_new_n14785_; 
wire u2__abc_52138_new_n14786_; 
wire u2__abc_52138_new_n14787_; 
wire u2__abc_52138_new_n14788_; 
wire u2__abc_52138_new_n14790_; 
wire u2__abc_52138_new_n14791_; 
wire u2__abc_52138_new_n14792_; 
wire u2__abc_52138_new_n14793_; 
wire u2__abc_52138_new_n14794_; 
wire u2__abc_52138_new_n14795_; 
wire u2__abc_52138_new_n14797_; 
wire u2__abc_52138_new_n14798_; 
wire u2__abc_52138_new_n14799_; 
wire u2__abc_52138_new_n14800_; 
wire u2__abc_52138_new_n14801_; 
wire u2__abc_52138_new_n14802_; 
wire u2__abc_52138_new_n14803_; 
wire u2__abc_52138_new_n14805_; 
wire u2__abc_52138_new_n14806_; 
wire u2__abc_52138_new_n14807_; 
wire u2__abc_52138_new_n14808_; 
wire u2__abc_52138_new_n14809_; 
wire u2__abc_52138_new_n14810_; 
wire u2__abc_52138_new_n14811_; 
wire u2__abc_52138_new_n14813_; 
wire u2__abc_52138_new_n14814_; 
wire u2__abc_52138_new_n14815_; 
wire u2__abc_52138_new_n14816_; 
wire u2__abc_52138_new_n14817_; 
wire u2__abc_52138_new_n14818_; 
wire u2__abc_52138_new_n14819_; 
wire u2__abc_52138_new_n14821_; 
wire u2__abc_52138_new_n14822_; 
wire u2__abc_52138_new_n14823_; 
wire u2__abc_52138_new_n14824_; 
wire u2__abc_52138_new_n14825_; 
wire u2__abc_52138_new_n14826_; 
wire u2__abc_52138_new_n14828_; 
wire u2__abc_52138_new_n14829_; 
wire u2__abc_52138_new_n14830_; 
wire u2__abc_52138_new_n14831_; 
wire u2__abc_52138_new_n14832_; 
wire u2__abc_52138_new_n14833_; 
wire u2__abc_52138_new_n14834_; 
wire u2__abc_52138_new_n14836_; 
wire u2__abc_52138_new_n14837_; 
wire u2__abc_52138_new_n14838_; 
wire u2__abc_52138_new_n14839_; 
wire u2__abc_52138_new_n14840_; 
wire u2__abc_52138_new_n14841_; 
wire u2__abc_52138_new_n14842_; 
wire u2__abc_52138_new_n14844_; 
wire u2__abc_52138_new_n14845_; 
wire u2__abc_52138_new_n14846_; 
wire u2__abc_52138_new_n14847_; 
wire u2__abc_52138_new_n14848_; 
wire u2__abc_52138_new_n14849_; 
wire u2__abc_52138_new_n14850_; 
wire u2__abc_52138_new_n14852_; 
wire u2__abc_52138_new_n14853_; 
wire u2__abc_52138_new_n14854_; 
wire u2__abc_52138_new_n14855_; 
wire u2__abc_52138_new_n14856_; 
wire u2__abc_52138_new_n14857_; 
wire u2__abc_52138_new_n14859_; 
wire u2__abc_52138_new_n14860_; 
wire u2__abc_52138_new_n14861_; 
wire u2__abc_52138_new_n14862_; 
wire u2__abc_52138_new_n14863_; 
wire u2__abc_52138_new_n14864_; 
wire u2__abc_52138_new_n14865_; 
wire u2__abc_52138_new_n14867_; 
wire u2__abc_52138_new_n14868_; 
wire u2__abc_52138_new_n14869_; 
wire u2__abc_52138_new_n14870_; 
wire u2__abc_52138_new_n14871_; 
wire u2__abc_52138_new_n14872_; 
wire u2__abc_52138_new_n14873_; 
wire u2__abc_52138_new_n14875_; 
wire u2__abc_52138_new_n14876_; 
wire u2__abc_52138_new_n14877_; 
wire u2__abc_52138_new_n14878_; 
wire u2__abc_52138_new_n14879_; 
wire u2__abc_52138_new_n14880_; 
wire u2__abc_52138_new_n14881_; 
wire u2__abc_52138_new_n14883_; 
wire u2__abc_52138_new_n14884_; 
wire u2__abc_52138_new_n14885_; 
wire u2__abc_52138_new_n14886_; 
wire u2__abc_52138_new_n14887_; 
wire u2__abc_52138_new_n14888_; 
wire u2__abc_52138_new_n14890_; 
wire u2__abc_52138_new_n14891_; 
wire u2__abc_52138_new_n14892_; 
wire u2__abc_52138_new_n14893_; 
wire u2__abc_52138_new_n14894_; 
wire u2__abc_52138_new_n14895_; 
wire u2__abc_52138_new_n14896_; 
wire u2__abc_52138_new_n14898_; 
wire u2__abc_52138_new_n14899_; 
wire u2__abc_52138_new_n14900_; 
wire u2__abc_52138_new_n14901_; 
wire u2__abc_52138_new_n14902_; 
wire u2__abc_52138_new_n14903_; 
wire u2__abc_52138_new_n14904_; 
wire u2__abc_52138_new_n14906_; 
wire u2__abc_52138_new_n14907_; 
wire u2__abc_52138_new_n14908_; 
wire u2__abc_52138_new_n14909_; 
wire u2__abc_52138_new_n14910_; 
wire u2__abc_52138_new_n14911_; 
wire u2__abc_52138_new_n14912_; 
wire u2__abc_52138_new_n14914_; 
wire u2__abc_52138_new_n14915_; 
wire u2__abc_52138_new_n14916_; 
wire u2__abc_52138_new_n14917_; 
wire u2__abc_52138_new_n14918_; 
wire u2__abc_52138_new_n14919_; 
wire u2__abc_52138_new_n14921_; 
wire u2__abc_52138_new_n14922_; 
wire u2__abc_52138_new_n14923_; 
wire u2__abc_52138_new_n14924_; 
wire u2__abc_52138_new_n14925_; 
wire u2__abc_52138_new_n14926_; 
wire u2__abc_52138_new_n14927_; 
wire u2__abc_52138_new_n14929_; 
wire u2__abc_52138_new_n14930_; 
wire u2__abc_52138_new_n14931_; 
wire u2__abc_52138_new_n14932_; 
wire u2__abc_52138_new_n14933_; 
wire u2__abc_52138_new_n14934_; 
wire u2__abc_52138_new_n14935_; 
wire u2__abc_52138_new_n14937_; 
wire u2__abc_52138_new_n14938_; 
wire u2__abc_52138_new_n14939_; 
wire u2__abc_52138_new_n14940_; 
wire u2__abc_52138_new_n14941_; 
wire u2__abc_52138_new_n14942_; 
wire u2__abc_52138_new_n14943_; 
wire u2__abc_52138_new_n14945_; 
wire u2__abc_52138_new_n14946_; 
wire u2__abc_52138_new_n14947_; 
wire u2__abc_52138_new_n14948_; 
wire u2__abc_52138_new_n14949_; 
wire u2__abc_52138_new_n14950_; 
wire u2__abc_52138_new_n14952_; 
wire u2__abc_52138_new_n14953_; 
wire u2__abc_52138_new_n14954_; 
wire u2__abc_52138_new_n14955_; 
wire u2__abc_52138_new_n14956_; 
wire u2__abc_52138_new_n14957_; 
wire u2__abc_52138_new_n14958_; 
wire u2__abc_52138_new_n14960_; 
wire u2__abc_52138_new_n14961_; 
wire u2__abc_52138_new_n14962_; 
wire u2__abc_52138_new_n14963_; 
wire u2__abc_52138_new_n14964_; 
wire u2__abc_52138_new_n14965_; 
wire u2__abc_52138_new_n14966_; 
wire u2__abc_52138_new_n14968_; 
wire u2__abc_52138_new_n14969_; 
wire u2__abc_52138_new_n14970_; 
wire u2__abc_52138_new_n14971_; 
wire u2__abc_52138_new_n14972_; 
wire u2__abc_52138_new_n14973_; 
wire u2__abc_52138_new_n14974_; 
wire u2__abc_52138_new_n14976_; 
wire u2__abc_52138_new_n14977_; 
wire u2__abc_52138_new_n14978_; 
wire u2__abc_52138_new_n14979_; 
wire u2__abc_52138_new_n14980_; 
wire u2__abc_52138_new_n14981_; 
wire u2__abc_52138_new_n14983_; 
wire u2__abc_52138_new_n14984_; 
wire u2__abc_52138_new_n14985_; 
wire u2__abc_52138_new_n14986_; 
wire u2__abc_52138_new_n14987_; 
wire u2__abc_52138_new_n14988_; 
wire u2__abc_52138_new_n14989_; 
wire u2__abc_52138_new_n14991_; 
wire u2__abc_52138_new_n14992_; 
wire u2__abc_52138_new_n14993_; 
wire u2__abc_52138_new_n14994_; 
wire u2__abc_52138_new_n14995_; 
wire u2__abc_52138_new_n14996_; 
wire u2__abc_52138_new_n14997_; 
wire u2__abc_52138_new_n14999_; 
wire u2__abc_52138_new_n15000_; 
wire u2__abc_52138_new_n15001_; 
wire u2__abc_52138_new_n15002_; 
wire u2__abc_52138_new_n15003_; 
wire u2__abc_52138_new_n15004_; 
wire u2__abc_52138_new_n15005_; 
wire u2__abc_52138_new_n15007_; 
wire u2__abc_52138_new_n15008_; 
wire u2__abc_52138_new_n15009_; 
wire u2__abc_52138_new_n15010_; 
wire u2__abc_52138_new_n15011_; 
wire u2__abc_52138_new_n15012_; 
wire u2__abc_52138_new_n15014_; 
wire u2__abc_52138_new_n15015_; 
wire u2__abc_52138_new_n15016_; 
wire u2__abc_52138_new_n15017_; 
wire u2__abc_52138_new_n15018_; 
wire u2__abc_52138_new_n15019_; 
wire u2__abc_52138_new_n15020_; 
wire u2__abc_52138_new_n15022_; 
wire u2__abc_52138_new_n15023_; 
wire u2__abc_52138_new_n15024_; 
wire u2__abc_52138_new_n15025_; 
wire u2__abc_52138_new_n15026_; 
wire u2__abc_52138_new_n15027_; 
wire u2__abc_52138_new_n15028_; 
wire u2__abc_52138_new_n15030_; 
wire u2__abc_52138_new_n15031_; 
wire u2__abc_52138_new_n15032_; 
wire u2__abc_52138_new_n15033_; 
wire u2__abc_52138_new_n15034_; 
wire u2__abc_52138_new_n15035_; 
wire u2__abc_52138_new_n15036_; 
wire u2__abc_52138_new_n15038_; 
wire u2__abc_52138_new_n15039_; 
wire u2__abc_52138_new_n15040_; 
wire u2__abc_52138_new_n15041_; 
wire u2__abc_52138_new_n15042_; 
wire u2__abc_52138_new_n15043_; 
wire u2__abc_52138_new_n15045_; 
wire u2__abc_52138_new_n15046_; 
wire u2__abc_52138_new_n15047_; 
wire u2__abc_52138_new_n15048_; 
wire u2__abc_52138_new_n15049_; 
wire u2__abc_52138_new_n15050_; 
wire u2__abc_52138_new_n15051_; 
wire u2__abc_52138_new_n15053_; 
wire u2__abc_52138_new_n15054_; 
wire u2__abc_52138_new_n15055_; 
wire u2__abc_52138_new_n15056_; 
wire u2__abc_52138_new_n15057_; 
wire u2__abc_52138_new_n15058_; 
wire u2__abc_52138_new_n15059_; 
wire u2__abc_52138_new_n15061_; 
wire u2__abc_52138_new_n15062_; 
wire u2__abc_52138_new_n15063_; 
wire u2__abc_52138_new_n15064_; 
wire u2__abc_52138_new_n15065_; 
wire u2__abc_52138_new_n15066_; 
wire u2__abc_52138_new_n15067_; 
wire u2__abc_52138_new_n15069_; 
wire u2__abc_52138_new_n15070_; 
wire u2__abc_52138_new_n15071_; 
wire u2__abc_52138_new_n15072_; 
wire u2__abc_52138_new_n15073_; 
wire u2__abc_52138_new_n15074_; 
wire u2__abc_52138_new_n15076_; 
wire u2__abc_52138_new_n15077_; 
wire u2__abc_52138_new_n15078_; 
wire u2__abc_52138_new_n15079_; 
wire u2__abc_52138_new_n15080_; 
wire u2__abc_52138_new_n15081_; 
wire u2__abc_52138_new_n15082_; 
wire u2__abc_52138_new_n15084_; 
wire u2__abc_52138_new_n15085_; 
wire u2__abc_52138_new_n15086_; 
wire u2__abc_52138_new_n15087_; 
wire u2__abc_52138_new_n15088_; 
wire u2__abc_52138_new_n15089_; 
wire u2__abc_52138_new_n15090_; 
wire u2__abc_52138_new_n15092_; 
wire u2__abc_52138_new_n15093_; 
wire u2__abc_52138_new_n15094_; 
wire u2__abc_52138_new_n15095_; 
wire u2__abc_52138_new_n15096_; 
wire u2__abc_52138_new_n15097_; 
wire u2__abc_52138_new_n15098_; 
wire u2__abc_52138_new_n15100_; 
wire u2__abc_52138_new_n15101_; 
wire u2__abc_52138_new_n15102_; 
wire u2__abc_52138_new_n15103_; 
wire u2__abc_52138_new_n15104_; 
wire u2__abc_52138_new_n15105_; 
wire u2__abc_52138_new_n15107_; 
wire u2__abc_52138_new_n15108_; 
wire u2__abc_52138_new_n15109_; 
wire u2__abc_52138_new_n15110_; 
wire u2__abc_52138_new_n15111_; 
wire u2__abc_52138_new_n15112_; 
wire u2__abc_52138_new_n15113_; 
wire u2__abc_52138_new_n15115_; 
wire u2__abc_52138_new_n15116_; 
wire u2__abc_52138_new_n15117_; 
wire u2__abc_52138_new_n15118_; 
wire u2__abc_52138_new_n15119_; 
wire u2__abc_52138_new_n15120_; 
wire u2__abc_52138_new_n15121_; 
wire u2__abc_52138_new_n15123_; 
wire u2__abc_52138_new_n15124_; 
wire u2__abc_52138_new_n15125_; 
wire u2__abc_52138_new_n15126_; 
wire u2__abc_52138_new_n15127_; 
wire u2__abc_52138_new_n15128_; 
wire u2__abc_52138_new_n15129_; 
wire u2__abc_52138_new_n15131_; 
wire u2__abc_52138_new_n15132_; 
wire u2__abc_52138_new_n15133_; 
wire u2__abc_52138_new_n15134_; 
wire u2__abc_52138_new_n15135_; 
wire u2__abc_52138_new_n15136_; 
wire u2__abc_52138_new_n15138_; 
wire u2__abc_52138_new_n15139_; 
wire u2__abc_52138_new_n15140_; 
wire u2__abc_52138_new_n15141_; 
wire u2__abc_52138_new_n15142_; 
wire u2__abc_52138_new_n15143_; 
wire u2__abc_52138_new_n15144_; 
wire u2__abc_52138_new_n15146_; 
wire u2__abc_52138_new_n15147_; 
wire u2__abc_52138_new_n15148_; 
wire u2__abc_52138_new_n15149_; 
wire u2__abc_52138_new_n15150_; 
wire u2__abc_52138_new_n15151_; 
wire u2__abc_52138_new_n15152_; 
wire u2__abc_52138_new_n15154_; 
wire u2__abc_52138_new_n15155_; 
wire u2__abc_52138_new_n15156_; 
wire u2__abc_52138_new_n15157_; 
wire u2__abc_52138_new_n15158_; 
wire u2__abc_52138_new_n15159_; 
wire u2__abc_52138_new_n15160_; 
wire u2__abc_52138_new_n15162_; 
wire u2__abc_52138_new_n15163_; 
wire u2__abc_52138_new_n15164_; 
wire u2__abc_52138_new_n15165_; 
wire u2__abc_52138_new_n15166_; 
wire u2__abc_52138_new_n15167_; 
wire u2__abc_52138_new_n15169_; 
wire u2__abc_52138_new_n15170_; 
wire u2__abc_52138_new_n15171_; 
wire u2__abc_52138_new_n15172_; 
wire u2__abc_52138_new_n15173_; 
wire u2__abc_52138_new_n15174_; 
wire u2__abc_52138_new_n15175_; 
wire u2__abc_52138_new_n15177_; 
wire u2__abc_52138_new_n15178_; 
wire u2__abc_52138_new_n15179_; 
wire u2__abc_52138_new_n15180_; 
wire u2__abc_52138_new_n15181_; 
wire u2__abc_52138_new_n15182_; 
wire u2__abc_52138_new_n15183_; 
wire u2__abc_52138_new_n15185_; 
wire u2__abc_52138_new_n15186_; 
wire u2__abc_52138_new_n15187_; 
wire u2__abc_52138_new_n15188_; 
wire u2__abc_52138_new_n15189_; 
wire u2__abc_52138_new_n15190_; 
wire u2__abc_52138_new_n15191_; 
wire u2__abc_52138_new_n15193_; 
wire u2__abc_52138_new_n15194_; 
wire u2__abc_52138_new_n15195_; 
wire u2__abc_52138_new_n15196_; 
wire u2__abc_52138_new_n15197_; 
wire u2__abc_52138_new_n15198_; 
wire u2__abc_52138_new_n15200_; 
wire u2__abc_52138_new_n15201_; 
wire u2__abc_52138_new_n15202_; 
wire u2__abc_52138_new_n15203_; 
wire u2__abc_52138_new_n15204_; 
wire u2__abc_52138_new_n15205_; 
wire u2__abc_52138_new_n15206_; 
wire u2__abc_52138_new_n15208_; 
wire u2__abc_52138_new_n15209_; 
wire u2__abc_52138_new_n15210_; 
wire u2__abc_52138_new_n15211_; 
wire u2__abc_52138_new_n15212_; 
wire u2__abc_52138_new_n15213_; 
wire u2__abc_52138_new_n15214_; 
wire u2__abc_52138_new_n15216_; 
wire u2__abc_52138_new_n15217_; 
wire u2__abc_52138_new_n15218_; 
wire u2__abc_52138_new_n15219_; 
wire u2__abc_52138_new_n15220_; 
wire u2__abc_52138_new_n15221_; 
wire u2__abc_52138_new_n15222_; 
wire u2__abc_52138_new_n15224_; 
wire u2__abc_52138_new_n15225_; 
wire u2__abc_52138_new_n15226_; 
wire u2__abc_52138_new_n15227_; 
wire u2__abc_52138_new_n15228_; 
wire u2__abc_52138_new_n15229_; 
wire u2__abc_52138_new_n15231_; 
wire u2__abc_52138_new_n15232_; 
wire u2__abc_52138_new_n15233_; 
wire u2__abc_52138_new_n15234_; 
wire u2__abc_52138_new_n15235_; 
wire u2__abc_52138_new_n15236_; 
wire u2__abc_52138_new_n15237_; 
wire u2__abc_52138_new_n15239_; 
wire u2__abc_52138_new_n15240_; 
wire u2__abc_52138_new_n15241_; 
wire u2__abc_52138_new_n15242_; 
wire u2__abc_52138_new_n15243_; 
wire u2__abc_52138_new_n15244_; 
wire u2__abc_52138_new_n15245_; 
wire u2__abc_52138_new_n15247_; 
wire u2__abc_52138_new_n15248_; 
wire u2__abc_52138_new_n15249_; 
wire u2__abc_52138_new_n15250_; 
wire u2__abc_52138_new_n15251_; 
wire u2__abc_52138_new_n15252_; 
wire u2__abc_52138_new_n15253_; 
wire u2__abc_52138_new_n15255_; 
wire u2__abc_52138_new_n15256_; 
wire u2__abc_52138_new_n15257_; 
wire u2__abc_52138_new_n15258_; 
wire u2__abc_52138_new_n15259_; 
wire u2__abc_52138_new_n15260_; 
wire u2__abc_52138_new_n15262_; 
wire u2__abc_52138_new_n15263_; 
wire u2__abc_52138_new_n15264_; 
wire u2__abc_52138_new_n15265_; 
wire u2__abc_52138_new_n15266_; 
wire u2__abc_52138_new_n15267_; 
wire u2__abc_52138_new_n15268_; 
wire u2__abc_52138_new_n15270_; 
wire u2__abc_52138_new_n15271_; 
wire u2__abc_52138_new_n15272_; 
wire u2__abc_52138_new_n15273_; 
wire u2__abc_52138_new_n15274_; 
wire u2__abc_52138_new_n15275_; 
wire u2__abc_52138_new_n15276_; 
wire u2__abc_52138_new_n15278_; 
wire u2__abc_52138_new_n15279_; 
wire u2__abc_52138_new_n15280_; 
wire u2__abc_52138_new_n15281_; 
wire u2__abc_52138_new_n15282_; 
wire u2__abc_52138_new_n15283_; 
wire u2__abc_52138_new_n15284_; 
wire u2__abc_52138_new_n15286_; 
wire u2__abc_52138_new_n15287_; 
wire u2__abc_52138_new_n15288_; 
wire u2__abc_52138_new_n15289_; 
wire u2__abc_52138_new_n15290_; 
wire u2__abc_52138_new_n15291_; 
wire u2__abc_52138_new_n15293_; 
wire u2__abc_52138_new_n15294_; 
wire u2__abc_52138_new_n15295_; 
wire u2__abc_52138_new_n15296_; 
wire u2__abc_52138_new_n15297_; 
wire u2__abc_52138_new_n15298_; 
wire u2__abc_52138_new_n15299_; 
wire u2__abc_52138_new_n15301_; 
wire u2__abc_52138_new_n15302_; 
wire u2__abc_52138_new_n15303_; 
wire u2__abc_52138_new_n15304_; 
wire u2__abc_52138_new_n15305_; 
wire u2__abc_52138_new_n15306_; 
wire u2__abc_52138_new_n15307_; 
wire u2__abc_52138_new_n15309_; 
wire u2__abc_52138_new_n15310_; 
wire u2__abc_52138_new_n15311_; 
wire u2__abc_52138_new_n15312_; 
wire u2__abc_52138_new_n15313_; 
wire u2__abc_52138_new_n15314_; 
wire u2__abc_52138_new_n15315_; 
wire u2__abc_52138_new_n15317_; 
wire u2__abc_52138_new_n15318_; 
wire u2__abc_52138_new_n15319_; 
wire u2__abc_52138_new_n15320_; 
wire u2__abc_52138_new_n15321_; 
wire u2__abc_52138_new_n15322_; 
wire u2__abc_52138_new_n15324_; 
wire u2__abc_52138_new_n15325_; 
wire u2__abc_52138_new_n15326_; 
wire u2__abc_52138_new_n15327_; 
wire u2__abc_52138_new_n15328_; 
wire u2__abc_52138_new_n15329_; 
wire u2__abc_52138_new_n15330_; 
wire u2__abc_52138_new_n15332_; 
wire u2__abc_52138_new_n15333_; 
wire u2__abc_52138_new_n15334_; 
wire u2__abc_52138_new_n15335_; 
wire u2__abc_52138_new_n15336_; 
wire u2__abc_52138_new_n15337_; 
wire u2__abc_52138_new_n15338_; 
wire u2__abc_52138_new_n15340_; 
wire u2__abc_52138_new_n15341_; 
wire u2__abc_52138_new_n15342_; 
wire u2__abc_52138_new_n15343_; 
wire u2__abc_52138_new_n15344_; 
wire u2__abc_52138_new_n15345_; 
wire u2__abc_52138_new_n15346_; 
wire u2__abc_52138_new_n15348_; 
wire u2__abc_52138_new_n15349_; 
wire u2__abc_52138_new_n15350_; 
wire u2__abc_52138_new_n15351_; 
wire u2__abc_52138_new_n15352_; 
wire u2__abc_52138_new_n15353_; 
wire u2__abc_52138_new_n15355_; 
wire u2__abc_52138_new_n15356_; 
wire u2__abc_52138_new_n15357_; 
wire u2__abc_52138_new_n15358_; 
wire u2__abc_52138_new_n15359_; 
wire u2__abc_52138_new_n15360_; 
wire u2__abc_52138_new_n15361_; 
wire u2__abc_52138_new_n15363_; 
wire u2__abc_52138_new_n15364_; 
wire u2__abc_52138_new_n15365_; 
wire u2__abc_52138_new_n15366_; 
wire u2__abc_52138_new_n15367_; 
wire u2__abc_52138_new_n15368_; 
wire u2__abc_52138_new_n15369_; 
wire u2__abc_52138_new_n15371_; 
wire u2__abc_52138_new_n15372_; 
wire u2__abc_52138_new_n15373_; 
wire u2__abc_52138_new_n15374_; 
wire u2__abc_52138_new_n15375_; 
wire u2__abc_52138_new_n15376_; 
wire u2__abc_52138_new_n15377_; 
wire u2__abc_52138_new_n15379_; 
wire u2__abc_52138_new_n15380_; 
wire u2__abc_52138_new_n15381_; 
wire u2__abc_52138_new_n15382_; 
wire u2__abc_52138_new_n15383_; 
wire u2__abc_52138_new_n15384_; 
wire u2__abc_52138_new_n15386_; 
wire u2__abc_52138_new_n15387_; 
wire u2__abc_52138_new_n15388_; 
wire u2__abc_52138_new_n15389_; 
wire u2__abc_52138_new_n15390_; 
wire u2__abc_52138_new_n15391_; 
wire u2__abc_52138_new_n15392_; 
wire u2__abc_52138_new_n15394_; 
wire u2__abc_52138_new_n15395_; 
wire u2__abc_52138_new_n15396_; 
wire u2__abc_52138_new_n15397_; 
wire u2__abc_52138_new_n15398_; 
wire u2__abc_52138_new_n15399_; 
wire u2__abc_52138_new_n15400_; 
wire u2__abc_52138_new_n15402_; 
wire u2__abc_52138_new_n15403_; 
wire u2__abc_52138_new_n15404_; 
wire u2__abc_52138_new_n15405_; 
wire u2__abc_52138_new_n15406_; 
wire u2__abc_52138_new_n15407_; 
wire u2__abc_52138_new_n15408_; 
wire u2__abc_52138_new_n15410_; 
wire u2__abc_52138_new_n15411_; 
wire u2__abc_52138_new_n15412_; 
wire u2__abc_52138_new_n15413_; 
wire u2__abc_52138_new_n15414_; 
wire u2__abc_52138_new_n15415_; 
wire u2__abc_52138_new_n15417_; 
wire u2__abc_52138_new_n15418_; 
wire u2__abc_52138_new_n15419_; 
wire u2__abc_52138_new_n15420_; 
wire u2__abc_52138_new_n15421_; 
wire u2__abc_52138_new_n15422_; 
wire u2__abc_52138_new_n15423_; 
wire u2__abc_52138_new_n15425_; 
wire u2__abc_52138_new_n15426_; 
wire u2__abc_52138_new_n15427_; 
wire u2__abc_52138_new_n15428_; 
wire u2__abc_52138_new_n15429_; 
wire u2__abc_52138_new_n15430_; 
wire u2__abc_52138_new_n15431_; 
wire u2__abc_52138_new_n15433_; 
wire u2__abc_52138_new_n15434_; 
wire u2__abc_52138_new_n15435_; 
wire u2__abc_52138_new_n15436_; 
wire u2__abc_52138_new_n15437_; 
wire u2__abc_52138_new_n15438_; 
wire u2__abc_52138_new_n15439_; 
wire u2__abc_52138_new_n15441_; 
wire u2__abc_52138_new_n15442_; 
wire u2__abc_52138_new_n15443_; 
wire u2__abc_52138_new_n15444_; 
wire u2__abc_52138_new_n15445_; 
wire u2__abc_52138_new_n15446_; 
wire u2__abc_52138_new_n15448_; 
wire u2__abc_52138_new_n15449_; 
wire u2__abc_52138_new_n15450_; 
wire u2__abc_52138_new_n15451_; 
wire u2__abc_52138_new_n15452_; 
wire u2__abc_52138_new_n15453_; 
wire u2__abc_52138_new_n15454_; 
wire u2__abc_52138_new_n15456_; 
wire u2__abc_52138_new_n15457_; 
wire u2__abc_52138_new_n15458_; 
wire u2__abc_52138_new_n15459_; 
wire u2__abc_52138_new_n15460_; 
wire u2__abc_52138_new_n15461_; 
wire u2__abc_52138_new_n15462_; 
wire u2__abc_52138_new_n15464_; 
wire u2__abc_52138_new_n15465_; 
wire u2__abc_52138_new_n15466_; 
wire u2__abc_52138_new_n15467_; 
wire u2__abc_52138_new_n15468_; 
wire u2__abc_52138_new_n15469_; 
wire u2__abc_52138_new_n15470_; 
wire u2__abc_52138_new_n15472_; 
wire u2__abc_52138_new_n15473_; 
wire u2__abc_52138_new_n15474_; 
wire u2__abc_52138_new_n15475_; 
wire u2__abc_52138_new_n15476_; 
wire u2__abc_52138_new_n15477_; 
wire u2__abc_52138_new_n15479_; 
wire u2__abc_52138_new_n15480_; 
wire u2__abc_52138_new_n15481_; 
wire u2__abc_52138_new_n15482_; 
wire u2__abc_52138_new_n15483_; 
wire u2__abc_52138_new_n15484_; 
wire u2__abc_52138_new_n15485_; 
wire u2__abc_52138_new_n15486_; 
wire u2__abc_52138_new_n15488_; 
wire u2__abc_52138_new_n15489_; 
wire u2__abc_52138_new_n15490_; 
wire u2__abc_52138_new_n15491_; 
wire u2__abc_52138_new_n15492_; 
wire u2__abc_52138_new_n15493_; 
wire u2__abc_52138_new_n15494_; 
wire u2__abc_52138_new_n15496_; 
wire u2__abc_52138_new_n15497_; 
wire u2__abc_52138_new_n15498_; 
wire u2__abc_52138_new_n15499_; 
wire u2__abc_52138_new_n15500_; 
wire u2__abc_52138_new_n15501_; 
wire u2__abc_52138_new_n15502_; 
wire u2__abc_52138_new_n15504_; 
wire u2__abc_52138_new_n15505_; 
wire u2__abc_52138_new_n15506_; 
wire u2__abc_52138_new_n15507_; 
wire u2__abc_52138_new_n15508_; 
wire u2__abc_52138_new_n15509_; 
wire u2__abc_52138_new_n15511_; 
wire u2__abc_52138_new_n15512_; 
wire u2__abc_52138_new_n15513_; 
wire u2__abc_52138_new_n15514_; 
wire u2__abc_52138_new_n15515_; 
wire u2__abc_52138_new_n15516_; 
wire u2__abc_52138_new_n15517_; 
wire u2__abc_52138_new_n15519_; 
wire u2__abc_52138_new_n15520_; 
wire u2__abc_52138_new_n15521_; 
wire u2__abc_52138_new_n15522_; 
wire u2__abc_52138_new_n15523_; 
wire u2__abc_52138_new_n15524_; 
wire u2__abc_52138_new_n15525_; 
wire u2__abc_52138_new_n15527_; 
wire u2__abc_52138_new_n15528_; 
wire u2__abc_52138_new_n15529_; 
wire u2__abc_52138_new_n15530_; 
wire u2__abc_52138_new_n15531_; 
wire u2__abc_52138_new_n15532_; 
wire u2__abc_52138_new_n15533_; 
wire u2__abc_52138_new_n15535_; 
wire u2__abc_52138_new_n15536_; 
wire u2__abc_52138_new_n15537_; 
wire u2__abc_52138_new_n15538_; 
wire u2__abc_52138_new_n15539_; 
wire u2__abc_52138_new_n15540_; 
wire u2__abc_52138_new_n15542_; 
wire u2__abc_52138_new_n15543_; 
wire u2__abc_52138_new_n15544_; 
wire u2__abc_52138_new_n15545_; 
wire u2__abc_52138_new_n15546_; 
wire u2__abc_52138_new_n15547_; 
wire u2__abc_52138_new_n15548_; 
wire u2__abc_52138_new_n15550_; 
wire u2__abc_52138_new_n15551_; 
wire u2__abc_52138_new_n15552_; 
wire u2__abc_52138_new_n15553_; 
wire u2__abc_52138_new_n15554_; 
wire u2__abc_52138_new_n15555_; 
wire u2__abc_52138_new_n15556_; 
wire u2__abc_52138_new_n15558_; 
wire u2__abc_52138_new_n15559_; 
wire u2__abc_52138_new_n15560_; 
wire u2__abc_52138_new_n15561_; 
wire u2__abc_52138_new_n15562_; 
wire u2__abc_52138_new_n15563_; 
wire u2__abc_52138_new_n15564_; 
wire u2__abc_52138_new_n15566_; 
wire u2__abc_52138_new_n15567_; 
wire u2__abc_52138_new_n15568_; 
wire u2__abc_52138_new_n15569_; 
wire u2__abc_52138_new_n15570_; 
wire u2__abc_52138_new_n15571_; 
wire u2__abc_52138_new_n15573_; 
wire u2__abc_52138_new_n15574_; 
wire u2__abc_52138_new_n15575_; 
wire u2__abc_52138_new_n15576_; 
wire u2__abc_52138_new_n15577_; 
wire u2__abc_52138_new_n15578_; 
wire u2__abc_52138_new_n15579_; 
wire u2__abc_52138_new_n15581_; 
wire u2__abc_52138_new_n15582_; 
wire u2__abc_52138_new_n15583_; 
wire u2__abc_52138_new_n15584_; 
wire u2__abc_52138_new_n15585_; 
wire u2__abc_52138_new_n15586_; 
wire u2__abc_52138_new_n15587_; 
wire u2__abc_52138_new_n15589_; 
wire u2__abc_52138_new_n15590_; 
wire u2__abc_52138_new_n15591_; 
wire u2__abc_52138_new_n15592_; 
wire u2__abc_52138_new_n15593_; 
wire u2__abc_52138_new_n15594_; 
wire u2__abc_52138_new_n15595_; 
wire u2__abc_52138_new_n15597_; 
wire u2__abc_52138_new_n15598_; 
wire u2__abc_52138_new_n15599_; 
wire u2__abc_52138_new_n15600_; 
wire u2__abc_52138_new_n15601_; 
wire u2__abc_52138_new_n15602_; 
wire u2__abc_52138_new_n15604_; 
wire u2__abc_52138_new_n15605_; 
wire u2__abc_52138_new_n15606_; 
wire u2__abc_52138_new_n15607_; 
wire u2__abc_52138_new_n15608_; 
wire u2__abc_52138_new_n15609_; 
wire u2__abc_52138_new_n15610_; 
wire u2__abc_52138_new_n15612_; 
wire u2__abc_52138_new_n15613_; 
wire u2__abc_52138_new_n15614_; 
wire u2__abc_52138_new_n15615_; 
wire u2__abc_52138_new_n15616_; 
wire u2__abc_52138_new_n15617_; 
wire u2__abc_52138_new_n15618_; 
wire u2__abc_52138_new_n15620_; 
wire u2__abc_52138_new_n15621_; 
wire u2__abc_52138_new_n15622_; 
wire u2__abc_52138_new_n15623_; 
wire u2__abc_52138_new_n15624_; 
wire u2__abc_52138_new_n15625_; 
wire u2__abc_52138_new_n15626_; 
wire u2__abc_52138_new_n15628_; 
wire u2__abc_52138_new_n15629_; 
wire u2__abc_52138_new_n15630_; 
wire u2__abc_52138_new_n15631_; 
wire u2__abc_52138_new_n15632_; 
wire u2__abc_52138_new_n15633_; 
wire u2__abc_52138_new_n15635_; 
wire u2__abc_52138_new_n15636_; 
wire u2__abc_52138_new_n15637_; 
wire u2__abc_52138_new_n15638_; 
wire u2__abc_52138_new_n15639_; 
wire u2__abc_52138_new_n15640_; 
wire u2__abc_52138_new_n15641_; 
wire u2__abc_52138_new_n15642_; 
wire u2__abc_52138_new_n15644_; 
wire u2__abc_52138_new_n15645_; 
wire u2__abc_52138_new_n15646_; 
wire u2__abc_52138_new_n15647_; 
wire u2__abc_52138_new_n15648_; 
wire u2__abc_52138_new_n15649_; 
wire u2__abc_52138_new_n15650_; 
wire u2__abc_52138_new_n15652_; 
wire u2__abc_52138_new_n15653_; 
wire u2__abc_52138_new_n15654_; 
wire u2__abc_52138_new_n15655_; 
wire u2__abc_52138_new_n15656_; 
wire u2__abc_52138_new_n15657_; 
wire u2__abc_52138_new_n15658_; 
wire u2__abc_52138_new_n15660_; 
wire u2__abc_52138_new_n15661_; 
wire u2__abc_52138_new_n15662_; 
wire u2__abc_52138_new_n15663_; 
wire u2__abc_52138_new_n15664_; 
wire u2__abc_52138_new_n15665_; 
wire u2__abc_52138_new_n15667_; 
wire u2__abc_52138_new_n15668_; 
wire u2__abc_52138_new_n15669_; 
wire u2__abc_52138_new_n15670_; 
wire u2__abc_52138_new_n15671_; 
wire u2__abc_52138_new_n15672_; 
wire u2__abc_52138_new_n15673_; 
wire u2__abc_52138_new_n15674_; 
wire u2__abc_52138_new_n15676_; 
wire u2__abc_52138_new_n15677_; 
wire u2__abc_52138_new_n15678_; 
wire u2__abc_52138_new_n15679_; 
wire u2__abc_52138_new_n15680_; 
wire u2__abc_52138_new_n15681_; 
wire u2__abc_52138_new_n15682_; 
wire u2__abc_52138_new_n15684_; 
wire u2__abc_52138_new_n15685_; 
wire u2__abc_52138_new_n15686_; 
wire u2__abc_52138_new_n15687_; 
wire u2__abc_52138_new_n15688_; 
wire u2__abc_52138_new_n15689_; 
wire u2__abc_52138_new_n15690_; 
wire u2__abc_52138_new_n15692_; 
wire u2__abc_52138_new_n15693_; 
wire u2__abc_52138_new_n15694_; 
wire u2__abc_52138_new_n15695_; 
wire u2__abc_52138_new_n15696_; 
wire u2__abc_52138_new_n15697_; 
wire u2__abc_52138_new_n15699_; 
wire u2__abc_52138_new_n15700_; 
wire u2__abc_52138_new_n15701_; 
wire u2__abc_52138_new_n15702_; 
wire u2__abc_52138_new_n15703_; 
wire u2__abc_52138_new_n15704_; 
wire u2__abc_52138_new_n15705_; 
wire u2__abc_52138_new_n15707_; 
wire u2__abc_52138_new_n15708_; 
wire u2__abc_52138_new_n15709_; 
wire u2__abc_52138_new_n15710_; 
wire u2__abc_52138_new_n15711_; 
wire u2__abc_52138_new_n15712_; 
wire u2__abc_52138_new_n15713_; 
wire u2__abc_52138_new_n15715_; 
wire u2__abc_52138_new_n15716_; 
wire u2__abc_52138_new_n15717_; 
wire u2__abc_52138_new_n15718_; 
wire u2__abc_52138_new_n15719_; 
wire u2__abc_52138_new_n15720_; 
wire u2__abc_52138_new_n15721_; 
wire u2__abc_52138_new_n15723_; 
wire u2__abc_52138_new_n15724_; 
wire u2__abc_52138_new_n15725_; 
wire u2__abc_52138_new_n15726_; 
wire u2__abc_52138_new_n15727_; 
wire u2__abc_52138_new_n15728_; 
wire u2__abc_52138_new_n15730_; 
wire u2__abc_52138_new_n15731_; 
wire u2__abc_52138_new_n15732_; 
wire u2__abc_52138_new_n15733_; 
wire u2__abc_52138_new_n15734_; 
wire u2__abc_52138_new_n15735_; 
wire u2__abc_52138_new_n15736_; 
wire u2__abc_52138_new_n15738_; 
wire u2__abc_52138_new_n15739_; 
wire u2__abc_52138_new_n15740_; 
wire u2__abc_52138_new_n15741_; 
wire u2__abc_52138_new_n15742_; 
wire u2__abc_52138_new_n15743_; 
wire u2__abc_52138_new_n15744_; 
wire u2__abc_52138_new_n15746_; 
wire u2__abc_52138_new_n15747_; 
wire u2__abc_52138_new_n15748_; 
wire u2__abc_52138_new_n15749_; 
wire u2__abc_52138_new_n15750_; 
wire u2__abc_52138_new_n15751_; 
wire u2__abc_52138_new_n15752_; 
wire u2__abc_52138_new_n15754_; 
wire u2__abc_52138_new_n15755_; 
wire u2__abc_52138_new_n15756_; 
wire u2__abc_52138_new_n15757_; 
wire u2__abc_52138_new_n15758_; 
wire u2__abc_52138_new_n15759_; 
wire u2__abc_52138_new_n15761_; 
wire u2__abc_52138_new_n15762_; 
wire u2__abc_52138_new_n15763_; 
wire u2__abc_52138_new_n15764_; 
wire u2__abc_52138_new_n15765_; 
wire u2__abc_52138_new_n15766_; 
wire u2__abc_52138_new_n15767_; 
wire u2__abc_52138_new_n15769_; 
wire u2__abc_52138_new_n15770_; 
wire u2__abc_52138_new_n15771_; 
wire u2__abc_52138_new_n15772_; 
wire u2__abc_52138_new_n15773_; 
wire u2__abc_52138_new_n15774_; 
wire u2__abc_52138_new_n15775_; 
wire u2__abc_52138_new_n15777_; 
wire u2__abc_52138_new_n15778_; 
wire u2__abc_52138_new_n15779_; 
wire u2__abc_52138_new_n15780_; 
wire u2__abc_52138_new_n15781_; 
wire u2__abc_52138_new_n15782_; 
wire u2__abc_52138_new_n15783_; 
wire u2__abc_52138_new_n15785_; 
wire u2__abc_52138_new_n15786_; 
wire u2__abc_52138_new_n15787_; 
wire u2__abc_52138_new_n15788_; 
wire u2__abc_52138_new_n15789_; 
wire u2__abc_52138_new_n15790_; 
wire u2__abc_52138_new_n15792_; 
wire u2__abc_52138_new_n15793_; 
wire u2__abc_52138_new_n15794_; 
wire u2__abc_52138_new_n15795_; 
wire u2__abc_52138_new_n15796_; 
wire u2__abc_52138_new_n15797_; 
wire u2__abc_52138_new_n15798_; 
wire u2__abc_52138_new_n15800_; 
wire u2__abc_52138_new_n15801_; 
wire u2__abc_52138_new_n15802_; 
wire u2__abc_52138_new_n15803_; 
wire u2__abc_52138_new_n15804_; 
wire u2__abc_52138_new_n15805_; 
wire u2__abc_52138_new_n15806_; 
wire u2__abc_52138_new_n15808_; 
wire u2__abc_52138_new_n15809_; 
wire u2__abc_52138_new_n15810_; 
wire u2__abc_52138_new_n15811_; 
wire u2__abc_52138_new_n15812_; 
wire u2__abc_52138_new_n15813_; 
wire u2__abc_52138_new_n15814_; 
wire u2__abc_52138_new_n15816_; 
wire u2__abc_52138_new_n15817_; 
wire u2__abc_52138_new_n15818_; 
wire u2__abc_52138_new_n15819_; 
wire u2__abc_52138_new_n15820_; 
wire u2__abc_52138_new_n15821_; 
wire u2__abc_52138_new_n15823_; 
wire u2__abc_52138_new_n15824_; 
wire u2__abc_52138_new_n15825_; 
wire u2__abc_52138_new_n15826_; 
wire u2__abc_52138_new_n15827_; 
wire u2__abc_52138_new_n15828_; 
wire u2__abc_52138_new_n15829_; 
wire u2__abc_52138_new_n15831_; 
wire u2__abc_52138_new_n15832_; 
wire u2__abc_52138_new_n15833_; 
wire u2__abc_52138_new_n15834_; 
wire u2__abc_52138_new_n15835_; 
wire u2__abc_52138_new_n15836_; 
wire u2__abc_52138_new_n15837_; 
wire u2__abc_52138_new_n15839_; 
wire u2__abc_52138_new_n15840_; 
wire u2__abc_52138_new_n15841_; 
wire u2__abc_52138_new_n15842_; 
wire u2__abc_52138_new_n15843_; 
wire u2__abc_52138_new_n15844_; 
wire u2__abc_52138_new_n15845_; 
wire u2__abc_52138_new_n15847_; 
wire u2__abc_52138_new_n15848_; 
wire u2__abc_52138_new_n15849_; 
wire u2__abc_52138_new_n15850_; 
wire u2__abc_52138_new_n15851_; 
wire u2__abc_52138_new_n15852_; 
wire u2__abc_52138_new_n15854_; 
wire u2__abc_52138_new_n15855_; 
wire u2__abc_52138_new_n15856_; 
wire u2__abc_52138_new_n15857_; 
wire u2__abc_52138_new_n15858_; 
wire u2__abc_52138_new_n15859_; 
wire u2__abc_52138_new_n15860_; 
wire u2__abc_52138_new_n15862_; 
wire u2__abc_52138_new_n15863_; 
wire u2__abc_52138_new_n15864_; 
wire u2__abc_52138_new_n15865_; 
wire u2__abc_52138_new_n15866_; 
wire u2__abc_52138_new_n15867_; 
wire u2__abc_52138_new_n15868_; 
wire u2__abc_52138_new_n15870_; 
wire u2__abc_52138_new_n15871_; 
wire u2__abc_52138_new_n15872_; 
wire u2__abc_52138_new_n15873_; 
wire u2__abc_52138_new_n15874_; 
wire u2__abc_52138_new_n15875_; 
wire u2__abc_52138_new_n15876_; 
wire u2__abc_52138_new_n15878_; 
wire u2__abc_52138_new_n15879_; 
wire u2__abc_52138_new_n15880_; 
wire u2__abc_52138_new_n15881_; 
wire u2__abc_52138_new_n15882_; 
wire u2__abc_52138_new_n15883_; 
wire u2__abc_52138_new_n15885_; 
wire u2__abc_52138_new_n15886_; 
wire u2__abc_52138_new_n15887_; 
wire u2__abc_52138_new_n15888_; 
wire u2__abc_52138_new_n15889_; 
wire u2__abc_52138_new_n15890_; 
wire u2__abc_52138_new_n15891_; 
wire u2__abc_52138_new_n15893_; 
wire u2__abc_52138_new_n15894_; 
wire u2__abc_52138_new_n15895_; 
wire u2__abc_52138_new_n15896_; 
wire u2__abc_52138_new_n15897_; 
wire u2__abc_52138_new_n15898_; 
wire u2__abc_52138_new_n15899_; 
wire u2__abc_52138_new_n15901_; 
wire u2__abc_52138_new_n15902_; 
wire u2__abc_52138_new_n15903_; 
wire u2__abc_52138_new_n15904_; 
wire u2__abc_52138_new_n15905_; 
wire u2__abc_52138_new_n15906_; 
wire u2__abc_52138_new_n15907_; 
wire u2__abc_52138_new_n15909_; 
wire u2__abc_52138_new_n15910_; 
wire u2__abc_52138_new_n15911_; 
wire u2__abc_52138_new_n15912_; 
wire u2__abc_52138_new_n15913_; 
wire u2__abc_52138_new_n15914_; 
wire u2__abc_52138_new_n15915_; 
wire u2__abc_52138_new_n15917_; 
wire u2__abc_52138_new_n15918_; 
wire u2__abc_52138_new_n15919_; 
wire u2__abc_52138_new_n15920_; 
wire u2__abc_52138_new_n15921_; 
wire u2__abc_52138_new_n15922_; 
wire u2__abc_52138_new_n15923_; 
wire u2__abc_52138_new_n15925_; 
wire u2__abc_52138_new_n15926_; 
wire u2__abc_52138_new_n15927_; 
wire u2__abc_52138_new_n15928_; 
wire u2__abc_52138_new_n15929_; 
wire u2__abc_52138_new_n15930_; 
wire u2__abc_52138_new_n15931_; 
wire u2__abc_52138_new_n15933_; 
wire u2__abc_52138_new_n15934_; 
wire u2__abc_52138_new_n15935_; 
wire u2__abc_52138_new_n15936_; 
wire u2__abc_52138_new_n15937_; 
wire u2__abc_52138_new_n15938_; 
wire u2__abc_52138_new_n15939_; 
wire u2__abc_52138_new_n15941_; 
wire u2__abc_52138_new_n15942_; 
wire u2__abc_52138_new_n15943_; 
wire u2__abc_52138_new_n15944_; 
wire u2__abc_52138_new_n15945_; 
wire u2__abc_52138_new_n15946_; 
wire u2__abc_52138_new_n15948_; 
wire u2__abc_52138_new_n15949_; 
wire u2__abc_52138_new_n15950_; 
wire u2__abc_52138_new_n15951_; 
wire u2__abc_52138_new_n15952_; 
wire u2__abc_52138_new_n15953_; 
wire u2__abc_52138_new_n15954_; 
wire u2__abc_52138_new_n15956_; 
wire u2__abc_52138_new_n15957_; 
wire u2__abc_52138_new_n15958_; 
wire u2__abc_52138_new_n15959_; 
wire u2__abc_52138_new_n15960_; 
wire u2__abc_52138_new_n15961_; 
wire u2__abc_52138_new_n15962_; 
wire u2__abc_52138_new_n15964_; 
wire u2__abc_52138_new_n15965_; 
wire u2__abc_52138_new_n15966_; 
wire u2__abc_52138_new_n15967_; 
wire u2__abc_52138_new_n15968_; 
wire u2__abc_52138_new_n15969_; 
wire u2__abc_52138_new_n15970_; 
wire u2__abc_52138_new_n15972_; 
wire u2__abc_52138_new_n15973_; 
wire u2__abc_52138_new_n15974_; 
wire u2__abc_52138_new_n15975_; 
wire u2__abc_52138_new_n15976_; 
wire u2__abc_52138_new_n15977_; 
wire u2__abc_52138_new_n15979_; 
wire u2__abc_52138_new_n15980_; 
wire u2__abc_52138_new_n15981_; 
wire u2__abc_52138_new_n15982_; 
wire u2__abc_52138_new_n15983_; 
wire u2__abc_52138_new_n15984_; 
wire u2__abc_52138_new_n15985_; 
wire u2__abc_52138_new_n15987_; 
wire u2__abc_52138_new_n15988_; 
wire u2__abc_52138_new_n15989_; 
wire u2__abc_52138_new_n15990_; 
wire u2__abc_52138_new_n15991_; 
wire u2__abc_52138_new_n15992_; 
wire u2__abc_52138_new_n15993_; 
wire u2__abc_52138_new_n15995_; 
wire u2__abc_52138_new_n15996_; 
wire u2__abc_52138_new_n15997_; 
wire u2__abc_52138_new_n15998_; 
wire u2__abc_52138_new_n15999_; 
wire u2__abc_52138_new_n16000_; 
wire u2__abc_52138_new_n16001_; 
wire u2__abc_52138_new_n16003_; 
wire u2__abc_52138_new_n16004_; 
wire u2__abc_52138_new_n16005_; 
wire u2__abc_52138_new_n16006_; 
wire u2__abc_52138_new_n16007_; 
wire u2__abc_52138_new_n16008_; 
wire u2__abc_52138_new_n16010_; 
wire u2__abc_52138_new_n16011_; 
wire u2__abc_52138_new_n16012_; 
wire u2__abc_52138_new_n16013_; 
wire u2__abc_52138_new_n16014_; 
wire u2__abc_52138_new_n16015_; 
wire u2__abc_52138_new_n16016_; 
wire u2__abc_52138_new_n16018_; 
wire u2__abc_52138_new_n16019_; 
wire u2__abc_52138_new_n16020_; 
wire u2__abc_52138_new_n16021_; 
wire u2__abc_52138_new_n16022_; 
wire u2__abc_52138_new_n16023_; 
wire u2__abc_52138_new_n16024_; 
wire u2__abc_52138_new_n16026_; 
wire u2__abc_52138_new_n16027_; 
wire u2__abc_52138_new_n16028_; 
wire u2__abc_52138_new_n16029_; 
wire u2__abc_52138_new_n16030_; 
wire u2__abc_52138_new_n16031_; 
wire u2__abc_52138_new_n16032_; 
wire u2__abc_52138_new_n16034_; 
wire u2__abc_52138_new_n16035_; 
wire u2__abc_52138_new_n16036_; 
wire u2__abc_52138_new_n16037_; 
wire u2__abc_52138_new_n16038_; 
wire u2__abc_52138_new_n16039_; 
wire u2__abc_52138_new_n16041_; 
wire u2__abc_52138_new_n16042_; 
wire u2__abc_52138_new_n16043_; 
wire u2__abc_52138_new_n16044_; 
wire u2__abc_52138_new_n16045_; 
wire u2__abc_52138_new_n16046_; 
wire u2__abc_52138_new_n16047_; 
wire u2__abc_52138_new_n16049_; 
wire u2__abc_52138_new_n16050_; 
wire u2__abc_52138_new_n16051_; 
wire u2__abc_52138_new_n16052_; 
wire u2__abc_52138_new_n16053_; 
wire u2__abc_52138_new_n16054_; 
wire u2__abc_52138_new_n16055_; 
wire u2__abc_52138_new_n16057_; 
wire u2__abc_52138_new_n16058_; 
wire u2__abc_52138_new_n16059_; 
wire u2__abc_52138_new_n16060_; 
wire u2__abc_52138_new_n16061_; 
wire u2__abc_52138_new_n16062_; 
wire u2__abc_52138_new_n16063_; 
wire u2__abc_52138_new_n16065_; 
wire u2__abc_52138_new_n16066_; 
wire u2__abc_52138_new_n16067_; 
wire u2__abc_52138_new_n16068_; 
wire u2__abc_52138_new_n16069_; 
wire u2__abc_52138_new_n16070_; 
wire u2__abc_52138_new_n16072_; 
wire u2__abc_52138_new_n16073_; 
wire u2__abc_52138_new_n16074_; 
wire u2__abc_52138_new_n16075_; 
wire u2__abc_52138_new_n16076_; 
wire u2__abc_52138_new_n16077_; 
wire u2__abc_52138_new_n16078_; 
wire u2__abc_52138_new_n16079_; 
wire u2__abc_52138_new_n16081_; 
wire u2__abc_52138_new_n16082_; 
wire u2__abc_52138_new_n16083_; 
wire u2__abc_52138_new_n16084_; 
wire u2__abc_52138_new_n16085_; 
wire u2__abc_52138_new_n16086_; 
wire u2__abc_52138_new_n16087_; 
wire u2__abc_52138_new_n16088_; 
wire u2__abc_52138_new_n16090_; 
wire u2__abc_52138_new_n16091_; 
wire u2__abc_52138_new_n16092_; 
wire u2__abc_52138_new_n16093_; 
wire u2__abc_52138_new_n16094_; 
wire u2__abc_52138_new_n16095_; 
wire u2__abc_52138_new_n16096_; 
wire u2__abc_52138_new_n16098_; 
wire u2__abc_52138_new_n16099_; 
wire u2__abc_52138_new_n16100_; 
wire u2__abc_52138_new_n16101_; 
wire u2__abc_52138_new_n16102_; 
wire u2__abc_52138_new_n16103_; 
wire u2__abc_52138_new_n16105_; 
wire u2__abc_52138_new_n16106_; 
wire u2__abc_52138_new_n16107_; 
wire u2__abc_52138_new_n16108_; 
wire u2__abc_52138_new_n16109_; 
wire u2__abc_52138_new_n16110_; 
wire u2__abc_52138_new_n16111_; 
wire u2__abc_52138_new_n16112_; 
wire u2__abc_52138_new_n16114_; 
wire u2__abc_52138_new_n16115_; 
wire u2__abc_52138_new_n16116_; 
wire u2__abc_52138_new_n16117_; 
wire u2__abc_52138_new_n16118_; 
wire u2__abc_52138_new_n16119_; 
wire u2__abc_52138_new_n16120_; 
wire u2__abc_52138_new_n16122_; 
wire u2__abc_52138_new_n16123_; 
wire u2__abc_52138_new_n16124_; 
wire u2__abc_52138_new_n16125_; 
wire u2__abc_52138_new_n16126_; 
wire u2__abc_52138_new_n16127_; 
wire u2__abc_52138_new_n16128_; 
wire u2__abc_52138_new_n16130_; 
wire u2__abc_52138_new_n16131_; 
wire u2__abc_52138_new_n16132_; 
wire u2__abc_52138_new_n16133_; 
wire u2__abc_52138_new_n16134_; 
wire u2__abc_52138_new_n16135_; 
wire u2__abc_52138_new_n16137_; 
wire u2__abc_52138_new_n16138_; 
wire u2__abc_52138_new_n16139_; 
wire u2__abc_52138_new_n16140_; 
wire u2__abc_52138_new_n16141_; 
wire u2__abc_52138_new_n16142_; 
wire u2__abc_52138_new_n16143_; 
wire u2__abc_52138_new_n16145_; 
wire u2__abc_52138_new_n16146_; 
wire u2__abc_52138_new_n16147_; 
wire u2__abc_52138_new_n16148_; 
wire u2__abc_52138_new_n16149_; 
wire u2__abc_52138_new_n16150_; 
wire u2__abc_52138_new_n16151_; 
wire u2__abc_52138_new_n16153_; 
wire u2__abc_52138_new_n16154_; 
wire u2__abc_52138_new_n16155_; 
wire u2__abc_52138_new_n16156_; 
wire u2__abc_52138_new_n16157_; 
wire u2__abc_52138_new_n16158_; 
wire u2__abc_52138_new_n16159_; 
wire u2__abc_52138_new_n16161_; 
wire u2__abc_52138_new_n16162_; 
wire u2__abc_52138_new_n16163_; 
wire u2__abc_52138_new_n16164_; 
wire u2__abc_52138_new_n16165_; 
wire u2__abc_52138_new_n16166_; 
wire u2__abc_52138_new_n16168_; 
wire u2__abc_52138_new_n16169_; 
wire u2__abc_52138_new_n16170_; 
wire u2__abc_52138_new_n16171_; 
wire u2__abc_52138_new_n16172_; 
wire u2__abc_52138_new_n16173_; 
wire u2__abc_52138_new_n16174_; 
wire u2__abc_52138_new_n16176_; 
wire u2__abc_52138_new_n16177_; 
wire u2__abc_52138_new_n16178_; 
wire u2__abc_52138_new_n16179_; 
wire u2__abc_52138_new_n16180_; 
wire u2__abc_52138_new_n16181_; 
wire u2__abc_52138_new_n16182_; 
wire u2__abc_52138_new_n16184_; 
wire u2__abc_52138_new_n16185_; 
wire u2__abc_52138_new_n16186_; 
wire u2__abc_52138_new_n16187_; 
wire u2__abc_52138_new_n16188_; 
wire u2__abc_52138_new_n16189_; 
wire u2__abc_52138_new_n16190_; 
wire u2__abc_52138_new_n16192_; 
wire u2__abc_52138_new_n16193_; 
wire u2__abc_52138_new_n16194_; 
wire u2__abc_52138_new_n16195_; 
wire u2__abc_52138_new_n16196_; 
wire u2__abc_52138_new_n16197_; 
wire u2__abc_52138_new_n16199_; 
wire u2__abc_52138_new_n16200_; 
wire u2__abc_52138_new_n16201_; 
wire u2__abc_52138_new_n16202_; 
wire u2__abc_52138_new_n16203_; 
wire u2__abc_52138_new_n16204_; 
wire u2__abc_52138_new_n16205_; 
wire u2__abc_52138_new_n16207_; 
wire u2__abc_52138_new_n16208_; 
wire u2__abc_52138_new_n16209_; 
wire u2__abc_52138_new_n16210_; 
wire u2__abc_52138_new_n16211_; 
wire u2__abc_52138_new_n16212_; 
wire u2__abc_52138_new_n16213_; 
wire u2__abc_52138_new_n16215_; 
wire u2__abc_52138_new_n16216_; 
wire u2__abc_52138_new_n16217_; 
wire u2__abc_52138_new_n16218_; 
wire u2__abc_52138_new_n16219_; 
wire u2__abc_52138_new_n16220_; 
wire u2__abc_52138_new_n16221_; 
wire u2__abc_52138_new_n16223_; 
wire u2__abc_52138_new_n16224_; 
wire u2__abc_52138_new_n16225_; 
wire u2__abc_52138_new_n16226_; 
wire u2__abc_52138_new_n16227_; 
wire u2__abc_52138_new_n16228_; 
wire u2__abc_52138_new_n16230_; 
wire u2__abc_52138_new_n16231_; 
wire u2__abc_52138_new_n16232_; 
wire u2__abc_52138_new_n16233_; 
wire u2__abc_52138_new_n16234_; 
wire u2__abc_52138_new_n16235_; 
wire u2__abc_52138_new_n16236_; 
wire u2__abc_52138_new_n16238_; 
wire u2__abc_52138_new_n16239_; 
wire u2__abc_52138_new_n16240_; 
wire u2__abc_52138_new_n16241_; 
wire u2__abc_52138_new_n16242_; 
wire u2__abc_52138_new_n16243_; 
wire u2__abc_52138_new_n16244_; 
wire u2__abc_52138_new_n16246_; 
wire u2__abc_52138_new_n16247_; 
wire u2__abc_52138_new_n16248_; 
wire u2__abc_52138_new_n16249_; 
wire u2__abc_52138_new_n16250_; 
wire u2__abc_52138_new_n16251_; 
wire u2__abc_52138_new_n16252_; 
wire u2__abc_52138_new_n16254_; 
wire u2__abc_52138_new_n16255_; 
wire u2__abc_52138_new_n16256_; 
wire u2__abc_52138_new_n16257_; 
wire u2__abc_52138_new_n16258_; 
wire u2__abc_52138_new_n16259_; 
wire u2__abc_52138_new_n16261_; 
wire u2__abc_52138_new_n16262_; 
wire u2__abc_52138_new_n16263_; 
wire u2__abc_52138_new_n16264_; 
wire u2__abc_52138_new_n16265_; 
wire u2__abc_52138_new_n16266_; 
wire u2__abc_52138_new_n16267_; 
wire u2__abc_52138_new_n16269_; 
wire u2__abc_52138_new_n16270_; 
wire u2__abc_52138_new_n16271_; 
wire u2__abc_52138_new_n16272_; 
wire u2__abc_52138_new_n16273_; 
wire u2__abc_52138_new_n16274_; 
wire u2__abc_52138_new_n16275_; 
wire u2__abc_52138_new_n16277_; 
wire u2__abc_52138_new_n16278_; 
wire u2__abc_52138_new_n16279_; 
wire u2__abc_52138_new_n16280_; 
wire u2__abc_52138_new_n16281_; 
wire u2__abc_52138_new_n16282_; 
wire u2__abc_52138_new_n16283_; 
wire u2__abc_52138_new_n16285_; 
wire u2__abc_52138_new_n16286_; 
wire u2__abc_52138_new_n16287_; 
wire u2__abc_52138_new_n16288_; 
wire u2__abc_52138_new_n16289_; 
wire u2__abc_52138_new_n16290_; 
wire u2__abc_52138_new_n16292_; 
wire u2__abc_52138_new_n16293_; 
wire u2__abc_52138_new_n16294_; 
wire u2__abc_52138_new_n16295_; 
wire u2__abc_52138_new_n16296_; 
wire u2__abc_52138_new_n16297_; 
wire u2__abc_52138_new_n16298_; 
wire u2__abc_52138_new_n16300_; 
wire u2__abc_52138_new_n16301_; 
wire u2__abc_52138_new_n16302_; 
wire u2__abc_52138_new_n16303_; 
wire u2__abc_52138_new_n16304_; 
wire u2__abc_52138_new_n16305_; 
wire u2__abc_52138_new_n16306_; 
wire u2__abc_52138_new_n16308_; 
wire u2__abc_52138_new_n16309_; 
wire u2__abc_52138_new_n16310_; 
wire u2__abc_52138_new_n16311_; 
wire u2__abc_52138_new_n16312_; 
wire u2__abc_52138_new_n16313_; 
wire u2__abc_52138_new_n16314_; 
wire u2__abc_52138_new_n16316_; 
wire u2__abc_52138_new_n16317_; 
wire u2__abc_52138_new_n16318_; 
wire u2__abc_52138_new_n16319_; 
wire u2__abc_52138_new_n16320_; 
wire u2__abc_52138_new_n16321_; 
wire u2__abc_52138_new_n16323_; 
wire u2__abc_52138_new_n16324_; 
wire u2__abc_52138_new_n16325_; 
wire u2__abc_52138_new_n16326_; 
wire u2__abc_52138_new_n16327_; 
wire u2__abc_52138_new_n16328_; 
wire u2__abc_52138_new_n16329_; 
wire u2__abc_52138_new_n16331_; 
wire u2__abc_52138_new_n16332_; 
wire u2__abc_52138_new_n16333_; 
wire u2__abc_52138_new_n16334_; 
wire u2__abc_52138_new_n16335_; 
wire u2__abc_52138_new_n16336_; 
wire u2__abc_52138_new_n16337_; 
wire u2__abc_52138_new_n16339_; 
wire u2__abc_52138_new_n16340_; 
wire u2__abc_52138_new_n16341_; 
wire u2__abc_52138_new_n16342_; 
wire u2__abc_52138_new_n16343_; 
wire u2__abc_52138_new_n16344_; 
wire u2__abc_52138_new_n16345_; 
wire u2__abc_52138_new_n16347_; 
wire u2__abc_52138_new_n16348_; 
wire u2__abc_52138_new_n16349_; 
wire u2__abc_52138_new_n16350_; 
wire u2__abc_52138_new_n16351_; 
wire u2__abc_52138_new_n16352_; 
wire u2__abc_52138_new_n16354_; 
wire u2__abc_52138_new_n16355_; 
wire u2__abc_52138_new_n16356_; 
wire u2__abc_52138_new_n16357_; 
wire u2__abc_52138_new_n16358_; 
wire u2__abc_52138_new_n16359_; 
wire u2__abc_52138_new_n16360_; 
wire u2__abc_52138_new_n16362_; 
wire u2__abc_52138_new_n16363_; 
wire u2__abc_52138_new_n16364_; 
wire u2__abc_52138_new_n16365_; 
wire u2__abc_52138_new_n16366_; 
wire u2__abc_52138_new_n16367_; 
wire u2__abc_52138_new_n16368_; 
wire u2__abc_52138_new_n16370_; 
wire u2__abc_52138_new_n16371_; 
wire u2__abc_52138_new_n16372_; 
wire u2__abc_52138_new_n16373_; 
wire u2__abc_52138_new_n16374_; 
wire u2__abc_52138_new_n16375_; 
wire u2__abc_52138_new_n16376_; 
wire u2__abc_52138_new_n16378_; 
wire u2__abc_52138_new_n16379_; 
wire u2__abc_52138_new_n16380_; 
wire u2__abc_52138_new_n16381_; 
wire u2__abc_52138_new_n16382_; 
wire u2__abc_52138_new_n16383_; 
wire u2__abc_52138_new_n16385_; 
wire u2__abc_52138_new_n16386_; 
wire u2__abc_52138_new_n16387_; 
wire u2__abc_52138_new_n16388_; 
wire u2__abc_52138_new_n16389_; 
wire u2__abc_52138_new_n16390_; 
wire u2__abc_52138_new_n16391_; 
wire u2__abc_52138_new_n16393_; 
wire u2__abc_52138_new_n16394_; 
wire u2__abc_52138_new_n16395_; 
wire u2__abc_52138_new_n16396_; 
wire u2__abc_52138_new_n16397_; 
wire u2__abc_52138_new_n16398_; 
wire u2__abc_52138_new_n16399_; 
wire u2__abc_52138_new_n16401_; 
wire u2__abc_52138_new_n16402_; 
wire u2__abc_52138_new_n16403_; 
wire u2__abc_52138_new_n16404_; 
wire u2__abc_52138_new_n16405_; 
wire u2__abc_52138_new_n16406_; 
wire u2__abc_52138_new_n16407_; 
wire u2__abc_52138_new_n16409_; 
wire u2__abc_52138_new_n16410_; 
wire u2__abc_52138_new_n16411_; 
wire u2__abc_52138_new_n16412_; 
wire u2__abc_52138_new_n16413_; 
wire u2__abc_52138_new_n16414_; 
wire u2__abc_52138_new_n16416_; 
wire u2__abc_52138_new_n16417_; 
wire u2__abc_52138_new_n16418_; 
wire u2__abc_52138_new_n16419_; 
wire u2__abc_52138_new_n16420_; 
wire u2__abc_52138_new_n16421_; 
wire u2__abc_52138_new_n16422_; 
wire u2__abc_52138_new_n16424_; 
wire u2__abc_52138_new_n16425_; 
wire u2__abc_52138_new_n16426_; 
wire u2__abc_52138_new_n16427_; 
wire u2__abc_52138_new_n16428_; 
wire u2__abc_52138_new_n16429_; 
wire u2__abc_52138_new_n16430_; 
wire u2__abc_52138_new_n16432_; 
wire u2__abc_52138_new_n16433_; 
wire u2__abc_52138_new_n16434_; 
wire u2__abc_52138_new_n16435_; 
wire u2__abc_52138_new_n16436_; 
wire u2__abc_52138_new_n16437_; 
wire u2__abc_52138_new_n16438_; 
wire u2__abc_52138_new_n16440_; 
wire u2__abc_52138_new_n16441_; 
wire u2__abc_52138_new_n16442_; 
wire u2__abc_52138_new_n16443_; 
wire u2__abc_52138_new_n16444_; 
wire u2__abc_52138_new_n16445_; 
wire u2__abc_52138_new_n16447_; 
wire u2__abc_52138_new_n16448_; 
wire u2__abc_52138_new_n16449_; 
wire u2__abc_52138_new_n16450_; 
wire u2__abc_52138_new_n16451_; 
wire u2__abc_52138_new_n16452_; 
wire u2__abc_52138_new_n16453_; 
wire u2__abc_52138_new_n16455_; 
wire u2__abc_52138_new_n16456_; 
wire u2__abc_52138_new_n16457_; 
wire u2__abc_52138_new_n16458_; 
wire u2__abc_52138_new_n16459_; 
wire u2__abc_52138_new_n16460_; 
wire u2__abc_52138_new_n16461_; 
wire u2__abc_52138_new_n16463_; 
wire u2__abc_52138_new_n16464_; 
wire u2__abc_52138_new_n16465_; 
wire u2__abc_52138_new_n16466_; 
wire u2__abc_52138_new_n16467_; 
wire u2__abc_52138_new_n16468_; 
wire u2__abc_52138_new_n16469_; 
wire u2__abc_52138_new_n16471_; 
wire u2__abc_52138_new_n16472_; 
wire u2__abc_52138_new_n16473_; 
wire u2__abc_52138_new_n16474_; 
wire u2__abc_52138_new_n16475_; 
wire u2__abc_52138_new_n16476_; 
wire u2__abc_52138_new_n16478_; 
wire u2__abc_52138_new_n16479_; 
wire u2__abc_52138_new_n16480_; 
wire u2__abc_52138_new_n16481_; 
wire u2__abc_52138_new_n16482_; 
wire u2__abc_52138_new_n16483_; 
wire u2__abc_52138_new_n16484_; 
wire u2__abc_52138_new_n16486_; 
wire u2__abc_52138_new_n16487_; 
wire u2__abc_52138_new_n16488_; 
wire u2__abc_52138_new_n16489_; 
wire u2__abc_52138_new_n16490_; 
wire u2__abc_52138_new_n16491_; 
wire u2__abc_52138_new_n16492_; 
wire u2__abc_52138_new_n16494_; 
wire u2__abc_52138_new_n16495_; 
wire u2__abc_52138_new_n16496_; 
wire u2__abc_52138_new_n16497_; 
wire u2__abc_52138_new_n16498_; 
wire u2__abc_52138_new_n16499_; 
wire u2__abc_52138_new_n16500_; 
wire u2__abc_52138_new_n16502_; 
wire u2__abc_52138_new_n16503_; 
wire u2__abc_52138_new_n16504_; 
wire u2__abc_52138_new_n16505_; 
wire u2__abc_52138_new_n16506_; 
wire u2__abc_52138_new_n16507_; 
wire u2__abc_52138_new_n16509_; 
wire u2__abc_52138_new_n16510_; 
wire u2__abc_52138_new_n16511_; 
wire u2__abc_52138_new_n16512_; 
wire u2__abc_52138_new_n16513_; 
wire u2__abc_52138_new_n16514_; 
wire u2__abc_52138_new_n16515_; 
wire u2__abc_52138_new_n16517_; 
wire u2__abc_52138_new_n16518_; 
wire u2__abc_52138_new_n16519_; 
wire u2__abc_52138_new_n16520_; 
wire u2__abc_52138_new_n16521_; 
wire u2__abc_52138_new_n16522_; 
wire u2__abc_52138_new_n16523_; 
wire u2__abc_52138_new_n16525_; 
wire u2__abc_52138_new_n16526_; 
wire u2__abc_52138_new_n16527_; 
wire u2__abc_52138_new_n16528_; 
wire u2__abc_52138_new_n16529_; 
wire u2__abc_52138_new_n16530_; 
wire u2__abc_52138_new_n16531_; 
wire u2__abc_52138_new_n16533_; 
wire u2__abc_52138_new_n16534_; 
wire u2__abc_52138_new_n16535_; 
wire u2__abc_52138_new_n16536_; 
wire u2__abc_52138_new_n16537_; 
wire u2__abc_52138_new_n16538_; 
wire u2__abc_52138_new_n2962_; 
wire u2__abc_52138_new_n2963_; 
wire u2__abc_52138_new_n2964_; 
wire u2__abc_52138_new_n2965_; 
wire u2__abc_52138_new_n2966_; 
wire u2__abc_52138_new_n2967_; 
wire u2__abc_52138_new_n2968_; 
wire u2__abc_52138_new_n2969_; 
wire u2__abc_52138_new_n2970_; 
wire u2__abc_52138_new_n2971_; 
wire u2__abc_52138_new_n2972_; 
wire u2__abc_52138_new_n2973_; 
wire u2__abc_52138_new_n2974_; 
wire u2__abc_52138_new_n2975_; 
wire u2__abc_52138_new_n2976_; 
wire u2__abc_52138_new_n2977_; 
wire u2__abc_52138_new_n2978_; 
wire u2__abc_52138_new_n2979_; 
wire u2__abc_52138_new_n2981_; 
wire u2__abc_52138_new_n2982_; 
wire u2__abc_52138_new_n2983_; 
wire u2__abc_52138_new_n2984_; 
wire u2__abc_52138_new_n2986_; 
wire u2__abc_52138_new_n2987_; 
wire u2__abc_52138_new_n2988_; 
wire u2__abc_52138_new_n2989_; 
wire u2__abc_52138_new_n2990_; 
wire u2__abc_52138_new_n2991_; 
wire u2__abc_52138_new_n2992_; 
wire u2__abc_52138_new_n2994_; 
wire u2__abc_52138_new_n2995_; 
wire u2__abc_52138_new_n2996_; 
wire u2__abc_52138_new_n2997_; 
wire u2__abc_52138_new_n2998_; 
wire u2__abc_52138_new_n2999_; 
wire u2__abc_52138_new_n3000_; 
wire u2__abc_52138_new_n3001_; 
wire u2__abc_52138_new_n3002_; 
wire u2__abc_52138_new_n3003_; 
wire u2__abc_52138_new_n3004_; 
wire u2__abc_52138_new_n3005_; 
wire u2__abc_52138_new_n3006_; 
wire u2__abc_52138_new_n3007_; 
wire u2__abc_52138_new_n3008_; 
wire u2__abc_52138_new_n3009_; 
wire u2__abc_52138_new_n3010_; 
wire u2__abc_52138_new_n3011_; 
wire u2__abc_52138_new_n3012_; 
wire u2__abc_52138_new_n3013_; 
wire u2__abc_52138_new_n3014_; 
wire u2__abc_52138_new_n3015_; 
wire u2__abc_52138_new_n3016_; 
wire u2__abc_52138_new_n3017_; 
wire u2__abc_52138_new_n3018_; 
wire u2__abc_52138_new_n3019_; 
wire u2__abc_52138_new_n3020_; 
wire u2__abc_52138_new_n3021_; 
wire u2__abc_52138_new_n3022_; 
wire u2__abc_52138_new_n3023_; 
wire u2__abc_52138_new_n3024_; 
wire u2__abc_52138_new_n3025_; 
wire u2__abc_52138_new_n3026_; 
wire u2__abc_52138_new_n3027_; 
wire u2__abc_52138_new_n3028_; 
wire u2__abc_52138_new_n3029_; 
wire u2__abc_52138_new_n3030_; 
wire u2__abc_52138_new_n3031_; 
wire u2__abc_52138_new_n3032_; 
wire u2__abc_52138_new_n3033_; 
wire u2__abc_52138_new_n3034_; 
wire u2__abc_52138_new_n3035_; 
wire u2__abc_52138_new_n3036_; 
wire u2__abc_52138_new_n3037_; 
wire u2__abc_52138_new_n3038_; 
wire u2__abc_52138_new_n3039_; 
wire u2__abc_52138_new_n3040_; 
wire u2__abc_52138_new_n3041_; 
wire u2__abc_52138_new_n3042_; 
wire u2__abc_52138_new_n3043_; 
wire u2__abc_52138_new_n3044_; 
wire u2__abc_52138_new_n3045_; 
wire u2__abc_52138_new_n3046_; 
wire u2__abc_52138_new_n3047_; 
wire u2__abc_52138_new_n3048_; 
wire u2__abc_52138_new_n3049_; 
wire u2__abc_52138_new_n3050_; 
wire u2__abc_52138_new_n3051_; 
wire u2__abc_52138_new_n3052_; 
wire u2__abc_52138_new_n3053_; 
wire u2__abc_52138_new_n3054_; 
wire u2__abc_52138_new_n3055_; 
wire u2__abc_52138_new_n3056_; 
wire u2__abc_52138_new_n3057_; 
wire u2__abc_52138_new_n3058_; 
wire u2__abc_52138_new_n3059_; 
wire u2__abc_52138_new_n3060_; 
wire u2__abc_52138_new_n3061_; 
wire u2__abc_52138_new_n3062_; 
wire u2__abc_52138_new_n3063_; 
wire u2__abc_52138_new_n3064_; 
wire u2__abc_52138_new_n3065_; 
wire u2__abc_52138_new_n3066_; 
wire u2__abc_52138_new_n3067_; 
wire u2__abc_52138_new_n3068_; 
wire u2__abc_52138_new_n3069_; 
wire u2__abc_52138_new_n3070_; 
wire u2__abc_52138_new_n3071_; 
wire u2__abc_52138_new_n3072_; 
wire u2__abc_52138_new_n3073_; 
wire u2__abc_52138_new_n3074_; 
wire u2__abc_52138_new_n3075_; 
wire u2__abc_52138_new_n3076_; 
wire u2__abc_52138_new_n3077_; 
wire u2__abc_52138_new_n3078_; 
wire u2__abc_52138_new_n3079_; 
wire u2__abc_52138_new_n3080_; 
wire u2__abc_52138_new_n3081_; 
wire u2__abc_52138_new_n3082_; 
wire u2__abc_52138_new_n3083_; 
wire u2__abc_52138_new_n3084_; 
wire u2__abc_52138_new_n3085_; 
wire u2__abc_52138_new_n3086_; 
wire u2__abc_52138_new_n3087_; 
wire u2__abc_52138_new_n3088_; 
wire u2__abc_52138_new_n3089_; 
wire u2__abc_52138_new_n3090_; 
wire u2__abc_52138_new_n3091_; 
wire u2__abc_52138_new_n3092_; 
wire u2__abc_52138_new_n3093_; 
wire u2__abc_52138_new_n3094_; 
wire u2__abc_52138_new_n3095_; 
wire u2__abc_52138_new_n3096_; 
wire u2__abc_52138_new_n3097_; 
wire u2__abc_52138_new_n3098_; 
wire u2__abc_52138_new_n3099_; 
wire u2__abc_52138_new_n3100_; 
wire u2__abc_52138_new_n3101_; 
wire u2__abc_52138_new_n3102_; 
wire u2__abc_52138_new_n3103_; 
wire u2__abc_52138_new_n3104_; 
wire u2__abc_52138_new_n3105_; 
wire u2__abc_52138_new_n3106_; 
wire u2__abc_52138_new_n3107_; 
wire u2__abc_52138_new_n3108_; 
wire u2__abc_52138_new_n3109_; 
wire u2__abc_52138_new_n3110_; 
wire u2__abc_52138_new_n3111_; 
wire u2__abc_52138_new_n3112_; 
wire u2__abc_52138_new_n3113_; 
wire u2__abc_52138_new_n3114_; 
wire u2__abc_52138_new_n3115_; 
wire u2__abc_52138_new_n3116_; 
wire u2__abc_52138_new_n3117_; 
wire u2__abc_52138_new_n3118_; 
wire u2__abc_52138_new_n3119_; 
wire u2__abc_52138_new_n3120_; 
wire u2__abc_52138_new_n3121_; 
wire u2__abc_52138_new_n3122_; 
wire u2__abc_52138_new_n3123_; 
wire u2__abc_52138_new_n3124_; 
wire u2__abc_52138_new_n3125_; 
wire u2__abc_52138_new_n3126_; 
wire u2__abc_52138_new_n3127_; 
wire u2__abc_52138_new_n3128_; 
wire u2__abc_52138_new_n3129_; 
wire u2__abc_52138_new_n3130_; 
wire u2__abc_52138_new_n3131_; 
wire u2__abc_52138_new_n3132_; 
wire u2__abc_52138_new_n3133_; 
wire u2__abc_52138_new_n3134_; 
wire u2__abc_52138_new_n3135_; 
wire u2__abc_52138_new_n3136_; 
wire u2__abc_52138_new_n3137_; 
wire u2__abc_52138_new_n3138_; 
wire u2__abc_52138_new_n3139_; 
wire u2__abc_52138_new_n3140_; 
wire u2__abc_52138_new_n3141_; 
wire u2__abc_52138_new_n3142_; 
wire u2__abc_52138_new_n3143_; 
wire u2__abc_52138_new_n3144_; 
wire u2__abc_52138_new_n3145_; 
wire u2__abc_52138_new_n3146_; 
wire u2__abc_52138_new_n3147_; 
wire u2__abc_52138_new_n3148_; 
wire u2__abc_52138_new_n3149_; 
wire u2__abc_52138_new_n3150_; 
wire u2__abc_52138_new_n3151_; 
wire u2__abc_52138_new_n3152_; 
wire u2__abc_52138_new_n3153_; 
wire u2__abc_52138_new_n3154_; 
wire u2__abc_52138_new_n3155_; 
wire u2__abc_52138_new_n3156_; 
wire u2__abc_52138_new_n3157_; 
wire u2__abc_52138_new_n3158_; 
wire u2__abc_52138_new_n3159_; 
wire u2__abc_52138_new_n3160_; 
wire u2__abc_52138_new_n3161_; 
wire u2__abc_52138_new_n3162_; 
wire u2__abc_52138_new_n3163_; 
wire u2__abc_52138_new_n3164_; 
wire u2__abc_52138_new_n3165_; 
wire u2__abc_52138_new_n3166_; 
wire u2__abc_52138_new_n3167_; 
wire u2__abc_52138_new_n3168_; 
wire u2__abc_52138_new_n3169_; 
wire u2__abc_52138_new_n3170_; 
wire u2__abc_52138_new_n3171_; 
wire u2__abc_52138_new_n3172_; 
wire u2__abc_52138_new_n3173_; 
wire u2__abc_52138_new_n3174_; 
wire u2__abc_52138_new_n3175_; 
wire u2__abc_52138_new_n3176_; 
wire u2__abc_52138_new_n3177_; 
wire u2__abc_52138_new_n3178_; 
wire u2__abc_52138_new_n3179_; 
wire u2__abc_52138_new_n3180_; 
wire u2__abc_52138_new_n3181_; 
wire u2__abc_52138_new_n3182_; 
wire u2__abc_52138_new_n3183_; 
wire u2__abc_52138_new_n3184_; 
wire u2__abc_52138_new_n3185_; 
wire u2__abc_52138_new_n3186_; 
wire u2__abc_52138_new_n3187_; 
wire u2__abc_52138_new_n3188_; 
wire u2__abc_52138_new_n3189_; 
wire u2__abc_52138_new_n3190_; 
wire u2__abc_52138_new_n3191_; 
wire u2__abc_52138_new_n3192_; 
wire u2__abc_52138_new_n3193_; 
wire u2__abc_52138_new_n3194_; 
wire u2__abc_52138_new_n3195_; 
wire u2__abc_52138_new_n3196_; 
wire u2__abc_52138_new_n3197_; 
wire u2__abc_52138_new_n3198_; 
wire u2__abc_52138_new_n3199_; 
wire u2__abc_52138_new_n3200_; 
wire u2__abc_52138_new_n3201_; 
wire u2__abc_52138_new_n3202_; 
wire u2__abc_52138_new_n3203_; 
wire u2__abc_52138_new_n3204_; 
wire u2__abc_52138_new_n3205_; 
wire u2__abc_52138_new_n3206_; 
wire u2__abc_52138_new_n3207_; 
wire u2__abc_52138_new_n3208_; 
wire u2__abc_52138_new_n3209_; 
wire u2__abc_52138_new_n3210_; 
wire u2__abc_52138_new_n3211_; 
wire u2__abc_52138_new_n3212_; 
wire u2__abc_52138_new_n3213_; 
wire u2__abc_52138_new_n3214_; 
wire u2__abc_52138_new_n3215_; 
wire u2__abc_52138_new_n3216_; 
wire u2__abc_52138_new_n3217_; 
wire u2__abc_52138_new_n3218_; 
wire u2__abc_52138_new_n3219_; 
wire u2__abc_52138_new_n3220_; 
wire u2__abc_52138_new_n3221_; 
wire u2__abc_52138_new_n3222_; 
wire u2__abc_52138_new_n3223_; 
wire u2__abc_52138_new_n3224_; 
wire u2__abc_52138_new_n3225_; 
wire u2__abc_52138_new_n3226_; 
wire u2__abc_52138_new_n3227_; 
wire u2__abc_52138_new_n3228_; 
wire u2__abc_52138_new_n3229_; 
wire u2__abc_52138_new_n3230_; 
wire u2__abc_52138_new_n3231_; 
wire u2__abc_52138_new_n3232_; 
wire u2__abc_52138_new_n3233_; 
wire u2__abc_52138_new_n3234_; 
wire u2__abc_52138_new_n3235_; 
wire u2__abc_52138_new_n3236_; 
wire u2__abc_52138_new_n3237_; 
wire u2__abc_52138_new_n3238_; 
wire u2__abc_52138_new_n3239_; 
wire u2__abc_52138_new_n3240_; 
wire u2__abc_52138_new_n3241_; 
wire u2__abc_52138_new_n3242_; 
wire u2__abc_52138_new_n3243_; 
wire u2__abc_52138_new_n3244_; 
wire u2__abc_52138_new_n3245_; 
wire u2__abc_52138_new_n3246_; 
wire u2__abc_52138_new_n3247_; 
wire u2__abc_52138_new_n3248_; 
wire u2__abc_52138_new_n3249_; 
wire u2__abc_52138_new_n3250_; 
wire u2__abc_52138_new_n3251_; 
wire u2__abc_52138_new_n3252_; 
wire u2__abc_52138_new_n3253_; 
wire u2__abc_52138_new_n3254_; 
wire u2__abc_52138_new_n3255_; 
wire u2__abc_52138_new_n3256_; 
wire u2__abc_52138_new_n3257_; 
wire u2__abc_52138_new_n3258_; 
wire u2__abc_52138_new_n3259_; 
wire u2__abc_52138_new_n3260_; 
wire u2__abc_52138_new_n3261_; 
wire u2__abc_52138_new_n3262_; 
wire u2__abc_52138_new_n3263_; 
wire u2__abc_52138_new_n3264_; 
wire u2__abc_52138_new_n3265_; 
wire u2__abc_52138_new_n3266_; 
wire u2__abc_52138_new_n3267_; 
wire u2__abc_52138_new_n3268_; 
wire u2__abc_52138_new_n3269_; 
wire u2__abc_52138_new_n3270_; 
wire u2__abc_52138_new_n3271_; 
wire u2__abc_52138_new_n3272_; 
wire u2__abc_52138_new_n3273_; 
wire u2__abc_52138_new_n3274_; 
wire u2__abc_52138_new_n3275_; 
wire u2__abc_52138_new_n3276_; 
wire u2__abc_52138_new_n3277_; 
wire u2__abc_52138_new_n3278_; 
wire u2__abc_52138_new_n3279_; 
wire u2__abc_52138_new_n3280_; 
wire u2__abc_52138_new_n3281_; 
wire u2__abc_52138_new_n3282_; 
wire u2__abc_52138_new_n3283_; 
wire u2__abc_52138_new_n3284_; 
wire u2__abc_52138_new_n3285_; 
wire u2__abc_52138_new_n3286_; 
wire u2__abc_52138_new_n3287_; 
wire u2__abc_52138_new_n3288_; 
wire u2__abc_52138_new_n3289_; 
wire u2__abc_52138_new_n3290_; 
wire u2__abc_52138_new_n3291_; 
wire u2__abc_52138_new_n3292_; 
wire u2__abc_52138_new_n3293_; 
wire u2__abc_52138_new_n3294_; 
wire u2__abc_52138_new_n3295_; 
wire u2__abc_52138_new_n3296_; 
wire u2__abc_52138_new_n3297_; 
wire u2__abc_52138_new_n3298_; 
wire u2__abc_52138_new_n3299_; 
wire u2__abc_52138_new_n3300_; 
wire u2__abc_52138_new_n3301_; 
wire u2__abc_52138_new_n3302_; 
wire u2__abc_52138_new_n3303_; 
wire u2__abc_52138_new_n3304_; 
wire u2__abc_52138_new_n3305_; 
wire u2__abc_52138_new_n3306_; 
wire u2__abc_52138_new_n3307_; 
wire u2__abc_52138_new_n3308_; 
wire u2__abc_52138_new_n3309_; 
wire u2__abc_52138_new_n3310_; 
wire u2__abc_52138_new_n3311_; 
wire u2__abc_52138_new_n3312_; 
wire u2__abc_52138_new_n3313_; 
wire u2__abc_52138_new_n3314_; 
wire u2__abc_52138_new_n3315_; 
wire u2__abc_52138_new_n3316_; 
wire u2__abc_52138_new_n3317_; 
wire u2__abc_52138_new_n3318_; 
wire u2__abc_52138_new_n3319_; 
wire u2__abc_52138_new_n3320_; 
wire u2__abc_52138_new_n3321_; 
wire u2__abc_52138_new_n3322_; 
wire u2__abc_52138_new_n3323_; 
wire u2__abc_52138_new_n3324_; 
wire u2__abc_52138_new_n3325_; 
wire u2__abc_52138_new_n3326_; 
wire u2__abc_52138_new_n3327_; 
wire u2__abc_52138_new_n3328_; 
wire u2__abc_52138_new_n3329_; 
wire u2__abc_52138_new_n3330_; 
wire u2__abc_52138_new_n3331_; 
wire u2__abc_52138_new_n3332_; 
wire u2__abc_52138_new_n3333_; 
wire u2__abc_52138_new_n3334_; 
wire u2__abc_52138_new_n3335_; 
wire u2__abc_52138_new_n3336_; 
wire u2__abc_52138_new_n3337_; 
wire u2__abc_52138_new_n3338_; 
wire u2__abc_52138_new_n3339_; 
wire u2__abc_52138_new_n3340_; 
wire u2__abc_52138_new_n3341_; 
wire u2__abc_52138_new_n3342_; 
wire u2__abc_52138_new_n3343_; 
wire u2__abc_52138_new_n3344_; 
wire u2__abc_52138_new_n3345_; 
wire u2__abc_52138_new_n3346_; 
wire u2__abc_52138_new_n3347_; 
wire u2__abc_52138_new_n3348_; 
wire u2__abc_52138_new_n3349_; 
wire u2__abc_52138_new_n3350_; 
wire u2__abc_52138_new_n3351_; 
wire u2__abc_52138_new_n3352_; 
wire u2__abc_52138_new_n3353_; 
wire u2__abc_52138_new_n3354_; 
wire u2__abc_52138_new_n3355_; 
wire u2__abc_52138_new_n3356_; 
wire u2__abc_52138_new_n3357_; 
wire u2__abc_52138_new_n3358_; 
wire u2__abc_52138_new_n3359_; 
wire u2__abc_52138_new_n3360_; 
wire u2__abc_52138_new_n3361_; 
wire u2__abc_52138_new_n3362_; 
wire u2__abc_52138_new_n3363_; 
wire u2__abc_52138_new_n3364_; 
wire u2__abc_52138_new_n3365_; 
wire u2__abc_52138_new_n3366_; 
wire u2__abc_52138_new_n3367_; 
wire u2__abc_52138_new_n3368_; 
wire u2__abc_52138_new_n3369_; 
wire u2__abc_52138_new_n3370_; 
wire u2__abc_52138_new_n3371_; 
wire u2__abc_52138_new_n3372_; 
wire u2__abc_52138_new_n3373_; 
wire u2__abc_52138_new_n3374_; 
wire u2__abc_52138_new_n3375_; 
wire u2__abc_52138_new_n3376_; 
wire u2__abc_52138_new_n3377_; 
wire u2__abc_52138_new_n3378_; 
wire u2__abc_52138_new_n3379_; 
wire u2__abc_52138_new_n3380_; 
wire u2__abc_52138_new_n3381_; 
wire u2__abc_52138_new_n3382_; 
wire u2__abc_52138_new_n3383_; 
wire u2__abc_52138_new_n3384_; 
wire u2__abc_52138_new_n3385_; 
wire u2__abc_52138_new_n3386_; 
wire u2__abc_52138_new_n3387_; 
wire u2__abc_52138_new_n3388_; 
wire u2__abc_52138_new_n3389_; 
wire u2__abc_52138_new_n3390_; 
wire u2__abc_52138_new_n3391_; 
wire u2__abc_52138_new_n3392_; 
wire u2__abc_52138_new_n3393_; 
wire u2__abc_52138_new_n3394_; 
wire u2__abc_52138_new_n3395_; 
wire u2__abc_52138_new_n3396_; 
wire u2__abc_52138_new_n3397_; 
wire u2__abc_52138_new_n3398_; 
wire u2__abc_52138_new_n3399_; 
wire u2__abc_52138_new_n3400_; 
wire u2__abc_52138_new_n3401_; 
wire u2__abc_52138_new_n3402_; 
wire u2__abc_52138_new_n3403_; 
wire u2__abc_52138_new_n3404_; 
wire u2__abc_52138_new_n3405_; 
wire u2__abc_52138_new_n3406_; 
wire u2__abc_52138_new_n3407_; 
wire u2__abc_52138_new_n3408_; 
wire u2__abc_52138_new_n3409_; 
wire u2__abc_52138_new_n3410_; 
wire u2__abc_52138_new_n3411_; 
wire u2__abc_52138_new_n3412_; 
wire u2__abc_52138_new_n3413_; 
wire u2__abc_52138_new_n3414_; 
wire u2__abc_52138_new_n3415_; 
wire u2__abc_52138_new_n3416_; 
wire u2__abc_52138_new_n3417_; 
wire u2__abc_52138_new_n3418_; 
wire u2__abc_52138_new_n3419_; 
wire u2__abc_52138_new_n3420_; 
wire u2__abc_52138_new_n3421_; 
wire u2__abc_52138_new_n3422_; 
wire u2__abc_52138_new_n3423_; 
wire u2__abc_52138_new_n3424_; 
wire u2__abc_52138_new_n3425_; 
wire u2__abc_52138_new_n3426_; 
wire u2__abc_52138_new_n3427_; 
wire u2__abc_52138_new_n3428_; 
wire u2__abc_52138_new_n3429_; 
wire u2__abc_52138_new_n3430_; 
wire u2__abc_52138_new_n3431_; 
wire u2__abc_52138_new_n3432_; 
wire u2__abc_52138_new_n3433_; 
wire u2__abc_52138_new_n3434_; 
wire u2__abc_52138_new_n3435_; 
wire u2__abc_52138_new_n3436_; 
wire u2__abc_52138_new_n3437_; 
wire u2__abc_52138_new_n3438_; 
wire u2__abc_52138_new_n3439_; 
wire u2__abc_52138_new_n3440_; 
wire u2__abc_52138_new_n3441_; 
wire u2__abc_52138_new_n3442_; 
wire u2__abc_52138_new_n3443_; 
wire u2__abc_52138_new_n3444_; 
wire u2__abc_52138_new_n3445_; 
wire u2__abc_52138_new_n3446_; 
wire u2__abc_52138_new_n3447_; 
wire u2__abc_52138_new_n3448_; 
wire u2__abc_52138_new_n3449_; 
wire u2__abc_52138_new_n3450_; 
wire u2__abc_52138_new_n3451_; 
wire u2__abc_52138_new_n3452_; 
wire u2__abc_52138_new_n3453_; 
wire u2__abc_52138_new_n3454_; 
wire u2__abc_52138_new_n3455_; 
wire u2__abc_52138_new_n3456_; 
wire u2__abc_52138_new_n3457_; 
wire u2__abc_52138_new_n3458_; 
wire u2__abc_52138_new_n3459_; 
wire u2__abc_52138_new_n3460_; 
wire u2__abc_52138_new_n3461_; 
wire u2__abc_52138_new_n3462_; 
wire u2__abc_52138_new_n3463_; 
wire u2__abc_52138_new_n3464_; 
wire u2__abc_52138_new_n3465_; 
wire u2__abc_52138_new_n3466_; 
wire u2__abc_52138_new_n3467_; 
wire u2__abc_52138_new_n3468_; 
wire u2__abc_52138_new_n3469_; 
wire u2__abc_52138_new_n3470_; 
wire u2__abc_52138_new_n3471_; 
wire u2__abc_52138_new_n3472_; 
wire u2__abc_52138_new_n3473_; 
wire u2__abc_52138_new_n3474_; 
wire u2__abc_52138_new_n3475_; 
wire u2__abc_52138_new_n3476_; 
wire u2__abc_52138_new_n3477_; 
wire u2__abc_52138_new_n3478_; 
wire u2__abc_52138_new_n3479_; 
wire u2__abc_52138_new_n3480_; 
wire u2__abc_52138_new_n3481_; 
wire u2__abc_52138_new_n3482_; 
wire u2__abc_52138_new_n3483_; 
wire u2__abc_52138_new_n3484_; 
wire u2__abc_52138_new_n3485_; 
wire u2__abc_52138_new_n3486_; 
wire u2__abc_52138_new_n3487_; 
wire u2__abc_52138_new_n3488_; 
wire u2__abc_52138_new_n3489_; 
wire u2__abc_52138_new_n3490_; 
wire u2__abc_52138_new_n3491_; 
wire u2__abc_52138_new_n3492_; 
wire u2__abc_52138_new_n3493_; 
wire u2__abc_52138_new_n3494_; 
wire u2__abc_52138_new_n3495_; 
wire u2__abc_52138_new_n3496_; 
wire u2__abc_52138_new_n3497_; 
wire u2__abc_52138_new_n3498_; 
wire u2__abc_52138_new_n3499_; 
wire u2__abc_52138_new_n3500_; 
wire u2__abc_52138_new_n3501_; 
wire u2__abc_52138_new_n3502_; 
wire u2__abc_52138_new_n3503_; 
wire u2__abc_52138_new_n3504_; 
wire u2__abc_52138_new_n3505_; 
wire u2__abc_52138_new_n3506_; 
wire u2__abc_52138_new_n3507_; 
wire u2__abc_52138_new_n3508_; 
wire u2__abc_52138_new_n3509_; 
wire u2__abc_52138_new_n3510_; 
wire u2__abc_52138_new_n3511_; 
wire u2__abc_52138_new_n3512_; 
wire u2__abc_52138_new_n3513_; 
wire u2__abc_52138_new_n3514_; 
wire u2__abc_52138_new_n3515_; 
wire u2__abc_52138_new_n3516_; 
wire u2__abc_52138_new_n3517_; 
wire u2__abc_52138_new_n3518_; 
wire u2__abc_52138_new_n3519_; 
wire u2__abc_52138_new_n3520_; 
wire u2__abc_52138_new_n3521_; 
wire u2__abc_52138_new_n3522_; 
wire u2__abc_52138_new_n3523_; 
wire u2__abc_52138_new_n3524_; 
wire u2__abc_52138_new_n3525_; 
wire u2__abc_52138_new_n3526_; 
wire u2__abc_52138_new_n3527_; 
wire u2__abc_52138_new_n3528_; 
wire u2__abc_52138_new_n3529_; 
wire u2__abc_52138_new_n3530_; 
wire u2__abc_52138_new_n3531_; 
wire u2__abc_52138_new_n3532_; 
wire u2__abc_52138_new_n3533_; 
wire u2__abc_52138_new_n3534_; 
wire u2__abc_52138_new_n3535_; 
wire u2__abc_52138_new_n3536_; 
wire u2__abc_52138_new_n3537_; 
wire u2__abc_52138_new_n3538_; 
wire u2__abc_52138_new_n3539_; 
wire u2__abc_52138_new_n3540_; 
wire u2__abc_52138_new_n3541_; 
wire u2__abc_52138_new_n3542_; 
wire u2__abc_52138_new_n3543_; 
wire u2__abc_52138_new_n3544_; 
wire u2__abc_52138_new_n3545_; 
wire u2__abc_52138_new_n3546_; 
wire u2__abc_52138_new_n3547_; 
wire u2__abc_52138_new_n3548_; 
wire u2__abc_52138_new_n3549_; 
wire u2__abc_52138_new_n3550_; 
wire u2__abc_52138_new_n3551_; 
wire u2__abc_52138_new_n3552_; 
wire u2__abc_52138_new_n3553_; 
wire u2__abc_52138_new_n3554_; 
wire u2__abc_52138_new_n3555_; 
wire u2__abc_52138_new_n3556_; 
wire u2__abc_52138_new_n3557_; 
wire u2__abc_52138_new_n3558_; 
wire u2__abc_52138_new_n3559_; 
wire u2__abc_52138_new_n3560_; 
wire u2__abc_52138_new_n3561_; 
wire u2__abc_52138_new_n3562_; 
wire u2__abc_52138_new_n3563_; 
wire u2__abc_52138_new_n3564_; 
wire u2__abc_52138_new_n3565_; 
wire u2__abc_52138_new_n3566_; 
wire u2__abc_52138_new_n3567_; 
wire u2__abc_52138_new_n3568_; 
wire u2__abc_52138_new_n3569_; 
wire u2__abc_52138_new_n3570_; 
wire u2__abc_52138_new_n3571_; 
wire u2__abc_52138_new_n3572_; 
wire u2__abc_52138_new_n3573_; 
wire u2__abc_52138_new_n3574_; 
wire u2__abc_52138_new_n3575_; 
wire u2__abc_52138_new_n3576_; 
wire u2__abc_52138_new_n3577_; 
wire u2__abc_52138_new_n3578_; 
wire u2__abc_52138_new_n3579_; 
wire u2__abc_52138_new_n3580_; 
wire u2__abc_52138_new_n3581_; 
wire u2__abc_52138_new_n3582_; 
wire u2__abc_52138_new_n3583_; 
wire u2__abc_52138_new_n3584_; 
wire u2__abc_52138_new_n3585_; 
wire u2__abc_52138_new_n3586_; 
wire u2__abc_52138_new_n3587_; 
wire u2__abc_52138_new_n3588_; 
wire u2__abc_52138_new_n3589_; 
wire u2__abc_52138_new_n3590_; 
wire u2__abc_52138_new_n3591_; 
wire u2__abc_52138_new_n3592_; 
wire u2__abc_52138_new_n3593_; 
wire u2__abc_52138_new_n3594_; 
wire u2__abc_52138_new_n3595_; 
wire u2__abc_52138_new_n3596_; 
wire u2__abc_52138_new_n3597_; 
wire u2__abc_52138_new_n3598_; 
wire u2__abc_52138_new_n3599_; 
wire u2__abc_52138_new_n3600_; 
wire u2__abc_52138_new_n3601_; 
wire u2__abc_52138_new_n3602_; 
wire u2__abc_52138_new_n3603_; 
wire u2__abc_52138_new_n3604_; 
wire u2__abc_52138_new_n3605_; 
wire u2__abc_52138_new_n3606_; 
wire u2__abc_52138_new_n3607_; 
wire u2__abc_52138_new_n3608_; 
wire u2__abc_52138_new_n3609_; 
wire u2__abc_52138_new_n3610_; 
wire u2__abc_52138_new_n3611_; 
wire u2__abc_52138_new_n3612_; 
wire u2__abc_52138_new_n3613_; 
wire u2__abc_52138_new_n3614_; 
wire u2__abc_52138_new_n3615_; 
wire u2__abc_52138_new_n3616_; 
wire u2__abc_52138_new_n3617_; 
wire u2__abc_52138_new_n3618_; 
wire u2__abc_52138_new_n3619_; 
wire u2__abc_52138_new_n3620_; 
wire u2__abc_52138_new_n3621_; 
wire u2__abc_52138_new_n3622_; 
wire u2__abc_52138_new_n3623_; 
wire u2__abc_52138_new_n3624_; 
wire u2__abc_52138_new_n3625_; 
wire u2__abc_52138_new_n3626_; 
wire u2__abc_52138_new_n3627_; 
wire u2__abc_52138_new_n3628_; 
wire u2__abc_52138_new_n3629_; 
wire u2__abc_52138_new_n3630_; 
wire u2__abc_52138_new_n3631_; 
wire u2__abc_52138_new_n3632_; 
wire u2__abc_52138_new_n3633_; 
wire u2__abc_52138_new_n3634_; 
wire u2__abc_52138_new_n3635_; 
wire u2__abc_52138_new_n3636_; 
wire u2__abc_52138_new_n3637_; 
wire u2__abc_52138_new_n3638_; 
wire u2__abc_52138_new_n3639_; 
wire u2__abc_52138_new_n3640_; 
wire u2__abc_52138_new_n3641_; 
wire u2__abc_52138_new_n3642_; 
wire u2__abc_52138_new_n3643_; 
wire u2__abc_52138_new_n3644_; 
wire u2__abc_52138_new_n3645_; 
wire u2__abc_52138_new_n3646_; 
wire u2__abc_52138_new_n3647_; 
wire u2__abc_52138_new_n3648_; 
wire u2__abc_52138_new_n3649_; 
wire u2__abc_52138_new_n3650_; 
wire u2__abc_52138_new_n3651_; 
wire u2__abc_52138_new_n3652_; 
wire u2__abc_52138_new_n3653_; 
wire u2__abc_52138_new_n3654_; 
wire u2__abc_52138_new_n3655_; 
wire u2__abc_52138_new_n3656_; 
wire u2__abc_52138_new_n3657_; 
wire u2__abc_52138_new_n3658_; 
wire u2__abc_52138_new_n3659_; 
wire u2__abc_52138_new_n3660_; 
wire u2__abc_52138_new_n3661_; 
wire u2__abc_52138_new_n3662_; 
wire u2__abc_52138_new_n3663_; 
wire u2__abc_52138_new_n3664_; 
wire u2__abc_52138_new_n3665_; 
wire u2__abc_52138_new_n3666_; 
wire u2__abc_52138_new_n3667_; 
wire u2__abc_52138_new_n3668_; 
wire u2__abc_52138_new_n3669_; 
wire u2__abc_52138_new_n3670_; 
wire u2__abc_52138_new_n3671_; 
wire u2__abc_52138_new_n3672_; 
wire u2__abc_52138_new_n3673_; 
wire u2__abc_52138_new_n3674_; 
wire u2__abc_52138_new_n3675_; 
wire u2__abc_52138_new_n3676_; 
wire u2__abc_52138_new_n3677_; 
wire u2__abc_52138_new_n3678_; 
wire u2__abc_52138_new_n3679_; 
wire u2__abc_52138_new_n3680_; 
wire u2__abc_52138_new_n3681_; 
wire u2__abc_52138_new_n3682_; 
wire u2__abc_52138_new_n3683_; 
wire u2__abc_52138_new_n3684_; 
wire u2__abc_52138_new_n3685_; 
wire u2__abc_52138_new_n3686_; 
wire u2__abc_52138_new_n3687_; 
wire u2__abc_52138_new_n3688_; 
wire u2__abc_52138_new_n3689_; 
wire u2__abc_52138_new_n3690_; 
wire u2__abc_52138_new_n3691_; 
wire u2__abc_52138_new_n3692_; 
wire u2__abc_52138_new_n3693_; 
wire u2__abc_52138_new_n3694_; 
wire u2__abc_52138_new_n3695_; 
wire u2__abc_52138_new_n3696_; 
wire u2__abc_52138_new_n3697_; 
wire u2__abc_52138_new_n3698_; 
wire u2__abc_52138_new_n3699_; 
wire u2__abc_52138_new_n3700_; 
wire u2__abc_52138_new_n3701_; 
wire u2__abc_52138_new_n3702_; 
wire u2__abc_52138_new_n3703_; 
wire u2__abc_52138_new_n3704_; 
wire u2__abc_52138_new_n3705_; 
wire u2__abc_52138_new_n3706_; 
wire u2__abc_52138_new_n3707_; 
wire u2__abc_52138_new_n3708_; 
wire u2__abc_52138_new_n3709_; 
wire u2__abc_52138_new_n3710_; 
wire u2__abc_52138_new_n3711_; 
wire u2__abc_52138_new_n3712_; 
wire u2__abc_52138_new_n3713_; 
wire u2__abc_52138_new_n3714_; 
wire u2__abc_52138_new_n3715_; 
wire u2__abc_52138_new_n3716_; 
wire u2__abc_52138_new_n3717_; 
wire u2__abc_52138_new_n3718_; 
wire u2__abc_52138_new_n3719_; 
wire u2__abc_52138_new_n3720_; 
wire u2__abc_52138_new_n3721_; 
wire u2__abc_52138_new_n3722_; 
wire u2__abc_52138_new_n3723_; 
wire u2__abc_52138_new_n3724_; 
wire u2__abc_52138_new_n3725_; 
wire u2__abc_52138_new_n3726_; 
wire u2__abc_52138_new_n3727_; 
wire u2__abc_52138_new_n3728_; 
wire u2__abc_52138_new_n3729_; 
wire u2__abc_52138_new_n3730_; 
wire u2__abc_52138_new_n3731_; 
wire u2__abc_52138_new_n3732_; 
wire u2__abc_52138_new_n3733_; 
wire u2__abc_52138_new_n3734_; 
wire u2__abc_52138_new_n3735_; 
wire u2__abc_52138_new_n3736_; 
wire u2__abc_52138_new_n3737_; 
wire u2__abc_52138_new_n3738_; 
wire u2__abc_52138_new_n3739_; 
wire u2__abc_52138_new_n3740_; 
wire u2__abc_52138_new_n3741_; 
wire u2__abc_52138_new_n3742_; 
wire u2__abc_52138_new_n3743_; 
wire u2__abc_52138_new_n3744_; 
wire u2__abc_52138_new_n3745_; 
wire u2__abc_52138_new_n3746_; 
wire u2__abc_52138_new_n3747_; 
wire u2__abc_52138_new_n3748_; 
wire u2__abc_52138_new_n3749_; 
wire u2__abc_52138_new_n3750_; 
wire u2__abc_52138_new_n3751_; 
wire u2__abc_52138_new_n3752_; 
wire u2__abc_52138_new_n3753_; 
wire u2__abc_52138_new_n3754_; 
wire u2__abc_52138_new_n3755_; 
wire u2__abc_52138_new_n3756_; 
wire u2__abc_52138_new_n3757_; 
wire u2__abc_52138_new_n3758_; 
wire u2__abc_52138_new_n3759_; 
wire u2__abc_52138_new_n3760_; 
wire u2__abc_52138_new_n3761_; 
wire u2__abc_52138_new_n3762_; 
wire u2__abc_52138_new_n3763_; 
wire u2__abc_52138_new_n3764_; 
wire u2__abc_52138_new_n3765_; 
wire u2__abc_52138_new_n3766_; 
wire u2__abc_52138_new_n3767_; 
wire u2__abc_52138_new_n3768_; 
wire u2__abc_52138_new_n3769_; 
wire u2__abc_52138_new_n3770_; 
wire u2__abc_52138_new_n3771_; 
wire u2__abc_52138_new_n3772_; 
wire u2__abc_52138_new_n3773_; 
wire u2__abc_52138_new_n3774_; 
wire u2__abc_52138_new_n3775_; 
wire u2__abc_52138_new_n3776_; 
wire u2__abc_52138_new_n3777_; 
wire u2__abc_52138_new_n3778_; 
wire u2__abc_52138_new_n3779_; 
wire u2__abc_52138_new_n3780_; 
wire u2__abc_52138_new_n3781_; 
wire u2__abc_52138_new_n3782_; 
wire u2__abc_52138_new_n3783_; 
wire u2__abc_52138_new_n3784_; 
wire u2__abc_52138_new_n3785_; 
wire u2__abc_52138_new_n3786_; 
wire u2__abc_52138_new_n3787_; 
wire u2__abc_52138_new_n3788_; 
wire u2__abc_52138_new_n3789_; 
wire u2__abc_52138_new_n3790_; 
wire u2__abc_52138_new_n3791_; 
wire u2__abc_52138_new_n3792_; 
wire u2__abc_52138_new_n3793_; 
wire u2__abc_52138_new_n3794_; 
wire u2__abc_52138_new_n3795_; 
wire u2__abc_52138_new_n3796_; 
wire u2__abc_52138_new_n3797_; 
wire u2__abc_52138_new_n3798_; 
wire u2__abc_52138_new_n3799_; 
wire u2__abc_52138_new_n3800_; 
wire u2__abc_52138_new_n3801_; 
wire u2__abc_52138_new_n3802_; 
wire u2__abc_52138_new_n3803_; 
wire u2__abc_52138_new_n3804_; 
wire u2__abc_52138_new_n3805_; 
wire u2__abc_52138_new_n3806_; 
wire u2__abc_52138_new_n3807_; 
wire u2__abc_52138_new_n3808_; 
wire u2__abc_52138_new_n3809_; 
wire u2__abc_52138_new_n3810_; 
wire u2__abc_52138_new_n3811_; 
wire u2__abc_52138_new_n3812_; 
wire u2__abc_52138_new_n3813_; 
wire u2__abc_52138_new_n3814_; 
wire u2__abc_52138_new_n3815_; 
wire u2__abc_52138_new_n3816_; 
wire u2__abc_52138_new_n3817_; 
wire u2__abc_52138_new_n3818_; 
wire u2__abc_52138_new_n3819_; 
wire u2__abc_52138_new_n3820_; 
wire u2__abc_52138_new_n3821_; 
wire u2__abc_52138_new_n3822_; 
wire u2__abc_52138_new_n3823_; 
wire u2__abc_52138_new_n3824_; 
wire u2__abc_52138_new_n3825_; 
wire u2__abc_52138_new_n3826_; 
wire u2__abc_52138_new_n3827_; 
wire u2__abc_52138_new_n3828_; 
wire u2__abc_52138_new_n3829_; 
wire u2__abc_52138_new_n3830_; 
wire u2__abc_52138_new_n3831_; 
wire u2__abc_52138_new_n3832_; 
wire u2__abc_52138_new_n3833_; 
wire u2__abc_52138_new_n3834_; 
wire u2__abc_52138_new_n3835_; 
wire u2__abc_52138_new_n3836_; 
wire u2__abc_52138_new_n3837_; 
wire u2__abc_52138_new_n3838_; 
wire u2__abc_52138_new_n3839_; 
wire u2__abc_52138_new_n3840_; 
wire u2__abc_52138_new_n3841_; 
wire u2__abc_52138_new_n3842_; 
wire u2__abc_52138_new_n3843_; 
wire u2__abc_52138_new_n3844_; 
wire u2__abc_52138_new_n3845_; 
wire u2__abc_52138_new_n3846_; 
wire u2__abc_52138_new_n3847_; 
wire u2__abc_52138_new_n3848_; 
wire u2__abc_52138_new_n3849_; 
wire u2__abc_52138_new_n3850_; 
wire u2__abc_52138_new_n3851_; 
wire u2__abc_52138_new_n3852_; 
wire u2__abc_52138_new_n3853_; 
wire u2__abc_52138_new_n3854_; 
wire u2__abc_52138_new_n3855_; 
wire u2__abc_52138_new_n3856_; 
wire u2__abc_52138_new_n3857_; 
wire u2__abc_52138_new_n3858_; 
wire u2__abc_52138_new_n3859_; 
wire u2__abc_52138_new_n3860_; 
wire u2__abc_52138_new_n3861_; 
wire u2__abc_52138_new_n3862_; 
wire u2__abc_52138_new_n3863_; 
wire u2__abc_52138_new_n3864_; 
wire u2__abc_52138_new_n3865_; 
wire u2__abc_52138_new_n3866_; 
wire u2__abc_52138_new_n3867_; 
wire u2__abc_52138_new_n3868_; 
wire u2__abc_52138_new_n3869_; 
wire u2__abc_52138_new_n3870_; 
wire u2__abc_52138_new_n3871_; 
wire u2__abc_52138_new_n3872_; 
wire u2__abc_52138_new_n3873_; 
wire u2__abc_52138_new_n3874_; 
wire u2__abc_52138_new_n3875_; 
wire u2__abc_52138_new_n3876_; 
wire u2__abc_52138_new_n3877_; 
wire u2__abc_52138_new_n3878_; 
wire u2__abc_52138_new_n3879_; 
wire u2__abc_52138_new_n3880_; 
wire u2__abc_52138_new_n3881_; 
wire u2__abc_52138_new_n3882_; 
wire u2__abc_52138_new_n3883_; 
wire u2__abc_52138_new_n3884_; 
wire u2__abc_52138_new_n3885_; 
wire u2__abc_52138_new_n3886_; 
wire u2__abc_52138_new_n3887_; 
wire u2__abc_52138_new_n3888_; 
wire u2__abc_52138_new_n3889_; 
wire u2__abc_52138_new_n3890_; 
wire u2__abc_52138_new_n3891_; 
wire u2__abc_52138_new_n3892_; 
wire u2__abc_52138_new_n3893_; 
wire u2__abc_52138_new_n3894_; 
wire u2__abc_52138_new_n3895_; 
wire u2__abc_52138_new_n3896_; 
wire u2__abc_52138_new_n3897_; 
wire u2__abc_52138_new_n3898_; 
wire u2__abc_52138_new_n3899_; 
wire u2__abc_52138_new_n3900_; 
wire u2__abc_52138_new_n3901_; 
wire u2__abc_52138_new_n3902_; 
wire u2__abc_52138_new_n3903_; 
wire u2__abc_52138_new_n3904_; 
wire u2__abc_52138_new_n3905_; 
wire u2__abc_52138_new_n3906_; 
wire u2__abc_52138_new_n3907_; 
wire u2__abc_52138_new_n3908_; 
wire u2__abc_52138_new_n3909_; 
wire u2__abc_52138_new_n3910_; 
wire u2__abc_52138_new_n3911_; 
wire u2__abc_52138_new_n3912_; 
wire u2__abc_52138_new_n3913_; 
wire u2__abc_52138_new_n3914_; 
wire u2__abc_52138_new_n3915_; 
wire u2__abc_52138_new_n3916_; 
wire u2__abc_52138_new_n3917_; 
wire u2__abc_52138_new_n3918_; 
wire u2__abc_52138_new_n3919_; 
wire u2__abc_52138_new_n3920_; 
wire u2__abc_52138_new_n3921_; 
wire u2__abc_52138_new_n3922_; 
wire u2__abc_52138_new_n3923_; 
wire u2__abc_52138_new_n3924_; 
wire u2__abc_52138_new_n3925_; 
wire u2__abc_52138_new_n3926_; 
wire u2__abc_52138_new_n3927_; 
wire u2__abc_52138_new_n3928_; 
wire u2__abc_52138_new_n3929_; 
wire u2__abc_52138_new_n3930_; 
wire u2__abc_52138_new_n3931_; 
wire u2__abc_52138_new_n3932_; 
wire u2__abc_52138_new_n3933_; 
wire u2__abc_52138_new_n3934_; 
wire u2__abc_52138_new_n3935_; 
wire u2__abc_52138_new_n3936_; 
wire u2__abc_52138_new_n3937_; 
wire u2__abc_52138_new_n3938_; 
wire u2__abc_52138_new_n3939_; 
wire u2__abc_52138_new_n3940_; 
wire u2__abc_52138_new_n3941_; 
wire u2__abc_52138_new_n3942_; 
wire u2__abc_52138_new_n3943_; 
wire u2__abc_52138_new_n3944_; 
wire u2__abc_52138_new_n3945_; 
wire u2__abc_52138_new_n3946_; 
wire u2__abc_52138_new_n3947_; 
wire u2__abc_52138_new_n3948_; 
wire u2__abc_52138_new_n3949_; 
wire u2__abc_52138_new_n3950_; 
wire u2__abc_52138_new_n3951_; 
wire u2__abc_52138_new_n3952_; 
wire u2__abc_52138_new_n3953_; 
wire u2__abc_52138_new_n3954_; 
wire u2__abc_52138_new_n3955_; 
wire u2__abc_52138_new_n3956_; 
wire u2__abc_52138_new_n3957_; 
wire u2__abc_52138_new_n3958_; 
wire u2__abc_52138_new_n3959_; 
wire u2__abc_52138_new_n3960_; 
wire u2__abc_52138_new_n3961_; 
wire u2__abc_52138_new_n3962_; 
wire u2__abc_52138_new_n3963_; 
wire u2__abc_52138_new_n3964_; 
wire u2__abc_52138_new_n3965_; 
wire u2__abc_52138_new_n3966_; 
wire u2__abc_52138_new_n3967_; 
wire u2__abc_52138_new_n3968_; 
wire u2__abc_52138_new_n3969_; 
wire u2__abc_52138_new_n3970_; 
wire u2__abc_52138_new_n3971_; 
wire u2__abc_52138_new_n3972_; 
wire u2__abc_52138_new_n3973_; 
wire u2__abc_52138_new_n3974_; 
wire u2__abc_52138_new_n3975_; 
wire u2__abc_52138_new_n3976_; 
wire u2__abc_52138_new_n3977_; 
wire u2__abc_52138_new_n3978_; 
wire u2__abc_52138_new_n3979_; 
wire u2__abc_52138_new_n3980_; 
wire u2__abc_52138_new_n3981_; 
wire u2__abc_52138_new_n3982_; 
wire u2__abc_52138_new_n3983_; 
wire u2__abc_52138_new_n3984_; 
wire u2__abc_52138_new_n3985_; 
wire u2__abc_52138_new_n3986_; 
wire u2__abc_52138_new_n3987_; 
wire u2__abc_52138_new_n3988_; 
wire u2__abc_52138_new_n3989_; 
wire u2__abc_52138_new_n3990_; 
wire u2__abc_52138_new_n3991_; 
wire u2__abc_52138_new_n3992_; 
wire u2__abc_52138_new_n3993_; 
wire u2__abc_52138_new_n3994_; 
wire u2__abc_52138_new_n3995_; 
wire u2__abc_52138_new_n3996_; 
wire u2__abc_52138_new_n3997_; 
wire u2__abc_52138_new_n3998_; 
wire u2__abc_52138_new_n3999_; 
wire u2__abc_52138_new_n4000_; 
wire u2__abc_52138_new_n4001_; 
wire u2__abc_52138_new_n4002_; 
wire u2__abc_52138_new_n4003_; 
wire u2__abc_52138_new_n4004_; 
wire u2__abc_52138_new_n4005_; 
wire u2__abc_52138_new_n4006_; 
wire u2__abc_52138_new_n4007_; 
wire u2__abc_52138_new_n4008_; 
wire u2__abc_52138_new_n4009_; 
wire u2__abc_52138_new_n4010_; 
wire u2__abc_52138_new_n4011_; 
wire u2__abc_52138_new_n4012_; 
wire u2__abc_52138_new_n4013_; 
wire u2__abc_52138_new_n4014_; 
wire u2__abc_52138_new_n4015_; 
wire u2__abc_52138_new_n4016_; 
wire u2__abc_52138_new_n4017_; 
wire u2__abc_52138_new_n4018_; 
wire u2__abc_52138_new_n4019_; 
wire u2__abc_52138_new_n4020_; 
wire u2__abc_52138_new_n4021_; 
wire u2__abc_52138_new_n4022_; 
wire u2__abc_52138_new_n4023_; 
wire u2__abc_52138_new_n4024_; 
wire u2__abc_52138_new_n4025_; 
wire u2__abc_52138_new_n4026_; 
wire u2__abc_52138_new_n4027_; 
wire u2__abc_52138_new_n4028_; 
wire u2__abc_52138_new_n4029_; 
wire u2__abc_52138_new_n4030_; 
wire u2__abc_52138_new_n4031_; 
wire u2__abc_52138_new_n4032_; 
wire u2__abc_52138_new_n4033_; 
wire u2__abc_52138_new_n4034_; 
wire u2__abc_52138_new_n4035_; 
wire u2__abc_52138_new_n4036_; 
wire u2__abc_52138_new_n4037_; 
wire u2__abc_52138_new_n4038_; 
wire u2__abc_52138_new_n4039_; 
wire u2__abc_52138_new_n4040_; 
wire u2__abc_52138_new_n4041_; 
wire u2__abc_52138_new_n4042_; 
wire u2__abc_52138_new_n4043_; 
wire u2__abc_52138_new_n4044_; 
wire u2__abc_52138_new_n4045_; 
wire u2__abc_52138_new_n4046_; 
wire u2__abc_52138_new_n4047_; 
wire u2__abc_52138_new_n4048_; 
wire u2__abc_52138_new_n4049_; 
wire u2__abc_52138_new_n4050_; 
wire u2__abc_52138_new_n4051_; 
wire u2__abc_52138_new_n4052_; 
wire u2__abc_52138_new_n4053_; 
wire u2__abc_52138_new_n4054_; 
wire u2__abc_52138_new_n4055_; 
wire u2__abc_52138_new_n4056_; 
wire u2__abc_52138_new_n4057_; 
wire u2__abc_52138_new_n4058_; 
wire u2__abc_52138_new_n4059_; 
wire u2__abc_52138_new_n4060_; 
wire u2__abc_52138_new_n4061_; 
wire u2__abc_52138_new_n4062_; 
wire u2__abc_52138_new_n4063_; 
wire u2__abc_52138_new_n4064_; 
wire u2__abc_52138_new_n4065_; 
wire u2__abc_52138_new_n4066_; 
wire u2__abc_52138_new_n4067_; 
wire u2__abc_52138_new_n4068_; 
wire u2__abc_52138_new_n4069_; 
wire u2__abc_52138_new_n4070_; 
wire u2__abc_52138_new_n4071_; 
wire u2__abc_52138_new_n4072_; 
wire u2__abc_52138_new_n4073_; 
wire u2__abc_52138_new_n4074_; 
wire u2__abc_52138_new_n4075_; 
wire u2__abc_52138_new_n4076_; 
wire u2__abc_52138_new_n4077_; 
wire u2__abc_52138_new_n4078_; 
wire u2__abc_52138_new_n4079_; 
wire u2__abc_52138_new_n4080_; 
wire u2__abc_52138_new_n4081_; 
wire u2__abc_52138_new_n4082_; 
wire u2__abc_52138_new_n4083_; 
wire u2__abc_52138_new_n4084_; 
wire u2__abc_52138_new_n4085_; 
wire u2__abc_52138_new_n4086_; 
wire u2__abc_52138_new_n4087_; 
wire u2__abc_52138_new_n4088_; 
wire u2__abc_52138_new_n4089_; 
wire u2__abc_52138_new_n4090_; 
wire u2__abc_52138_new_n4091_; 
wire u2__abc_52138_new_n4092_; 
wire u2__abc_52138_new_n4093_; 
wire u2__abc_52138_new_n4094_; 
wire u2__abc_52138_new_n4095_; 
wire u2__abc_52138_new_n4096_; 
wire u2__abc_52138_new_n4097_; 
wire u2__abc_52138_new_n4098_; 
wire u2__abc_52138_new_n4099_; 
wire u2__abc_52138_new_n4100_; 
wire u2__abc_52138_new_n4101_; 
wire u2__abc_52138_new_n4102_; 
wire u2__abc_52138_new_n4103_; 
wire u2__abc_52138_new_n4104_; 
wire u2__abc_52138_new_n4105_; 
wire u2__abc_52138_new_n4106_; 
wire u2__abc_52138_new_n4107_; 
wire u2__abc_52138_new_n4108_; 
wire u2__abc_52138_new_n4109_; 
wire u2__abc_52138_new_n4110_; 
wire u2__abc_52138_new_n4111_; 
wire u2__abc_52138_new_n4112_; 
wire u2__abc_52138_new_n4113_; 
wire u2__abc_52138_new_n4114_; 
wire u2__abc_52138_new_n4115_; 
wire u2__abc_52138_new_n4116_; 
wire u2__abc_52138_new_n4117_; 
wire u2__abc_52138_new_n4118_; 
wire u2__abc_52138_new_n4119_; 
wire u2__abc_52138_new_n4120_; 
wire u2__abc_52138_new_n4121_; 
wire u2__abc_52138_new_n4122_; 
wire u2__abc_52138_new_n4123_; 
wire u2__abc_52138_new_n4124_; 
wire u2__abc_52138_new_n4125_; 
wire u2__abc_52138_new_n4126_; 
wire u2__abc_52138_new_n4127_; 
wire u2__abc_52138_new_n4128_; 
wire u2__abc_52138_new_n4129_; 
wire u2__abc_52138_new_n4130_; 
wire u2__abc_52138_new_n4131_; 
wire u2__abc_52138_new_n4132_; 
wire u2__abc_52138_new_n4133_; 
wire u2__abc_52138_new_n4134_; 
wire u2__abc_52138_new_n4135_; 
wire u2__abc_52138_new_n4136_; 
wire u2__abc_52138_new_n4137_; 
wire u2__abc_52138_new_n4138_; 
wire u2__abc_52138_new_n4139_; 
wire u2__abc_52138_new_n4140_; 
wire u2__abc_52138_new_n4141_; 
wire u2__abc_52138_new_n4142_; 
wire u2__abc_52138_new_n4143_; 
wire u2__abc_52138_new_n4144_; 
wire u2__abc_52138_new_n4145_; 
wire u2__abc_52138_new_n4146_; 
wire u2__abc_52138_new_n4147_; 
wire u2__abc_52138_new_n4148_; 
wire u2__abc_52138_new_n4149_; 
wire u2__abc_52138_new_n4150_; 
wire u2__abc_52138_new_n4151_; 
wire u2__abc_52138_new_n4152_; 
wire u2__abc_52138_new_n4153_; 
wire u2__abc_52138_new_n4154_; 
wire u2__abc_52138_new_n4155_; 
wire u2__abc_52138_new_n4156_; 
wire u2__abc_52138_new_n4157_; 
wire u2__abc_52138_new_n4158_; 
wire u2__abc_52138_new_n4159_; 
wire u2__abc_52138_new_n4160_; 
wire u2__abc_52138_new_n4161_; 
wire u2__abc_52138_new_n4162_; 
wire u2__abc_52138_new_n4163_; 
wire u2__abc_52138_new_n4164_; 
wire u2__abc_52138_new_n4165_; 
wire u2__abc_52138_new_n4166_; 
wire u2__abc_52138_new_n4167_; 
wire u2__abc_52138_new_n4168_; 
wire u2__abc_52138_new_n4169_; 
wire u2__abc_52138_new_n4170_; 
wire u2__abc_52138_new_n4171_; 
wire u2__abc_52138_new_n4172_; 
wire u2__abc_52138_new_n4173_; 
wire u2__abc_52138_new_n4174_; 
wire u2__abc_52138_new_n4175_; 
wire u2__abc_52138_new_n4176_; 
wire u2__abc_52138_new_n4177_; 
wire u2__abc_52138_new_n4178_; 
wire u2__abc_52138_new_n4179_; 
wire u2__abc_52138_new_n4180_; 
wire u2__abc_52138_new_n4181_; 
wire u2__abc_52138_new_n4182_; 
wire u2__abc_52138_new_n4183_; 
wire u2__abc_52138_new_n4184_; 
wire u2__abc_52138_new_n4185_; 
wire u2__abc_52138_new_n4186_; 
wire u2__abc_52138_new_n4187_; 
wire u2__abc_52138_new_n4188_; 
wire u2__abc_52138_new_n4189_; 
wire u2__abc_52138_new_n4190_; 
wire u2__abc_52138_new_n4191_; 
wire u2__abc_52138_new_n4192_; 
wire u2__abc_52138_new_n4193_; 
wire u2__abc_52138_new_n4194_; 
wire u2__abc_52138_new_n4195_; 
wire u2__abc_52138_new_n4196_; 
wire u2__abc_52138_new_n4197_; 
wire u2__abc_52138_new_n4198_; 
wire u2__abc_52138_new_n4199_; 
wire u2__abc_52138_new_n4200_; 
wire u2__abc_52138_new_n4201_; 
wire u2__abc_52138_new_n4202_; 
wire u2__abc_52138_new_n4203_; 
wire u2__abc_52138_new_n4204_; 
wire u2__abc_52138_new_n4205_; 
wire u2__abc_52138_new_n4206_; 
wire u2__abc_52138_new_n4207_; 
wire u2__abc_52138_new_n4208_; 
wire u2__abc_52138_new_n4209_; 
wire u2__abc_52138_new_n4210_; 
wire u2__abc_52138_new_n4211_; 
wire u2__abc_52138_new_n4212_; 
wire u2__abc_52138_new_n4213_; 
wire u2__abc_52138_new_n4214_; 
wire u2__abc_52138_new_n4215_; 
wire u2__abc_52138_new_n4216_; 
wire u2__abc_52138_new_n4217_; 
wire u2__abc_52138_new_n4218_; 
wire u2__abc_52138_new_n4219_; 
wire u2__abc_52138_new_n4220_; 
wire u2__abc_52138_new_n4221_; 
wire u2__abc_52138_new_n4222_; 
wire u2__abc_52138_new_n4223_; 
wire u2__abc_52138_new_n4224_; 
wire u2__abc_52138_new_n4225_; 
wire u2__abc_52138_new_n4226_; 
wire u2__abc_52138_new_n4227_; 
wire u2__abc_52138_new_n4228_; 
wire u2__abc_52138_new_n4229_; 
wire u2__abc_52138_new_n4230_; 
wire u2__abc_52138_new_n4231_; 
wire u2__abc_52138_new_n4232_; 
wire u2__abc_52138_new_n4233_; 
wire u2__abc_52138_new_n4234_; 
wire u2__abc_52138_new_n4235_; 
wire u2__abc_52138_new_n4236_; 
wire u2__abc_52138_new_n4237_; 
wire u2__abc_52138_new_n4238_; 
wire u2__abc_52138_new_n4239_; 
wire u2__abc_52138_new_n4240_; 
wire u2__abc_52138_new_n4241_; 
wire u2__abc_52138_new_n4242_; 
wire u2__abc_52138_new_n4243_; 
wire u2__abc_52138_new_n4244_; 
wire u2__abc_52138_new_n4245_; 
wire u2__abc_52138_new_n4246_; 
wire u2__abc_52138_new_n4247_; 
wire u2__abc_52138_new_n4248_; 
wire u2__abc_52138_new_n4249_; 
wire u2__abc_52138_new_n4250_; 
wire u2__abc_52138_new_n4251_; 
wire u2__abc_52138_new_n4252_; 
wire u2__abc_52138_new_n4253_; 
wire u2__abc_52138_new_n4254_; 
wire u2__abc_52138_new_n4255_; 
wire u2__abc_52138_new_n4256_; 
wire u2__abc_52138_new_n4257_; 
wire u2__abc_52138_new_n4258_; 
wire u2__abc_52138_new_n4259_; 
wire u2__abc_52138_new_n4260_; 
wire u2__abc_52138_new_n4261_; 
wire u2__abc_52138_new_n4262_; 
wire u2__abc_52138_new_n4263_; 
wire u2__abc_52138_new_n4264_; 
wire u2__abc_52138_new_n4265_; 
wire u2__abc_52138_new_n4266_; 
wire u2__abc_52138_new_n4267_; 
wire u2__abc_52138_new_n4268_; 
wire u2__abc_52138_new_n4269_; 
wire u2__abc_52138_new_n4270_; 
wire u2__abc_52138_new_n4271_; 
wire u2__abc_52138_new_n4272_; 
wire u2__abc_52138_new_n4273_; 
wire u2__abc_52138_new_n4274_; 
wire u2__abc_52138_new_n4275_; 
wire u2__abc_52138_new_n4276_; 
wire u2__abc_52138_new_n4277_; 
wire u2__abc_52138_new_n4278_; 
wire u2__abc_52138_new_n4279_; 
wire u2__abc_52138_new_n4280_; 
wire u2__abc_52138_new_n4281_; 
wire u2__abc_52138_new_n4282_; 
wire u2__abc_52138_new_n4283_; 
wire u2__abc_52138_new_n4284_; 
wire u2__abc_52138_new_n4285_; 
wire u2__abc_52138_new_n4286_; 
wire u2__abc_52138_new_n4287_; 
wire u2__abc_52138_new_n4288_; 
wire u2__abc_52138_new_n4289_; 
wire u2__abc_52138_new_n4290_; 
wire u2__abc_52138_new_n4291_; 
wire u2__abc_52138_new_n4292_; 
wire u2__abc_52138_new_n4293_; 
wire u2__abc_52138_new_n4294_; 
wire u2__abc_52138_new_n4295_; 
wire u2__abc_52138_new_n4296_; 
wire u2__abc_52138_new_n4297_; 
wire u2__abc_52138_new_n4298_; 
wire u2__abc_52138_new_n4299_; 
wire u2__abc_52138_new_n4300_; 
wire u2__abc_52138_new_n4301_; 
wire u2__abc_52138_new_n4302_; 
wire u2__abc_52138_new_n4303_; 
wire u2__abc_52138_new_n4304_; 
wire u2__abc_52138_new_n4305_; 
wire u2__abc_52138_new_n4306_; 
wire u2__abc_52138_new_n4307_; 
wire u2__abc_52138_new_n4308_; 
wire u2__abc_52138_new_n4309_; 
wire u2__abc_52138_new_n4310_; 
wire u2__abc_52138_new_n4311_; 
wire u2__abc_52138_new_n4312_; 
wire u2__abc_52138_new_n4313_; 
wire u2__abc_52138_new_n4314_; 
wire u2__abc_52138_new_n4315_; 
wire u2__abc_52138_new_n4316_; 
wire u2__abc_52138_new_n4317_; 
wire u2__abc_52138_new_n4318_; 
wire u2__abc_52138_new_n4319_; 
wire u2__abc_52138_new_n4320_; 
wire u2__abc_52138_new_n4321_; 
wire u2__abc_52138_new_n4322_; 
wire u2__abc_52138_new_n4323_; 
wire u2__abc_52138_new_n4324_; 
wire u2__abc_52138_new_n4325_; 
wire u2__abc_52138_new_n4326_; 
wire u2__abc_52138_new_n4327_; 
wire u2__abc_52138_new_n4328_; 
wire u2__abc_52138_new_n4329_; 
wire u2__abc_52138_new_n4330_; 
wire u2__abc_52138_new_n4331_; 
wire u2__abc_52138_new_n4332_; 
wire u2__abc_52138_new_n4333_; 
wire u2__abc_52138_new_n4334_; 
wire u2__abc_52138_new_n4335_; 
wire u2__abc_52138_new_n4336_; 
wire u2__abc_52138_new_n4337_; 
wire u2__abc_52138_new_n4338_; 
wire u2__abc_52138_new_n4339_; 
wire u2__abc_52138_new_n4340_; 
wire u2__abc_52138_new_n4341_; 
wire u2__abc_52138_new_n4342_; 
wire u2__abc_52138_new_n4343_; 
wire u2__abc_52138_new_n4344_; 
wire u2__abc_52138_new_n4345_; 
wire u2__abc_52138_new_n4346_; 
wire u2__abc_52138_new_n4347_; 
wire u2__abc_52138_new_n4348_; 
wire u2__abc_52138_new_n4349_; 
wire u2__abc_52138_new_n4350_; 
wire u2__abc_52138_new_n4351_; 
wire u2__abc_52138_new_n4352_; 
wire u2__abc_52138_new_n4353_; 
wire u2__abc_52138_new_n4354_; 
wire u2__abc_52138_new_n4355_; 
wire u2__abc_52138_new_n4356_; 
wire u2__abc_52138_new_n4357_; 
wire u2__abc_52138_new_n4358_; 
wire u2__abc_52138_new_n4359_; 
wire u2__abc_52138_new_n4360_; 
wire u2__abc_52138_new_n4361_; 
wire u2__abc_52138_new_n4362_; 
wire u2__abc_52138_new_n4363_; 
wire u2__abc_52138_new_n4364_; 
wire u2__abc_52138_new_n4365_; 
wire u2__abc_52138_new_n4366_; 
wire u2__abc_52138_new_n4367_; 
wire u2__abc_52138_new_n4368_; 
wire u2__abc_52138_new_n4369_; 
wire u2__abc_52138_new_n4370_; 
wire u2__abc_52138_new_n4371_; 
wire u2__abc_52138_new_n4372_; 
wire u2__abc_52138_new_n4373_; 
wire u2__abc_52138_new_n4374_; 
wire u2__abc_52138_new_n4375_; 
wire u2__abc_52138_new_n4376_; 
wire u2__abc_52138_new_n4377_; 
wire u2__abc_52138_new_n4378_; 
wire u2__abc_52138_new_n4379_; 
wire u2__abc_52138_new_n4380_; 
wire u2__abc_52138_new_n4381_; 
wire u2__abc_52138_new_n4382_; 
wire u2__abc_52138_new_n4383_; 
wire u2__abc_52138_new_n4384_; 
wire u2__abc_52138_new_n4385_; 
wire u2__abc_52138_new_n4386_; 
wire u2__abc_52138_new_n4387_; 
wire u2__abc_52138_new_n4388_; 
wire u2__abc_52138_new_n4389_; 
wire u2__abc_52138_new_n4390_; 
wire u2__abc_52138_new_n4391_; 
wire u2__abc_52138_new_n4392_; 
wire u2__abc_52138_new_n4393_; 
wire u2__abc_52138_new_n4394_; 
wire u2__abc_52138_new_n4395_; 
wire u2__abc_52138_new_n4396_; 
wire u2__abc_52138_new_n4397_; 
wire u2__abc_52138_new_n4398_; 
wire u2__abc_52138_new_n4399_; 
wire u2__abc_52138_new_n4400_; 
wire u2__abc_52138_new_n4401_; 
wire u2__abc_52138_new_n4402_; 
wire u2__abc_52138_new_n4403_; 
wire u2__abc_52138_new_n4404_; 
wire u2__abc_52138_new_n4405_; 
wire u2__abc_52138_new_n4406_; 
wire u2__abc_52138_new_n4407_; 
wire u2__abc_52138_new_n4408_; 
wire u2__abc_52138_new_n4409_; 
wire u2__abc_52138_new_n4410_; 
wire u2__abc_52138_new_n4411_; 
wire u2__abc_52138_new_n4412_; 
wire u2__abc_52138_new_n4413_; 
wire u2__abc_52138_new_n4414_; 
wire u2__abc_52138_new_n4415_; 
wire u2__abc_52138_new_n4416_; 
wire u2__abc_52138_new_n4417_; 
wire u2__abc_52138_new_n4418_; 
wire u2__abc_52138_new_n4419_; 
wire u2__abc_52138_new_n4420_; 
wire u2__abc_52138_new_n4421_; 
wire u2__abc_52138_new_n4422_; 
wire u2__abc_52138_new_n4423_; 
wire u2__abc_52138_new_n4424_; 
wire u2__abc_52138_new_n4425_; 
wire u2__abc_52138_new_n4426_; 
wire u2__abc_52138_new_n4427_; 
wire u2__abc_52138_new_n4428_; 
wire u2__abc_52138_new_n4429_; 
wire u2__abc_52138_new_n4430_; 
wire u2__abc_52138_new_n4431_; 
wire u2__abc_52138_new_n4432_; 
wire u2__abc_52138_new_n4433_; 
wire u2__abc_52138_new_n4434_; 
wire u2__abc_52138_new_n4435_; 
wire u2__abc_52138_new_n4436_; 
wire u2__abc_52138_new_n4437_; 
wire u2__abc_52138_new_n4438_; 
wire u2__abc_52138_new_n4439_; 
wire u2__abc_52138_new_n4440_; 
wire u2__abc_52138_new_n4441_; 
wire u2__abc_52138_new_n4442_; 
wire u2__abc_52138_new_n4443_; 
wire u2__abc_52138_new_n4444_; 
wire u2__abc_52138_new_n4445_; 
wire u2__abc_52138_new_n4446_; 
wire u2__abc_52138_new_n4447_; 
wire u2__abc_52138_new_n4448_; 
wire u2__abc_52138_new_n4449_; 
wire u2__abc_52138_new_n4450_; 
wire u2__abc_52138_new_n4451_; 
wire u2__abc_52138_new_n4452_; 
wire u2__abc_52138_new_n4453_; 
wire u2__abc_52138_new_n4454_; 
wire u2__abc_52138_new_n4455_; 
wire u2__abc_52138_new_n4456_; 
wire u2__abc_52138_new_n4457_; 
wire u2__abc_52138_new_n4458_; 
wire u2__abc_52138_new_n4459_; 
wire u2__abc_52138_new_n4460_; 
wire u2__abc_52138_new_n4461_; 
wire u2__abc_52138_new_n4462_; 
wire u2__abc_52138_new_n4463_; 
wire u2__abc_52138_new_n4464_; 
wire u2__abc_52138_new_n4465_; 
wire u2__abc_52138_new_n4466_; 
wire u2__abc_52138_new_n4467_; 
wire u2__abc_52138_new_n4468_; 
wire u2__abc_52138_new_n4469_; 
wire u2__abc_52138_new_n4470_; 
wire u2__abc_52138_new_n4471_; 
wire u2__abc_52138_new_n4472_; 
wire u2__abc_52138_new_n4473_; 
wire u2__abc_52138_new_n4474_; 
wire u2__abc_52138_new_n4475_; 
wire u2__abc_52138_new_n4476_; 
wire u2__abc_52138_new_n4477_; 
wire u2__abc_52138_new_n4478_; 
wire u2__abc_52138_new_n4479_; 
wire u2__abc_52138_new_n4480_; 
wire u2__abc_52138_new_n4481_; 
wire u2__abc_52138_new_n4482_; 
wire u2__abc_52138_new_n4483_; 
wire u2__abc_52138_new_n4484_; 
wire u2__abc_52138_new_n4485_; 
wire u2__abc_52138_new_n4486_; 
wire u2__abc_52138_new_n4487_; 
wire u2__abc_52138_new_n4488_; 
wire u2__abc_52138_new_n4489_; 
wire u2__abc_52138_new_n4490_; 
wire u2__abc_52138_new_n4491_; 
wire u2__abc_52138_new_n4492_; 
wire u2__abc_52138_new_n4493_; 
wire u2__abc_52138_new_n4494_; 
wire u2__abc_52138_new_n4495_; 
wire u2__abc_52138_new_n4496_; 
wire u2__abc_52138_new_n4497_; 
wire u2__abc_52138_new_n4498_; 
wire u2__abc_52138_new_n4499_; 
wire u2__abc_52138_new_n4500_; 
wire u2__abc_52138_new_n4501_; 
wire u2__abc_52138_new_n4502_; 
wire u2__abc_52138_new_n4503_; 
wire u2__abc_52138_new_n4504_; 
wire u2__abc_52138_new_n4505_; 
wire u2__abc_52138_new_n4506_; 
wire u2__abc_52138_new_n4507_; 
wire u2__abc_52138_new_n4508_; 
wire u2__abc_52138_new_n4509_; 
wire u2__abc_52138_new_n4510_; 
wire u2__abc_52138_new_n4511_; 
wire u2__abc_52138_new_n4512_; 
wire u2__abc_52138_new_n4513_; 
wire u2__abc_52138_new_n4514_; 
wire u2__abc_52138_new_n4515_; 
wire u2__abc_52138_new_n4516_; 
wire u2__abc_52138_new_n4517_; 
wire u2__abc_52138_new_n4518_; 
wire u2__abc_52138_new_n4519_; 
wire u2__abc_52138_new_n4520_; 
wire u2__abc_52138_new_n4521_; 
wire u2__abc_52138_new_n4522_; 
wire u2__abc_52138_new_n4523_; 
wire u2__abc_52138_new_n4524_; 
wire u2__abc_52138_new_n4525_; 
wire u2__abc_52138_new_n4526_; 
wire u2__abc_52138_new_n4527_; 
wire u2__abc_52138_new_n4528_; 
wire u2__abc_52138_new_n4529_; 
wire u2__abc_52138_new_n4530_; 
wire u2__abc_52138_new_n4531_; 
wire u2__abc_52138_new_n4532_; 
wire u2__abc_52138_new_n4533_; 
wire u2__abc_52138_new_n4534_; 
wire u2__abc_52138_new_n4535_; 
wire u2__abc_52138_new_n4536_; 
wire u2__abc_52138_new_n4537_; 
wire u2__abc_52138_new_n4538_; 
wire u2__abc_52138_new_n4539_; 
wire u2__abc_52138_new_n4540_; 
wire u2__abc_52138_new_n4541_; 
wire u2__abc_52138_new_n4542_; 
wire u2__abc_52138_new_n4543_; 
wire u2__abc_52138_new_n4544_; 
wire u2__abc_52138_new_n4545_; 
wire u2__abc_52138_new_n4546_; 
wire u2__abc_52138_new_n4547_; 
wire u2__abc_52138_new_n4548_; 
wire u2__abc_52138_new_n4549_; 
wire u2__abc_52138_new_n4550_; 
wire u2__abc_52138_new_n4551_; 
wire u2__abc_52138_new_n4552_; 
wire u2__abc_52138_new_n4553_; 
wire u2__abc_52138_new_n4554_; 
wire u2__abc_52138_new_n4555_; 
wire u2__abc_52138_new_n4556_; 
wire u2__abc_52138_new_n4557_; 
wire u2__abc_52138_new_n4558_; 
wire u2__abc_52138_new_n4559_; 
wire u2__abc_52138_new_n4560_; 
wire u2__abc_52138_new_n4561_; 
wire u2__abc_52138_new_n4562_; 
wire u2__abc_52138_new_n4563_; 
wire u2__abc_52138_new_n4564_; 
wire u2__abc_52138_new_n4565_; 
wire u2__abc_52138_new_n4566_; 
wire u2__abc_52138_new_n4567_; 
wire u2__abc_52138_new_n4568_; 
wire u2__abc_52138_new_n4569_; 
wire u2__abc_52138_new_n4570_; 
wire u2__abc_52138_new_n4571_; 
wire u2__abc_52138_new_n4572_; 
wire u2__abc_52138_new_n4573_; 
wire u2__abc_52138_new_n4574_; 
wire u2__abc_52138_new_n4575_; 
wire u2__abc_52138_new_n4576_; 
wire u2__abc_52138_new_n4577_; 
wire u2__abc_52138_new_n4578_; 
wire u2__abc_52138_new_n4579_; 
wire u2__abc_52138_new_n4580_; 
wire u2__abc_52138_new_n4581_; 
wire u2__abc_52138_new_n4582_; 
wire u2__abc_52138_new_n4583_; 
wire u2__abc_52138_new_n4584_; 
wire u2__abc_52138_new_n4585_; 
wire u2__abc_52138_new_n4586_; 
wire u2__abc_52138_new_n4587_; 
wire u2__abc_52138_new_n4588_; 
wire u2__abc_52138_new_n4589_; 
wire u2__abc_52138_new_n4590_; 
wire u2__abc_52138_new_n4591_; 
wire u2__abc_52138_new_n4592_; 
wire u2__abc_52138_new_n4593_; 
wire u2__abc_52138_new_n4594_; 
wire u2__abc_52138_new_n4595_; 
wire u2__abc_52138_new_n4596_; 
wire u2__abc_52138_new_n4597_; 
wire u2__abc_52138_new_n4598_; 
wire u2__abc_52138_new_n4599_; 
wire u2__abc_52138_new_n4600_; 
wire u2__abc_52138_new_n4601_; 
wire u2__abc_52138_new_n4602_; 
wire u2__abc_52138_new_n4603_; 
wire u2__abc_52138_new_n4604_; 
wire u2__abc_52138_new_n4605_; 
wire u2__abc_52138_new_n4606_; 
wire u2__abc_52138_new_n4607_; 
wire u2__abc_52138_new_n4608_; 
wire u2__abc_52138_new_n4609_; 
wire u2__abc_52138_new_n4610_; 
wire u2__abc_52138_new_n4611_; 
wire u2__abc_52138_new_n4612_; 
wire u2__abc_52138_new_n4613_; 
wire u2__abc_52138_new_n4614_; 
wire u2__abc_52138_new_n4615_; 
wire u2__abc_52138_new_n4616_; 
wire u2__abc_52138_new_n4617_; 
wire u2__abc_52138_new_n4618_; 
wire u2__abc_52138_new_n4619_; 
wire u2__abc_52138_new_n4620_; 
wire u2__abc_52138_new_n4621_; 
wire u2__abc_52138_new_n4622_; 
wire u2__abc_52138_new_n4623_; 
wire u2__abc_52138_new_n4624_; 
wire u2__abc_52138_new_n4625_; 
wire u2__abc_52138_new_n4626_; 
wire u2__abc_52138_new_n4627_; 
wire u2__abc_52138_new_n4628_; 
wire u2__abc_52138_new_n4629_; 
wire u2__abc_52138_new_n4630_; 
wire u2__abc_52138_new_n4631_; 
wire u2__abc_52138_new_n4632_; 
wire u2__abc_52138_new_n4633_; 
wire u2__abc_52138_new_n4634_; 
wire u2__abc_52138_new_n4635_; 
wire u2__abc_52138_new_n4636_; 
wire u2__abc_52138_new_n4637_; 
wire u2__abc_52138_new_n4638_; 
wire u2__abc_52138_new_n4639_; 
wire u2__abc_52138_new_n4640_; 
wire u2__abc_52138_new_n4641_; 
wire u2__abc_52138_new_n4642_; 
wire u2__abc_52138_new_n4643_; 
wire u2__abc_52138_new_n4644_; 
wire u2__abc_52138_new_n4645_; 
wire u2__abc_52138_new_n4646_; 
wire u2__abc_52138_new_n4647_; 
wire u2__abc_52138_new_n4648_; 
wire u2__abc_52138_new_n4649_; 
wire u2__abc_52138_new_n4650_; 
wire u2__abc_52138_new_n4651_; 
wire u2__abc_52138_new_n4652_; 
wire u2__abc_52138_new_n4653_; 
wire u2__abc_52138_new_n4654_; 
wire u2__abc_52138_new_n4655_; 
wire u2__abc_52138_new_n4656_; 
wire u2__abc_52138_new_n4657_; 
wire u2__abc_52138_new_n4658_; 
wire u2__abc_52138_new_n4659_; 
wire u2__abc_52138_new_n4660_; 
wire u2__abc_52138_new_n4661_; 
wire u2__abc_52138_new_n4662_; 
wire u2__abc_52138_new_n4663_; 
wire u2__abc_52138_new_n4664_; 
wire u2__abc_52138_new_n4665_; 
wire u2__abc_52138_new_n4666_; 
wire u2__abc_52138_new_n4667_; 
wire u2__abc_52138_new_n4668_; 
wire u2__abc_52138_new_n4669_; 
wire u2__abc_52138_new_n4670_; 
wire u2__abc_52138_new_n4671_; 
wire u2__abc_52138_new_n4672_; 
wire u2__abc_52138_new_n4673_; 
wire u2__abc_52138_new_n4674_; 
wire u2__abc_52138_new_n4675_; 
wire u2__abc_52138_new_n4676_; 
wire u2__abc_52138_new_n4677_; 
wire u2__abc_52138_new_n4678_; 
wire u2__abc_52138_new_n4679_; 
wire u2__abc_52138_new_n4680_; 
wire u2__abc_52138_new_n4681_; 
wire u2__abc_52138_new_n4682_; 
wire u2__abc_52138_new_n4683_; 
wire u2__abc_52138_new_n4684_; 
wire u2__abc_52138_new_n4685_; 
wire u2__abc_52138_new_n4686_; 
wire u2__abc_52138_new_n4687_; 
wire u2__abc_52138_new_n4688_; 
wire u2__abc_52138_new_n4689_; 
wire u2__abc_52138_new_n4690_; 
wire u2__abc_52138_new_n4691_; 
wire u2__abc_52138_new_n4692_; 
wire u2__abc_52138_new_n4693_; 
wire u2__abc_52138_new_n4694_; 
wire u2__abc_52138_new_n4695_; 
wire u2__abc_52138_new_n4696_; 
wire u2__abc_52138_new_n4697_; 
wire u2__abc_52138_new_n4698_; 
wire u2__abc_52138_new_n4699_; 
wire u2__abc_52138_new_n4700_; 
wire u2__abc_52138_new_n4701_; 
wire u2__abc_52138_new_n4702_; 
wire u2__abc_52138_new_n4703_; 
wire u2__abc_52138_new_n4704_; 
wire u2__abc_52138_new_n4705_; 
wire u2__abc_52138_new_n4706_; 
wire u2__abc_52138_new_n4707_; 
wire u2__abc_52138_new_n4708_; 
wire u2__abc_52138_new_n4709_; 
wire u2__abc_52138_new_n4710_; 
wire u2__abc_52138_new_n4711_; 
wire u2__abc_52138_new_n4712_; 
wire u2__abc_52138_new_n4713_; 
wire u2__abc_52138_new_n4714_; 
wire u2__abc_52138_new_n4715_; 
wire u2__abc_52138_new_n4716_; 
wire u2__abc_52138_new_n4717_; 
wire u2__abc_52138_new_n4718_; 
wire u2__abc_52138_new_n4719_; 
wire u2__abc_52138_new_n4720_; 
wire u2__abc_52138_new_n4721_; 
wire u2__abc_52138_new_n4722_; 
wire u2__abc_52138_new_n4723_; 
wire u2__abc_52138_new_n4724_; 
wire u2__abc_52138_new_n4725_; 
wire u2__abc_52138_new_n4726_; 
wire u2__abc_52138_new_n4727_; 
wire u2__abc_52138_new_n4728_; 
wire u2__abc_52138_new_n4729_; 
wire u2__abc_52138_new_n4730_; 
wire u2__abc_52138_new_n4731_; 
wire u2__abc_52138_new_n4732_; 
wire u2__abc_52138_new_n4733_; 
wire u2__abc_52138_new_n4734_; 
wire u2__abc_52138_new_n4735_; 
wire u2__abc_52138_new_n4736_; 
wire u2__abc_52138_new_n4737_; 
wire u2__abc_52138_new_n4738_; 
wire u2__abc_52138_new_n4739_; 
wire u2__abc_52138_new_n4740_; 
wire u2__abc_52138_new_n4741_; 
wire u2__abc_52138_new_n4742_; 
wire u2__abc_52138_new_n4743_; 
wire u2__abc_52138_new_n4744_; 
wire u2__abc_52138_new_n4745_; 
wire u2__abc_52138_new_n4746_; 
wire u2__abc_52138_new_n4747_; 
wire u2__abc_52138_new_n4748_; 
wire u2__abc_52138_new_n4749_; 
wire u2__abc_52138_new_n4750_; 
wire u2__abc_52138_new_n4751_; 
wire u2__abc_52138_new_n4752_; 
wire u2__abc_52138_new_n4753_; 
wire u2__abc_52138_new_n4754_; 
wire u2__abc_52138_new_n4755_; 
wire u2__abc_52138_new_n4756_; 
wire u2__abc_52138_new_n4757_; 
wire u2__abc_52138_new_n4758_; 
wire u2__abc_52138_new_n4759_; 
wire u2__abc_52138_new_n4760_; 
wire u2__abc_52138_new_n4761_; 
wire u2__abc_52138_new_n4762_; 
wire u2__abc_52138_new_n4763_; 
wire u2__abc_52138_new_n4764_; 
wire u2__abc_52138_new_n4765_; 
wire u2__abc_52138_new_n4766_; 
wire u2__abc_52138_new_n4767_; 
wire u2__abc_52138_new_n4768_; 
wire u2__abc_52138_new_n4769_; 
wire u2__abc_52138_new_n4770_; 
wire u2__abc_52138_new_n4771_; 
wire u2__abc_52138_new_n4772_; 
wire u2__abc_52138_new_n4773_; 
wire u2__abc_52138_new_n4774_; 
wire u2__abc_52138_new_n4775_; 
wire u2__abc_52138_new_n4776_; 
wire u2__abc_52138_new_n4777_; 
wire u2__abc_52138_new_n4778_; 
wire u2__abc_52138_new_n4779_; 
wire u2__abc_52138_new_n4780_; 
wire u2__abc_52138_new_n4781_; 
wire u2__abc_52138_new_n4782_; 
wire u2__abc_52138_new_n4783_; 
wire u2__abc_52138_new_n4784_; 
wire u2__abc_52138_new_n4785_; 
wire u2__abc_52138_new_n4786_; 
wire u2__abc_52138_new_n4787_; 
wire u2__abc_52138_new_n4788_; 
wire u2__abc_52138_new_n4789_; 
wire u2__abc_52138_new_n4790_; 
wire u2__abc_52138_new_n4791_; 
wire u2__abc_52138_new_n4792_; 
wire u2__abc_52138_new_n4793_; 
wire u2__abc_52138_new_n4794_; 
wire u2__abc_52138_new_n4795_; 
wire u2__abc_52138_new_n4796_; 
wire u2__abc_52138_new_n4797_; 
wire u2__abc_52138_new_n4798_; 
wire u2__abc_52138_new_n4799_; 
wire u2__abc_52138_new_n4800_; 
wire u2__abc_52138_new_n4801_; 
wire u2__abc_52138_new_n4802_; 
wire u2__abc_52138_new_n4803_; 
wire u2__abc_52138_new_n4804_; 
wire u2__abc_52138_new_n4805_; 
wire u2__abc_52138_new_n4806_; 
wire u2__abc_52138_new_n4807_; 
wire u2__abc_52138_new_n4808_; 
wire u2__abc_52138_new_n4809_; 
wire u2__abc_52138_new_n4810_; 
wire u2__abc_52138_new_n4811_; 
wire u2__abc_52138_new_n4812_; 
wire u2__abc_52138_new_n4813_; 
wire u2__abc_52138_new_n4814_; 
wire u2__abc_52138_new_n4815_; 
wire u2__abc_52138_new_n4816_; 
wire u2__abc_52138_new_n4817_; 
wire u2__abc_52138_new_n4818_; 
wire u2__abc_52138_new_n4819_; 
wire u2__abc_52138_new_n4820_; 
wire u2__abc_52138_new_n4821_; 
wire u2__abc_52138_new_n4822_; 
wire u2__abc_52138_new_n4823_; 
wire u2__abc_52138_new_n4824_; 
wire u2__abc_52138_new_n4825_; 
wire u2__abc_52138_new_n4826_; 
wire u2__abc_52138_new_n4827_; 
wire u2__abc_52138_new_n4828_; 
wire u2__abc_52138_new_n4829_; 
wire u2__abc_52138_new_n4830_; 
wire u2__abc_52138_new_n4831_; 
wire u2__abc_52138_new_n4832_; 
wire u2__abc_52138_new_n4833_; 
wire u2__abc_52138_new_n4834_; 
wire u2__abc_52138_new_n4835_; 
wire u2__abc_52138_new_n4836_; 
wire u2__abc_52138_new_n4837_; 
wire u2__abc_52138_new_n4838_; 
wire u2__abc_52138_new_n4839_; 
wire u2__abc_52138_new_n4840_; 
wire u2__abc_52138_new_n4841_; 
wire u2__abc_52138_new_n4842_; 
wire u2__abc_52138_new_n4843_; 
wire u2__abc_52138_new_n4844_; 
wire u2__abc_52138_new_n4845_; 
wire u2__abc_52138_new_n4846_; 
wire u2__abc_52138_new_n4847_; 
wire u2__abc_52138_new_n4848_; 
wire u2__abc_52138_new_n4849_; 
wire u2__abc_52138_new_n4850_; 
wire u2__abc_52138_new_n4851_; 
wire u2__abc_52138_new_n4852_; 
wire u2__abc_52138_new_n4853_; 
wire u2__abc_52138_new_n4854_; 
wire u2__abc_52138_new_n4855_; 
wire u2__abc_52138_new_n4856_; 
wire u2__abc_52138_new_n4857_; 
wire u2__abc_52138_new_n4858_; 
wire u2__abc_52138_new_n4859_; 
wire u2__abc_52138_new_n4860_; 
wire u2__abc_52138_new_n4861_; 
wire u2__abc_52138_new_n4862_; 
wire u2__abc_52138_new_n4863_; 
wire u2__abc_52138_new_n4864_; 
wire u2__abc_52138_new_n4865_; 
wire u2__abc_52138_new_n4866_; 
wire u2__abc_52138_new_n4867_; 
wire u2__abc_52138_new_n4868_; 
wire u2__abc_52138_new_n4869_; 
wire u2__abc_52138_new_n4870_; 
wire u2__abc_52138_new_n4871_; 
wire u2__abc_52138_new_n4872_; 
wire u2__abc_52138_new_n4873_; 
wire u2__abc_52138_new_n4874_; 
wire u2__abc_52138_new_n4875_; 
wire u2__abc_52138_new_n4876_; 
wire u2__abc_52138_new_n4877_; 
wire u2__abc_52138_new_n4878_; 
wire u2__abc_52138_new_n4879_; 
wire u2__abc_52138_new_n4880_; 
wire u2__abc_52138_new_n4881_; 
wire u2__abc_52138_new_n4882_; 
wire u2__abc_52138_new_n4883_; 
wire u2__abc_52138_new_n4884_; 
wire u2__abc_52138_new_n4885_; 
wire u2__abc_52138_new_n4886_; 
wire u2__abc_52138_new_n4887_; 
wire u2__abc_52138_new_n4888_; 
wire u2__abc_52138_new_n4889_; 
wire u2__abc_52138_new_n4890_; 
wire u2__abc_52138_new_n4891_; 
wire u2__abc_52138_new_n4892_; 
wire u2__abc_52138_new_n4893_; 
wire u2__abc_52138_new_n4894_; 
wire u2__abc_52138_new_n4895_; 
wire u2__abc_52138_new_n4896_; 
wire u2__abc_52138_new_n4897_; 
wire u2__abc_52138_new_n4898_; 
wire u2__abc_52138_new_n4899_; 
wire u2__abc_52138_new_n4900_; 
wire u2__abc_52138_new_n4901_; 
wire u2__abc_52138_new_n4902_; 
wire u2__abc_52138_new_n4903_; 
wire u2__abc_52138_new_n4904_; 
wire u2__abc_52138_new_n4905_; 
wire u2__abc_52138_new_n4906_; 
wire u2__abc_52138_new_n4907_; 
wire u2__abc_52138_new_n4908_; 
wire u2__abc_52138_new_n4909_; 
wire u2__abc_52138_new_n4910_; 
wire u2__abc_52138_new_n4911_; 
wire u2__abc_52138_new_n4912_; 
wire u2__abc_52138_new_n4913_; 
wire u2__abc_52138_new_n4914_; 
wire u2__abc_52138_new_n4915_; 
wire u2__abc_52138_new_n4916_; 
wire u2__abc_52138_new_n4917_; 
wire u2__abc_52138_new_n4918_; 
wire u2__abc_52138_new_n4919_; 
wire u2__abc_52138_new_n4920_; 
wire u2__abc_52138_new_n4921_; 
wire u2__abc_52138_new_n4922_; 
wire u2__abc_52138_new_n4923_; 
wire u2__abc_52138_new_n4924_; 
wire u2__abc_52138_new_n4925_; 
wire u2__abc_52138_new_n4926_; 
wire u2__abc_52138_new_n4927_; 
wire u2__abc_52138_new_n4928_; 
wire u2__abc_52138_new_n4929_; 
wire u2__abc_52138_new_n4930_; 
wire u2__abc_52138_new_n4931_; 
wire u2__abc_52138_new_n4932_; 
wire u2__abc_52138_new_n4933_; 
wire u2__abc_52138_new_n4934_; 
wire u2__abc_52138_new_n4935_; 
wire u2__abc_52138_new_n4936_; 
wire u2__abc_52138_new_n4937_; 
wire u2__abc_52138_new_n4938_; 
wire u2__abc_52138_new_n4939_; 
wire u2__abc_52138_new_n4940_; 
wire u2__abc_52138_new_n4941_; 
wire u2__abc_52138_new_n4942_; 
wire u2__abc_52138_new_n4943_; 
wire u2__abc_52138_new_n4944_; 
wire u2__abc_52138_new_n4945_; 
wire u2__abc_52138_new_n4946_; 
wire u2__abc_52138_new_n4947_; 
wire u2__abc_52138_new_n4948_; 
wire u2__abc_52138_new_n4949_; 
wire u2__abc_52138_new_n4950_; 
wire u2__abc_52138_new_n4951_; 
wire u2__abc_52138_new_n4952_; 
wire u2__abc_52138_new_n4953_; 
wire u2__abc_52138_new_n4954_; 
wire u2__abc_52138_new_n4955_; 
wire u2__abc_52138_new_n4956_; 
wire u2__abc_52138_new_n4957_; 
wire u2__abc_52138_new_n4958_; 
wire u2__abc_52138_new_n4959_; 
wire u2__abc_52138_new_n4960_; 
wire u2__abc_52138_new_n4961_; 
wire u2__abc_52138_new_n4962_; 
wire u2__abc_52138_new_n4963_; 
wire u2__abc_52138_new_n4964_; 
wire u2__abc_52138_new_n4965_; 
wire u2__abc_52138_new_n4966_; 
wire u2__abc_52138_new_n4967_; 
wire u2__abc_52138_new_n4968_; 
wire u2__abc_52138_new_n4969_; 
wire u2__abc_52138_new_n4970_; 
wire u2__abc_52138_new_n4971_; 
wire u2__abc_52138_new_n4972_; 
wire u2__abc_52138_new_n4973_; 
wire u2__abc_52138_new_n4974_; 
wire u2__abc_52138_new_n4975_; 
wire u2__abc_52138_new_n4976_; 
wire u2__abc_52138_new_n4977_; 
wire u2__abc_52138_new_n4978_; 
wire u2__abc_52138_new_n4979_; 
wire u2__abc_52138_new_n4980_; 
wire u2__abc_52138_new_n4981_; 
wire u2__abc_52138_new_n4982_; 
wire u2__abc_52138_new_n4983_; 
wire u2__abc_52138_new_n4984_; 
wire u2__abc_52138_new_n4985_; 
wire u2__abc_52138_new_n4986_; 
wire u2__abc_52138_new_n4987_; 
wire u2__abc_52138_new_n4988_; 
wire u2__abc_52138_new_n4989_; 
wire u2__abc_52138_new_n4990_; 
wire u2__abc_52138_new_n4991_; 
wire u2__abc_52138_new_n4992_; 
wire u2__abc_52138_new_n4993_; 
wire u2__abc_52138_new_n4994_; 
wire u2__abc_52138_new_n4995_; 
wire u2__abc_52138_new_n4996_; 
wire u2__abc_52138_new_n4997_; 
wire u2__abc_52138_new_n4998_; 
wire u2__abc_52138_new_n4999_; 
wire u2__abc_52138_new_n5000_; 
wire u2__abc_52138_new_n5001_; 
wire u2__abc_52138_new_n5002_; 
wire u2__abc_52138_new_n5003_; 
wire u2__abc_52138_new_n5004_; 
wire u2__abc_52138_new_n5005_; 
wire u2__abc_52138_new_n5006_; 
wire u2__abc_52138_new_n5007_; 
wire u2__abc_52138_new_n5008_; 
wire u2__abc_52138_new_n5009_; 
wire u2__abc_52138_new_n5010_; 
wire u2__abc_52138_new_n5011_; 
wire u2__abc_52138_new_n5012_; 
wire u2__abc_52138_new_n5013_; 
wire u2__abc_52138_new_n5014_; 
wire u2__abc_52138_new_n5015_; 
wire u2__abc_52138_new_n5016_; 
wire u2__abc_52138_new_n5017_; 
wire u2__abc_52138_new_n5018_; 
wire u2__abc_52138_new_n5019_; 
wire u2__abc_52138_new_n5020_; 
wire u2__abc_52138_new_n5021_; 
wire u2__abc_52138_new_n5022_; 
wire u2__abc_52138_new_n5023_; 
wire u2__abc_52138_new_n5024_; 
wire u2__abc_52138_new_n5025_; 
wire u2__abc_52138_new_n5026_; 
wire u2__abc_52138_new_n5027_; 
wire u2__abc_52138_new_n5028_; 
wire u2__abc_52138_new_n5029_; 
wire u2__abc_52138_new_n5030_; 
wire u2__abc_52138_new_n5031_; 
wire u2__abc_52138_new_n5032_; 
wire u2__abc_52138_new_n5033_; 
wire u2__abc_52138_new_n5034_; 
wire u2__abc_52138_new_n5035_; 
wire u2__abc_52138_new_n5036_; 
wire u2__abc_52138_new_n5037_; 
wire u2__abc_52138_new_n5038_; 
wire u2__abc_52138_new_n5039_; 
wire u2__abc_52138_new_n5040_; 
wire u2__abc_52138_new_n5041_; 
wire u2__abc_52138_new_n5042_; 
wire u2__abc_52138_new_n5043_; 
wire u2__abc_52138_new_n5044_; 
wire u2__abc_52138_new_n5045_; 
wire u2__abc_52138_new_n5046_; 
wire u2__abc_52138_new_n5047_; 
wire u2__abc_52138_new_n5048_; 
wire u2__abc_52138_new_n5049_; 
wire u2__abc_52138_new_n5050_; 
wire u2__abc_52138_new_n5051_; 
wire u2__abc_52138_new_n5052_; 
wire u2__abc_52138_new_n5053_; 
wire u2__abc_52138_new_n5054_; 
wire u2__abc_52138_new_n5055_; 
wire u2__abc_52138_new_n5056_; 
wire u2__abc_52138_new_n5057_; 
wire u2__abc_52138_new_n5058_; 
wire u2__abc_52138_new_n5059_; 
wire u2__abc_52138_new_n5060_; 
wire u2__abc_52138_new_n5061_; 
wire u2__abc_52138_new_n5062_; 
wire u2__abc_52138_new_n5063_; 
wire u2__abc_52138_new_n5064_; 
wire u2__abc_52138_new_n5065_; 
wire u2__abc_52138_new_n5066_; 
wire u2__abc_52138_new_n5067_; 
wire u2__abc_52138_new_n5068_; 
wire u2__abc_52138_new_n5069_; 
wire u2__abc_52138_new_n5070_; 
wire u2__abc_52138_new_n5071_; 
wire u2__abc_52138_new_n5072_; 
wire u2__abc_52138_new_n5073_; 
wire u2__abc_52138_new_n5074_; 
wire u2__abc_52138_new_n5075_; 
wire u2__abc_52138_new_n5076_; 
wire u2__abc_52138_new_n5077_; 
wire u2__abc_52138_new_n5078_; 
wire u2__abc_52138_new_n5079_; 
wire u2__abc_52138_new_n5080_; 
wire u2__abc_52138_new_n5081_; 
wire u2__abc_52138_new_n5082_; 
wire u2__abc_52138_new_n5083_; 
wire u2__abc_52138_new_n5084_; 
wire u2__abc_52138_new_n5085_; 
wire u2__abc_52138_new_n5086_; 
wire u2__abc_52138_new_n5087_; 
wire u2__abc_52138_new_n5088_; 
wire u2__abc_52138_new_n5089_; 
wire u2__abc_52138_new_n5090_; 
wire u2__abc_52138_new_n5091_; 
wire u2__abc_52138_new_n5092_; 
wire u2__abc_52138_new_n5093_; 
wire u2__abc_52138_new_n5094_; 
wire u2__abc_52138_new_n5095_; 
wire u2__abc_52138_new_n5096_; 
wire u2__abc_52138_new_n5097_; 
wire u2__abc_52138_new_n5098_; 
wire u2__abc_52138_new_n5099_; 
wire u2__abc_52138_new_n5100_; 
wire u2__abc_52138_new_n5101_; 
wire u2__abc_52138_new_n5102_; 
wire u2__abc_52138_new_n5103_; 
wire u2__abc_52138_new_n5104_; 
wire u2__abc_52138_new_n5105_; 
wire u2__abc_52138_new_n5106_; 
wire u2__abc_52138_new_n5107_; 
wire u2__abc_52138_new_n5108_; 
wire u2__abc_52138_new_n5109_; 
wire u2__abc_52138_new_n5110_; 
wire u2__abc_52138_new_n5111_; 
wire u2__abc_52138_new_n5112_; 
wire u2__abc_52138_new_n5113_; 
wire u2__abc_52138_new_n5114_; 
wire u2__abc_52138_new_n5115_; 
wire u2__abc_52138_new_n5116_; 
wire u2__abc_52138_new_n5117_; 
wire u2__abc_52138_new_n5118_; 
wire u2__abc_52138_new_n5119_; 
wire u2__abc_52138_new_n5120_; 
wire u2__abc_52138_new_n5121_; 
wire u2__abc_52138_new_n5122_; 
wire u2__abc_52138_new_n5123_; 
wire u2__abc_52138_new_n5124_; 
wire u2__abc_52138_new_n5125_; 
wire u2__abc_52138_new_n5126_; 
wire u2__abc_52138_new_n5127_; 
wire u2__abc_52138_new_n5128_; 
wire u2__abc_52138_new_n5129_; 
wire u2__abc_52138_new_n5130_; 
wire u2__abc_52138_new_n5131_; 
wire u2__abc_52138_new_n5132_; 
wire u2__abc_52138_new_n5133_; 
wire u2__abc_52138_new_n5134_; 
wire u2__abc_52138_new_n5135_; 
wire u2__abc_52138_new_n5136_; 
wire u2__abc_52138_new_n5137_; 
wire u2__abc_52138_new_n5138_; 
wire u2__abc_52138_new_n5139_; 
wire u2__abc_52138_new_n5140_; 
wire u2__abc_52138_new_n5141_; 
wire u2__abc_52138_new_n5142_; 
wire u2__abc_52138_new_n5143_; 
wire u2__abc_52138_new_n5144_; 
wire u2__abc_52138_new_n5145_; 
wire u2__abc_52138_new_n5146_; 
wire u2__abc_52138_new_n5147_; 
wire u2__abc_52138_new_n5148_; 
wire u2__abc_52138_new_n5149_; 
wire u2__abc_52138_new_n5150_; 
wire u2__abc_52138_new_n5151_; 
wire u2__abc_52138_new_n5152_; 
wire u2__abc_52138_new_n5153_; 
wire u2__abc_52138_new_n5154_; 
wire u2__abc_52138_new_n5155_; 
wire u2__abc_52138_new_n5156_; 
wire u2__abc_52138_new_n5157_; 
wire u2__abc_52138_new_n5158_; 
wire u2__abc_52138_new_n5159_; 
wire u2__abc_52138_new_n5160_; 
wire u2__abc_52138_new_n5161_; 
wire u2__abc_52138_new_n5162_; 
wire u2__abc_52138_new_n5163_; 
wire u2__abc_52138_new_n5164_; 
wire u2__abc_52138_new_n5165_; 
wire u2__abc_52138_new_n5166_; 
wire u2__abc_52138_new_n5167_; 
wire u2__abc_52138_new_n5168_; 
wire u2__abc_52138_new_n5169_; 
wire u2__abc_52138_new_n5170_; 
wire u2__abc_52138_new_n5171_; 
wire u2__abc_52138_new_n5172_; 
wire u2__abc_52138_new_n5173_; 
wire u2__abc_52138_new_n5174_; 
wire u2__abc_52138_new_n5175_; 
wire u2__abc_52138_new_n5176_; 
wire u2__abc_52138_new_n5177_; 
wire u2__abc_52138_new_n5178_; 
wire u2__abc_52138_new_n5179_; 
wire u2__abc_52138_new_n5180_; 
wire u2__abc_52138_new_n5181_; 
wire u2__abc_52138_new_n5182_; 
wire u2__abc_52138_new_n5183_; 
wire u2__abc_52138_new_n5184_; 
wire u2__abc_52138_new_n5185_; 
wire u2__abc_52138_new_n5186_; 
wire u2__abc_52138_new_n5187_; 
wire u2__abc_52138_new_n5188_; 
wire u2__abc_52138_new_n5189_; 
wire u2__abc_52138_new_n5190_; 
wire u2__abc_52138_new_n5191_; 
wire u2__abc_52138_new_n5192_; 
wire u2__abc_52138_new_n5193_; 
wire u2__abc_52138_new_n5194_; 
wire u2__abc_52138_new_n5195_; 
wire u2__abc_52138_new_n5196_; 
wire u2__abc_52138_new_n5197_; 
wire u2__abc_52138_new_n5198_; 
wire u2__abc_52138_new_n5199_; 
wire u2__abc_52138_new_n5200_; 
wire u2__abc_52138_new_n5201_; 
wire u2__abc_52138_new_n5202_; 
wire u2__abc_52138_new_n5203_; 
wire u2__abc_52138_new_n5204_; 
wire u2__abc_52138_new_n5205_; 
wire u2__abc_52138_new_n5206_; 
wire u2__abc_52138_new_n5207_; 
wire u2__abc_52138_new_n5208_; 
wire u2__abc_52138_new_n5209_; 
wire u2__abc_52138_new_n5210_; 
wire u2__abc_52138_new_n5211_; 
wire u2__abc_52138_new_n5212_; 
wire u2__abc_52138_new_n5213_; 
wire u2__abc_52138_new_n5214_; 
wire u2__abc_52138_new_n5215_; 
wire u2__abc_52138_new_n5216_; 
wire u2__abc_52138_new_n5217_; 
wire u2__abc_52138_new_n5218_; 
wire u2__abc_52138_new_n5219_; 
wire u2__abc_52138_new_n5220_; 
wire u2__abc_52138_new_n5221_; 
wire u2__abc_52138_new_n5222_; 
wire u2__abc_52138_new_n5223_; 
wire u2__abc_52138_new_n5224_; 
wire u2__abc_52138_new_n5225_; 
wire u2__abc_52138_new_n5226_; 
wire u2__abc_52138_new_n5227_; 
wire u2__abc_52138_new_n5228_; 
wire u2__abc_52138_new_n5229_; 
wire u2__abc_52138_new_n5230_; 
wire u2__abc_52138_new_n5231_; 
wire u2__abc_52138_new_n5232_; 
wire u2__abc_52138_new_n5233_; 
wire u2__abc_52138_new_n5234_; 
wire u2__abc_52138_new_n5235_; 
wire u2__abc_52138_new_n5236_; 
wire u2__abc_52138_new_n5237_; 
wire u2__abc_52138_new_n5238_; 
wire u2__abc_52138_new_n5239_; 
wire u2__abc_52138_new_n5240_; 
wire u2__abc_52138_new_n5241_; 
wire u2__abc_52138_new_n5242_; 
wire u2__abc_52138_new_n5243_; 
wire u2__abc_52138_new_n5244_; 
wire u2__abc_52138_new_n5245_; 
wire u2__abc_52138_new_n5246_; 
wire u2__abc_52138_new_n5247_; 
wire u2__abc_52138_new_n5248_; 
wire u2__abc_52138_new_n5249_; 
wire u2__abc_52138_new_n5250_; 
wire u2__abc_52138_new_n5251_; 
wire u2__abc_52138_new_n5252_; 
wire u2__abc_52138_new_n5253_; 
wire u2__abc_52138_new_n5254_; 
wire u2__abc_52138_new_n5255_; 
wire u2__abc_52138_new_n5256_; 
wire u2__abc_52138_new_n5257_; 
wire u2__abc_52138_new_n5258_; 
wire u2__abc_52138_new_n5259_; 
wire u2__abc_52138_new_n5260_; 
wire u2__abc_52138_new_n5261_; 
wire u2__abc_52138_new_n5262_; 
wire u2__abc_52138_new_n5263_; 
wire u2__abc_52138_new_n5264_; 
wire u2__abc_52138_new_n5265_; 
wire u2__abc_52138_new_n5266_; 
wire u2__abc_52138_new_n5267_; 
wire u2__abc_52138_new_n5268_; 
wire u2__abc_52138_new_n5269_; 
wire u2__abc_52138_new_n5270_; 
wire u2__abc_52138_new_n5271_; 
wire u2__abc_52138_new_n5272_; 
wire u2__abc_52138_new_n5273_; 
wire u2__abc_52138_new_n5274_; 
wire u2__abc_52138_new_n5275_; 
wire u2__abc_52138_new_n5276_; 
wire u2__abc_52138_new_n5277_; 
wire u2__abc_52138_new_n5278_; 
wire u2__abc_52138_new_n5279_; 
wire u2__abc_52138_new_n5280_; 
wire u2__abc_52138_new_n5281_; 
wire u2__abc_52138_new_n5282_; 
wire u2__abc_52138_new_n5283_; 
wire u2__abc_52138_new_n5284_; 
wire u2__abc_52138_new_n5285_; 
wire u2__abc_52138_new_n5286_; 
wire u2__abc_52138_new_n5287_; 
wire u2__abc_52138_new_n5288_; 
wire u2__abc_52138_new_n5289_; 
wire u2__abc_52138_new_n5290_; 
wire u2__abc_52138_new_n5291_; 
wire u2__abc_52138_new_n5292_; 
wire u2__abc_52138_new_n5293_; 
wire u2__abc_52138_new_n5294_; 
wire u2__abc_52138_new_n5295_; 
wire u2__abc_52138_new_n5296_; 
wire u2__abc_52138_new_n5297_; 
wire u2__abc_52138_new_n5298_; 
wire u2__abc_52138_new_n5299_; 
wire u2__abc_52138_new_n5300_; 
wire u2__abc_52138_new_n5301_; 
wire u2__abc_52138_new_n5302_; 
wire u2__abc_52138_new_n5303_; 
wire u2__abc_52138_new_n5304_; 
wire u2__abc_52138_new_n5305_; 
wire u2__abc_52138_new_n5306_; 
wire u2__abc_52138_new_n5307_; 
wire u2__abc_52138_new_n5308_; 
wire u2__abc_52138_new_n5309_; 
wire u2__abc_52138_new_n5310_; 
wire u2__abc_52138_new_n5311_; 
wire u2__abc_52138_new_n5312_; 
wire u2__abc_52138_new_n5313_; 
wire u2__abc_52138_new_n5314_; 
wire u2__abc_52138_new_n5315_; 
wire u2__abc_52138_new_n5316_; 
wire u2__abc_52138_new_n5317_; 
wire u2__abc_52138_new_n5318_; 
wire u2__abc_52138_new_n5319_; 
wire u2__abc_52138_new_n5320_; 
wire u2__abc_52138_new_n5321_; 
wire u2__abc_52138_new_n5322_; 
wire u2__abc_52138_new_n5323_; 
wire u2__abc_52138_new_n5324_; 
wire u2__abc_52138_new_n5325_; 
wire u2__abc_52138_new_n5326_; 
wire u2__abc_52138_new_n5327_; 
wire u2__abc_52138_new_n5328_; 
wire u2__abc_52138_new_n5329_; 
wire u2__abc_52138_new_n5330_; 
wire u2__abc_52138_new_n5331_; 
wire u2__abc_52138_new_n5332_; 
wire u2__abc_52138_new_n5333_; 
wire u2__abc_52138_new_n5334_; 
wire u2__abc_52138_new_n5335_; 
wire u2__abc_52138_new_n5336_; 
wire u2__abc_52138_new_n5337_; 
wire u2__abc_52138_new_n5338_; 
wire u2__abc_52138_new_n5339_; 
wire u2__abc_52138_new_n5340_; 
wire u2__abc_52138_new_n5341_; 
wire u2__abc_52138_new_n5342_; 
wire u2__abc_52138_new_n5343_; 
wire u2__abc_52138_new_n5344_; 
wire u2__abc_52138_new_n5345_; 
wire u2__abc_52138_new_n5346_; 
wire u2__abc_52138_new_n5347_; 
wire u2__abc_52138_new_n5348_; 
wire u2__abc_52138_new_n5349_; 
wire u2__abc_52138_new_n5350_; 
wire u2__abc_52138_new_n5351_; 
wire u2__abc_52138_new_n5352_; 
wire u2__abc_52138_new_n5353_; 
wire u2__abc_52138_new_n5354_; 
wire u2__abc_52138_new_n5355_; 
wire u2__abc_52138_new_n5356_; 
wire u2__abc_52138_new_n5357_; 
wire u2__abc_52138_new_n5358_; 
wire u2__abc_52138_new_n5359_; 
wire u2__abc_52138_new_n5360_; 
wire u2__abc_52138_new_n5361_; 
wire u2__abc_52138_new_n5362_; 
wire u2__abc_52138_new_n5363_; 
wire u2__abc_52138_new_n5364_; 
wire u2__abc_52138_new_n5365_; 
wire u2__abc_52138_new_n5366_; 
wire u2__abc_52138_new_n5367_; 
wire u2__abc_52138_new_n5368_; 
wire u2__abc_52138_new_n5369_; 
wire u2__abc_52138_new_n5370_; 
wire u2__abc_52138_new_n5371_; 
wire u2__abc_52138_new_n5372_; 
wire u2__abc_52138_new_n5373_; 
wire u2__abc_52138_new_n5374_; 
wire u2__abc_52138_new_n5375_; 
wire u2__abc_52138_new_n5376_; 
wire u2__abc_52138_new_n5377_; 
wire u2__abc_52138_new_n5378_; 
wire u2__abc_52138_new_n5379_; 
wire u2__abc_52138_new_n5380_; 
wire u2__abc_52138_new_n5381_; 
wire u2__abc_52138_new_n5382_; 
wire u2__abc_52138_new_n5383_; 
wire u2__abc_52138_new_n5384_; 
wire u2__abc_52138_new_n5385_; 
wire u2__abc_52138_new_n5386_; 
wire u2__abc_52138_new_n5387_; 
wire u2__abc_52138_new_n5388_; 
wire u2__abc_52138_new_n5389_; 
wire u2__abc_52138_new_n5390_; 
wire u2__abc_52138_new_n5391_; 
wire u2__abc_52138_new_n5392_; 
wire u2__abc_52138_new_n5393_; 
wire u2__abc_52138_new_n5394_; 
wire u2__abc_52138_new_n5395_; 
wire u2__abc_52138_new_n5396_; 
wire u2__abc_52138_new_n5397_; 
wire u2__abc_52138_new_n5398_; 
wire u2__abc_52138_new_n5399_; 
wire u2__abc_52138_new_n5400_; 
wire u2__abc_52138_new_n5401_; 
wire u2__abc_52138_new_n5402_; 
wire u2__abc_52138_new_n5403_; 
wire u2__abc_52138_new_n5404_; 
wire u2__abc_52138_new_n5405_; 
wire u2__abc_52138_new_n5406_; 
wire u2__abc_52138_new_n5407_; 
wire u2__abc_52138_new_n5408_; 
wire u2__abc_52138_new_n5409_; 
wire u2__abc_52138_new_n5410_; 
wire u2__abc_52138_new_n5411_; 
wire u2__abc_52138_new_n5412_; 
wire u2__abc_52138_new_n5413_; 
wire u2__abc_52138_new_n5414_; 
wire u2__abc_52138_new_n5415_; 
wire u2__abc_52138_new_n5416_; 
wire u2__abc_52138_new_n5417_; 
wire u2__abc_52138_new_n5418_; 
wire u2__abc_52138_new_n5419_; 
wire u2__abc_52138_new_n5420_; 
wire u2__abc_52138_new_n5421_; 
wire u2__abc_52138_new_n5422_; 
wire u2__abc_52138_new_n5423_; 
wire u2__abc_52138_new_n5424_; 
wire u2__abc_52138_new_n5425_; 
wire u2__abc_52138_new_n5426_; 
wire u2__abc_52138_new_n5427_; 
wire u2__abc_52138_new_n5428_; 
wire u2__abc_52138_new_n5429_; 
wire u2__abc_52138_new_n5430_; 
wire u2__abc_52138_new_n5431_; 
wire u2__abc_52138_new_n5432_; 
wire u2__abc_52138_new_n5433_; 
wire u2__abc_52138_new_n5434_; 
wire u2__abc_52138_new_n5435_; 
wire u2__abc_52138_new_n5436_; 
wire u2__abc_52138_new_n5437_; 
wire u2__abc_52138_new_n5438_; 
wire u2__abc_52138_new_n5439_; 
wire u2__abc_52138_new_n5440_; 
wire u2__abc_52138_new_n5441_; 
wire u2__abc_52138_new_n5442_; 
wire u2__abc_52138_new_n5443_; 
wire u2__abc_52138_new_n5444_; 
wire u2__abc_52138_new_n5445_; 
wire u2__abc_52138_new_n5446_; 
wire u2__abc_52138_new_n5447_; 
wire u2__abc_52138_new_n5448_; 
wire u2__abc_52138_new_n5449_; 
wire u2__abc_52138_new_n5450_; 
wire u2__abc_52138_new_n5451_; 
wire u2__abc_52138_new_n5452_; 
wire u2__abc_52138_new_n5453_; 
wire u2__abc_52138_new_n5454_; 
wire u2__abc_52138_new_n5455_; 
wire u2__abc_52138_new_n5456_; 
wire u2__abc_52138_new_n5457_; 
wire u2__abc_52138_new_n5458_; 
wire u2__abc_52138_new_n5459_; 
wire u2__abc_52138_new_n5460_; 
wire u2__abc_52138_new_n5461_; 
wire u2__abc_52138_new_n5462_; 
wire u2__abc_52138_new_n5463_; 
wire u2__abc_52138_new_n5464_; 
wire u2__abc_52138_new_n5465_; 
wire u2__abc_52138_new_n5466_; 
wire u2__abc_52138_new_n5467_; 
wire u2__abc_52138_new_n5468_; 
wire u2__abc_52138_new_n5469_; 
wire u2__abc_52138_new_n5470_; 
wire u2__abc_52138_new_n5471_; 
wire u2__abc_52138_new_n5472_; 
wire u2__abc_52138_new_n5473_; 
wire u2__abc_52138_new_n5474_; 
wire u2__abc_52138_new_n5475_; 
wire u2__abc_52138_new_n5476_; 
wire u2__abc_52138_new_n5477_; 
wire u2__abc_52138_new_n5478_; 
wire u2__abc_52138_new_n5479_; 
wire u2__abc_52138_new_n5480_; 
wire u2__abc_52138_new_n5481_; 
wire u2__abc_52138_new_n5482_; 
wire u2__abc_52138_new_n5483_; 
wire u2__abc_52138_new_n5484_; 
wire u2__abc_52138_new_n5485_; 
wire u2__abc_52138_new_n5486_; 
wire u2__abc_52138_new_n5487_; 
wire u2__abc_52138_new_n5488_; 
wire u2__abc_52138_new_n5489_; 
wire u2__abc_52138_new_n5490_; 
wire u2__abc_52138_new_n5491_; 
wire u2__abc_52138_new_n5492_; 
wire u2__abc_52138_new_n5493_; 
wire u2__abc_52138_new_n5494_; 
wire u2__abc_52138_new_n5495_; 
wire u2__abc_52138_new_n5496_; 
wire u2__abc_52138_new_n5497_; 
wire u2__abc_52138_new_n5498_; 
wire u2__abc_52138_new_n5499_; 
wire u2__abc_52138_new_n5500_; 
wire u2__abc_52138_new_n5501_; 
wire u2__abc_52138_new_n5502_; 
wire u2__abc_52138_new_n5503_; 
wire u2__abc_52138_new_n5504_; 
wire u2__abc_52138_new_n5505_; 
wire u2__abc_52138_new_n5506_; 
wire u2__abc_52138_new_n5507_; 
wire u2__abc_52138_new_n5508_; 
wire u2__abc_52138_new_n5509_; 
wire u2__abc_52138_new_n5510_; 
wire u2__abc_52138_new_n5511_; 
wire u2__abc_52138_new_n5512_; 
wire u2__abc_52138_new_n5513_; 
wire u2__abc_52138_new_n5514_; 
wire u2__abc_52138_new_n5515_; 
wire u2__abc_52138_new_n5516_; 
wire u2__abc_52138_new_n5517_; 
wire u2__abc_52138_new_n5518_; 
wire u2__abc_52138_new_n5519_; 
wire u2__abc_52138_new_n5520_; 
wire u2__abc_52138_new_n5521_; 
wire u2__abc_52138_new_n5522_; 
wire u2__abc_52138_new_n5523_; 
wire u2__abc_52138_new_n5524_; 
wire u2__abc_52138_new_n5525_; 
wire u2__abc_52138_new_n5526_; 
wire u2__abc_52138_new_n5527_; 
wire u2__abc_52138_new_n5528_; 
wire u2__abc_52138_new_n5529_; 
wire u2__abc_52138_new_n5530_; 
wire u2__abc_52138_new_n5531_; 
wire u2__abc_52138_new_n5532_; 
wire u2__abc_52138_new_n5533_; 
wire u2__abc_52138_new_n5534_; 
wire u2__abc_52138_new_n5535_; 
wire u2__abc_52138_new_n5536_; 
wire u2__abc_52138_new_n5537_; 
wire u2__abc_52138_new_n5538_; 
wire u2__abc_52138_new_n5539_; 
wire u2__abc_52138_new_n5540_; 
wire u2__abc_52138_new_n5541_; 
wire u2__abc_52138_new_n5542_; 
wire u2__abc_52138_new_n5543_; 
wire u2__abc_52138_new_n5544_; 
wire u2__abc_52138_new_n5545_; 
wire u2__abc_52138_new_n5546_; 
wire u2__abc_52138_new_n5547_; 
wire u2__abc_52138_new_n5548_; 
wire u2__abc_52138_new_n5549_; 
wire u2__abc_52138_new_n5550_; 
wire u2__abc_52138_new_n5551_; 
wire u2__abc_52138_new_n5552_; 
wire u2__abc_52138_new_n5553_; 
wire u2__abc_52138_new_n5554_; 
wire u2__abc_52138_new_n5555_; 
wire u2__abc_52138_new_n5556_; 
wire u2__abc_52138_new_n5557_; 
wire u2__abc_52138_new_n5558_; 
wire u2__abc_52138_new_n5559_; 
wire u2__abc_52138_new_n5560_; 
wire u2__abc_52138_new_n5561_; 
wire u2__abc_52138_new_n5562_; 
wire u2__abc_52138_new_n5563_; 
wire u2__abc_52138_new_n5564_; 
wire u2__abc_52138_new_n5565_; 
wire u2__abc_52138_new_n5566_; 
wire u2__abc_52138_new_n5567_; 
wire u2__abc_52138_new_n5568_; 
wire u2__abc_52138_new_n5569_; 
wire u2__abc_52138_new_n5570_; 
wire u2__abc_52138_new_n5571_; 
wire u2__abc_52138_new_n5572_; 
wire u2__abc_52138_new_n5573_; 
wire u2__abc_52138_new_n5574_; 
wire u2__abc_52138_new_n5575_; 
wire u2__abc_52138_new_n5576_; 
wire u2__abc_52138_new_n5577_; 
wire u2__abc_52138_new_n5578_; 
wire u2__abc_52138_new_n5579_; 
wire u2__abc_52138_new_n5580_; 
wire u2__abc_52138_new_n5581_; 
wire u2__abc_52138_new_n5582_; 
wire u2__abc_52138_new_n5583_; 
wire u2__abc_52138_new_n5584_; 
wire u2__abc_52138_new_n5585_; 
wire u2__abc_52138_new_n5586_; 
wire u2__abc_52138_new_n5587_; 
wire u2__abc_52138_new_n5588_; 
wire u2__abc_52138_new_n5589_; 
wire u2__abc_52138_new_n5590_; 
wire u2__abc_52138_new_n5591_; 
wire u2__abc_52138_new_n5592_; 
wire u2__abc_52138_new_n5593_; 
wire u2__abc_52138_new_n5594_; 
wire u2__abc_52138_new_n5595_; 
wire u2__abc_52138_new_n5596_; 
wire u2__abc_52138_new_n5597_; 
wire u2__abc_52138_new_n5598_; 
wire u2__abc_52138_new_n5599_; 
wire u2__abc_52138_new_n5600_; 
wire u2__abc_52138_new_n5601_; 
wire u2__abc_52138_new_n5602_; 
wire u2__abc_52138_new_n5603_; 
wire u2__abc_52138_new_n5604_; 
wire u2__abc_52138_new_n5605_; 
wire u2__abc_52138_new_n5606_; 
wire u2__abc_52138_new_n5607_; 
wire u2__abc_52138_new_n5608_; 
wire u2__abc_52138_new_n5609_; 
wire u2__abc_52138_new_n5610_; 
wire u2__abc_52138_new_n5611_; 
wire u2__abc_52138_new_n5612_; 
wire u2__abc_52138_new_n5613_; 
wire u2__abc_52138_new_n5614_; 
wire u2__abc_52138_new_n5615_; 
wire u2__abc_52138_new_n5616_; 
wire u2__abc_52138_new_n5617_; 
wire u2__abc_52138_new_n5618_; 
wire u2__abc_52138_new_n5619_; 
wire u2__abc_52138_new_n5620_; 
wire u2__abc_52138_new_n5621_; 
wire u2__abc_52138_new_n5622_; 
wire u2__abc_52138_new_n5623_; 
wire u2__abc_52138_new_n5624_; 
wire u2__abc_52138_new_n5625_; 
wire u2__abc_52138_new_n5626_; 
wire u2__abc_52138_new_n5627_; 
wire u2__abc_52138_new_n5628_; 
wire u2__abc_52138_new_n5629_; 
wire u2__abc_52138_new_n5630_; 
wire u2__abc_52138_new_n5631_; 
wire u2__abc_52138_new_n5632_; 
wire u2__abc_52138_new_n5633_; 
wire u2__abc_52138_new_n5634_; 
wire u2__abc_52138_new_n5635_; 
wire u2__abc_52138_new_n5636_; 
wire u2__abc_52138_new_n5637_; 
wire u2__abc_52138_new_n5638_; 
wire u2__abc_52138_new_n5639_; 
wire u2__abc_52138_new_n5640_; 
wire u2__abc_52138_new_n5641_; 
wire u2__abc_52138_new_n5642_; 
wire u2__abc_52138_new_n5643_; 
wire u2__abc_52138_new_n5644_; 
wire u2__abc_52138_new_n5645_; 
wire u2__abc_52138_new_n5646_; 
wire u2__abc_52138_new_n5647_; 
wire u2__abc_52138_new_n5648_; 
wire u2__abc_52138_new_n5649_; 
wire u2__abc_52138_new_n5650_; 
wire u2__abc_52138_new_n5651_; 
wire u2__abc_52138_new_n5652_; 
wire u2__abc_52138_new_n5653_; 
wire u2__abc_52138_new_n5654_; 
wire u2__abc_52138_new_n5655_; 
wire u2__abc_52138_new_n5656_; 
wire u2__abc_52138_new_n5657_; 
wire u2__abc_52138_new_n5658_; 
wire u2__abc_52138_new_n5659_; 
wire u2__abc_52138_new_n5660_; 
wire u2__abc_52138_new_n5661_; 
wire u2__abc_52138_new_n5662_; 
wire u2__abc_52138_new_n5663_; 
wire u2__abc_52138_new_n5664_; 
wire u2__abc_52138_new_n5665_; 
wire u2__abc_52138_new_n5666_; 
wire u2__abc_52138_new_n5667_; 
wire u2__abc_52138_new_n5668_; 
wire u2__abc_52138_new_n5669_; 
wire u2__abc_52138_new_n5670_; 
wire u2__abc_52138_new_n5671_; 
wire u2__abc_52138_new_n5672_; 
wire u2__abc_52138_new_n5673_; 
wire u2__abc_52138_new_n5674_; 
wire u2__abc_52138_new_n5675_; 
wire u2__abc_52138_new_n5676_; 
wire u2__abc_52138_new_n5677_; 
wire u2__abc_52138_new_n5678_; 
wire u2__abc_52138_new_n5679_; 
wire u2__abc_52138_new_n5680_; 
wire u2__abc_52138_new_n5681_; 
wire u2__abc_52138_new_n5682_; 
wire u2__abc_52138_new_n5683_; 
wire u2__abc_52138_new_n5684_; 
wire u2__abc_52138_new_n5685_; 
wire u2__abc_52138_new_n5686_; 
wire u2__abc_52138_new_n5687_; 
wire u2__abc_52138_new_n5688_; 
wire u2__abc_52138_new_n5689_; 
wire u2__abc_52138_new_n5690_; 
wire u2__abc_52138_new_n5691_; 
wire u2__abc_52138_new_n5692_; 
wire u2__abc_52138_new_n5693_; 
wire u2__abc_52138_new_n5694_; 
wire u2__abc_52138_new_n5695_; 
wire u2__abc_52138_new_n5696_; 
wire u2__abc_52138_new_n5697_; 
wire u2__abc_52138_new_n5698_; 
wire u2__abc_52138_new_n5699_; 
wire u2__abc_52138_new_n5700_; 
wire u2__abc_52138_new_n5701_; 
wire u2__abc_52138_new_n5702_; 
wire u2__abc_52138_new_n5703_; 
wire u2__abc_52138_new_n5704_; 
wire u2__abc_52138_new_n5705_; 
wire u2__abc_52138_new_n5706_; 
wire u2__abc_52138_new_n5707_; 
wire u2__abc_52138_new_n5708_; 
wire u2__abc_52138_new_n5709_; 
wire u2__abc_52138_new_n5710_; 
wire u2__abc_52138_new_n5711_; 
wire u2__abc_52138_new_n5712_; 
wire u2__abc_52138_new_n5713_; 
wire u2__abc_52138_new_n5714_; 
wire u2__abc_52138_new_n5715_; 
wire u2__abc_52138_new_n5716_; 
wire u2__abc_52138_new_n5717_; 
wire u2__abc_52138_new_n5718_; 
wire u2__abc_52138_new_n5719_; 
wire u2__abc_52138_new_n5720_; 
wire u2__abc_52138_new_n5721_; 
wire u2__abc_52138_new_n5722_; 
wire u2__abc_52138_new_n5723_; 
wire u2__abc_52138_new_n5724_; 
wire u2__abc_52138_new_n5725_; 
wire u2__abc_52138_new_n5726_; 
wire u2__abc_52138_new_n5727_; 
wire u2__abc_52138_new_n5728_; 
wire u2__abc_52138_new_n5729_; 
wire u2__abc_52138_new_n5730_; 
wire u2__abc_52138_new_n5731_; 
wire u2__abc_52138_new_n5732_; 
wire u2__abc_52138_new_n5733_; 
wire u2__abc_52138_new_n5734_; 
wire u2__abc_52138_new_n5735_; 
wire u2__abc_52138_new_n5736_; 
wire u2__abc_52138_new_n5737_; 
wire u2__abc_52138_new_n5738_; 
wire u2__abc_52138_new_n5739_; 
wire u2__abc_52138_new_n5740_; 
wire u2__abc_52138_new_n5741_; 
wire u2__abc_52138_new_n5742_; 
wire u2__abc_52138_new_n5743_; 
wire u2__abc_52138_new_n5744_; 
wire u2__abc_52138_new_n5745_; 
wire u2__abc_52138_new_n5746_; 
wire u2__abc_52138_new_n5747_; 
wire u2__abc_52138_new_n5748_; 
wire u2__abc_52138_new_n5749_; 
wire u2__abc_52138_new_n5750_; 
wire u2__abc_52138_new_n5751_; 
wire u2__abc_52138_new_n5752_; 
wire u2__abc_52138_new_n5753_; 
wire u2__abc_52138_new_n5754_; 
wire u2__abc_52138_new_n5755_; 
wire u2__abc_52138_new_n5756_; 
wire u2__abc_52138_new_n5757_; 
wire u2__abc_52138_new_n5758_; 
wire u2__abc_52138_new_n5759_; 
wire u2__abc_52138_new_n5760_; 
wire u2__abc_52138_new_n5761_; 
wire u2__abc_52138_new_n5762_; 
wire u2__abc_52138_new_n5763_; 
wire u2__abc_52138_new_n5764_; 
wire u2__abc_52138_new_n5765_; 
wire u2__abc_52138_new_n5766_; 
wire u2__abc_52138_new_n5767_; 
wire u2__abc_52138_new_n5768_; 
wire u2__abc_52138_new_n5769_; 
wire u2__abc_52138_new_n5770_; 
wire u2__abc_52138_new_n5771_; 
wire u2__abc_52138_new_n5772_; 
wire u2__abc_52138_new_n5773_; 
wire u2__abc_52138_new_n5774_; 
wire u2__abc_52138_new_n5775_; 
wire u2__abc_52138_new_n5776_; 
wire u2__abc_52138_new_n5777_; 
wire u2__abc_52138_new_n5778_; 
wire u2__abc_52138_new_n5779_; 
wire u2__abc_52138_new_n5780_; 
wire u2__abc_52138_new_n5781_; 
wire u2__abc_52138_new_n5782_; 
wire u2__abc_52138_new_n5783_; 
wire u2__abc_52138_new_n5784_; 
wire u2__abc_52138_new_n5785_; 
wire u2__abc_52138_new_n5786_; 
wire u2__abc_52138_new_n5787_; 
wire u2__abc_52138_new_n5788_; 
wire u2__abc_52138_new_n5789_; 
wire u2__abc_52138_new_n5790_; 
wire u2__abc_52138_new_n5791_; 
wire u2__abc_52138_new_n5792_; 
wire u2__abc_52138_new_n5793_; 
wire u2__abc_52138_new_n5794_; 
wire u2__abc_52138_new_n5795_; 
wire u2__abc_52138_new_n5796_; 
wire u2__abc_52138_new_n5797_; 
wire u2__abc_52138_new_n5798_; 
wire u2__abc_52138_new_n5799_; 
wire u2__abc_52138_new_n5800_; 
wire u2__abc_52138_new_n5801_; 
wire u2__abc_52138_new_n5802_; 
wire u2__abc_52138_new_n5803_; 
wire u2__abc_52138_new_n5804_; 
wire u2__abc_52138_new_n5805_; 
wire u2__abc_52138_new_n5806_; 
wire u2__abc_52138_new_n5807_; 
wire u2__abc_52138_new_n5808_; 
wire u2__abc_52138_new_n5809_; 
wire u2__abc_52138_new_n5810_; 
wire u2__abc_52138_new_n5811_; 
wire u2__abc_52138_new_n5812_; 
wire u2__abc_52138_new_n5813_; 
wire u2__abc_52138_new_n5814_; 
wire u2__abc_52138_new_n5815_; 
wire u2__abc_52138_new_n5816_; 
wire u2__abc_52138_new_n5817_; 
wire u2__abc_52138_new_n5818_; 
wire u2__abc_52138_new_n5819_; 
wire u2__abc_52138_new_n5820_; 
wire u2__abc_52138_new_n5821_; 
wire u2__abc_52138_new_n5822_; 
wire u2__abc_52138_new_n5823_; 
wire u2__abc_52138_new_n5824_; 
wire u2__abc_52138_new_n5825_; 
wire u2__abc_52138_new_n5826_; 
wire u2__abc_52138_new_n5827_; 
wire u2__abc_52138_new_n5828_; 
wire u2__abc_52138_new_n5829_; 
wire u2__abc_52138_new_n5830_; 
wire u2__abc_52138_new_n5831_; 
wire u2__abc_52138_new_n5832_; 
wire u2__abc_52138_new_n5833_; 
wire u2__abc_52138_new_n5834_; 
wire u2__abc_52138_new_n5835_; 
wire u2__abc_52138_new_n5836_; 
wire u2__abc_52138_new_n5837_; 
wire u2__abc_52138_new_n5838_; 
wire u2__abc_52138_new_n5839_; 
wire u2__abc_52138_new_n5840_; 
wire u2__abc_52138_new_n5841_; 
wire u2__abc_52138_new_n5842_; 
wire u2__abc_52138_new_n5843_; 
wire u2__abc_52138_new_n5844_; 
wire u2__abc_52138_new_n5845_; 
wire u2__abc_52138_new_n5846_; 
wire u2__abc_52138_new_n5847_; 
wire u2__abc_52138_new_n5848_; 
wire u2__abc_52138_new_n5849_; 
wire u2__abc_52138_new_n5850_; 
wire u2__abc_52138_new_n5851_; 
wire u2__abc_52138_new_n5852_; 
wire u2__abc_52138_new_n5853_; 
wire u2__abc_52138_new_n5854_; 
wire u2__abc_52138_new_n5855_; 
wire u2__abc_52138_new_n5856_; 
wire u2__abc_52138_new_n5857_; 
wire u2__abc_52138_new_n5858_; 
wire u2__abc_52138_new_n5859_; 
wire u2__abc_52138_new_n5860_; 
wire u2__abc_52138_new_n5861_; 
wire u2__abc_52138_new_n5862_; 
wire u2__abc_52138_new_n5863_; 
wire u2__abc_52138_new_n5864_; 
wire u2__abc_52138_new_n5865_; 
wire u2__abc_52138_new_n5866_; 
wire u2__abc_52138_new_n5867_; 
wire u2__abc_52138_new_n5868_; 
wire u2__abc_52138_new_n5869_; 
wire u2__abc_52138_new_n5870_; 
wire u2__abc_52138_new_n5871_; 
wire u2__abc_52138_new_n5872_; 
wire u2__abc_52138_new_n5873_; 
wire u2__abc_52138_new_n5874_; 
wire u2__abc_52138_new_n5875_; 
wire u2__abc_52138_new_n5876_; 
wire u2__abc_52138_new_n5877_; 
wire u2__abc_52138_new_n5878_; 
wire u2__abc_52138_new_n5879_; 
wire u2__abc_52138_new_n5880_; 
wire u2__abc_52138_new_n5881_; 
wire u2__abc_52138_new_n5882_; 
wire u2__abc_52138_new_n5883_; 
wire u2__abc_52138_new_n5884_; 
wire u2__abc_52138_new_n5885_; 
wire u2__abc_52138_new_n5886_; 
wire u2__abc_52138_new_n5887_; 
wire u2__abc_52138_new_n5888_; 
wire u2__abc_52138_new_n5889_; 
wire u2__abc_52138_new_n5890_; 
wire u2__abc_52138_new_n5891_; 
wire u2__abc_52138_new_n5892_; 
wire u2__abc_52138_new_n5893_; 
wire u2__abc_52138_new_n5894_; 
wire u2__abc_52138_new_n5895_; 
wire u2__abc_52138_new_n5896_; 
wire u2__abc_52138_new_n5897_; 
wire u2__abc_52138_new_n5898_; 
wire u2__abc_52138_new_n5899_; 
wire u2__abc_52138_new_n5900_; 
wire u2__abc_52138_new_n5901_; 
wire u2__abc_52138_new_n5902_; 
wire u2__abc_52138_new_n5903_; 
wire u2__abc_52138_new_n5904_; 
wire u2__abc_52138_new_n5905_; 
wire u2__abc_52138_new_n5906_; 
wire u2__abc_52138_new_n5907_; 
wire u2__abc_52138_new_n5908_; 
wire u2__abc_52138_new_n5909_; 
wire u2__abc_52138_new_n5910_; 
wire u2__abc_52138_new_n5911_; 
wire u2__abc_52138_new_n5912_; 
wire u2__abc_52138_new_n5913_; 
wire u2__abc_52138_new_n5914_; 
wire u2__abc_52138_new_n5915_; 
wire u2__abc_52138_new_n5916_; 
wire u2__abc_52138_new_n5917_; 
wire u2__abc_52138_new_n5918_; 
wire u2__abc_52138_new_n5919_; 
wire u2__abc_52138_new_n5920_; 
wire u2__abc_52138_new_n5921_; 
wire u2__abc_52138_new_n5922_; 
wire u2__abc_52138_new_n5923_; 
wire u2__abc_52138_new_n5924_; 
wire u2__abc_52138_new_n5925_; 
wire u2__abc_52138_new_n5926_; 
wire u2__abc_52138_new_n5927_; 
wire u2__abc_52138_new_n5928_; 
wire u2__abc_52138_new_n5929_; 
wire u2__abc_52138_new_n5930_; 
wire u2__abc_52138_new_n5931_; 
wire u2__abc_52138_new_n5932_; 
wire u2__abc_52138_new_n5933_; 
wire u2__abc_52138_new_n5934_; 
wire u2__abc_52138_new_n5935_; 
wire u2__abc_52138_new_n5936_; 
wire u2__abc_52138_new_n5937_; 
wire u2__abc_52138_new_n5938_; 
wire u2__abc_52138_new_n5939_; 
wire u2__abc_52138_new_n5940_; 
wire u2__abc_52138_new_n5941_; 
wire u2__abc_52138_new_n5942_; 
wire u2__abc_52138_new_n5943_; 
wire u2__abc_52138_new_n5944_; 
wire u2__abc_52138_new_n5945_; 
wire u2__abc_52138_new_n5946_; 
wire u2__abc_52138_new_n5947_; 
wire u2__abc_52138_new_n5948_; 
wire u2__abc_52138_new_n5949_; 
wire u2__abc_52138_new_n5950_; 
wire u2__abc_52138_new_n5951_; 
wire u2__abc_52138_new_n5952_; 
wire u2__abc_52138_new_n5953_; 
wire u2__abc_52138_new_n5954_; 
wire u2__abc_52138_new_n5955_; 
wire u2__abc_52138_new_n5956_; 
wire u2__abc_52138_new_n5957_; 
wire u2__abc_52138_new_n5958_; 
wire u2__abc_52138_new_n5959_; 
wire u2__abc_52138_new_n5960_; 
wire u2__abc_52138_new_n5961_; 
wire u2__abc_52138_new_n5962_; 
wire u2__abc_52138_new_n5963_; 
wire u2__abc_52138_new_n5964_; 
wire u2__abc_52138_new_n5965_; 
wire u2__abc_52138_new_n5966_; 
wire u2__abc_52138_new_n5967_; 
wire u2__abc_52138_new_n5968_; 
wire u2__abc_52138_new_n5969_; 
wire u2__abc_52138_new_n5970_; 
wire u2__abc_52138_new_n5971_; 
wire u2__abc_52138_new_n5972_; 
wire u2__abc_52138_new_n5973_; 
wire u2__abc_52138_new_n5974_; 
wire u2__abc_52138_new_n5975_; 
wire u2__abc_52138_new_n5976_; 
wire u2__abc_52138_new_n5977_; 
wire u2__abc_52138_new_n5978_; 
wire u2__abc_52138_new_n5979_; 
wire u2__abc_52138_new_n5980_; 
wire u2__abc_52138_new_n5981_; 
wire u2__abc_52138_new_n5982_; 
wire u2__abc_52138_new_n5983_; 
wire u2__abc_52138_new_n5984_; 
wire u2__abc_52138_new_n5985_; 
wire u2__abc_52138_new_n5986_; 
wire u2__abc_52138_new_n5987_; 
wire u2__abc_52138_new_n5988_; 
wire u2__abc_52138_new_n5989_; 
wire u2__abc_52138_new_n5990_; 
wire u2__abc_52138_new_n5991_; 
wire u2__abc_52138_new_n5992_; 
wire u2__abc_52138_new_n5993_; 
wire u2__abc_52138_new_n5994_; 
wire u2__abc_52138_new_n5995_; 
wire u2__abc_52138_new_n5996_; 
wire u2__abc_52138_new_n5997_; 
wire u2__abc_52138_new_n5998_; 
wire u2__abc_52138_new_n5999_; 
wire u2__abc_52138_new_n6000_; 
wire u2__abc_52138_new_n6001_; 
wire u2__abc_52138_new_n6002_; 
wire u2__abc_52138_new_n6003_; 
wire u2__abc_52138_new_n6004_; 
wire u2__abc_52138_new_n6005_; 
wire u2__abc_52138_new_n6006_; 
wire u2__abc_52138_new_n6007_; 
wire u2__abc_52138_new_n6008_; 
wire u2__abc_52138_new_n6009_; 
wire u2__abc_52138_new_n6010_; 
wire u2__abc_52138_new_n6011_; 
wire u2__abc_52138_new_n6012_; 
wire u2__abc_52138_new_n6013_; 
wire u2__abc_52138_new_n6014_; 
wire u2__abc_52138_new_n6015_; 
wire u2__abc_52138_new_n6016_; 
wire u2__abc_52138_new_n6017_; 
wire u2__abc_52138_new_n6018_; 
wire u2__abc_52138_new_n6019_; 
wire u2__abc_52138_new_n6020_; 
wire u2__abc_52138_new_n6021_; 
wire u2__abc_52138_new_n6022_; 
wire u2__abc_52138_new_n6023_; 
wire u2__abc_52138_new_n6024_; 
wire u2__abc_52138_new_n6025_; 
wire u2__abc_52138_new_n6026_; 
wire u2__abc_52138_new_n6027_; 
wire u2__abc_52138_new_n6028_; 
wire u2__abc_52138_new_n6029_; 
wire u2__abc_52138_new_n6030_; 
wire u2__abc_52138_new_n6031_; 
wire u2__abc_52138_new_n6032_; 
wire u2__abc_52138_new_n6033_; 
wire u2__abc_52138_new_n6034_; 
wire u2__abc_52138_new_n6035_; 
wire u2__abc_52138_new_n6036_; 
wire u2__abc_52138_new_n6037_; 
wire u2__abc_52138_new_n6038_; 
wire u2__abc_52138_new_n6039_; 
wire u2__abc_52138_new_n6040_; 
wire u2__abc_52138_new_n6041_; 
wire u2__abc_52138_new_n6042_; 
wire u2__abc_52138_new_n6043_; 
wire u2__abc_52138_new_n6044_; 
wire u2__abc_52138_new_n6045_; 
wire u2__abc_52138_new_n6046_; 
wire u2__abc_52138_new_n6047_; 
wire u2__abc_52138_new_n6048_; 
wire u2__abc_52138_new_n6049_; 
wire u2__abc_52138_new_n6050_; 
wire u2__abc_52138_new_n6051_; 
wire u2__abc_52138_new_n6052_; 
wire u2__abc_52138_new_n6053_; 
wire u2__abc_52138_new_n6054_; 
wire u2__abc_52138_new_n6055_; 
wire u2__abc_52138_new_n6056_; 
wire u2__abc_52138_new_n6057_; 
wire u2__abc_52138_new_n6058_; 
wire u2__abc_52138_new_n6059_; 
wire u2__abc_52138_new_n6060_; 
wire u2__abc_52138_new_n6061_; 
wire u2__abc_52138_new_n6062_; 
wire u2__abc_52138_new_n6063_; 
wire u2__abc_52138_new_n6064_; 
wire u2__abc_52138_new_n6065_; 
wire u2__abc_52138_new_n6066_; 
wire u2__abc_52138_new_n6067_; 
wire u2__abc_52138_new_n6068_; 
wire u2__abc_52138_new_n6069_; 
wire u2__abc_52138_new_n6070_; 
wire u2__abc_52138_new_n6071_; 
wire u2__abc_52138_new_n6072_; 
wire u2__abc_52138_new_n6073_; 
wire u2__abc_52138_new_n6074_; 
wire u2__abc_52138_new_n6075_; 
wire u2__abc_52138_new_n6076_; 
wire u2__abc_52138_new_n6077_; 
wire u2__abc_52138_new_n6078_; 
wire u2__abc_52138_new_n6079_; 
wire u2__abc_52138_new_n6080_; 
wire u2__abc_52138_new_n6081_; 
wire u2__abc_52138_new_n6082_; 
wire u2__abc_52138_new_n6083_; 
wire u2__abc_52138_new_n6084_; 
wire u2__abc_52138_new_n6085_; 
wire u2__abc_52138_new_n6086_; 
wire u2__abc_52138_new_n6087_; 
wire u2__abc_52138_new_n6088_; 
wire u2__abc_52138_new_n6089_; 
wire u2__abc_52138_new_n6090_; 
wire u2__abc_52138_new_n6091_; 
wire u2__abc_52138_new_n6092_; 
wire u2__abc_52138_new_n6093_; 
wire u2__abc_52138_new_n6094_; 
wire u2__abc_52138_new_n6095_; 
wire u2__abc_52138_new_n6096_; 
wire u2__abc_52138_new_n6097_; 
wire u2__abc_52138_new_n6098_; 
wire u2__abc_52138_new_n6099_; 
wire u2__abc_52138_new_n6100_; 
wire u2__abc_52138_new_n6101_; 
wire u2__abc_52138_new_n6102_; 
wire u2__abc_52138_new_n6103_; 
wire u2__abc_52138_new_n6104_; 
wire u2__abc_52138_new_n6105_; 
wire u2__abc_52138_new_n6106_; 
wire u2__abc_52138_new_n6107_; 
wire u2__abc_52138_new_n6108_; 
wire u2__abc_52138_new_n6109_; 
wire u2__abc_52138_new_n6110_; 
wire u2__abc_52138_new_n6111_; 
wire u2__abc_52138_new_n6112_; 
wire u2__abc_52138_new_n6113_; 
wire u2__abc_52138_new_n6114_; 
wire u2__abc_52138_new_n6115_; 
wire u2__abc_52138_new_n6116_; 
wire u2__abc_52138_new_n6117_; 
wire u2__abc_52138_new_n6118_; 
wire u2__abc_52138_new_n6119_; 
wire u2__abc_52138_new_n6120_; 
wire u2__abc_52138_new_n6121_; 
wire u2__abc_52138_new_n6122_; 
wire u2__abc_52138_new_n6123_; 
wire u2__abc_52138_new_n6124_; 
wire u2__abc_52138_new_n6125_; 
wire u2__abc_52138_new_n6126_; 
wire u2__abc_52138_new_n6127_; 
wire u2__abc_52138_new_n6128_; 
wire u2__abc_52138_new_n6129_; 
wire u2__abc_52138_new_n6130_; 
wire u2__abc_52138_new_n6131_; 
wire u2__abc_52138_new_n6132_; 
wire u2__abc_52138_new_n6133_; 
wire u2__abc_52138_new_n6134_; 
wire u2__abc_52138_new_n6135_; 
wire u2__abc_52138_new_n6136_; 
wire u2__abc_52138_new_n6137_; 
wire u2__abc_52138_new_n6138_; 
wire u2__abc_52138_new_n6139_; 
wire u2__abc_52138_new_n6140_; 
wire u2__abc_52138_new_n6141_; 
wire u2__abc_52138_new_n6142_; 
wire u2__abc_52138_new_n6143_; 
wire u2__abc_52138_new_n6144_; 
wire u2__abc_52138_new_n6145_; 
wire u2__abc_52138_new_n6146_; 
wire u2__abc_52138_new_n6147_; 
wire u2__abc_52138_new_n6148_; 
wire u2__abc_52138_new_n6149_; 
wire u2__abc_52138_new_n6150_; 
wire u2__abc_52138_new_n6151_; 
wire u2__abc_52138_new_n6152_; 
wire u2__abc_52138_new_n6153_; 
wire u2__abc_52138_new_n6154_; 
wire u2__abc_52138_new_n6155_; 
wire u2__abc_52138_new_n6156_; 
wire u2__abc_52138_new_n6157_; 
wire u2__abc_52138_new_n6158_; 
wire u2__abc_52138_new_n6159_; 
wire u2__abc_52138_new_n6160_; 
wire u2__abc_52138_new_n6161_; 
wire u2__abc_52138_new_n6162_; 
wire u2__abc_52138_new_n6163_; 
wire u2__abc_52138_new_n6164_; 
wire u2__abc_52138_new_n6165_; 
wire u2__abc_52138_new_n6166_; 
wire u2__abc_52138_new_n6167_; 
wire u2__abc_52138_new_n6168_; 
wire u2__abc_52138_new_n6169_; 
wire u2__abc_52138_new_n6170_; 
wire u2__abc_52138_new_n6171_; 
wire u2__abc_52138_new_n6172_; 
wire u2__abc_52138_new_n6173_; 
wire u2__abc_52138_new_n6174_; 
wire u2__abc_52138_new_n6175_; 
wire u2__abc_52138_new_n6176_; 
wire u2__abc_52138_new_n6177_; 
wire u2__abc_52138_new_n6178_; 
wire u2__abc_52138_new_n6179_; 
wire u2__abc_52138_new_n6180_; 
wire u2__abc_52138_new_n6181_; 
wire u2__abc_52138_new_n6182_; 
wire u2__abc_52138_new_n6183_; 
wire u2__abc_52138_new_n6184_; 
wire u2__abc_52138_new_n6185_; 
wire u2__abc_52138_new_n6186_; 
wire u2__abc_52138_new_n6187_; 
wire u2__abc_52138_new_n6188_; 
wire u2__abc_52138_new_n6189_; 
wire u2__abc_52138_new_n6190_; 
wire u2__abc_52138_new_n6191_; 
wire u2__abc_52138_new_n6192_; 
wire u2__abc_52138_new_n6193_; 
wire u2__abc_52138_new_n6194_; 
wire u2__abc_52138_new_n6195_; 
wire u2__abc_52138_new_n6196_; 
wire u2__abc_52138_new_n6197_; 
wire u2__abc_52138_new_n6198_; 
wire u2__abc_52138_new_n6199_; 
wire u2__abc_52138_new_n6200_; 
wire u2__abc_52138_new_n6201_; 
wire u2__abc_52138_new_n6202_; 
wire u2__abc_52138_new_n6203_; 
wire u2__abc_52138_new_n6204_; 
wire u2__abc_52138_new_n6205_; 
wire u2__abc_52138_new_n6206_; 
wire u2__abc_52138_new_n6207_; 
wire u2__abc_52138_new_n6208_; 
wire u2__abc_52138_new_n6209_; 
wire u2__abc_52138_new_n6210_; 
wire u2__abc_52138_new_n6211_; 
wire u2__abc_52138_new_n6212_; 
wire u2__abc_52138_new_n6213_; 
wire u2__abc_52138_new_n6214_; 
wire u2__abc_52138_new_n6215_; 
wire u2__abc_52138_new_n6216_; 
wire u2__abc_52138_new_n6217_; 
wire u2__abc_52138_new_n6218_; 
wire u2__abc_52138_new_n6219_; 
wire u2__abc_52138_new_n6220_; 
wire u2__abc_52138_new_n6221_; 
wire u2__abc_52138_new_n6222_; 
wire u2__abc_52138_new_n6223_; 
wire u2__abc_52138_new_n6224_; 
wire u2__abc_52138_new_n6225_; 
wire u2__abc_52138_new_n6226_; 
wire u2__abc_52138_new_n6227_; 
wire u2__abc_52138_new_n6228_; 
wire u2__abc_52138_new_n6229_; 
wire u2__abc_52138_new_n6230_; 
wire u2__abc_52138_new_n6231_; 
wire u2__abc_52138_new_n6232_; 
wire u2__abc_52138_new_n6233_; 
wire u2__abc_52138_new_n6234_; 
wire u2__abc_52138_new_n6235_; 
wire u2__abc_52138_new_n6236_; 
wire u2__abc_52138_new_n6237_; 
wire u2__abc_52138_new_n6238_; 
wire u2__abc_52138_new_n6239_; 
wire u2__abc_52138_new_n6240_; 
wire u2__abc_52138_new_n6241_; 
wire u2__abc_52138_new_n6242_; 
wire u2__abc_52138_new_n6243_; 
wire u2__abc_52138_new_n6244_; 
wire u2__abc_52138_new_n6245_; 
wire u2__abc_52138_new_n6246_; 
wire u2__abc_52138_new_n6247_; 
wire u2__abc_52138_new_n6248_; 
wire u2__abc_52138_new_n6249_; 
wire u2__abc_52138_new_n6250_; 
wire u2__abc_52138_new_n6251_; 
wire u2__abc_52138_new_n6252_; 
wire u2__abc_52138_new_n6253_; 
wire u2__abc_52138_new_n6254_; 
wire u2__abc_52138_new_n6255_; 
wire u2__abc_52138_new_n6256_; 
wire u2__abc_52138_new_n6257_; 
wire u2__abc_52138_new_n6258_; 
wire u2__abc_52138_new_n6259_; 
wire u2__abc_52138_new_n6260_; 
wire u2__abc_52138_new_n6261_; 
wire u2__abc_52138_new_n6262_; 
wire u2__abc_52138_new_n6263_; 
wire u2__abc_52138_new_n6264_; 
wire u2__abc_52138_new_n6265_; 
wire u2__abc_52138_new_n6266_; 
wire u2__abc_52138_new_n6267_; 
wire u2__abc_52138_new_n6268_; 
wire u2__abc_52138_new_n6269_; 
wire u2__abc_52138_new_n6270_; 
wire u2__abc_52138_new_n6271_; 
wire u2__abc_52138_new_n6272_; 
wire u2__abc_52138_new_n6273_; 
wire u2__abc_52138_new_n6274_; 
wire u2__abc_52138_new_n6275_; 
wire u2__abc_52138_new_n6276_; 
wire u2__abc_52138_new_n6277_; 
wire u2__abc_52138_new_n6278_; 
wire u2__abc_52138_new_n6279_; 
wire u2__abc_52138_new_n6280_; 
wire u2__abc_52138_new_n6281_; 
wire u2__abc_52138_new_n6282_; 
wire u2__abc_52138_new_n6283_; 
wire u2__abc_52138_new_n6284_; 
wire u2__abc_52138_new_n6285_; 
wire u2__abc_52138_new_n6286_; 
wire u2__abc_52138_new_n6287_; 
wire u2__abc_52138_new_n6288_; 
wire u2__abc_52138_new_n6289_; 
wire u2__abc_52138_new_n6290_; 
wire u2__abc_52138_new_n6291_; 
wire u2__abc_52138_new_n6292_; 
wire u2__abc_52138_new_n6293_; 
wire u2__abc_52138_new_n6294_; 
wire u2__abc_52138_new_n6295_; 
wire u2__abc_52138_new_n6296_; 
wire u2__abc_52138_new_n6297_; 
wire u2__abc_52138_new_n6298_; 
wire u2__abc_52138_new_n6299_; 
wire u2__abc_52138_new_n6300_; 
wire u2__abc_52138_new_n6301_; 
wire u2__abc_52138_new_n6302_; 
wire u2__abc_52138_new_n6303_; 
wire u2__abc_52138_new_n6304_; 
wire u2__abc_52138_new_n6305_; 
wire u2__abc_52138_new_n6306_; 
wire u2__abc_52138_new_n6307_; 
wire u2__abc_52138_new_n6308_; 
wire u2__abc_52138_new_n6309_; 
wire u2__abc_52138_new_n6310_; 
wire u2__abc_52138_new_n6311_; 
wire u2__abc_52138_new_n6312_; 
wire u2__abc_52138_new_n6313_; 
wire u2__abc_52138_new_n6314_; 
wire u2__abc_52138_new_n6315_; 
wire u2__abc_52138_new_n6316_; 
wire u2__abc_52138_new_n6317_; 
wire u2__abc_52138_new_n6318_; 
wire u2__abc_52138_new_n6319_; 
wire u2__abc_52138_new_n6320_; 
wire u2__abc_52138_new_n6321_; 
wire u2__abc_52138_new_n6322_; 
wire u2__abc_52138_new_n6323_; 
wire u2__abc_52138_new_n6324_; 
wire u2__abc_52138_new_n6325_; 
wire u2__abc_52138_new_n6326_; 
wire u2__abc_52138_new_n6327_; 
wire u2__abc_52138_new_n6328_; 
wire u2__abc_52138_new_n6329_; 
wire u2__abc_52138_new_n6330_; 
wire u2__abc_52138_new_n6331_; 
wire u2__abc_52138_new_n6332_; 
wire u2__abc_52138_new_n6333_; 
wire u2__abc_52138_new_n6334_; 
wire u2__abc_52138_new_n6335_; 
wire u2__abc_52138_new_n6336_; 
wire u2__abc_52138_new_n6337_; 
wire u2__abc_52138_new_n6338_; 
wire u2__abc_52138_new_n6339_; 
wire u2__abc_52138_new_n6340_; 
wire u2__abc_52138_new_n6341_; 
wire u2__abc_52138_new_n6342_; 
wire u2__abc_52138_new_n6343_; 
wire u2__abc_52138_new_n6344_; 
wire u2__abc_52138_new_n6345_; 
wire u2__abc_52138_new_n6346_; 
wire u2__abc_52138_new_n6347_; 
wire u2__abc_52138_new_n6348_; 
wire u2__abc_52138_new_n6349_; 
wire u2__abc_52138_new_n6350_; 
wire u2__abc_52138_new_n6351_; 
wire u2__abc_52138_new_n6352_; 
wire u2__abc_52138_new_n6353_; 
wire u2__abc_52138_new_n6354_; 
wire u2__abc_52138_new_n6355_; 
wire u2__abc_52138_new_n6356_; 
wire u2__abc_52138_new_n6357_; 
wire u2__abc_52138_new_n6358_; 
wire u2__abc_52138_new_n6359_; 
wire u2__abc_52138_new_n6360_; 
wire u2__abc_52138_new_n6361_; 
wire u2__abc_52138_new_n6362_; 
wire u2__abc_52138_new_n6363_; 
wire u2__abc_52138_new_n6364_; 
wire u2__abc_52138_new_n6365_; 
wire u2__abc_52138_new_n6366_; 
wire u2__abc_52138_new_n6367_; 
wire u2__abc_52138_new_n6368_; 
wire u2__abc_52138_new_n6369_; 
wire u2__abc_52138_new_n6370_; 
wire u2__abc_52138_new_n6371_; 
wire u2__abc_52138_new_n6372_; 
wire u2__abc_52138_new_n6373_; 
wire u2__abc_52138_new_n6374_; 
wire u2__abc_52138_new_n6375_; 
wire u2__abc_52138_new_n6376_; 
wire u2__abc_52138_new_n6377_; 
wire u2__abc_52138_new_n6378_; 
wire u2__abc_52138_new_n6379_; 
wire u2__abc_52138_new_n6380_; 
wire u2__abc_52138_new_n6381_; 
wire u2__abc_52138_new_n6382_; 
wire u2__abc_52138_new_n6383_; 
wire u2__abc_52138_new_n6384_; 
wire u2__abc_52138_new_n6385_; 
wire u2__abc_52138_new_n6386_; 
wire u2__abc_52138_new_n6387_; 
wire u2__abc_52138_new_n6388_; 
wire u2__abc_52138_new_n6389_; 
wire u2__abc_52138_new_n6390_; 
wire u2__abc_52138_new_n6391_; 
wire u2__abc_52138_new_n6392_; 
wire u2__abc_52138_new_n6393_; 
wire u2__abc_52138_new_n6394_; 
wire u2__abc_52138_new_n6395_; 
wire u2__abc_52138_new_n6396_; 
wire u2__abc_52138_new_n6397_; 
wire u2__abc_52138_new_n6398_; 
wire u2__abc_52138_new_n6399_; 
wire u2__abc_52138_new_n6400_; 
wire u2__abc_52138_new_n6401_; 
wire u2__abc_52138_new_n6402_; 
wire u2__abc_52138_new_n6403_; 
wire u2__abc_52138_new_n6404_; 
wire u2__abc_52138_new_n6405_; 
wire u2__abc_52138_new_n6406_; 
wire u2__abc_52138_new_n6407_; 
wire u2__abc_52138_new_n6408_; 
wire u2__abc_52138_new_n6409_; 
wire u2__abc_52138_new_n6410_; 
wire u2__abc_52138_new_n6411_; 
wire u2__abc_52138_new_n6412_; 
wire u2__abc_52138_new_n6413_; 
wire u2__abc_52138_new_n6414_; 
wire u2__abc_52138_new_n6415_; 
wire u2__abc_52138_new_n6416_; 
wire u2__abc_52138_new_n6417_; 
wire u2__abc_52138_new_n6418_; 
wire u2__abc_52138_new_n6419_; 
wire u2__abc_52138_new_n6420_; 
wire u2__abc_52138_new_n6421_; 
wire u2__abc_52138_new_n6422_; 
wire u2__abc_52138_new_n6423_; 
wire u2__abc_52138_new_n6424_; 
wire u2__abc_52138_new_n6425_; 
wire u2__abc_52138_new_n6426_; 
wire u2__abc_52138_new_n6427_; 
wire u2__abc_52138_new_n6428_; 
wire u2__abc_52138_new_n6429_; 
wire u2__abc_52138_new_n6430_; 
wire u2__abc_52138_new_n6431_; 
wire u2__abc_52138_new_n6432_; 
wire u2__abc_52138_new_n6433_; 
wire u2__abc_52138_new_n6434_; 
wire u2__abc_52138_new_n6435_; 
wire u2__abc_52138_new_n6436_; 
wire u2__abc_52138_new_n6437_; 
wire u2__abc_52138_new_n6438_; 
wire u2__abc_52138_new_n6439_; 
wire u2__abc_52138_new_n6440_; 
wire u2__abc_52138_new_n6441_; 
wire u2__abc_52138_new_n6442_; 
wire u2__abc_52138_new_n6443_; 
wire u2__abc_52138_new_n6444_; 
wire u2__abc_52138_new_n6445_; 
wire u2__abc_52138_new_n6446_; 
wire u2__abc_52138_new_n6447_; 
wire u2__abc_52138_new_n6448_; 
wire u2__abc_52138_new_n6449_; 
wire u2__abc_52138_new_n6450_; 
wire u2__abc_52138_new_n6451_; 
wire u2__abc_52138_new_n6452_; 
wire u2__abc_52138_new_n6453_; 
wire u2__abc_52138_new_n6454_; 
wire u2__abc_52138_new_n6455_; 
wire u2__abc_52138_new_n6456_; 
wire u2__abc_52138_new_n6457_; 
wire u2__abc_52138_new_n6458_; 
wire u2__abc_52138_new_n6459_; 
wire u2__abc_52138_new_n6460_; 
wire u2__abc_52138_new_n6461_; 
wire u2__abc_52138_new_n6462_; 
wire u2__abc_52138_new_n6463_; 
wire u2__abc_52138_new_n6464_; 
wire u2__abc_52138_new_n6465_; 
wire u2__abc_52138_new_n6466_; 
wire u2__abc_52138_new_n6467_; 
wire u2__abc_52138_new_n6468_; 
wire u2__abc_52138_new_n6469_; 
wire u2__abc_52138_new_n6470_; 
wire u2__abc_52138_new_n6471_; 
wire u2__abc_52138_new_n6472_; 
wire u2__abc_52138_new_n6473_; 
wire u2__abc_52138_new_n6474_; 
wire u2__abc_52138_new_n6475_; 
wire u2__abc_52138_new_n6476_; 
wire u2__abc_52138_new_n6477_; 
wire u2__abc_52138_new_n6478_; 
wire u2__abc_52138_new_n6479_; 
wire u2__abc_52138_new_n6480_; 
wire u2__abc_52138_new_n6481_; 
wire u2__abc_52138_new_n6482_; 
wire u2__abc_52138_new_n6483_; 
wire u2__abc_52138_new_n6484_; 
wire u2__abc_52138_new_n6485_; 
wire u2__abc_52138_new_n6486_; 
wire u2__abc_52138_new_n6487_; 
wire u2__abc_52138_new_n6488_; 
wire u2__abc_52138_new_n6489_; 
wire u2__abc_52138_new_n6490_; 
wire u2__abc_52138_new_n6491_; 
wire u2__abc_52138_new_n6492_; 
wire u2__abc_52138_new_n6493_; 
wire u2__abc_52138_new_n6494_; 
wire u2__abc_52138_new_n6495_; 
wire u2__abc_52138_new_n6496_; 
wire u2__abc_52138_new_n6497_; 
wire u2__abc_52138_new_n6498_; 
wire u2__abc_52138_new_n6499_; 
wire u2__abc_52138_new_n6500_; 
wire u2__abc_52138_new_n6501_; 
wire u2__abc_52138_new_n6502_; 
wire u2__abc_52138_new_n6503_; 
wire u2__abc_52138_new_n6504_; 
wire u2__abc_52138_new_n6505_; 
wire u2__abc_52138_new_n6506_; 
wire u2__abc_52138_new_n6507_; 
wire u2__abc_52138_new_n6509_; 
wire u2__abc_52138_new_n6510_; 
wire u2__abc_52138_new_n6511_; 
wire u2__abc_52138_new_n6512_; 
wire u2__abc_52138_new_n6513_; 
wire u2__abc_52138_new_n6514_; 
wire u2__abc_52138_new_n6515_; 
wire u2__abc_52138_new_n6516_; 
wire u2__abc_52138_new_n6517_; 
wire u2__abc_52138_new_n6519_; 
wire u2__abc_52138_new_n6520_; 
wire u2__abc_52138_new_n6521_; 
wire u2__abc_52138_new_n6522_; 
wire u2__abc_52138_new_n6523_; 
wire u2__abc_52138_new_n6524_; 
wire u2__abc_52138_new_n6525_; 
wire u2__abc_52138_new_n6526_; 
wire u2__abc_52138_new_n6528_; 
wire u2__abc_52138_new_n6529_; 
wire u2__abc_52138_new_n6530_; 
wire u2__abc_52138_new_n6531_; 
wire u2__abc_52138_new_n6532_; 
wire u2__abc_52138_new_n6533_; 
wire u2__abc_52138_new_n6534_; 
wire u2__abc_52138_new_n6535_; 
wire u2__abc_52138_new_n6537_; 
wire u2__abc_52138_new_n6538_; 
wire u2__abc_52138_new_n6539_; 
wire u2__abc_52138_new_n6540_; 
wire u2__abc_52138_new_n6541_; 
wire u2__abc_52138_new_n6542_; 
wire u2__abc_52138_new_n6543_; 
wire u2__abc_52138_new_n6544_; 
wire u2__abc_52138_new_n6545_; 
wire u2__abc_52138_new_n6546_; 
wire u2__abc_52138_new_n6547_; 
wire u2__abc_52138_new_n6549_; 
wire u2__abc_52138_new_n6550_; 
wire u2__abc_52138_new_n6551_; 
wire u2__abc_52138_new_n6552_; 
wire u2__abc_52138_new_n6553_; 
wire u2__abc_52138_new_n6554_; 
wire u2__abc_52138_new_n6555_; 
wire u2__abc_52138_new_n6556_; 
wire u2__abc_52138_new_n6558_; 
wire u2__abc_52138_new_n6559_; 
wire u2__abc_52138_new_n6560_; 
wire u2__abc_52138_new_n6561_; 
wire u2__abc_52138_new_n6562_; 
wire u2__abc_52138_new_n6563_; 
wire u2__abc_52138_new_n6564_; 
wire u2__abc_52138_new_n6565_; 
wire u2__abc_52138_new_n6567_; 
wire u2__abc_52138_new_n6568_; 
wire u2__abc_52138_new_n6569_; 
wire u2__abc_52138_new_n6570_; 
wire u2__abc_52138_new_n6571_; 
wire u2__abc_52138_new_n6572_; 
wire u2__abc_52138_new_n6573_; 
wire u2__abc_52138_new_n6575_; 
wire u2__abc_52138_new_n6576_; 
wire u2__abc_52138_new_n6577_; 
wire u2__abc_52138_new_n6578_; 
wire u2__abc_52138_new_n6579_; 
wire u2__abc_52138_new_n6580_; 
wire u2__abc_52138_new_n6581_; 
wire u2__abc_52138_new_n6582_; 
wire u2__abc_52138_new_n6583_; 
wire u2__abc_52138_new_n6584_; 
wire u2__abc_52138_new_n6585_; 
wire u2__abc_52138_new_n6586_; 
wire u2__abc_52138_new_n6587_; 
wire u2__abc_52138_new_n6588_; 
wire u2__abc_52138_new_n6590_; 
wire u2__abc_52138_new_n6591_; 
wire u2__abc_52138_new_n6592_; 
wire u2__abc_52138_new_n6593_; 
wire u2__abc_52138_new_n6594_; 
wire u2__abc_52138_new_n6595_; 
wire u2__abc_52138_new_n6596_; 
wire u2__abc_52138_new_n6598_; 
wire u2__abc_52138_new_n6599_; 
wire u2__abc_52138_new_n6600_; 
wire u2__abc_52138_new_n6601_; 
wire u2__abc_52138_new_n6602_; 
wire u2__abc_52138_new_n6603_; 
wire u2__abc_52138_new_n6604_; 
wire u2__abc_52138_new_n6605_; 
wire u2__abc_52138_new_n6606_; 
wire u2__abc_52138_new_n6607_; 
wire u2__abc_52138_new_n6608_; 
wire u2__abc_52138_new_n6609_; 
wire u2__abc_52138_new_n6610_; 
wire u2__abc_52138_new_n6611_; 
wire u2__abc_52138_new_n6613_; 
wire u2__abc_52138_new_n6614_; 
wire u2__abc_52138_new_n6615_; 
wire u2__abc_52138_new_n6616_; 
wire u2__abc_52138_new_n6617_; 
wire u2__abc_52138_new_n6618_; 
wire u2__abc_52138_new_n6619_; 
wire u2__abc_52138_new_n6620_; 
wire u2__abc_52138_new_n6621_; 
wire u2__abc_52138_new_n6623_; 
wire u2__abc_52138_new_n6624_; 
wire u2__abc_52138_new_n6625_; 
wire u2__abc_52138_new_n6626_; 
wire u2__abc_52138_new_n6627_; 
wire u2__abc_52138_new_n6628_; 
wire u2__abc_52138_new_n6629_; 
wire u2__abc_52138_new_n6630_; 
wire u2__abc_52138_new_n6631_; 
wire u2__abc_52138_new_n6632_; 
wire u2__abc_52138_new_n6634_; 
wire u2__abc_52138_new_n6635_; 
wire u2__abc_52138_new_n6636_; 
wire u2__abc_52138_new_n6637_; 
wire u2__abc_52138_new_n6638_; 
wire u2__abc_52138_new_n6639_; 
wire u2__abc_52138_new_n6640_; 
wire u2__abc_52138_new_n6642_; 
wire u2__abc_52138_new_n6643_; 
wire u2__abc_52138_new_n6644_; 
wire u2__abc_52138_new_n6645_; 
wire u2__abc_52138_new_n6646_; 
wire u2__abc_52138_new_n6647_; 
wire u2__abc_52138_new_n6648_; 
wire u2__abc_52138_new_n6649_; 
wire u2__abc_52138_new_n6650_; 
wire u2__abc_52138_new_n6652_; 
wire u2__abc_52138_new_n6653_; 
wire u2__abc_52138_new_n6654_; 
wire u2__abc_52138_new_n6655_; 
wire u2__abc_52138_new_n6656_; 
wire u2__abc_52138_new_n6657_; 
wire u2__abc_52138_new_n6658_; 
wire u2__abc_52138_new_n6659_; 
wire u2__abc_52138_new_n6660_; 
wire u2__abc_52138_new_n6661_; 
wire u2__abc_52138_new_n6663_; 
wire u2__abc_52138_new_n6664_; 
wire u2__abc_52138_new_n6665_; 
wire u2__abc_52138_new_n6666_; 
wire u2__abc_52138_new_n6667_; 
wire u2__abc_52138_new_n6668_; 
wire u2__abc_52138_new_n6669_; 
wire u2__abc_52138_new_n6670_; 
wire u2__abc_52138_new_n6671_; 
wire u2__abc_52138_new_n6672_; 
wire u2__abc_52138_new_n6673_; 
wire u2__abc_52138_new_n6674_; 
wire u2__abc_52138_new_n6675_; 
wire u2__abc_52138_new_n6676_; 
wire u2__abc_52138_new_n6677_; 
wire u2__abc_52138_new_n6678_; 
wire u2__abc_52138_new_n6679_; 
wire u2__abc_52138_new_n6680_; 
wire u2__abc_52138_new_n6682_; 
wire u2__abc_52138_new_n6683_; 
wire u2__abc_52138_new_n6684_; 
wire u2__abc_52138_new_n6685_; 
wire u2__abc_52138_new_n6686_; 
wire u2__abc_52138_new_n6687_; 
wire u2__abc_52138_new_n6688_; 
wire u2__abc_52138_new_n6690_; 
wire u2__abc_52138_new_n6691_; 
wire u2__abc_52138_new_n6692_; 
wire u2__abc_52138_new_n6693_; 
wire u2__abc_52138_new_n6694_; 
wire u2__abc_52138_new_n6695_; 
wire u2__abc_52138_new_n6696_; 
wire u2__abc_52138_new_n6697_; 
wire u2__abc_52138_new_n6698_; 
wire u2__abc_52138_new_n6699_; 
wire u2__abc_52138_new_n6701_; 
wire u2__abc_52138_new_n6702_; 
wire u2__abc_52138_new_n6703_; 
wire u2__abc_52138_new_n6704_; 
wire u2__abc_52138_new_n6705_; 
wire u2__abc_52138_new_n6706_; 
wire u2__abc_52138_new_n6707_; 
wire u2__abc_52138_new_n6708_; 
wire u2__abc_52138_new_n6710_; 
wire u2__abc_52138_new_n6711_; 
wire u2__abc_52138_new_n6712_; 
wire u2__abc_52138_new_n6713_; 
wire u2__abc_52138_new_n6714_; 
wire u2__abc_52138_new_n6715_; 
wire u2__abc_52138_new_n6716_; 
wire u2__abc_52138_new_n6717_; 
wire u2__abc_52138_new_n6718_; 
wire u2__abc_52138_new_n6719_; 
wire u2__abc_52138_new_n6720_; 
wire u2__abc_52138_new_n6721_; 
wire u2__abc_52138_new_n6722_; 
wire u2__abc_52138_new_n6724_; 
wire u2__abc_52138_new_n6725_; 
wire u2__abc_52138_new_n6726_; 
wire u2__abc_52138_new_n6727_; 
wire u2__abc_52138_new_n6728_; 
wire u2__abc_52138_new_n6729_; 
wire u2__abc_52138_new_n6730_; 
wire u2__abc_52138_new_n6732_; 
wire u2__abc_52138_new_n6733_; 
wire u2__abc_52138_new_n6734_; 
wire u2__abc_52138_new_n6735_; 
wire u2__abc_52138_new_n6736_; 
wire u2__abc_52138_new_n6737_; 
wire u2__abc_52138_new_n6738_; 
wire u2__abc_52138_new_n6739_; 
wire u2__abc_52138_new_n6740_; 
wire u2__abc_52138_new_n6741_; 
wire u2__abc_52138_new_n6742_; 
wire u2__abc_52138_new_n6743_; 
wire u2__abc_52138_new_n6744_; 
wire u2__abc_52138_new_n6746_; 
wire u2__abc_52138_new_n6747_; 
wire u2__abc_52138_new_n6748_; 
wire u2__abc_52138_new_n6749_; 
wire u2__abc_52138_new_n6750_; 
wire u2__abc_52138_new_n6751_; 
wire u2__abc_52138_new_n6752_; 
wire u2__abc_52138_new_n6753_; 
wire u2__abc_52138_new_n6755_; 
wire u2__abc_52138_new_n6756_; 
wire u2__abc_52138_new_n6757_; 
wire u2__abc_52138_new_n6758_; 
wire u2__abc_52138_new_n6759_; 
wire u2__abc_52138_new_n6760_; 
wire u2__abc_52138_new_n6761_; 
wire u2__abc_52138_new_n6762_; 
wire u2__abc_52138_new_n6763_; 
wire u2__abc_52138_new_n6764_; 
wire u2__abc_52138_new_n6765_; 
wire u2__abc_52138_new_n6766_; 
wire u2__abc_52138_new_n6767_; 
wire u2__abc_52138_new_n6768_; 
wire u2__abc_52138_new_n6769_; 
wire u2__abc_52138_new_n6770_; 
wire u2__abc_52138_new_n6772_; 
wire u2__abc_52138_new_n6773_; 
wire u2__abc_52138_new_n6774_; 
wire u2__abc_52138_new_n6775_; 
wire u2__abc_52138_new_n6776_; 
wire u2__abc_52138_new_n6777_; 
wire u2__abc_52138_new_n6778_; 
wire u2__abc_52138_new_n6780_; 
wire u2__abc_52138_new_n6781_; 
wire u2__abc_52138_new_n6782_; 
wire u2__abc_52138_new_n6783_; 
wire u2__abc_52138_new_n6784_; 
wire u2__abc_52138_new_n6785_; 
wire u2__abc_52138_new_n6786_; 
wire u2__abc_52138_new_n6787_; 
wire u2__abc_52138_new_n6788_; 
wire u2__abc_52138_new_n6789_; 
wire u2__abc_52138_new_n6790_; 
wire u2__abc_52138_new_n6792_; 
wire u2__abc_52138_new_n6793_; 
wire u2__abc_52138_new_n6794_; 
wire u2__abc_52138_new_n6795_; 
wire u2__abc_52138_new_n6796_; 
wire u2__abc_52138_new_n6797_; 
wire u2__abc_52138_new_n6798_; 
wire u2__abc_52138_new_n6800_; 
wire u2__abc_52138_new_n6801_; 
wire u2__abc_52138_new_n6802_; 
wire u2__abc_52138_new_n6803_; 
wire u2__abc_52138_new_n6804_; 
wire u2__abc_52138_new_n6805_; 
wire u2__abc_52138_new_n6806_; 
wire u2__abc_52138_new_n6807_; 
wire u2__abc_52138_new_n6808_; 
wire u2__abc_52138_new_n6809_; 
wire u2__abc_52138_new_n6810_; 
wire u2__abc_52138_new_n6811_; 
wire u2__abc_52138_new_n6812_; 
wire u2__abc_52138_new_n6813_; 
wire u2__abc_52138_new_n6815_; 
wire u2__abc_52138_new_n6816_; 
wire u2__abc_52138_new_n6817_; 
wire u2__abc_52138_new_n6818_; 
wire u2__abc_52138_new_n6819_; 
wire u2__abc_52138_new_n6820_; 
wire u2__abc_52138_new_n6821_; 
wire u2__abc_52138_new_n6823_; 
wire u2__abc_52138_new_n6824_; 
wire u2__abc_52138_new_n6825_; 
wire u2__abc_52138_new_n6826_; 
wire u2__abc_52138_new_n6827_; 
wire u2__abc_52138_new_n6828_; 
wire u2__abc_52138_new_n6829_; 
wire u2__abc_52138_new_n6830_; 
wire u2__abc_52138_new_n6832_; 
wire u2__abc_52138_new_n6833_; 
wire u2__abc_52138_new_n6834_; 
wire u2__abc_52138_new_n6835_; 
wire u2__abc_52138_new_n6836_; 
wire u2__abc_52138_new_n6837_; 
wire u2__abc_52138_new_n6838_; 
wire u2__abc_52138_new_n6840_; 
wire u2__abc_52138_new_n6841_; 
wire u2__abc_52138_new_n6842_; 
wire u2__abc_52138_new_n6843_; 
wire u2__abc_52138_new_n6844_; 
wire u2__abc_52138_new_n6845_; 
wire u2__abc_52138_new_n6846_; 
wire u2__abc_52138_new_n6847_; 
wire u2__abc_52138_new_n6848_; 
wire u2__abc_52138_new_n6849_; 
wire u2__abc_52138_new_n6850_; 
wire u2__abc_52138_new_n6852_; 
wire u2__abc_52138_new_n6853_; 
wire u2__abc_52138_new_n6854_; 
wire u2__abc_52138_new_n6855_; 
wire u2__abc_52138_new_n6856_; 
wire u2__abc_52138_new_n6857_; 
wire u2__abc_52138_new_n6858_; 
wire u2__abc_52138_new_n6859_; 
wire u2__abc_52138_new_n6861_; 
wire u2__abc_52138_new_n6862_; 
wire u2__abc_52138_new_n6863_; 
wire u2__abc_52138_new_n6864_; 
wire u2__abc_52138_new_n6865_; 
wire u2__abc_52138_new_n6866_; 
wire u2__abc_52138_new_n6867_; 
wire u2__abc_52138_new_n6868_; 
wire u2__abc_52138_new_n6869_; 
wire u2__abc_52138_new_n6871_; 
wire u2__abc_52138_new_n6872_; 
wire u2__abc_52138_new_n6873_; 
wire u2__abc_52138_new_n6874_; 
wire u2__abc_52138_new_n6875_; 
wire u2__abc_52138_new_n6876_; 
wire u2__abc_52138_new_n6877_; 
wire u2__abc_52138_new_n6878_; 
wire u2__abc_52138_new_n6880_; 
wire u2__abc_52138_new_n6881_; 
wire u2__abc_52138_new_n6882_; 
wire u2__abc_52138_new_n6883_; 
wire u2__abc_52138_new_n6884_; 
wire u2__abc_52138_new_n6885_; 
wire u2__abc_52138_new_n6886_; 
wire u2__abc_52138_new_n6887_; 
wire u2__abc_52138_new_n6888_; 
wire u2__abc_52138_new_n6889_; 
wire u2__abc_52138_new_n6890_; 
wire u2__abc_52138_new_n6891_; 
wire u2__abc_52138_new_n6892_; 
wire u2__abc_52138_new_n6894_; 
wire u2__abc_52138_new_n6895_; 
wire u2__abc_52138_new_n6896_; 
wire u2__abc_52138_new_n6897_; 
wire u2__abc_52138_new_n6898_; 
wire u2__abc_52138_new_n6899_; 
wire u2__abc_52138_new_n6900_; 
wire u2__abc_52138_new_n6901_; 
wire u2__abc_52138_new_n6903_; 
wire u2__abc_52138_new_n6904_; 
wire u2__abc_52138_new_n6905_; 
wire u2__abc_52138_new_n6906_; 
wire u2__abc_52138_new_n6907_; 
wire u2__abc_52138_new_n6908_; 
wire u2__abc_52138_new_n6909_; 
wire u2__abc_52138_new_n6910_; 
wire u2__abc_52138_new_n6911_; 
wire u2__abc_52138_new_n6912_; 
wire u2__abc_52138_new_n6914_; 
wire u2__abc_52138_new_n6915_; 
wire u2__abc_52138_new_n6916_; 
wire u2__abc_52138_new_n6917_; 
wire u2__abc_52138_new_n6918_; 
wire u2__abc_52138_new_n6919_; 
wire u2__abc_52138_new_n6920_; 
wire u2__abc_52138_new_n6922_; 
wire u2__abc_52138_new_n6923_; 
wire u2__abc_52138_new_n6924_; 
wire u2__abc_52138_new_n6925_; 
wire u2__abc_52138_new_n6926_; 
wire u2__abc_52138_new_n6927_; 
wire u2__abc_52138_new_n6928_; 
wire u2__abc_52138_new_n6929_; 
wire u2__abc_52138_new_n6930_; 
wire u2__abc_52138_new_n6931_; 
wire u2__abc_52138_new_n6932_; 
wire u2__abc_52138_new_n6933_; 
wire u2__abc_52138_new_n6934_; 
wire u2__abc_52138_new_n6935_; 
wire u2__abc_52138_new_n6936_; 
wire u2__abc_52138_new_n6938_; 
wire u2__abc_52138_new_n6939_; 
wire u2__abc_52138_new_n6940_; 
wire u2__abc_52138_new_n6941_; 
wire u2__abc_52138_new_n6942_; 
wire u2__abc_52138_new_n6943_; 
wire u2__abc_52138_new_n6944_; 
wire u2__abc_52138_new_n6946_; 
wire u2__abc_52138_new_n6947_; 
wire u2__abc_52138_new_n6948_; 
wire u2__abc_52138_new_n6949_; 
wire u2__abc_52138_new_n6950_; 
wire u2__abc_52138_new_n6951_; 
wire u2__abc_52138_new_n6952_; 
wire u2__abc_52138_new_n6953_; 
wire u2__abc_52138_new_n6955_; 
wire u2__abc_52138_new_n6956_; 
wire u2__abc_52138_new_n6957_; 
wire u2__abc_52138_new_n6958_; 
wire u2__abc_52138_new_n6959_; 
wire u2__abc_52138_new_n6960_; 
wire u2__abc_52138_new_n6961_; 
wire u2__abc_52138_new_n6962_; 
wire u2__abc_52138_new_n6963_; 
wire u2__abc_52138_new_n6965_; 
wire u2__abc_52138_new_n6966_; 
wire u2__abc_52138_new_n6967_; 
wire u2__abc_52138_new_n6968_; 
wire u2__abc_52138_new_n6969_; 
wire u2__abc_52138_new_n6970_; 
wire u2__abc_52138_new_n6971_; 
wire u2__abc_52138_new_n6972_; 
wire u2__abc_52138_new_n6973_; 
wire u2__abc_52138_new_n6974_; 
wire u2__abc_52138_new_n6975_; 
wire u2__abc_52138_new_n6976_; 
wire u2__abc_52138_new_n6977_; 
wire u2__abc_52138_new_n6979_; 
wire u2__abc_52138_new_n6980_; 
wire u2__abc_52138_new_n6981_; 
wire u2__abc_52138_new_n6982_; 
wire u2__abc_52138_new_n6983_; 
wire u2__abc_52138_new_n6984_; 
wire u2__abc_52138_new_n6985_; 
wire u2__abc_52138_new_n6987_; 
wire u2__abc_52138_new_n6988_; 
wire u2__abc_52138_new_n6989_; 
wire u2__abc_52138_new_n6990_; 
wire u2__abc_52138_new_n6991_; 
wire u2__abc_52138_new_n6992_; 
wire u2__abc_52138_new_n6993_; 
wire u2__abc_52138_new_n6994_; 
wire u2__abc_52138_new_n6995_; 
wire u2__abc_52138_new_n6997_; 
wire u2__abc_52138_new_n6998_; 
wire u2__abc_52138_new_n6999_; 
wire u2__abc_52138_new_n7000_; 
wire u2__abc_52138_new_n7001_; 
wire u2__abc_52138_new_n7002_; 
wire u2__abc_52138_new_n7003_; 
wire u2__abc_52138_new_n7004_; 
wire u2__abc_52138_new_n7006_; 
wire u2__abc_52138_new_n7007_; 
wire u2__abc_52138_new_n7008_; 
wire u2__abc_52138_new_n7009_; 
wire u2__abc_52138_new_n7010_; 
wire u2__abc_52138_new_n7011_; 
wire u2__abc_52138_new_n7012_; 
wire u2__abc_52138_new_n7013_; 
wire u2__abc_52138_new_n7014_; 
wire u2__abc_52138_new_n7015_; 
wire u2__abc_52138_new_n7016_; 
wire u2__abc_52138_new_n7017_; 
wire u2__abc_52138_new_n7018_; 
wire u2__abc_52138_new_n7019_; 
wire u2__abc_52138_new_n7021_; 
wire u2__abc_52138_new_n7022_; 
wire u2__abc_52138_new_n7023_; 
wire u2__abc_52138_new_n7024_; 
wire u2__abc_52138_new_n7025_; 
wire u2__abc_52138_new_n7026_; 
wire u2__abc_52138_new_n7027_; 
wire u2__abc_52138_new_n7029_; 
wire u2__abc_52138_new_n7030_; 
wire u2__abc_52138_new_n7031_; 
wire u2__abc_52138_new_n7032_; 
wire u2__abc_52138_new_n7033_; 
wire u2__abc_52138_new_n7034_; 
wire u2__abc_52138_new_n7035_; 
wire u2__abc_52138_new_n7036_; 
wire u2__abc_52138_new_n7037_; 
wire u2__abc_52138_new_n7038_; 
wire u2__abc_52138_new_n7039_; 
wire u2__abc_52138_new_n7040_; 
wire u2__abc_52138_new_n7042_; 
wire u2__abc_52138_new_n7043_; 
wire u2__abc_52138_new_n7044_; 
wire u2__abc_52138_new_n7045_; 
wire u2__abc_52138_new_n7046_; 
wire u2__abc_52138_new_n7047_; 
wire u2__abc_52138_new_n7048_; 
wire u2__abc_52138_new_n7050_; 
wire u2__abc_52138_new_n7051_; 
wire u2__abc_52138_new_n7052_; 
wire u2__abc_52138_new_n7053_; 
wire u2__abc_52138_new_n7054_; 
wire u2__abc_52138_new_n7055_; 
wire u2__abc_52138_new_n7056_; 
wire u2__abc_52138_new_n7057_; 
wire u2__abc_52138_new_n7058_; 
wire u2__abc_52138_new_n7059_; 
wire u2__abc_52138_new_n7060_; 
wire u2__abc_52138_new_n7061_; 
wire u2__abc_52138_new_n7062_; 
wire u2__abc_52138_new_n7064_; 
wire u2__abc_52138_new_n7065_; 
wire u2__abc_52138_new_n7066_; 
wire u2__abc_52138_new_n7067_; 
wire u2__abc_52138_new_n7068_; 
wire u2__abc_52138_new_n7069_; 
wire u2__abc_52138_new_n7070_; 
wire u2__abc_52138_new_n7072_; 
wire u2__abc_52138_new_n7073_; 
wire u2__abc_52138_new_n7074_; 
wire u2__abc_52138_new_n7075_; 
wire u2__abc_52138_new_n7076_; 
wire u2__abc_52138_new_n7077_; 
wire u2__abc_52138_new_n7078_; 
wire u2__abc_52138_new_n7079_; 
wire u2__abc_52138_new_n7080_; 
wire u2__abc_52138_new_n7081_; 
wire u2__abc_52138_new_n7083_; 
wire u2__abc_52138_new_n7084_; 
wire u2__abc_52138_new_n7085_; 
wire u2__abc_52138_new_n7086_; 
wire u2__abc_52138_new_n7087_; 
wire u2__abc_52138_new_n7088_; 
wire u2__abc_52138_new_n7089_; 
wire u2__abc_52138_new_n7090_; 
wire u2__abc_52138_new_n7092_; 
wire u2__abc_52138_new_n7093_; 
wire u2__abc_52138_new_n7094_; 
wire u2__abc_52138_new_n7095_; 
wire u2__abc_52138_new_n7096_; 
wire u2__abc_52138_new_n7097_; 
wire u2__abc_52138_new_n7098_; 
wire u2__abc_52138_new_n7099_; 
wire u2__abc_52138_new_n7100_; 
wire u2__abc_52138_new_n7101_; 
wire u2__abc_52138_new_n7102_; 
wire u2__abc_52138_new_n7103_; 
wire u2__abc_52138_new_n7104_; 
wire u2__abc_52138_new_n7105_; 
wire u2__abc_52138_new_n7106_; 
wire u2__abc_52138_new_n7108_; 
wire u2__abc_52138_new_n7109_; 
wire u2__abc_52138_new_n7110_; 
wire u2__abc_52138_new_n7111_; 
wire u2__abc_52138_new_n7112_; 
wire u2__abc_52138_new_n7113_; 
wire u2__abc_52138_new_n7114_; 
wire u2__abc_52138_new_n7116_; 
wire u2__abc_52138_new_n7117_; 
wire u2__abc_52138_new_n7118_; 
wire u2__abc_52138_new_n7119_; 
wire u2__abc_52138_new_n7120_; 
wire u2__abc_52138_new_n7121_; 
wire u2__abc_52138_new_n7122_; 
wire u2__abc_52138_new_n7123_; 
wire u2__abc_52138_new_n7125_; 
wire u2__abc_52138_new_n7126_; 
wire u2__abc_52138_new_n7127_; 
wire u2__abc_52138_new_n7128_; 
wire u2__abc_52138_new_n7129_; 
wire u2__abc_52138_new_n7130_; 
wire u2__abc_52138_new_n7131_; 
wire u2__abc_52138_new_n7132_; 
wire u2__abc_52138_new_n7134_; 
wire u2__abc_52138_new_n7135_; 
wire u2__abc_52138_new_n7136_; 
wire u2__abc_52138_new_n7137_; 
wire u2__abc_52138_new_n7138_; 
wire u2__abc_52138_new_n7139_; 
wire u2__abc_52138_new_n7140_; 
wire u2__abc_52138_new_n7141_; 
wire u2__abc_52138_new_n7142_; 
wire u2__abc_52138_new_n7143_; 
wire u2__abc_52138_new_n7144_; 
wire u2__abc_52138_new_n7145_; 
wire u2__abc_52138_new_n7146_; 
wire u2__abc_52138_new_n7147_; 
wire u2__abc_52138_new_n7149_; 
wire u2__abc_52138_new_n7150_; 
wire u2__abc_52138_new_n7151_; 
wire u2__abc_52138_new_n7152_; 
wire u2__abc_52138_new_n7153_; 
wire u2__abc_52138_new_n7154_; 
wire u2__abc_52138_new_n7155_; 
wire u2__abc_52138_new_n7156_; 
wire u2__abc_52138_new_n7157_; 
wire u2__abc_52138_new_n7159_; 
wire u2__abc_52138_new_n7160_; 
wire u2__abc_52138_new_n7161_; 
wire u2__abc_52138_new_n7162_; 
wire u2__abc_52138_new_n7163_; 
wire u2__abc_52138_new_n7164_; 
wire u2__abc_52138_new_n7165_; 
wire u2__abc_52138_new_n7166_; 
wire u2__abc_52138_new_n7168_; 
wire u2__abc_52138_new_n7169_; 
wire u2__abc_52138_new_n7170_; 
wire u2__abc_52138_new_n7171_; 
wire u2__abc_52138_new_n7172_; 
wire u2__abc_52138_new_n7173_; 
wire u2__abc_52138_new_n7174_; 
wire u2__abc_52138_new_n7176_; 
wire u2__abc_52138_new_n7177_; 
wire u2__abc_52138_new_n7178_; 
wire u2__abc_52138_new_n7179_; 
wire u2__abc_52138_new_n7180_; 
wire u2__abc_52138_new_n7181_; 
wire u2__abc_52138_new_n7182_; 
wire u2__abc_52138_new_n7183_; 
wire u2__abc_52138_new_n7184_; 
wire u2__abc_52138_new_n7185_; 
wire u2__abc_52138_new_n7186_; 
wire u2__abc_52138_new_n7187_; 
wire u2__abc_52138_new_n7188_; 
wire u2__abc_52138_new_n7189_; 
wire u2__abc_52138_new_n7190_; 
wire u2__abc_52138_new_n7191_; 
wire u2__abc_52138_new_n7192_; 
wire u2__abc_52138_new_n7194_; 
wire u2__abc_52138_new_n7195_; 
wire u2__abc_52138_new_n7196_; 
wire u2__abc_52138_new_n7197_; 
wire u2__abc_52138_new_n7198_; 
wire u2__abc_52138_new_n7199_; 
wire u2__abc_52138_new_n7200_; 
wire u2__abc_52138_new_n7202_; 
wire u2__abc_52138_new_n7203_; 
wire u2__abc_52138_new_n7204_; 
wire u2__abc_52138_new_n7205_; 
wire u2__abc_52138_new_n7206_; 
wire u2__abc_52138_new_n7207_; 
wire u2__abc_52138_new_n7208_; 
wire u2__abc_52138_new_n7209_; 
wire u2__abc_52138_new_n7211_; 
wire u2__abc_52138_new_n7212_; 
wire u2__abc_52138_new_n7213_; 
wire u2__abc_52138_new_n7214_; 
wire u2__abc_52138_new_n7215_; 
wire u2__abc_52138_new_n7216_; 
wire u2__abc_52138_new_n7217_; 
wire u2__abc_52138_new_n7218_; 
wire u2__abc_52138_new_n7219_; 
wire u2__abc_52138_new_n7221_; 
wire u2__abc_52138_new_n7222_; 
wire u2__abc_52138_new_n7223_; 
wire u2__abc_52138_new_n7224_; 
wire u2__abc_52138_new_n7225_; 
wire u2__abc_52138_new_n7226_; 
wire u2__abc_52138_new_n7227_; 
wire u2__abc_52138_new_n7228_; 
wire u2__abc_52138_new_n7229_; 
wire u2__abc_52138_new_n7230_; 
wire u2__abc_52138_new_n7231_; 
wire u2__abc_52138_new_n7232_; 
wire u2__abc_52138_new_n7234_; 
wire u2__abc_52138_new_n7235_; 
wire u2__abc_52138_new_n7236_; 
wire u2__abc_52138_new_n7237_; 
wire u2__abc_52138_new_n7238_; 
wire u2__abc_52138_new_n7239_; 
wire u2__abc_52138_new_n7240_; 
wire u2__abc_52138_new_n7242_; 
wire u2__abc_52138_new_n7243_; 
wire u2__abc_52138_new_n7244_; 
wire u2__abc_52138_new_n7245_; 
wire u2__abc_52138_new_n7246_; 
wire u2__abc_52138_new_n7247_; 
wire u2__abc_52138_new_n7248_; 
wire u2__abc_52138_new_n7249_; 
wire u2__abc_52138_new_n7251_; 
wire u2__abc_52138_new_n7252_; 
wire u2__abc_52138_new_n7253_; 
wire u2__abc_52138_new_n7254_; 
wire u2__abc_52138_new_n7255_; 
wire u2__abc_52138_new_n7256_; 
wire u2__abc_52138_new_n7257_; 
wire u2__abc_52138_new_n7258_; 
wire u2__abc_52138_new_n7259_; 
wire u2__abc_52138_new_n7261_; 
wire u2__abc_52138_new_n7262_; 
wire u2__abc_52138_new_n7263_; 
wire u2__abc_52138_new_n7264_; 
wire u2__abc_52138_new_n7265_; 
wire u2__abc_52138_new_n7266_; 
wire u2__abc_52138_new_n7267_; 
wire u2__abc_52138_new_n7268_; 
wire u2__abc_52138_new_n7269_; 
wire u2__abc_52138_new_n7270_; 
wire u2__abc_52138_new_n7271_; 
wire u2__abc_52138_new_n7272_; 
wire u2__abc_52138_new_n7273_; 
wire u2__abc_52138_new_n7274_; 
wire u2__abc_52138_new_n7275_; 
wire u2__abc_52138_new_n7276_; 
wire u2__abc_52138_new_n7277_; 
wire u2__abc_52138_new_n7279_; 
wire u2__abc_52138_new_n7280_; 
wire u2__abc_52138_new_n7281_; 
wire u2__abc_52138_new_n7282_; 
wire u2__abc_52138_new_n7283_; 
wire u2__abc_52138_new_n7284_; 
wire u2__abc_52138_new_n7285_; 
wire u2__abc_52138_new_n7287_; 
wire u2__abc_52138_new_n7288_; 
wire u2__abc_52138_new_n7289_; 
wire u2__abc_52138_new_n7290_; 
wire u2__abc_52138_new_n7291_; 
wire u2__abc_52138_new_n7292_; 
wire u2__abc_52138_new_n7293_; 
wire u2__abc_52138_new_n7294_; 
wire u2__abc_52138_new_n7295_; 
wire u2__abc_52138_new_n7297_; 
wire u2__abc_52138_new_n7298_; 
wire u2__abc_52138_new_n7299_; 
wire u2__abc_52138_new_n7300_; 
wire u2__abc_52138_new_n7301_; 
wire u2__abc_52138_new_n7302_; 
wire u2__abc_52138_new_n7303_; 
wire u2__abc_52138_new_n7304_; 
wire u2__abc_52138_new_n7305_; 
wire u2__abc_52138_new_n7307_; 
wire u2__abc_52138_new_n7308_; 
wire u2__abc_52138_new_n7309_; 
wire u2__abc_52138_new_n7310_; 
wire u2__abc_52138_new_n7311_; 
wire u2__abc_52138_new_n7312_; 
wire u2__abc_52138_new_n7313_; 
wire u2__abc_52138_new_n7314_; 
wire u2__abc_52138_new_n7315_; 
wire u2__abc_52138_new_n7316_; 
wire u2__abc_52138_new_n7317_; 
wire u2__abc_52138_new_n7318_; 
wire u2__abc_52138_new_n7319_; 
wire u2__abc_52138_new_n7320_; 
wire u2__abc_52138_new_n7321_; 
wire u2__abc_52138_new_n7322_; 
wire u2__abc_52138_new_n7324_; 
wire u2__abc_52138_new_n7325_; 
wire u2__abc_52138_new_n7326_; 
wire u2__abc_52138_new_n7327_; 
wire u2__abc_52138_new_n7328_; 
wire u2__abc_52138_new_n7329_; 
wire u2__abc_52138_new_n7330_; 
wire u2__abc_52138_new_n7331_; 
wire u2__abc_52138_new_n7332_; 
wire u2__abc_52138_new_n7334_; 
wire u2__abc_52138_new_n7335_; 
wire u2__abc_52138_new_n7336_; 
wire u2__abc_52138_new_n7337_; 
wire u2__abc_52138_new_n7338_; 
wire u2__abc_52138_new_n7339_; 
wire u2__abc_52138_new_n7340_; 
wire u2__abc_52138_new_n7341_; 
wire u2__abc_52138_new_n7343_; 
wire u2__abc_52138_new_n7344_; 
wire u2__abc_52138_new_n7345_; 
wire u2__abc_52138_new_n7346_; 
wire u2__abc_52138_new_n7347_; 
wire u2__abc_52138_new_n7348_; 
wire u2__abc_52138_new_n7349_; 
wire u2__abc_52138_new_n7351_; 
wire u2__abc_52138_new_n7352_; 
wire u2__abc_52138_new_n7353_; 
wire u2__abc_52138_new_n7354_; 
wire u2__abc_52138_new_n7355_; 
wire u2__abc_52138_new_n7356_; 
wire u2__abc_52138_new_n7357_; 
wire u2__abc_52138_new_n7358_; 
wire u2__abc_52138_new_n7359_; 
wire u2__abc_52138_new_n7360_; 
wire u2__abc_52138_new_n7361_; 
wire u2__abc_52138_new_n7362_; 
wire u2__abc_52138_new_n7363_; 
wire u2__abc_52138_new_n7364_; 
wire u2__abc_52138_new_n7365_; 
wire u2__abc_52138_new_n7366_; 
wire u2__abc_52138_new_n7367_; 
wire u2__abc_52138_new_n7368_; 
wire u2__abc_52138_new_n7370_; 
wire u2__abc_52138_new_n7371_; 
wire u2__abc_52138_new_n7372_; 
wire u2__abc_52138_new_n7373_; 
wire u2__abc_52138_new_n7374_; 
wire u2__abc_52138_new_n7375_; 
wire u2__abc_52138_new_n7376_; 
wire u2__abc_52138_new_n7377_; 
wire u2__abc_52138_new_n7379_; 
wire u2__abc_52138_new_n7380_; 
wire u2__abc_52138_new_n7381_; 
wire u2__abc_52138_new_n7382_; 
wire u2__abc_52138_new_n7383_; 
wire u2__abc_52138_new_n7384_; 
wire u2__abc_52138_new_n7385_; 
wire u2__abc_52138_new_n7386_; 
wire u2__abc_52138_new_n7387_; 
wire u2__abc_52138_new_n7389_; 
wire u2__abc_52138_new_n7390_; 
wire u2__abc_52138_new_n7391_; 
wire u2__abc_52138_new_n7392_; 
wire u2__abc_52138_new_n7393_; 
wire u2__abc_52138_new_n7394_; 
wire u2__abc_52138_new_n7395_; 
wire u2__abc_52138_new_n7396_; 
wire u2__abc_52138_new_n7398_; 
wire u2__abc_52138_new_n7399_; 
wire u2__abc_52138_new_n7400_; 
wire u2__abc_52138_new_n7401_; 
wire u2__abc_52138_new_n7402_; 
wire u2__abc_52138_new_n7403_; 
wire u2__abc_52138_new_n7404_; 
wire u2__abc_52138_new_n7405_; 
wire u2__abc_52138_new_n7406_; 
wire u2__abc_52138_new_n7407_; 
wire u2__abc_52138_new_n7408_; 
wire u2__abc_52138_new_n7409_; 
wire u2__abc_52138_new_n7410_; 
wire u2__abc_52138_new_n7411_; 
wire u2__abc_52138_new_n7412_; 
wire u2__abc_52138_new_n7413_; 
wire u2__abc_52138_new_n7414_; 
wire u2__abc_52138_new_n7416_; 
wire u2__abc_52138_new_n7417_; 
wire u2__abc_52138_new_n7418_; 
wire u2__abc_52138_new_n7419_; 
wire u2__abc_52138_new_n7420_; 
wire u2__abc_52138_new_n7421_; 
wire u2__abc_52138_new_n7422_; 
wire u2__abc_52138_new_n7424_; 
wire u2__abc_52138_new_n7425_; 
wire u2__abc_52138_new_n7426_; 
wire u2__abc_52138_new_n7427_; 
wire u2__abc_52138_new_n7428_; 
wire u2__abc_52138_new_n7429_; 
wire u2__abc_52138_new_n7430_; 
wire u2__abc_52138_new_n7431_; 
wire u2__abc_52138_new_n7432_; 
wire u2__abc_52138_new_n7433_; 
wire u2__abc_52138_new_n7435_; 
wire u2__abc_52138_new_n7436_; 
wire u2__abc_52138_new_n7437_; 
wire u2__abc_52138_new_n7438_; 
wire u2__abc_52138_new_n7439_; 
wire u2__abc_52138_new_n7440_; 
wire u2__abc_52138_new_n7441_; 
wire u2__abc_52138_new_n7442_; 
wire u2__abc_52138_new_n7443_; 
wire u2__abc_52138_new_n7445_; 
wire u2__abc_52138_new_n7446_; 
wire u2__abc_52138_new_n7447_; 
wire u2__abc_52138_new_n7448_; 
wire u2__abc_52138_new_n7449_; 
wire u2__abc_52138_new_n7450_; 
wire u2__abc_52138_new_n7451_; 
wire u2__abc_52138_new_n7452_; 
wire u2__abc_52138_new_n7453_; 
wire u2__abc_52138_new_n7454_; 
wire u2__abc_52138_new_n7455_; 
wire u2__abc_52138_new_n7456_; 
wire u2__abc_52138_new_n7457_; 
wire u2__abc_52138_new_n7458_; 
wire u2__abc_52138_new_n7459_; 
wire u2__abc_52138_new_n7461_; 
wire u2__abc_52138_new_n7462_; 
wire u2__abc_52138_new_n7463_; 
wire u2__abc_52138_new_n7464_; 
wire u2__abc_52138_new_n7465_; 
wire u2__abc_52138_new_n7466_; 
wire u2__abc_52138_new_n7467_; 
wire u2__abc_52138_new_n7468_; 
wire u2__abc_52138_new_n7469_; 
wire u2__abc_52138_new_n7471_; 
wire u2__abc_52138_new_n7472_; 
wire u2__abc_52138_new_n7473_; 
wire u2__abc_52138_new_n7474_; 
wire u2__abc_52138_new_n7475_; 
wire u2__abc_52138_new_n7476_; 
wire u2__abc_52138_new_n7477_; 
wire u2__abc_52138_new_n7478_; 
wire u2__abc_52138_new_n7479_; 
wire u2__abc_52138_new_n7480_; 
wire u2__abc_52138_new_n7482_; 
wire u2__abc_52138_new_n7483_; 
wire u2__abc_52138_new_n7484_; 
wire u2__abc_52138_new_n7485_; 
wire u2__abc_52138_new_n7486_; 
wire u2__abc_52138_new_n7487_; 
wire u2__abc_52138_new_n7488_; 
wire u2__abc_52138_new_n7490_; 
wire u2__abc_52138_new_n7491_; 
wire u2__abc_52138_new_n7492_; 
wire u2__abc_52138_new_n7493_; 
wire u2__abc_52138_new_n7494_; 
wire u2__abc_52138_new_n7495_; 
wire u2__abc_52138_new_n7496_; 
wire u2__abc_52138_new_n7497_; 
wire u2__abc_52138_new_n7498_; 
wire u2__abc_52138_new_n7499_; 
wire u2__abc_52138_new_n7500_; 
wire u2__abc_52138_new_n7502_; 
wire u2__abc_52138_new_n7503_; 
wire u2__abc_52138_new_n7504_; 
wire u2__abc_52138_new_n7505_; 
wire u2__abc_52138_new_n7506_; 
wire u2__abc_52138_new_n7507_; 
wire u2__abc_52138_new_n7508_; 
wire u2__abc_52138_new_n7509_; 
wire u2__abc_52138_new_n7511_; 
wire u2__abc_52138_new_n7512_; 
wire u2__abc_52138_new_n7513_; 
wire u2__abc_52138_new_n7514_; 
wire u2__abc_52138_new_n7515_; 
wire u2__abc_52138_new_n7516_; 
wire u2__abc_52138_new_n7517_; 
wire u2__abc_52138_new_n7518_; 
wire u2__abc_52138_new_n7519_; 
wire u2__abc_52138_new_n7521_; 
wire u2__abc_52138_new_n7522_; 
wire u2__abc_52138_new_n7523_; 
wire u2__abc_52138_new_n7524_; 
wire u2__abc_52138_new_n7525_; 
wire u2__abc_52138_new_n7526_; 
wire u2__abc_52138_new_n7527_; 
wire u2__abc_52138_new_n7528_; 
wire u2__abc_52138_new_n7530_; 
wire u2__abc_52138_new_n7531_; 
wire u2__abc_52138_new_n7532_; 
wire u2__abc_52138_new_n7533_; 
wire u2__abc_52138_new_n7534_; 
wire u2__abc_52138_new_n7535_; 
wire u2__abc_52138_new_n7536_; 
wire u2__abc_52138_new_n7537_; 
wire u2__abc_52138_new_n7538_; 
wire u2__abc_52138_new_n7539_; 
wire u2__abc_52138_new_n7540_; 
wire u2__abc_52138_new_n7541_; 
wire u2__abc_52138_new_n7542_; 
wire u2__abc_52138_new_n7543_; 
wire u2__abc_52138_new_n7544_; 
wire u2__abc_52138_new_n7545_; 
wire u2__abc_52138_new_n7546_; 
wire u2__abc_52138_new_n7547_; 
wire u2__abc_52138_new_n7548_; 
wire u2__abc_52138_new_n7550_; 
wire u2__abc_52138_new_n7551_; 
wire u2__abc_52138_new_n7552_; 
wire u2__abc_52138_new_n7553_; 
wire u2__abc_52138_new_n7554_; 
wire u2__abc_52138_new_n7555_; 
wire u2__abc_52138_new_n7556_; 
wire u2__abc_52138_new_n7558_; 
wire u2__abc_52138_new_n7559_; 
wire u2__abc_52138_new_n7560_; 
wire u2__abc_52138_new_n7561_; 
wire u2__abc_52138_new_n7562_; 
wire u2__abc_52138_new_n7563_; 
wire u2__abc_52138_new_n7564_; 
wire u2__abc_52138_new_n7565_; 
wire u2__abc_52138_new_n7566_; 
wire u2__abc_52138_new_n7568_; 
wire u2__abc_52138_new_n7569_; 
wire u2__abc_52138_new_n7570_; 
wire u2__abc_52138_new_n7571_; 
wire u2__abc_52138_new_n7572_; 
wire u2__abc_52138_new_n7573_; 
wire u2__abc_52138_new_n7574_; 
wire u2__abc_52138_new_n7575_; 
wire u2__abc_52138_new_n7576_; 
wire u2__abc_52138_new_n7578_; 
wire u2__abc_52138_new_n7579_; 
wire u2__abc_52138_new_n7580_; 
wire u2__abc_52138_new_n7581_; 
wire u2__abc_52138_new_n7582_; 
wire u2__abc_52138_new_n7583_; 
wire u2__abc_52138_new_n7584_; 
wire u2__abc_52138_new_n7585_; 
wire u2__abc_52138_new_n7586_; 
wire u2__abc_52138_new_n7587_; 
wire u2__abc_52138_new_n7588_; 
wire u2__abc_52138_new_n7589_; 
wire u2__abc_52138_new_n7590_; 
wire u2__abc_52138_new_n7591_; 
wire u2__abc_52138_new_n7592_; 
wire u2__abc_52138_new_n7593_; 
wire u2__abc_52138_new_n7594_; 
wire u2__abc_52138_new_n7596_; 
wire u2__abc_52138_new_n7597_; 
wire u2__abc_52138_new_n7598_; 
wire u2__abc_52138_new_n7599_; 
wire u2__abc_52138_new_n7600_; 
wire u2__abc_52138_new_n7601_; 
wire u2__abc_52138_new_n7602_; 
wire u2__abc_52138_new_n7604_; 
wire u2__abc_52138_new_n7605_; 
wire u2__abc_52138_new_n7606_; 
wire u2__abc_52138_new_n7607_; 
wire u2__abc_52138_new_n7608_; 
wire u2__abc_52138_new_n7609_; 
wire u2__abc_52138_new_n7610_; 
wire u2__abc_52138_new_n7611_; 
wire u2__abc_52138_new_n7612_; 
wire u2__abc_52138_new_n7613_; 
wire u2__abc_52138_new_n7615_; 
wire u2__abc_52138_new_n7616_; 
wire u2__abc_52138_new_n7617_; 
wire u2__abc_52138_new_n7618_; 
wire u2__abc_52138_new_n7619_; 
wire u2__abc_52138_new_n7620_; 
wire u2__abc_52138_new_n7621_; 
wire u2__abc_52138_new_n7622_; 
wire u2__abc_52138_new_n7624_; 
wire u2__abc_52138_new_n7625_; 
wire u2__abc_52138_new_n7626_; 
wire u2__abc_52138_new_n7627_; 
wire u2__abc_52138_new_n7628_; 
wire u2__abc_52138_new_n7629_; 
wire u2__abc_52138_new_n7630_; 
wire u2__abc_52138_new_n7631_; 
wire u2__abc_52138_new_n7632_; 
wire u2__abc_52138_new_n7633_; 
wire u2__abc_52138_new_n7634_; 
wire u2__abc_52138_new_n7635_; 
wire u2__abc_52138_new_n7636_; 
wire u2__abc_52138_new_n7637_; 
wire u2__abc_52138_new_n7638_; 
wire u2__abc_52138_new_n7639_; 
wire u2__abc_52138_new_n7641_; 
wire u2__abc_52138_new_n7642_; 
wire u2__abc_52138_new_n7643_; 
wire u2__abc_52138_new_n7644_; 
wire u2__abc_52138_new_n7645_; 
wire u2__abc_52138_new_n7646_; 
wire u2__abc_52138_new_n7647_; 
wire u2__abc_52138_new_n7648_; 
wire u2__abc_52138_new_n7650_; 
wire u2__abc_52138_new_n7651_; 
wire u2__abc_52138_new_n7652_; 
wire u2__abc_52138_new_n7653_; 
wire u2__abc_52138_new_n7654_; 
wire u2__abc_52138_new_n7655_; 
wire u2__abc_52138_new_n7656_; 
wire u2__abc_52138_new_n7657_; 
wire u2__abc_52138_new_n7658_; 
wire u2__abc_52138_new_n7659_; 
wire u2__abc_52138_new_n7661_; 
wire u2__abc_52138_new_n7662_; 
wire u2__abc_52138_new_n7663_; 
wire u2__abc_52138_new_n7664_; 
wire u2__abc_52138_new_n7665_; 
wire u2__abc_52138_new_n7666_; 
wire u2__abc_52138_new_n7667_; 
wire u2__abc_52138_new_n7669_; 
wire u2__abc_52138_new_n7670_; 
wire u2__abc_52138_new_n7671_; 
wire u2__abc_52138_new_n7672_; 
wire u2__abc_52138_new_n7673_; 
wire u2__abc_52138_new_n7674_; 
wire u2__abc_52138_new_n7675_; 
wire u2__abc_52138_new_n7676_; 
wire u2__abc_52138_new_n7677_; 
wire u2__abc_52138_new_n7678_; 
wire u2__abc_52138_new_n7679_; 
wire u2__abc_52138_new_n7680_; 
wire u2__abc_52138_new_n7681_; 
wire u2__abc_52138_new_n7683_; 
wire u2__abc_52138_new_n7684_; 
wire u2__abc_52138_new_n7685_; 
wire u2__abc_52138_new_n7686_; 
wire u2__abc_52138_new_n7687_; 
wire u2__abc_52138_new_n7688_; 
wire u2__abc_52138_new_n7689_; 
wire u2__abc_52138_new_n7690_; 
wire u2__abc_52138_new_n7692_; 
wire u2__abc_52138_new_n7693_; 
wire u2__abc_52138_new_n7694_; 
wire u2__abc_52138_new_n7695_; 
wire u2__abc_52138_new_n7696_; 
wire u2__abc_52138_new_n7697_; 
wire u2__abc_52138_new_n7698_; 
wire u2__abc_52138_new_n7699_; 
wire u2__abc_52138_new_n7700_; 
wire u2__abc_52138_new_n7702_; 
wire u2__abc_52138_new_n7703_; 
wire u2__abc_52138_new_n7704_; 
wire u2__abc_52138_new_n7705_; 
wire u2__abc_52138_new_n7706_; 
wire u2__abc_52138_new_n7707_; 
wire u2__abc_52138_new_n7708_; 
wire u2__abc_52138_new_n7709_; 
wire u2__abc_52138_new_n7710_; 
wire u2__abc_52138_new_n7711_; 
wire u2__abc_52138_new_n7713_; 
wire u2__abc_52138_new_n7714_; 
wire u2__abc_52138_new_n7715_; 
wire u2__abc_52138_new_n7716_; 
wire u2__abc_52138_new_n7717_; 
wire u2__abc_52138_new_n7718_; 
wire u2__abc_52138_new_n7719_; 
wire u2__abc_52138_new_n7720_; 
wire u2__abc_52138_new_n7721_; 
wire u2__abc_52138_new_n7722_; 
wire u2__abc_52138_new_n7723_; 
wire u2__abc_52138_new_n7724_; 
wire u2__abc_52138_new_n7725_; 
wire u2__abc_52138_new_n7726_; 
wire u2__abc_52138_new_n7728_; 
wire u2__abc_52138_new_n7729_; 
wire u2__abc_52138_new_n7730_; 
wire u2__abc_52138_new_n7731_; 
wire u2__abc_52138_new_n7732_; 
wire u2__abc_52138_new_n7733_; 
wire u2__abc_52138_new_n7734_; 
wire u2__abc_52138_new_n7735_; 
wire u2__abc_52138_new_n7737_; 
wire u2__abc_52138_new_n7738_; 
wire u2__abc_52138_new_n7739_; 
wire u2__abc_52138_new_n7740_; 
wire u2__abc_52138_new_n7741_; 
wire u2__abc_52138_new_n7742_; 
wire u2__abc_52138_new_n7743_; 
wire u2__abc_52138_new_n7744_; 
wire u2__abc_52138_new_n7745_; 
wire u2__abc_52138_new_n7746_; 
wire u2__abc_52138_new_n7748_; 
wire u2__abc_52138_new_n7749_; 
wire u2__abc_52138_new_n7750_; 
wire u2__abc_52138_new_n7751_; 
wire u2__abc_52138_new_n7752_; 
wire u2__abc_52138_new_n7753_; 
wire u2__abc_52138_new_n7754_; 
wire u2__abc_52138_new_n7756_; 
wire u2__abc_52138_new_n7757_; 
wire u2__abc_52138_new_n7758_; 
wire u2__abc_52138_new_n7759_; 
wire u2__abc_52138_new_n7760_; 
wire u2__abc_52138_new_n7761_; 
wire u2__abc_52138_new_n7762_; 
wire u2__abc_52138_new_n7763_; 
wire u2__abc_52138_new_n7764_; 
wire u2__abc_52138_new_n7765_; 
wire u2__abc_52138_new_n7766_; 
wire u2__abc_52138_new_n7767_; 
wire u2__abc_52138_new_n7768_; 
wire u2__abc_52138_new_n7770_; 
wire u2__abc_52138_new_n7771_; 
wire u2__abc_52138_new_n7772_; 
wire u2__abc_52138_new_n7773_; 
wire u2__abc_52138_new_n7774_; 
wire u2__abc_52138_new_n7775_; 
wire u2__abc_52138_new_n7776_; 
wire u2__abc_52138_new_n7777_; 
wire u2__abc_52138_new_n7779_; 
wire u2__abc_52138_new_n7780_; 
wire u2__abc_52138_new_n7781_; 
wire u2__abc_52138_new_n7782_; 
wire u2__abc_52138_new_n7783_; 
wire u2__abc_52138_new_n7784_; 
wire u2__abc_52138_new_n7785_; 
wire u2__abc_52138_new_n7786_; 
wire u2__abc_52138_new_n7787_; 
wire u2__abc_52138_new_n7788_; 
wire u2__abc_52138_new_n7789_; 
wire u2__abc_52138_new_n7791_; 
wire u2__abc_52138_new_n7792_; 
wire u2__abc_52138_new_n7793_; 
wire u2__abc_52138_new_n7794_; 
wire u2__abc_52138_new_n7795_; 
wire u2__abc_52138_new_n7796_; 
wire u2__abc_52138_new_n7797_; 
wire u2__abc_52138_new_n7798_; 
wire u2__abc_52138_new_n7800_; 
wire u2__abc_52138_new_n7801_; 
wire u2__abc_52138_new_n7802_; 
wire u2__abc_52138_new_n7803_; 
wire u2__abc_52138_new_n7804_; 
wire u2__abc_52138_new_n7805_; 
wire u2__abc_52138_new_n7806_; 
wire u2__abc_52138_new_n7807_; 
wire u2__abc_52138_new_n7808_; 
wire u2__abc_52138_new_n7809_; 
wire u2__abc_52138_new_n7810_; 
wire u2__abc_52138_new_n7811_; 
wire u2__abc_52138_new_n7812_; 
wire u2__abc_52138_new_n7813_; 
wire u2__abc_52138_new_n7814_; 
wire u2__abc_52138_new_n7815_; 
wire u2__abc_52138_new_n7816_; 
wire u2__abc_52138_new_n7818_; 
wire u2__abc_52138_new_n7819_; 
wire u2__abc_52138_new_n7820_; 
wire u2__abc_52138_new_n7821_; 
wire u2__abc_52138_new_n7822_; 
wire u2__abc_52138_new_n7823_; 
wire u2__abc_52138_new_n7824_; 
wire u2__abc_52138_new_n7825_; 
wire u2__abc_52138_new_n7827_; 
wire u2__abc_52138_new_n7828_; 
wire u2__abc_52138_new_n7829_; 
wire u2__abc_52138_new_n7830_; 
wire u2__abc_52138_new_n7831_; 
wire u2__abc_52138_new_n7832_; 
wire u2__abc_52138_new_n7833_; 
wire u2__abc_52138_new_n7834_; 
wire u2__abc_52138_new_n7835_; 
wire u2__abc_52138_new_n7836_; 
wire u2__abc_52138_new_n7837_; 
wire u2__abc_52138_new_n7839_; 
wire u2__abc_52138_new_n7840_; 
wire u2__abc_52138_new_n7841_; 
wire u2__abc_52138_new_n7842_; 
wire u2__abc_52138_new_n7843_; 
wire u2__abc_52138_new_n7844_; 
wire u2__abc_52138_new_n7845_; 
wire u2__abc_52138_new_n7846_; 
wire u2__abc_52138_new_n7848_; 
wire u2__abc_52138_new_n7849_; 
wire u2__abc_52138_new_n7850_; 
wire u2__abc_52138_new_n7851_; 
wire u2__abc_52138_new_n7852_; 
wire u2__abc_52138_new_n7853_; 
wire u2__abc_52138_new_n7854_; 
wire u2__abc_52138_new_n7855_; 
wire u2__abc_52138_new_n7856_; 
wire u2__abc_52138_new_n7857_; 
wire u2__abc_52138_new_n7858_; 
wire u2__abc_52138_new_n7859_; 
wire u2__abc_52138_new_n7861_; 
wire u2__abc_52138_new_n7862_; 
wire u2__abc_52138_new_n7863_; 
wire u2__abc_52138_new_n7864_; 
wire u2__abc_52138_new_n7865_; 
wire u2__abc_52138_new_n7866_; 
wire u2__abc_52138_new_n7867_; 
wire u2__abc_52138_new_n7868_; 
wire u2__abc_52138_new_n7870_; 
wire u2__abc_52138_new_n7871_; 
wire u2__abc_52138_new_n7872_; 
wire u2__abc_52138_new_n7873_; 
wire u2__abc_52138_new_n7874_; 
wire u2__abc_52138_new_n7875_; 
wire u2__abc_52138_new_n7876_; 
wire u2__abc_52138_new_n7877_; 
wire u2__abc_52138_new_n7879_; 
wire u2__abc_52138_new_n7880_; 
wire u2__abc_52138_new_n7881_; 
wire u2__abc_52138_new_n7882_; 
wire u2__abc_52138_new_n7883_; 
wire u2__abc_52138_new_n7884_; 
wire u2__abc_52138_new_n7885_; 
wire u2__abc_52138_new_n7887_; 
wire u2__abc_52138_new_n7888_; 
wire u2__abc_52138_new_n7889_; 
wire u2__abc_52138_new_n7890_; 
wire u2__abc_52138_new_n7891_; 
wire u2__abc_52138_new_n7892_; 
wire u2__abc_52138_new_n7893_; 
wire u2__abc_52138_new_n7894_; 
wire u2__abc_52138_new_n7895_; 
wire u2__abc_52138_new_n7896_; 
wire u2__abc_52138_new_n7897_; 
wire u2__abc_52138_new_n7898_; 
wire u2__abc_52138_new_n7899_; 
wire u2__abc_52138_new_n7900_; 
wire u2__abc_52138_new_n7901_; 
wire u2__abc_52138_new_n7902_; 
wire u2__abc_52138_new_n7903_; 
wire u2__abc_52138_new_n7904_; 
wire u2__abc_52138_new_n7905_; 
wire u2__abc_52138_new_n7906_; 
wire u2__abc_52138_new_n7907_; 
wire u2__abc_52138_new_n7909_; 
wire u2__abc_52138_new_n7910_; 
wire u2__abc_52138_new_n7911_; 
wire u2__abc_52138_new_n7912_; 
wire u2__abc_52138_new_n7913_; 
wire u2__abc_52138_new_n7914_; 
wire u2__abc_52138_new_n7915_; 
wire u2__abc_52138_new_n7917_; 
wire u2__abc_52138_new_n7918_; 
wire u2__abc_52138_new_n7919_; 
wire u2__abc_52138_new_n7920_; 
wire u2__abc_52138_new_n7921_; 
wire u2__abc_52138_new_n7922_; 
wire u2__abc_52138_new_n7923_; 
wire u2__abc_52138_new_n7924_; 
wire u2__abc_52138_new_n7925_; 
wire u2__abc_52138_new_n7927_; 
wire u2__abc_52138_new_n7928_; 
wire u2__abc_52138_new_n7929_; 
wire u2__abc_52138_new_n7930_; 
wire u2__abc_52138_new_n7931_; 
wire u2__abc_52138_new_n7932_; 
wire u2__abc_52138_new_n7933_; 
wire u2__abc_52138_new_n7934_; 
wire u2__abc_52138_new_n7935_; 
wire u2__abc_52138_new_n7937_; 
wire u2__abc_52138_new_n7938_; 
wire u2__abc_52138_new_n7939_; 
wire u2__abc_52138_new_n7940_; 
wire u2__abc_52138_new_n7941_; 
wire u2__abc_52138_new_n7942_; 
wire u2__abc_52138_new_n7943_; 
wire u2__abc_52138_new_n7944_; 
wire u2__abc_52138_new_n7945_; 
wire u2__abc_52138_new_n7946_; 
wire u2__abc_52138_new_n7947_; 
wire u2__abc_52138_new_n7948_; 
wire u2__abc_52138_new_n7949_; 
wire u2__abc_52138_new_n7950_; 
wire u2__abc_52138_new_n7951_; 
wire u2__abc_52138_new_n7953_; 
wire u2__abc_52138_new_n7954_; 
wire u2__abc_52138_new_n7955_; 
wire u2__abc_52138_new_n7956_; 
wire u2__abc_52138_new_n7957_; 
wire u2__abc_52138_new_n7958_; 
wire u2__abc_52138_new_n7959_; 
wire u2__abc_52138_new_n7961_; 
wire u2__abc_52138_new_n7962_; 
wire u2__abc_52138_new_n7963_; 
wire u2__abc_52138_new_n7964_; 
wire u2__abc_52138_new_n7965_; 
wire u2__abc_52138_new_n7966_; 
wire u2__abc_52138_new_n7967_; 
wire u2__abc_52138_new_n7968_; 
wire u2__abc_52138_new_n7969_; 
wire u2__abc_52138_new_n7970_; 
wire u2__abc_52138_new_n7972_; 
wire u2__abc_52138_new_n7973_; 
wire u2__abc_52138_new_n7974_; 
wire u2__abc_52138_new_n7975_; 
wire u2__abc_52138_new_n7976_; 
wire u2__abc_52138_new_n7977_; 
wire u2__abc_52138_new_n7978_; 
wire u2__abc_52138_new_n7980_; 
wire u2__abc_52138_new_n7981_; 
wire u2__abc_52138_new_n7982_; 
wire u2__abc_52138_new_n7983_; 
wire u2__abc_52138_new_n7984_; 
wire u2__abc_52138_new_n7985_; 
wire u2__abc_52138_new_n7986_; 
wire u2__abc_52138_new_n7987_; 
wire u2__abc_52138_new_n7988_; 
wire u2__abc_52138_new_n7989_; 
wire u2__abc_52138_new_n7990_; 
wire u2__abc_52138_new_n7991_; 
wire u2__abc_52138_new_n7992_; 
wire u2__abc_52138_new_n7993_; 
wire u2__abc_52138_new_n7994_; 
wire u2__abc_52138_new_n7995_; 
wire u2__abc_52138_new_n7996_; 
wire u2__abc_52138_new_n7998_; 
wire u2__abc_52138_new_n7999_; 
wire u2__abc_52138_new_n8000_; 
wire u2__abc_52138_new_n8001_; 
wire u2__abc_52138_new_n8002_; 
wire u2__abc_52138_new_n8003_; 
wire u2__abc_52138_new_n8004_; 
wire u2__abc_52138_new_n8006_; 
wire u2__abc_52138_new_n8007_; 
wire u2__abc_52138_new_n8008_; 
wire u2__abc_52138_new_n8009_; 
wire u2__abc_52138_new_n8010_; 
wire u2__abc_52138_new_n8011_; 
wire u2__abc_52138_new_n8012_; 
wire u2__abc_52138_new_n8013_; 
wire u2__abc_52138_new_n8014_; 
wire u2__abc_52138_new_n8015_; 
wire u2__abc_52138_new_n8016_; 
wire u2__abc_52138_new_n8017_; 
wire u2__abc_52138_new_n8019_; 
wire u2__abc_52138_new_n8020_; 
wire u2__abc_52138_new_n8021_; 
wire u2__abc_52138_new_n8022_; 
wire u2__abc_52138_new_n8023_; 
wire u2__abc_52138_new_n8024_; 
wire u2__abc_52138_new_n8025_; 
wire u2__abc_52138_new_n8026_; 
wire u2__abc_52138_new_n8027_; 
wire u2__abc_52138_new_n8029_; 
wire u2__abc_52138_new_n8030_; 
wire u2__abc_52138_new_n8031_; 
wire u2__abc_52138_new_n8032_; 
wire u2__abc_52138_new_n8033_; 
wire u2__abc_52138_new_n8034_; 
wire u2__abc_52138_new_n8035_; 
wire u2__abc_52138_new_n8036_; 
wire u2__abc_52138_new_n8037_; 
wire u2__abc_52138_new_n8038_; 
wire u2__abc_52138_new_n8039_; 
wire u2__abc_52138_new_n8040_; 
wire u2__abc_52138_new_n8041_; 
wire u2__abc_52138_new_n8043_; 
wire u2__abc_52138_new_n8044_; 
wire u2__abc_52138_new_n8045_; 
wire u2__abc_52138_new_n8046_; 
wire u2__abc_52138_new_n8047_; 
wire u2__abc_52138_new_n8048_; 
wire u2__abc_52138_new_n8049_; 
wire u2__abc_52138_new_n8051_; 
wire u2__abc_52138_new_n8052_; 
wire u2__abc_52138_new_n8053_; 
wire u2__abc_52138_new_n8054_; 
wire u2__abc_52138_new_n8055_; 
wire u2__abc_52138_new_n8056_; 
wire u2__abc_52138_new_n8057_; 
wire u2__abc_52138_new_n8058_; 
wire u2__abc_52138_new_n8060_; 
wire u2__abc_52138_new_n8061_; 
wire u2__abc_52138_new_n8062_; 
wire u2__abc_52138_new_n8063_; 
wire u2__abc_52138_new_n8064_; 
wire u2__abc_52138_new_n8065_; 
wire u2__abc_52138_new_n8066_; 
wire u2__abc_52138_new_n8068_; 
wire u2__abc_52138_new_n8069_; 
wire u2__abc_52138_new_n8070_; 
wire u2__abc_52138_new_n8071_; 
wire u2__abc_52138_new_n8072_; 
wire u2__abc_52138_new_n8073_; 
wire u2__abc_52138_new_n8074_; 
wire u2__abc_52138_new_n8075_; 
wire u2__abc_52138_new_n8076_; 
wire u2__abc_52138_new_n8077_; 
wire u2__abc_52138_new_n8078_; 
wire u2__abc_52138_new_n8079_; 
wire u2__abc_52138_new_n8080_; 
wire u2__abc_52138_new_n8081_; 
wire u2__abc_52138_new_n8082_; 
wire u2__abc_52138_new_n8083_; 
wire u2__abc_52138_new_n8084_; 
wire u2__abc_52138_new_n8085_; 
wire u2__abc_52138_new_n8086_; 
wire u2__abc_52138_new_n8087_; 
wire u2__abc_52138_new_n8088_; 
wire u2__abc_52138_new_n8089_; 
wire u2__abc_52138_new_n8091_; 
wire u2__abc_52138_new_n8092_; 
wire u2__abc_52138_new_n8093_; 
wire u2__abc_52138_new_n8094_; 
wire u2__abc_52138_new_n8095_; 
wire u2__abc_52138_new_n8096_; 
wire u2__abc_52138_new_n8097_; 
wire u2__abc_52138_new_n8098_; 
wire u2__abc_52138_new_n8100_; 
wire u2__abc_52138_new_n8101_; 
wire u2__abc_52138_new_n8102_; 
wire u2__abc_52138_new_n8103_; 
wire u2__abc_52138_new_n8104_; 
wire u2__abc_52138_new_n8105_; 
wire u2__abc_52138_new_n8106_; 
wire u2__abc_52138_new_n8107_; 
wire u2__abc_52138_new_n8108_; 
wire u2__abc_52138_new_n8109_; 
wire u2__abc_52138_new_n8111_; 
wire u2__abc_52138_new_n8112_; 
wire u2__abc_52138_new_n8113_; 
wire u2__abc_52138_new_n8114_; 
wire u2__abc_52138_new_n8115_; 
wire u2__abc_52138_new_n8116_; 
wire u2__abc_52138_new_n8117_; 
wire u2__abc_52138_new_n8118_; 
wire u2__abc_52138_new_n8120_; 
wire u2__abc_52138_new_n8121_; 
wire u2__abc_52138_new_n8122_; 
wire u2__abc_52138_new_n8123_; 
wire u2__abc_52138_new_n8124_; 
wire u2__abc_52138_new_n8125_; 
wire u2__abc_52138_new_n8126_; 
wire u2__abc_52138_new_n8127_; 
wire u2__abc_52138_new_n8128_; 
wire u2__abc_52138_new_n8129_; 
wire u2__abc_52138_new_n8131_; 
wire u2__abc_52138_new_n8132_; 
wire u2__abc_52138_new_n8133_; 
wire u2__abc_52138_new_n8134_; 
wire u2__abc_52138_new_n8135_; 
wire u2__abc_52138_new_n8136_; 
wire u2__abc_52138_new_n8137_; 
wire u2__abc_52138_new_n8138_; 
wire u2__abc_52138_new_n8140_; 
wire u2__abc_52138_new_n8141_; 
wire u2__abc_52138_new_n8142_; 
wire u2__abc_52138_new_n8143_; 
wire u2__abc_52138_new_n8144_; 
wire u2__abc_52138_new_n8145_; 
wire u2__abc_52138_new_n8146_; 
wire u2__abc_52138_new_n8147_; 
wire u2__abc_52138_new_n8148_; 
wire u2__abc_52138_new_n8149_; 
wire u2__abc_52138_new_n8150_; 
wire u2__abc_52138_new_n8151_; 
wire u2__abc_52138_new_n8153_; 
wire u2__abc_52138_new_n8154_; 
wire u2__abc_52138_new_n8155_; 
wire u2__abc_52138_new_n8156_; 
wire u2__abc_52138_new_n8157_; 
wire u2__abc_52138_new_n8158_; 
wire u2__abc_52138_new_n8159_; 
wire u2__abc_52138_new_n8161_; 
wire u2__abc_52138_new_n8162_; 
wire u2__abc_52138_new_n8163_; 
wire u2__abc_52138_new_n8164_; 
wire u2__abc_52138_new_n8165_; 
wire u2__abc_52138_new_n8166_; 
wire u2__abc_52138_new_n8167_; 
wire u2__abc_52138_new_n8168_; 
wire u2__abc_52138_new_n8169_; 
wire u2__abc_52138_new_n8170_; 
wire u2__abc_52138_new_n8171_; 
wire u2__abc_52138_new_n8172_; 
wire u2__abc_52138_new_n8173_; 
wire u2__abc_52138_new_n8174_; 
wire u2__abc_52138_new_n8175_; 
wire u2__abc_52138_new_n8176_; 
wire u2__abc_52138_new_n8177_; 
wire u2__abc_52138_new_n8178_; 
wire u2__abc_52138_new_n8180_; 
wire u2__abc_52138_new_n8181_; 
wire u2__abc_52138_new_n8182_; 
wire u2__abc_52138_new_n8183_; 
wire u2__abc_52138_new_n8184_; 
wire u2__abc_52138_new_n8185_; 
wire u2__abc_52138_new_n8186_; 
wire u2__abc_52138_new_n8188_; 
wire u2__abc_52138_new_n8189_; 
wire u2__abc_52138_new_n8190_; 
wire u2__abc_52138_new_n8191_; 
wire u2__abc_52138_new_n8192_; 
wire u2__abc_52138_new_n8193_; 
wire u2__abc_52138_new_n8194_; 
wire u2__abc_52138_new_n8195_; 
wire u2__abc_52138_new_n8196_; 
wire u2__abc_52138_new_n8198_; 
wire u2__abc_52138_new_n8199_; 
wire u2__abc_52138_new_n8200_; 
wire u2__abc_52138_new_n8201_; 
wire u2__abc_52138_new_n8202_; 
wire u2__abc_52138_new_n8203_; 
wire u2__abc_52138_new_n8204_; 
wire u2__abc_52138_new_n8206_; 
wire u2__abc_52138_new_n8207_; 
wire u2__abc_52138_new_n8208_; 
wire u2__abc_52138_new_n8209_; 
wire u2__abc_52138_new_n8210_; 
wire u2__abc_52138_new_n8211_; 
wire u2__abc_52138_new_n8212_; 
wire u2__abc_52138_new_n8213_; 
wire u2__abc_52138_new_n8214_; 
wire u2__abc_52138_new_n8215_; 
wire u2__abc_52138_new_n8216_; 
wire u2__abc_52138_new_n8217_; 
wire u2__abc_52138_new_n8218_; 
wire u2__abc_52138_new_n8220_; 
wire u2__abc_52138_new_n8221_; 
wire u2__abc_52138_new_n8222_; 
wire u2__abc_52138_new_n8223_; 
wire u2__abc_52138_new_n8224_; 
wire u2__abc_52138_new_n8225_; 
wire u2__abc_52138_new_n8226_; 
wire u2__abc_52138_new_n8228_; 
wire u2__abc_52138_new_n8229_; 
wire u2__abc_52138_new_n8230_; 
wire u2__abc_52138_new_n8231_; 
wire u2__abc_52138_new_n8232_; 
wire u2__abc_52138_new_n8233_; 
wire u2__abc_52138_new_n8234_; 
wire u2__abc_52138_new_n8235_; 
wire u2__abc_52138_new_n8236_; 
wire u2__abc_52138_new_n8238_; 
wire u2__abc_52138_new_n8239_; 
wire u2__abc_52138_new_n8240_; 
wire u2__abc_52138_new_n8241_; 
wire u2__abc_52138_new_n8242_; 
wire u2__abc_52138_new_n8243_; 
wire u2__abc_52138_new_n8244_; 
wire u2__abc_52138_new_n8245_; 
wire u2__abc_52138_new_n8247_; 
wire u2__abc_52138_new_n8248_; 
wire u2__abc_52138_new_n8249_; 
wire u2__abc_52138_new_n8250_; 
wire u2__abc_52138_new_n8251_; 
wire u2__abc_52138_new_n8252_; 
wire u2__abc_52138_new_n8253_; 
wire u2__abc_52138_new_n8254_; 
wire u2__abc_52138_new_n8255_; 
wire u2__abc_52138_new_n8256_; 
wire u2__abc_52138_new_n8257_; 
wire u2__abc_52138_new_n8258_; 
wire u2__abc_52138_new_n8259_; 
wire u2__abc_52138_new_n8260_; 
wire u2__abc_52138_new_n8261_; 
wire u2__abc_52138_new_n8262_; 
wire u2__abc_52138_new_n8263_; 
wire u2__abc_52138_new_n8264_; 
wire u2__abc_52138_new_n8265_; 
wire u2__abc_52138_new_n8267_; 
wire u2__abc_52138_new_n8268_; 
wire u2__abc_52138_new_n8269_; 
wire u2__abc_52138_new_n8270_; 
wire u2__abc_52138_new_n8271_; 
wire u2__abc_52138_new_n8272_; 
wire u2__abc_52138_new_n8273_; 
wire u2__abc_52138_new_n8275_; 
wire u2__abc_52138_new_n8276_; 
wire u2__abc_52138_new_n8277_; 
wire u2__abc_52138_new_n8278_; 
wire u2__abc_52138_new_n8279_; 
wire u2__abc_52138_new_n8280_; 
wire u2__abc_52138_new_n8281_; 
wire u2__abc_52138_new_n8282_; 
wire u2__abc_52138_new_n8283_; 
wire u2__abc_52138_new_n8284_; 
wire u2__abc_52138_new_n8285_; 
wire u2__abc_52138_new_n8286_; 
wire u2__abc_52138_new_n8288_; 
wire u2__abc_52138_new_n8289_; 
wire u2__abc_52138_new_n8290_; 
wire u2__abc_52138_new_n8291_; 
wire u2__abc_52138_new_n8292_; 
wire u2__abc_52138_new_n8293_; 
wire u2__abc_52138_new_n8294_; 
wire u2__abc_52138_new_n8295_; 
wire u2__abc_52138_new_n8296_; 
wire u2__abc_52138_new_n8298_; 
wire u2__abc_52138_new_n8299_; 
wire u2__abc_52138_new_n8300_; 
wire u2__abc_52138_new_n8301_; 
wire u2__abc_52138_new_n8302_; 
wire u2__abc_52138_new_n8303_; 
wire u2__abc_52138_new_n8304_; 
wire u2__abc_52138_new_n8305_; 
wire u2__abc_52138_new_n8306_; 
wire u2__abc_52138_new_n8307_; 
wire u2__abc_52138_new_n8308_; 
wire u2__abc_52138_new_n8309_; 
wire u2__abc_52138_new_n8311_; 
wire u2__abc_52138_new_n8312_; 
wire u2__abc_52138_new_n8313_; 
wire u2__abc_52138_new_n8314_; 
wire u2__abc_52138_new_n8315_; 
wire u2__abc_52138_new_n8316_; 
wire u2__abc_52138_new_n8317_; 
wire u2__abc_52138_new_n8318_; 
wire u2__abc_52138_new_n8320_; 
wire u2__abc_52138_new_n8321_; 
wire u2__abc_52138_new_n8322_; 
wire u2__abc_52138_new_n8323_; 
wire u2__abc_52138_new_n8324_; 
wire u2__abc_52138_new_n8325_; 
wire u2__abc_52138_new_n8326_; 
wire u2__abc_52138_new_n8327_; 
wire u2__abc_52138_new_n8328_; 
wire u2__abc_52138_new_n8330_; 
wire u2__abc_52138_new_n8331_; 
wire u2__abc_52138_new_n8332_; 
wire u2__abc_52138_new_n8333_; 
wire u2__abc_52138_new_n8334_; 
wire u2__abc_52138_new_n8335_; 
wire u2__abc_52138_new_n8336_; 
wire u2__abc_52138_new_n8337_; 
wire u2__abc_52138_new_n8339_; 
wire u2__abc_52138_new_n8340_; 
wire u2__abc_52138_new_n8341_; 
wire u2__abc_52138_new_n8342_; 
wire u2__abc_52138_new_n8343_; 
wire u2__abc_52138_new_n8344_; 
wire u2__abc_52138_new_n8345_; 
wire u2__abc_52138_new_n8346_; 
wire u2__abc_52138_new_n8347_; 
wire u2__abc_52138_new_n8348_; 
wire u2__abc_52138_new_n8349_; 
wire u2__abc_52138_new_n8350_; 
wire u2__abc_52138_new_n8351_; 
wire u2__abc_52138_new_n8352_; 
wire u2__abc_52138_new_n8354_; 
wire u2__abc_52138_new_n8355_; 
wire u2__abc_52138_new_n8356_; 
wire u2__abc_52138_new_n8357_; 
wire u2__abc_52138_new_n8358_; 
wire u2__abc_52138_new_n8359_; 
wire u2__abc_52138_new_n8360_; 
wire u2__abc_52138_new_n8362_; 
wire u2__abc_52138_new_n8363_; 
wire u2__abc_52138_new_n8364_; 
wire u2__abc_52138_new_n8365_; 
wire u2__abc_52138_new_n8366_; 
wire u2__abc_52138_new_n8367_; 
wire u2__abc_52138_new_n8368_; 
wire u2__abc_52138_new_n8369_; 
wire u2__abc_52138_new_n8370_; 
wire u2__abc_52138_new_n8371_; 
wire u2__abc_52138_new_n8373_; 
wire u2__abc_52138_new_n8374_; 
wire u2__abc_52138_new_n8375_; 
wire u2__abc_52138_new_n8376_; 
wire u2__abc_52138_new_n8377_; 
wire u2__abc_52138_new_n8378_; 
wire u2__abc_52138_new_n8379_; 
wire u2__abc_52138_new_n8381_; 
wire u2__abc_52138_new_n8382_; 
wire u2__abc_52138_new_n8383_; 
wire u2__abc_52138_new_n8384_; 
wire u2__abc_52138_new_n8385_; 
wire u2__abc_52138_new_n8386_; 
wire u2__abc_52138_new_n8387_; 
wire u2__abc_52138_new_n8388_; 
wire u2__abc_52138_new_n8389_; 
wire u2__abc_52138_new_n8390_; 
wire u2__abc_52138_new_n8392_; 
wire u2__abc_52138_new_n8393_; 
wire u2__abc_52138_new_n8394_; 
wire u2__abc_52138_new_n8395_; 
wire u2__abc_52138_new_n8396_; 
wire u2__abc_52138_new_n8397_; 
wire u2__abc_52138_new_n8398_; 
wire u2__abc_52138_new_n8400_; 
wire u2__abc_52138_new_n8401_; 
wire u2__abc_52138_new_n8402_; 
wire u2__abc_52138_new_n8403_; 
wire u2__abc_52138_new_n8404_; 
wire u2__abc_52138_new_n8405_; 
wire u2__abc_52138_new_n8406_; 
wire u2__abc_52138_new_n8407_; 
wire u2__abc_52138_new_n8409_; 
wire u2__abc_52138_new_n8410_; 
wire u2__abc_52138_new_n8411_; 
wire u2__abc_52138_new_n8412_; 
wire u2__abc_52138_new_n8413_; 
wire u2__abc_52138_new_n8414_; 
wire u2__abc_52138_new_n8415_; 
wire u2__abc_52138_new_n8417_; 
wire u2__abc_52138_new_n8418_; 
wire u2__abc_52138_new_n8419_; 
wire u2__abc_52138_new_n8420_; 
wire u2__abc_52138_new_n8421_; 
wire u2__abc_52138_new_n8422_; 
wire u2__abc_52138_new_n8423_; 
wire u2__abc_52138_new_n8424_; 
wire u2__abc_52138_new_n8425_; 
wire u2__abc_52138_new_n8426_; 
wire u2__abc_52138_new_n8427_; 
wire u2__abc_52138_new_n8428_; 
wire u2__abc_52138_new_n8429_; 
wire u2__abc_52138_new_n8430_; 
wire u2__abc_52138_new_n8431_; 
wire u2__abc_52138_new_n8432_; 
wire u2__abc_52138_new_n8433_; 
wire u2__abc_52138_new_n8434_; 
wire u2__abc_52138_new_n8435_; 
wire u2__abc_52138_new_n8436_; 
wire u2__abc_52138_new_n8437_; 
wire u2__abc_52138_new_n8439_; 
wire u2__abc_52138_new_n8440_; 
wire u2__abc_52138_new_n8441_; 
wire u2__abc_52138_new_n8442_; 
wire u2__abc_52138_new_n8443_; 
wire u2__abc_52138_new_n8444_; 
wire u2__abc_52138_new_n8445_; 
wire u2__abc_52138_new_n8447_; 
wire u2__abc_52138_new_n8448_; 
wire u2__abc_52138_new_n8449_; 
wire u2__abc_52138_new_n8450_; 
wire u2__abc_52138_new_n8451_; 
wire u2__abc_52138_new_n8452_; 
wire u2__abc_52138_new_n8453_; 
wire u2__abc_52138_new_n8454_; 
wire u2__abc_52138_new_n8455_; 
wire u2__abc_52138_new_n8456_; 
wire u2__abc_52138_new_n8457_; 
wire u2__abc_52138_new_n8458_; 
wire u2__abc_52138_new_n8459_; 
wire u2__abc_52138_new_n8460_; 
wire u2__abc_52138_new_n8462_; 
wire u2__abc_52138_new_n8463_; 
wire u2__abc_52138_new_n8464_; 
wire u2__abc_52138_new_n8465_; 
wire u2__abc_52138_new_n8466_; 
wire u2__abc_52138_new_n8467_; 
wire u2__abc_52138_new_n8468_; 
wire u2__abc_52138_new_n8470_; 
wire u2__abc_52138_new_n8471_; 
wire u2__abc_52138_new_n8472_; 
wire u2__abc_52138_new_n8473_; 
wire u2__abc_52138_new_n8474_; 
wire u2__abc_52138_new_n8475_; 
wire u2__abc_52138_new_n8476_; 
wire u2__abc_52138_new_n8477_; 
wire u2__abc_52138_new_n8478_; 
wire u2__abc_52138_new_n8479_; 
wire u2__abc_52138_new_n8480_; 
wire u2__abc_52138_new_n8481_; 
wire u2__abc_52138_new_n8483_; 
wire u2__abc_52138_new_n8484_; 
wire u2__abc_52138_new_n8485_; 
wire u2__abc_52138_new_n8486_; 
wire u2__abc_52138_new_n8487_; 
wire u2__abc_52138_new_n8488_; 
wire u2__abc_52138_new_n8489_; 
wire u2__abc_52138_new_n8491_; 
wire u2__abc_52138_new_n8492_; 
wire u2__abc_52138_new_n8493_; 
wire u2__abc_52138_new_n8494_; 
wire u2__abc_52138_new_n8495_; 
wire u2__abc_52138_new_n8496_; 
wire u2__abc_52138_new_n8497_; 
wire u2__abc_52138_new_n8498_; 
wire u2__abc_52138_new_n8500_; 
wire u2__abc_52138_new_n8501_; 
wire u2__abc_52138_new_n8502_; 
wire u2__abc_52138_new_n8503_; 
wire u2__abc_52138_new_n8504_; 
wire u2__abc_52138_new_n8505_; 
wire u2__abc_52138_new_n8506_; 
wire u2__abc_52138_new_n8508_; 
wire u2__abc_52138_new_n8509_; 
wire u2__abc_52138_new_n8510_; 
wire u2__abc_52138_new_n8511_; 
wire u2__abc_52138_new_n8512_; 
wire u2__abc_52138_new_n8513_; 
wire u2__abc_52138_new_n8514_; 
wire u2__abc_52138_new_n8515_; 
wire u2__abc_52138_new_n8516_; 
wire u2__abc_52138_new_n8517_; 
wire u2__abc_52138_new_n8518_; 
wire u2__abc_52138_new_n8519_; 
wire u2__abc_52138_new_n8520_; 
wire u2__abc_52138_new_n8522_; 
wire u2__abc_52138_new_n8523_; 
wire u2__abc_52138_new_n8524_; 
wire u2__abc_52138_new_n8525_; 
wire u2__abc_52138_new_n8526_; 
wire u2__abc_52138_new_n8527_; 
wire u2__abc_52138_new_n8528_; 
wire u2__abc_52138_new_n8529_; 
wire u2__abc_52138_new_n8531_; 
wire u2__abc_52138_new_n8532_; 
wire u2__abc_52138_new_n8533_; 
wire u2__abc_52138_new_n8534_; 
wire u2__abc_52138_new_n8535_; 
wire u2__abc_52138_new_n8536_; 
wire u2__abc_52138_new_n8537_; 
wire u2__abc_52138_new_n8538_; 
wire u2__abc_52138_new_n8539_; 
wire u2__abc_52138_new_n8540_; 
wire u2__abc_52138_new_n8542_; 
wire u2__abc_52138_new_n8543_; 
wire u2__abc_52138_new_n8544_; 
wire u2__abc_52138_new_n8545_; 
wire u2__abc_52138_new_n8546_; 
wire u2__abc_52138_new_n8547_; 
wire u2__abc_52138_new_n8548_; 
wire u2__abc_52138_new_n8549_; 
wire u2__abc_52138_new_n8551_; 
wire u2__abc_52138_new_n8552_; 
wire u2__abc_52138_new_n8553_; 
wire u2__abc_52138_new_n8554_; 
wire u2__abc_52138_new_n8555_; 
wire u2__abc_52138_new_n8556_; 
wire u2__abc_52138_new_n8557_; 
wire u2__abc_52138_new_n8558_; 
wire u2__abc_52138_new_n8559_; 
wire u2__abc_52138_new_n8560_; 
wire u2__abc_52138_new_n8561_; 
wire u2__abc_52138_new_n8562_; 
wire u2__abc_52138_new_n8564_; 
wire u2__abc_52138_new_n8565_; 
wire u2__abc_52138_new_n8566_; 
wire u2__abc_52138_new_n8567_; 
wire u2__abc_52138_new_n8568_; 
wire u2__abc_52138_new_n8569_; 
wire u2__abc_52138_new_n8570_; 
wire u2__abc_52138_new_n8572_; 
wire u2__abc_52138_new_n8573_; 
wire u2__abc_52138_new_n8574_; 
wire u2__abc_52138_new_n8575_; 
wire u2__abc_52138_new_n8576_; 
wire u2__abc_52138_new_n8577_; 
wire u2__abc_52138_new_n8578_; 
wire u2__abc_52138_new_n8579_; 
wire u2__abc_52138_new_n8581_; 
wire u2__abc_52138_new_n8582_; 
wire u2__abc_52138_new_n8583_; 
wire u2__abc_52138_new_n8584_; 
wire u2__abc_52138_new_n8585_; 
wire u2__abc_52138_new_n8586_; 
wire u2__abc_52138_new_n8587_; 
wire u2__abc_52138_new_n8589_; 
wire u2__abc_52138_new_n8590_; 
wire u2__abc_52138_new_n8591_; 
wire u2__abc_52138_new_n8592_; 
wire u2__abc_52138_new_n8593_; 
wire u2__abc_52138_new_n8594_; 
wire u2__abc_52138_new_n8595_; 
wire u2__abc_52138_new_n8596_; 
wire u2__abc_52138_new_n8597_; 
wire u2__abc_52138_new_n8598_; 
wire u2__abc_52138_new_n8599_; 
wire u2__abc_52138_new_n8600_; 
wire u2__abc_52138_new_n8601_; 
wire u2__abc_52138_new_n8602_; 
wire u2__abc_52138_new_n8603_; 
wire u2__abc_52138_new_n8604_; 
wire u2__abc_52138_new_n8605_; 
wire u2__abc_52138_new_n8606_; 
wire u2__abc_52138_new_n8607_; 
wire u2__abc_52138_new_n8608_; 
wire u2__abc_52138_new_n8609_; 
wire u2__abc_52138_new_n8610_; 
wire u2__abc_52138_new_n8611_; 
wire u2__abc_52138_new_n8612_; 
wire u2__abc_52138_new_n8614_; 
wire u2__abc_52138_new_n8615_; 
wire u2__abc_52138_new_n8616_; 
wire u2__abc_52138_new_n8617_; 
wire u2__abc_52138_new_n8618_; 
wire u2__abc_52138_new_n8619_; 
wire u2__abc_52138_new_n8620_; 
wire u2__abc_52138_new_n8622_; 
wire u2__abc_52138_new_n8623_; 
wire u2__abc_52138_new_n8624_; 
wire u2__abc_52138_new_n8625_; 
wire u2__abc_52138_new_n8626_; 
wire u2__abc_52138_new_n8627_; 
wire u2__abc_52138_new_n8628_; 
wire u2__abc_52138_new_n8629_; 
wire u2__abc_52138_new_n8630_; 
wire u2__abc_52138_new_n8632_; 
wire u2__abc_52138_new_n8633_; 
wire u2__abc_52138_new_n8634_; 
wire u2__abc_52138_new_n8635_; 
wire u2__abc_52138_new_n8636_; 
wire u2__abc_52138_new_n8637_; 
wire u2__abc_52138_new_n8638_; 
wire u2__abc_52138_new_n8640_; 
wire u2__abc_52138_new_n8641_; 
wire u2__abc_52138_new_n8642_; 
wire u2__abc_52138_new_n8643_; 
wire u2__abc_52138_new_n8644_; 
wire u2__abc_52138_new_n8645_; 
wire u2__abc_52138_new_n8646_; 
wire u2__abc_52138_new_n8647_; 
wire u2__abc_52138_new_n8648_; 
wire u2__abc_52138_new_n8649_; 
wire u2__abc_52138_new_n8650_; 
wire u2__abc_52138_new_n8651_; 
wire u2__abc_52138_new_n8653_; 
wire u2__abc_52138_new_n8654_; 
wire u2__abc_52138_new_n8655_; 
wire u2__abc_52138_new_n8656_; 
wire u2__abc_52138_new_n8657_; 
wire u2__abc_52138_new_n8658_; 
wire u2__abc_52138_new_n8659_; 
wire u2__abc_52138_new_n8660_; 
wire u2__abc_52138_new_n8662_; 
wire u2__abc_52138_new_n8663_; 
wire u2__abc_52138_new_n8664_; 
wire u2__abc_52138_new_n8665_; 
wire u2__abc_52138_new_n8666_; 
wire u2__abc_52138_new_n8667_; 
wire u2__abc_52138_new_n8668_; 
wire u2__abc_52138_new_n8669_; 
wire u2__abc_52138_new_n8670_; 
wire u2__abc_52138_new_n8671_; 
wire u2__abc_52138_new_n8672_; 
wire u2__abc_52138_new_n8673_; 
wire u2__abc_52138_new_n8674_; 
wire u2__abc_52138_new_n8676_; 
wire u2__abc_52138_new_n8677_; 
wire u2__abc_52138_new_n8678_; 
wire u2__abc_52138_new_n8679_; 
wire u2__abc_52138_new_n8680_; 
wire u2__abc_52138_new_n8681_; 
wire u2__abc_52138_new_n8682_; 
wire u2__abc_52138_new_n8684_; 
wire u2__abc_52138_new_n8685_; 
wire u2__abc_52138_new_n8686_; 
wire u2__abc_52138_new_n8687_; 
wire u2__abc_52138_new_n8688_; 
wire u2__abc_52138_new_n8689_; 
wire u2__abc_52138_new_n8690_; 
wire u2__abc_52138_new_n8691_; 
wire u2__abc_52138_new_n8692_; 
wire u2__abc_52138_new_n8693_; 
wire u2__abc_52138_new_n8694_; 
wire u2__abc_52138_new_n8695_; 
wire u2__abc_52138_new_n8696_; 
wire u2__abc_52138_new_n8697_; 
wire u2__abc_52138_new_n8698_; 
wire u2__abc_52138_new_n8700_; 
wire u2__abc_52138_new_n8701_; 
wire u2__abc_52138_new_n8702_; 
wire u2__abc_52138_new_n8703_; 
wire u2__abc_52138_new_n8704_; 
wire u2__abc_52138_new_n8705_; 
wire u2__abc_52138_new_n8706_; 
wire u2__abc_52138_new_n8708_; 
wire u2__abc_52138_new_n8709_; 
wire u2__abc_52138_new_n8710_; 
wire u2__abc_52138_new_n8711_; 
wire u2__abc_52138_new_n8712_; 
wire u2__abc_52138_new_n8713_; 
wire u2__abc_52138_new_n8714_; 
wire u2__abc_52138_new_n8715_; 
wire u2__abc_52138_new_n8716_; 
wire u2__abc_52138_new_n8718_; 
wire u2__abc_52138_new_n8719_; 
wire u2__abc_52138_new_n8720_; 
wire u2__abc_52138_new_n8721_; 
wire u2__abc_52138_new_n8722_; 
wire u2__abc_52138_new_n8723_; 
wire u2__abc_52138_new_n8724_; 
wire u2__abc_52138_new_n8726_; 
wire u2__abc_52138_new_n8727_; 
wire u2__abc_52138_new_n8728_; 
wire u2__abc_52138_new_n8729_; 
wire u2__abc_52138_new_n8730_; 
wire u2__abc_52138_new_n8731_; 
wire u2__abc_52138_new_n8732_; 
wire u2__abc_52138_new_n8733_; 
wire u2__abc_52138_new_n8734_; 
wire u2__abc_52138_new_n8735_; 
wire u2__abc_52138_new_n8736_; 
wire u2__abc_52138_new_n8737_; 
wire u2__abc_52138_new_n8738_; 
wire u2__abc_52138_new_n8740_; 
wire u2__abc_52138_new_n8741_; 
wire u2__abc_52138_new_n8742_; 
wire u2__abc_52138_new_n8743_; 
wire u2__abc_52138_new_n8744_; 
wire u2__abc_52138_new_n8745_; 
wire u2__abc_52138_new_n8746_; 
wire u2__abc_52138_new_n8748_; 
wire u2__abc_52138_new_n8749_; 
wire u2__abc_52138_new_n8750_; 
wire u2__abc_52138_new_n8751_; 
wire u2__abc_52138_new_n8752_; 
wire u2__abc_52138_new_n8753_; 
wire u2__abc_52138_new_n8754_; 
wire u2__abc_52138_new_n8755_; 
wire u2__abc_52138_new_n8756_; 
wire u2__abc_52138_new_n8758_; 
wire u2__abc_52138_new_n8759_; 
wire u2__abc_52138_new_n8760_; 
wire u2__abc_52138_new_n8761_; 
wire u2__abc_52138_new_n8762_; 
wire u2__abc_52138_new_n8763_; 
wire u2__abc_52138_new_n8764_; 
wire u2__abc_52138_new_n8766_; 
wire u2__abc_52138_new_n8767_; 
wire u2__abc_52138_new_n8768_; 
wire u2__abc_52138_new_n8769_; 
wire u2__abc_52138_new_n8770_; 
wire u2__abc_52138_new_n8771_; 
wire u2__abc_52138_new_n8772_; 
wire u2__abc_52138_new_n8773_; 
wire u2__abc_52138_new_n8774_; 
wire u2__abc_52138_new_n8775_; 
wire u2__abc_52138_new_n8776_; 
wire u2__abc_52138_new_n8777_; 
wire u2__abc_52138_new_n8778_; 
wire u2__abc_52138_new_n8779_; 
wire u2__abc_52138_new_n8780_; 
wire u2__abc_52138_new_n8781_; 
wire u2__abc_52138_new_n8782_; 
wire u2__abc_52138_new_n8784_; 
wire u2__abc_52138_new_n8785_; 
wire u2__abc_52138_new_n8786_; 
wire u2__abc_52138_new_n8787_; 
wire u2__abc_52138_new_n8788_; 
wire u2__abc_52138_new_n8789_; 
wire u2__abc_52138_new_n8790_; 
wire u2__abc_52138_new_n8792_; 
wire u2__abc_52138_new_n8793_; 
wire u2__abc_52138_new_n8794_; 
wire u2__abc_52138_new_n8795_; 
wire u2__abc_52138_new_n8796_; 
wire u2__abc_52138_new_n8797_; 
wire u2__abc_52138_new_n8798_; 
wire u2__abc_52138_new_n8799_; 
wire u2__abc_52138_new_n8801_; 
wire u2__abc_52138_new_n8802_; 
wire u2__abc_52138_new_n8803_; 
wire u2__abc_52138_new_n8804_; 
wire u2__abc_52138_new_n8805_; 
wire u2__abc_52138_new_n8806_; 
wire u2__abc_52138_new_n8807_; 
wire u2__abc_52138_new_n8808_; 
wire u2__abc_52138_new_n8810_; 
wire u2__abc_52138_new_n8811_; 
wire u2__abc_52138_new_n8812_; 
wire u2__abc_52138_new_n8813_; 
wire u2__abc_52138_new_n8814_; 
wire u2__abc_52138_new_n8815_; 
wire u2__abc_52138_new_n8816_; 
wire u2__abc_52138_new_n8817_; 
wire u2__abc_52138_new_n8818_; 
wire u2__abc_52138_new_n8819_; 
wire u2__abc_52138_new_n8820_; 
wire u2__abc_52138_new_n8821_; 
wire u2__abc_52138_new_n8822_; 
wire u2__abc_52138_new_n8823_; 
wire u2__abc_52138_new_n8825_; 
wire u2__abc_52138_new_n8826_; 
wire u2__abc_52138_new_n8827_; 
wire u2__abc_52138_new_n8828_; 
wire u2__abc_52138_new_n8829_; 
wire u2__abc_52138_new_n8830_; 
wire u2__abc_52138_new_n8831_; 
wire u2__abc_52138_new_n8833_; 
wire u2__abc_52138_new_n8834_; 
wire u2__abc_52138_new_n8835_; 
wire u2__abc_52138_new_n8836_; 
wire u2__abc_52138_new_n8837_; 
wire u2__abc_52138_new_n8838_; 
wire u2__abc_52138_new_n8839_; 
wire u2__abc_52138_new_n8840_; 
wire u2__abc_52138_new_n8842_; 
wire u2__abc_52138_new_n8843_; 
wire u2__abc_52138_new_n8844_; 
wire u2__abc_52138_new_n8845_; 
wire u2__abc_52138_new_n8846_; 
wire u2__abc_52138_new_n8847_; 
wire u2__abc_52138_new_n8848_; 
wire u2__abc_52138_new_n8850_; 
wire u2__abc_52138_new_n8851_; 
wire u2__abc_52138_new_n8852_; 
wire u2__abc_52138_new_n8853_; 
wire u2__abc_52138_new_n8854_; 
wire u2__abc_52138_new_n8855_; 
wire u2__abc_52138_new_n8856_; 
wire u2__abc_52138_new_n8857_; 
wire u2__abc_52138_new_n8858_; 
wire u2__abc_52138_new_n8859_; 
wire u2__abc_52138_new_n8860_; 
wire u2__abc_52138_new_n8861_; 
wire u2__abc_52138_new_n8862_; 
wire u2__abc_52138_new_n8863_; 
wire u2__abc_52138_new_n8865_; 
wire u2__abc_52138_new_n8866_; 
wire u2__abc_52138_new_n8867_; 
wire u2__abc_52138_new_n8868_; 
wire u2__abc_52138_new_n8869_; 
wire u2__abc_52138_new_n8870_; 
wire u2__abc_52138_new_n8871_; 
wire u2__abc_52138_new_n8872_; 
wire u2__abc_52138_new_n8874_; 
wire u2__abc_52138_new_n8875_; 
wire u2__abc_52138_new_n8876_; 
wire u2__abc_52138_new_n8877_; 
wire u2__abc_52138_new_n8878_; 
wire u2__abc_52138_new_n8879_; 
wire u2__abc_52138_new_n8880_; 
wire u2__abc_52138_new_n8881_; 
wire u2__abc_52138_new_n8882_; 
wire u2__abc_52138_new_n8884_; 
wire u2__abc_52138_new_n8885_; 
wire u2__abc_52138_new_n8886_; 
wire u2__abc_52138_new_n8887_; 
wire u2__abc_52138_new_n8888_; 
wire u2__abc_52138_new_n8889_; 
wire u2__abc_52138_new_n8890_; 
wire u2__abc_52138_new_n8891_; 
wire u2__abc_52138_new_n8893_; 
wire u2__abc_52138_new_n8894_; 
wire u2__abc_52138_new_n8895_; 
wire u2__abc_52138_new_n8896_; 
wire u2__abc_52138_new_n8897_; 
wire u2__abc_52138_new_n8898_; 
wire u2__abc_52138_new_n8899_; 
wire u2__abc_52138_new_n8900_; 
wire u2__abc_52138_new_n8901_; 
wire u2__abc_52138_new_n8902_; 
wire u2__abc_52138_new_n8903_; 
wire u2__abc_52138_new_n8904_; 
wire u2__abc_52138_new_n8905_; 
wire u2__abc_52138_new_n8907_; 
wire u2__abc_52138_new_n8908_; 
wire u2__abc_52138_new_n8909_; 
wire u2__abc_52138_new_n8910_; 
wire u2__abc_52138_new_n8911_; 
wire u2__abc_52138_new_n8912_; 
wire u2__abc_52138_new_n8913_; 
wire u2__abc_52138_new_n8915_; 
wire u2__abc_52138_new_n8916_; 
wire u2__abc_52138_new_n8917_; 
wire u2__abc_52138_new_n8918_; 
wire u2__abc_52138_new_n8919_; 
wire u2__abc_52138_new_n8920_; 
wire u2__abc_52138_new_n8921_; 
wire u2__abc_52138_new_n8922_; 
wire u2__abc_52138_new_n8923_; 
wire u2__abc_52138_new_n8925_; 
wire u2__abc_52138_new_n8926_; 
wire u2__abc_52138_new_n8927_; 
wire u2__abc_52138_new_n8928_; 
wire u2__abc_52138_new_n8929_; 
wire u2__abc_52138_new_n8930_; 
wire u2__abc_52138_new_n8931_; 
wire u2__abc_52138_new_n8932_; 
wire u2__abc_52138_new_n8934_; 
wire u2__abc_52138_new_n8935_; 
wire u2__abc_52138_new_n8936_; 
wire u2__abc_52138_new_n8937_; 
wire u2__abc_52138_new_n8938_; 
wire u2__abc_52138_new_n8939_; 
wire u2__abc_52138_new_n8940_; 
wire u2__abc_52138_new_n8941_; 
wire u2__abc_52138_new_n8942_; 
wire u2__abc_52138_new_n8943_; 
wire u2__abc_52138_new_n8944_; 
wire u2__abc_52138_new_n8945_; 
wire u2__abc_52138_new_n8946_; 
wire u2__abc_52138_new_n8947_; 
wire u2__abc_52138_new_n8948_; 
wire u2__abc_52138_new_n8949_; 
wire u2__abc_52138_new_n8950_; 
wire u2__abc_52138_new_n8951_; 
wire u2__abc_52138_new_n8952_; 
wire u2__abc_52138_new_n8954_; 
wire u2__abc_52138_new_n8955_; 
wire u2__abc_52138_new_n8956_; 
wire u2__abc_52138_new_n8957_; 
wire u2__abc_52138_new_n8958_; 
wire u2__abc_52138_new_n8959_; 
wire u2__abc_52138_new_n8960_; 
wire u2__abc_52138_new_n8962_; 
wire u2__abc_52138_new_n8963_; 
wire u2__abc_52138_new_n8964_; 
wire u2__abc_52138_new_n8965_; 
wire u2__abc_52138_new_n8966_; 
wire u2__abc_52138_new_n8967_; 
wire u2__abc_52138_new_n8968_; 
wire u2__abc_52138_new_n8969_; 
wire u2__abc_52138_new_n8971_; 
wire u2__abc_52138_new_n8972_; 
wire u2__abc_52138_new_n8973_; 
wire u2__abc_52138_new_n8974_; 
wire u2__abc_52138_new_n8975_; 
wire u2__abc_52138_new_n8976_; 
wire u2__abc_52138_new_n8977_; 
wire u2__abc_52138_new_n8979_; 
wire u2__abc_52138_new_n8980_; 
wire u2__abc_52138_new_n8981_; 
wire u2__abc_52138_new_n8982_; 
wire u2__abc_52138_new_n8983_; 
wire u2__abc_52138_new_n8984_; 
wire u2__abc_52138_new_n8985_; 
wire u2__abc_52138_new_n8986_; 
wire u2__abc_52138_new_n8987_; 
wire u2__abc_52138_new_n8988_; 
wire u2__abc_52138_new_n8989_; 
wire u2__abc_52138_new_n8990_; 
wire u2__abc_52138_new_n8992_; 
wire u2__abc_52138_new_n8993_; 
wire u2__abc_52138_new_n8994_; 
wire u2__abc_52138_new_n8995_; 
wire u2__abc_52138_new_n8996_; 
wire u2__abc_52138_new_n8997_; 
wire u2__abc_52138_new_n8998_; 
wire u2__abc_52138_new_n9000_; 
wire u2__abc_52138_new_n9001_; 
wire u2__abc_52138_new_n9002_; 
wire u2__abc_52138_new_n9003_; 
wire u2__abc_52138_new_n9004_; 
wire u2__abc_52138_new_n9005_; 
wire u2__abc_52138_new_n9006_; 
wire u2__abc_52138_new_n9007_; 
wire u2__abc_52138_new_n9008_; 
wire u2__abc_52138_new_n9010_; 
wire u2__abc_52138_new_n9011_; 
wire u2__abc_52138_new_n9012_; 
wire u2__abc_52138_new_n9013_; 
wire u2__abc_52138_new_n9014_; 
wire u2__abc_52138_new_n9015_; 
wire u2__abc_52138_new_n9016_; 
wire u2__abc_52138_new_n9018_; 
wire u2__abc_52138_new_n9019_; 
wire u2__abc_52138_new_n9020_; 
wire u2__abc_52138_new_n9021_; 
wire u2__abc_52138_new_n9022_; 
wire u2__abc_52138_new_n9023_; 
wire u2__abc_52138_new_n9024_; 
wire u2__abc_52138_new_n9025_; 
wire u2__abc_52138_new_n9026_; 
wire u2__abc_52138_new_n9027_; 
wire u2__abc_52138_new_n9028_; 
wire u2__abc_52138_new_n9029_; 
wire u2__abc_52138_new_n9030_; 
wire u2__abc_52138_new_n9031_; 
wire u2__abc_52138_new_n9033_; 
wire u2__abc_52138_new_n9034_; 
wire u2__abc_52138_new_n9035_; 
wire u2__abc_52138_new_n9036_; 
wire u2__abc_52138_new_n9037_; 
wire u2__abc_52138_new_n9038_; 
wire u2__abc_52138_new_n9039_; 
wire u2__abc_52138_new_n9040_; 
wire u2__abc_52138_new_n9042_; 
wire u2__abc_52138_new_n9043_; 
wire u2__abc_52138_new_n9044_; 
wire u2__abc_52138_new_n9045_; 
wire u2__abc_52138_new_n9046_; 
wire u2__abc_52138_new_n9047_; 
wire u2__abc_52138_new_n9048_; 
wire u2__abc_52138_new_n9049_; 
wire u2__abc_52138_new_n9050_; 
wire u2__abc_52138_new_n9052_; 
wire u2__abc_52138_new_n9053_; 
wire u2__abc_52138_new_n9054_; 
wire u2__abc_52138_new_n9055_; 
wire u2__abc_52138_new_n9056_; 
wire u2__abc_52138_new_n9057_; 
wire u2__abc_52138_new_n9058_; 
wire u2__abc_52138_new_n9060_; 
wire u2__abc_52138_new_n9061_; 
wire u2__abc_52138_new_n9062_; 
wire u2__abc_52138_new_n9063_; 
wire u2__abc_52138_new_n9064_; 
wire u2__abc_52138_new_n9065_; 
wire u2__abc_52138_new_n9066_; 
wire u2__abc_52138_new_n9067_; 
wire u2__abc_52138_new_n9068_; 
wire u2__abc_52138_new_n9069_; 
wire u2__abc_52138_new_n9071_; 
wire u2__abc_52138_new_n9072_; 
wire u2__abc_52138_new_n9073_; 
wire u2__abc_52138_new_n9074_; 
wire u2__abc_52138_new_n9075_; 
wire u2__abc_52138_new_n9076_; 
wire u2__abc_52138_new_n9077_; 
wire u2__abc_52138_new_n9079_; 
wire u2__abc_52138_new_n9080_; 
wire u2__abc_52138_new_n9081_; 
wire u2__abc_52138_new_n9082_; 
wire u2__abc_52138_new_n9083_; 
wire u2__abc_52138_new_n9084_; 
wire u2__abc_52138_new_n9085_; 
wire u2__abc_52138_new_n9086_; 
wire u2__abc_52138_new_n9088_; 
wire u2__abc_52138_new_n9089_; 
wire u2__abc_52138_new_n9090_; 
wire u2__abc_52138_new_n9091_; 
wire u2__abc_52138_new_n9092_; 
wire u2__abc_52138_new_n9093_; 
wire u2__abc_52138_new_n9094_; 
wire u2__abc_52138_new_n9096_; 
wire u2__abc_52138_new_n9097_; 
wire u2__abc_52138_new_n9098_; 
wire u2__abc_52138_new_n9099_; 
wire u2__abc_52138_new_n9100_; 
wire u2__abc_52138_new_n9101_; 
wire u2__abc_52138_new_n9102_; 
wire u2__abc_52138_new_n9103_; 
wire u2__abc_52138_new_n9104_; 
wire u2__abc_52138_new_n9105_; 
wire u2__abc_52138_new_n9106_; 
wire u2__abc_52138_new_n9107_; 
wire u2__abc_52138_new_n9108_; 
wire u2__abc_52138_new_n9109_; 
wire u2__abc_52138_new_n9110_; 
wire u2__abc_52138_new_n9111_; 
wire u2__abc_52138_new_n9112_; 
wire u2__abc_52138_new_n9114_; 
wire u2__abc_52138_new_n9115_; 
wire u2__abc_52138_new_n9116_; 
wire u2__abc_52138_new_n9117_; 
wire u2__abc_52138_new_n9118_; 
wire u2__abc_52138_new_n9119_; 
wire u2__abc_52138_new_n9120_; 
wire u2__abc_52138_new_n9121_; 
wire u2__abc_52138_new_n9123_; 
wire u2__abc_52138_new_n9124_; 
wire u2__abc_52138_new_n9125_; 
wire u2__abc_52138_new_n9126_; 
wire u2__abc_52138_new_n9127_; 
wire u2__abc_52138_new_n9128_; 
wire u2__abc_52138_new_n9129_; 
wire u2__abc_52138_new_n9130_; 
wire u2__abc_52138_new_n9131_; 
wire u2__abc_52138_new_n9133_; 
wire u2__abc_52138_new_n9134_; 
wire u2__abc_52138_new_n9135_; 
wire u2__abc_52138_new_n9136_; 
wire u2__abc_52138_new_n9137_; 
wire u2__abc_52138_new_n9138_; 
wire u2__abc_52138_new_n9139_; 
wire u2__abc_52138_new_n9140_; 
wire u2__abc_52138_new_n9142_; 
wire u2__abc_52138_new_n9143_; 
wire u2__abc_52138_new_n9144_; 
wire u2__abc_52138_new_n9145_; 
wire u2__abc_52138_new_n9146_; 
wire u2__abc_52138_new_n9147_; 
wire u2__abc_52138_new_n9148_; 
wire u2__abc_52138_new_n9149_; 
wire u2__abc_52138_new_n9150_; 
wire u2__abc_52138_new_n9151_; 
wire u2__abc_52138_new_n9152_; 
wire u2__abc_52138_new_n9154_; 
wire u2__abc_52138_new_n9155_; 
wire u2__abc_52138_new_n9156_; 
wire u2__abc_52138_new_n9157_; 
wire u2__abc_52138_new_n9158_; 
wire u2__abc_52138_new_n9159_; 
wire u2__abc_52138_new_n9160_; 
wire u2__abc_52138_new_n9162_; 
wire u2__abc_52138_new_n9163_; 
wire u2__abc_52138_new_n9164_; 
wire u2__abc_52138_new_n9165_; 
wire u2__abc_52138_new_n9166_; 
wire u2__abc_52138_new_n9167_; 
wire u2__abc_52138_new_n9168_; 
wire u2__abc_52138_new_n9169_; 
wire u2__abc_52138_new_n9170_; 
wire u2__abc_52138_new_n9172_; 
wire u2__abc_52138_new_n9173_; 
wire u2__abc_52138_new_n9174_; 
wire u2__abc_52138_new_n9175_; 
wire u2__abc_52138_new_n9176_; 
wire u2__abc_52138_new_n9177_; 
wire u2__abc_52138_new_n9178_; 
wire u2__abc_52138_new_n9179_; 
wire u2__abc_52138_new_n9181_; 
wire u2__abc_52138_new_n9182_; 
wire u2__abc_52138_new_n9183_; 
wire u2__abc_52138_new_n9184_; 
wire u2__abc_52138_new_n9185_; 
wire u2__abc_52138_new_n9186_; 
wire u2__abc_52138_new_n9187_; 
wire u2__abc_52138_new_n9188_; 
wire u2__abc_52138_new_n9189_; 
wire u2__abc_52138_new_n9190_; 
wire u2__abc_52138_new_n9191_; 
wire u2__abc_52138_new_n9192_; 
wire u2__abc_52138_new_n9193_; 
wire u2__abc_52138_new_n9194_; 
wire u2__abc_52138_new_n9196_; 
wire u2__abc_52138_new_n9197_; 
wire u2__abc_52138_new_n9198_; 
wire u2__abc_52138_new_n9199_; 
wire u2__abc_52138_new_n9200_; 
wire u2__abc_52138_new_n9201_; 
wire u2__abc_52138_new_n9202_; 
wire u2__abc_52138_new_n9204_; 
wire u2__abc_52138_new_n9205_; 
wire u2__abc_52138_new_n9206_; 
wire u2__abc_52138_new_n9207_; 
wire u2__abc_52138_new_n9208_; 
wire u2__abc_52138_new_n9209_; 
wire u2__abc_52138_new_n9210_; 
wire u2__abc_52138_new_n9211_; 
wire u2__abc_52138_new_n9212_; 
wire u2__abc_52138_new_n9213_; 
wire u2__abc_52138_new_n9214_; 
wire u2__abc_52138_new_n9216_; 
wire u2__abc_52138_new_n9217_; 
wire u2__abc_52138_new_n9218_; 
wire u2__abc_52138_new_n9219_; 
wire u2__abc_52138_new_n9220_; 
wire u2__abc_52138_new_n9221_; 
wire u2__abc_52138_new_n9222_; 
wire u2__abc_52138_new_n9223_; 
wire u2__abc_52138_new_n9225_; 
wire u2__abc_52138_new_n9226_; 
wire u2__abc_52138_new_n9227_; 
wire u2__abc_52138_new_n9228_; 
wire u2__abc_52138_new_n9229_; 
wire u2__abc_52138_new_n9230_; 
wire u2__abc_52138_new_n9231_; 
wire u2__abc_52138_new_n9232_; 
wire u2__abc_52138_new_n9233_; 
wire u2__abc_52138_new_n9234_; 
wire u2__abc_52138_new_n9235_; 
wire u2__abc_52138_new_n9236_; 
wire u2__abc_52138_new_n9238_; 
wire u2__abc_52138_new_n9239_; 
wire u2__abc_52138_new_n9240_; 
wire u2__abc_52138_new_n9241_; 
wire u2__abc_52138_new_n9242_; 
wire u2__abc_52138_new_n9243_; 
wire u2__abc_52138_new_n9244_; 
wire u2__abc_52138_new_n9246_; 
wire u2__abc_52138_new_n9247_; 
wire u2__abc_52138_new_n9248_; 
wire u2__abc_52138_new_n9249_; 
wire u2__abc_52138_new_n9250_; 
wire u2__abc_52138_new_n9251_; 
wire u2__abc_52138_new_n9252_; 
wire u2__abc_52138_new_n9253_; 
wire u2__abc_52138_new_n9255_; 
wire u2__abc_52138_new_n9256_; 
wire u2__abc_52138_new_n9257_; 
wire u2__abc_52138_new_n9258_; 
wire u2__abc_52138_new_n9259_; 
wire u2__abc_52138_new_n9260_; 
wire u2__abc_52138_new_n9261_; 
wire u2__abc_52138_new_n9263_; 
wire u2__abc_52138_new_n9264_; 
wire u2__abc_52138_new_n9265_; 
wire u2__abc_52138_new_n9266_; 
wire u2__abc_52138_new_n9267_; 
wire u2__abc_52138_new_n9268_; 
wire u2__abc_52138_new_n9269_; 
wire u2__abc_52138_new_n9270_; 
wire u2__abc_52138_new_n9271_; 
wire u2__abc_52138_new_n9272_; 
wire u2__abc_52138_new_n9273_; 
wire u2__abc_52138_new_n9274_; 
wire u2__abc_52138_new_n9275_; 
wire u2__abc_52138_new_n9276_; 
wire u2__abc_52138_new_n9277_; 
wire u2__abc_52138_new_n9278_; 
wire u2__abc_52138_new_n9279_; 
wire u2__abc_52138_new_n9280_; 
wire u2__abc_52138_new_n9281_; 
wire u2__abc_52138_new_n9282_; 
wire u2__abc_52138_new_n9283_; 
wire u2__abc_52138_new_n9285_; 
wire u2__abc_52138_new_n9286_; 
wire u2__abc_52138_new_n9287_; 
wire u2__abc_52138_new_n9288_; 
wire u2__abc_52138_new_n9289_; 
wire u2__abc_52138_new_n9290_; 
wire u2__abc_52138_new_n9291_; 
wire u2__abc_52138_new_n9292_; 
wire u2__abc_52138_new_n9293_; 
wire u2__abc_52138_new_n9294_; 
wire u2__abc_52138_new_n9296_; 
wire u2__abc_52138_new_n9297_; 
wire u2__abc_52138_new_n9298_; 
wire u2__abc_52138_new_n9299_; 
wire u2__abc_52138_new_n9300_; 
wire u2__abc_52138_new_n9301_; 
wire u2__abc_52138_new_n9302_; 
wire u2__abc_52138_new_n9303_; 
wire u2__abc_52138_new_n9305_; 
wire u2__abc_52138_new_n9306_; 
wire u2__abc_52138_new_n9307_; 
wire u2__abc_52138_new_n9308_; 
wire u2__abc_52138_new_n9309_; 
wire u2__abc_52138_new_n9310_; 
wire u2__abc_52138_new_n9311_; 
wire u2__abc_52138_new_n9312_; 
wire u2__abc_52138_new_n9313_; 
wire u2__abc_52138_new_n9315_; 
wire u2__abc_52138_new_n9316_; 
wire u2__abc_52138_new_n9317_; 
wire u2__abc_52138_new_n9318_; 
wire u2__abc_52138_new_n9319_; 
wire u2__abc_52138_new_n9320_; 
wire u2__abc_52138_new_n9321_; 
wire u2__abc_52138_new_n9322_; 
wire u2__abc_52138_new_n9323_; 
wire u2__abc_52138_new_n9324_; 
wire u2__abc_52138_new_n9325_; 
wire u2__abc_52138_new_n9326_; 
wire u2__abc_52138_new_n9327_; 
wire u2__abc_52138_new_n9328_; 
wire u2__abc_52138_new_n9330_; 
wire u2__abc_52138_new_n9331_; 
wire u2__abc_52138_new_n9332_; 
wire u2__abc_52138_new_n9333_; 
wire u2__abc_52138_new_n9334_; 
wire u2__abc_52138_new_n9335_; 
wire u2__abc_52138_new_n9336_; 
wire u2__abc_52138_new_n9338_; 
wire u2__abc_52138_new_n9339_; 
wire u2__abc_52138_new_n9340_; 
wire u2__abc_52138_new_n9341_; 
wire u2__abc_52138_new_n9342_; 
wire u2__abc_52138_new_n9343_; 
wire u2__abc_52138_new_n9344_; 
wire u2__abc_52138_new_n9345_; 
wire u2__abc_52138_new_n9346_; 
wire u2__abc_52138_new_n9347_; 
wire u2__abc_52138_new_n9348_; 
wire u2__abc_52138_new_n9350_; 
wire u2__abc_52138_new_n9351_; 
wire u2__abc_52138_new_n9352_; 
wire u2__abc_52138_new_n9353_; 
wire u2__abc_52138_new_n9354_; 
wire u2__abc_52138_new_n9355_; 
wire u2__abc_52138_new_n9356_; 
wire u2__abc_52138_new_n9357_; 
wire u2__abc_52138_new_n9359_; 
wire u2__abc_52138_new_n9360_; 
wire u2__abc_52138_new_n9361_; 
wire u2__abc_52138_new_n9362_; 
wire u2__abc_52138_new_n9363_; 
wire u2__abc_52138_new_n9364_; 
wire u2__abc_52138_new_n9365_; 
wire u2__abc_52138_new_n9366_; 
wire u2__abc_52138_new_n9367_; 
wire u2__abc_52138_new_n9368_; 
wire u2__abc_52138_new_n9369_; 
wire u2__abc_52138_new_n9371_; 
wire u2__abc_52138_new_n9372_; 
wire u2__abc_52138_new_n9373_; 
wire u2__abc_52138_new_n9374_; 
wire u2__abc_52138_new_n9375_; 
wire u2__abc_52138_new_n9376_; 
wire u2__abc_52138_new_n9377_; 
wire u2__abc_52138_new_n9378_; 
wire u2__abc_52138_new_n9379_; 
wire u2__abc_52138_new_n9381_; 
wire u2__abc_52138_new_n9382_; 
wire u2__abc_52138_new_n9383_; 
wire u2__abc_52138_new_n9384_; 
wire u2__abc_52138_new_n9385_; 
wire u2__abc_52138_new_n9386_; 
wire u2__abc_52138_new_n9387_; 
wire u2__abc_52138_new_n9388_; 
wire u2__abc_52138_new_n9390_; 
wire u2__abc_52138_new_n9391_; 
wire u2__abc_52138_new_n9392_; 
wire u2__abc_52138_new_n9393_; 
wire u2__abc_52138_new_n9394_; 
wire u2__abc_52138_new_n9395_; 
wire u2__abc_52138_new_n9396_; 
wire u2__abc_52138_new_n9397_; 
wire u2__abc_52138_new_n9399_; 
wire u2__abc_52138_new_n9400_; 
wire u2__abc_52138_new_n9401_; 
wire u2__abc_52138_new_n9402_; 
wire u2__abc_52138_new_n9403_; 
wire u2__abc_52138_new_n9404_; 
wire u2__abc_52138_new_n9405_; 
wire u2__abc_52138_new_n9406_; 
wire u2__abc_52138_new_n9407_; 
wire u2__abc_52138_new_n9409_; 
wire u2__abc_52138_new_n9410_; 
wire u2__abc_52138_new_n9411_; 
wire u2__abc_52138_new_n9412_; 
wire u2__abc_52138_new_n9413_; 
wire u2__abc_52138_new_n9414_; 
wire u2__abc_52138_new_n9415_; 
wire u2__abc_52138_new_n9417_; 
wire u2__abc_52138_new_n9418_; 
wire u2__abc_52138_new_n9419_; 
wire u2__abc_52138_new_n9420_; 
wire u2__abc_52138_new_n9421_; 
wire u2__abc_52138_new_n9422_; 
wire u2__abc_52138_new_n9423_; 
wire u2__abc_52138_new_n9424_; 
wire u2__abc_52138_new_n9425_; 
wire u2__abc_52138_new_n9426_; 
wire u2__abc_52138_new_n9427_; 
wire u2__abc_52138_new_n9429_; 
wire u2__abc_52138_new_n9430_; 
wire u2__abc_52138_new_n9431_; 
wire u2__abc_52138_new_n9432_; 
wire u2__abc_52138_new_n9433_; 
wire u2__abc_52138_new_n9434_; 
wire u2__abc_52138_new_n9435_; 
wire u2__abc_52138_new_n9436_; 
wire u2__abc_52138_new_n9438_; 
wire u2__abc_52138_new_n9439_; 
wire u2__abc_52138_new_n9440_; 
wire u2__abc_52138_new_n9441_; 
wire u2__abc_52138_new_n9442_; 
wire u2__abc_52138_new_n9443_; 
wire u2__abc_52138_new_n9444_; 
wire u2__abc_52138_new_n9445_; 
wire u2__abc_52138_new_n9446_; 
wire u2__abc_52138_new_n9447_; 
wire u2__abc_52138_new_n9448_; 
wire u2__abc_52138_new_n9449_; 
wire u2__abc_52138_new_n9450_; 
wire u2__abc_52138_new_n9451_; 
wire u2__abc_52138_new_n9452_; 
wire u2__abc_52138_new_n9453_; 
wire u2__abc_52138_new_n9454_; 
wire u2__abc_52138_new_n9456_; 
wire u2__abc_52138_new_n9457_; 
wire u2__abc_52138_new_n9458_; 
wire u2__abc_52138_new_n9459_; 
wire u2__abc_52138_new_n9460_; 
wire u2__abc_52138_new_n9461_; 
wire u2__abc_52138_new_n9462_; 
wire u2__abc_52138_new_n9464_; 
wire u2__abc_52138_new_n9465_; 
wire u2__abc_52138_new_n9466_; 
wire u2__abc_52138_new_n9467_; 
wire u2__abc_52138_new_n9468_; 
wire u2__abc_52138_new_n9469_; 
wire u2__abc_52138_new_n9470_; 
wire u2__abc_52138_new_n9471_; 
wire u2__abc_52138_new_n9472_; 
wire u2__abc_52138_new_n9473_; 
wire u2__abc_52138_new_n9475_; 
wire u2__abc_52138_new_n9476_; 
wire u2__abc_52138_new_n9477_; 
wire u2__abc_52138_new_n9478_; 
wire u2__abc_52138_new_n9479_; 
wire u2__abc_52138_new_n9480_; 
wire u2__abc_52138_new_n9481_; 
wire u2__abc_52138_new_n9482_; 
wire u2__abc_52138_new_n9484_; 
wire u2__abc_52138_new_n9485_; 
wire u2__abc_52138_new_n9486_; 
wire u2__abc_52138_new_n9487_; 
wire u2__abc_52138_new_n9488_; 
wire u2__abc_52138_new_n9489_; 
wire u2__abc_52138_new_n9490_; 
wire u2__abc_52138_new_n9491_; 
wire u2__abc_52138_new_n9492_; 
wire u2__abc_52138_new_n9493_; 
wire u2__abc_52138_new_n9494_; 
wire u2__abc_52138_new_n9495_; 
wire u2__abc_52138_new_n9496_; 
wire u2__abc_52138_new_n9497_; 
wire u2__abc_52138_new_n9499_; 
wire u2__abc_52138_new_n9500_; 
wire u2__abc_52138_new_n9501_; 
wire u2__abc_52138_new_n9502_; 
wire u2__abc_52138_new_n9503_; 
wire u2__abc_52138_new_n9504_; 
wire u2__abc_52138_new_n9505_; 
wire u2__abc_52138_new_n9507_; 
wire u2__abc_52138_new_n9508_; 
wire u2__abc_52138_new_n9509_; 
wire u2__abc_52138_new_n9510_; 
wire u2__abc_52138_new_n9511_; 
wire u2__abc_52138_new_n9512_; 
wire u2__abc_52138_new_n9513_; 
wire u2__abc_52138_new_n9514_; 
wire u2__abc_52138_new_n9515_; 
wire u2__abc_52138_new_n9516_; 
wire u2__abc_52138_new_n9518_; 
wire u2__abc_52138_new_n9519_; 
wire u2__abc_52138_new_n9520_; 
wire u2__abc_52138_new_n9521_; 
wire u2__abc_52138_new_n9522_; 
wire u2__abc_52138_new_n9523_; 
wire u2__abc_52138_new_n9524_; 
wire u2__abc_52138_new_n9525_; 
wire u2__abc_52138_new_n9527_; 
wire u2__abc_52138_new_n9528_; 
wire u2__abc_52138_new_n9529_; 
wire u2__abc_52138_new_n9530_; 
wire u2__abc_52138_new_n9531_; 
wire u2__abc_52138_new_n9532_; 
wire u2__abc_52138_new_n9533_; 
wire u2__abc_52138_new_n9534_; 
wire u2__abc_52138_new_n9535_; 
wire u2__abc_52138_new_n9536_; 
wire u2__abc_52138_new_n9537_; 
wire u2__abc_52138_new_n9538_; 
wire u2__abc_52138_new_n9539_; 
wire u2__abc_52138_new_n9541_; 
wire u2__abc_52138_new_n9542_; 
wire u2__abc_52138_new_n9543_; 
wire u2__abc_52138_new_n9544_; 
wire u2__abc_52138_new_n9545_; 
wire u2__abc_52138_new_n9546_; 
wire u2__abc_52138_new_n9547_; 
wire u2__abc_52138_new_n9549_; 
wire u2__abc_52138_new_n9550_; 
wire u2__abc_52138_new_n9551_; 
wire u2__abc_52138_new_n9552_; 
wire u2__abc_52138_new_n9553_; 
wire u2__abc_52138_new_n9554_; 
wire u2__abc_52138_new_n9555_; 
wire u2__abc_52138_new_n9556_; 
wire u2__abc_52138_new_n9557_; 
wire u2__abc_52138_new_n9559_; 
wire u2__abc_52138_new_n9560_; 
wire u2__abc_52138_new_n9561_; 
wire u2__abc_52138_new_n9562_; 
wire u2__abc_52138_new_n9563_; 
wire u2__abc_52138_new_n9564_; 
wire u2__abc_52138_new_n9565_; 
wire u2__abc_52138_new_n9566_; 
wire u2__abc_52138_new_n9568_; 
wire u2__abc_52138_new_n9569_; 
wire u2__abc_52138_new_n9570_; 
wire u2__abc_52138_new_n9571_; 
wire u2__abc_52138_new_n9572_; 
wire u2__abc_52138_new_n9573_; 
wire u2__abc_52138_new_n9574_; 
wire u2__abc_52138_new_n9575_; 
wire u2__abc_52138_new_n9576_; 
wire u2__abc_52138_new_n9577_; 
wire u2__abc_52138_new_n9578_; 
wire u2__abc_52138_new_n9579_; 
wire u2__abc_52138_new_n9580_; 
wire u2__abc_52138_new_n9581_; 
wire u2__abc_52138_new_n9583_; 
wire u2__abc_52138_new_n9584_; 
wire u2__abc_52138_new_n9585_; 
wire u2__abc_52138_new_n9586_; 
wire u2__abc_52138_new_n9587_; 
wire u2__abc_52138_new_n9588_; 
wire u2__abc_52138_new_n9589_; 
wire u2__abc_52138_new_n9590_; 
wire u2__abc_52138_new_n9592_; 
wire u2__abc_52138_new_n9593_; 
wire u2__abc_52138_new_n9594_; 
wire u2__abc_52138_new_n9595_; 
wire u2__abc_52138_new_n9596_; 
wire u2__abc_52138_new_n9597_; 
wire u2__abc_52138_new_n9598_; 
wire u2__abc_52138_new_n9599_; 
wire u2__abc_52138_new_n9600_; 
wire u2__abc_52138_new_n9601_; 
wire u2__abc_52138_new_n9603_; 
wire u2__abc_52138_new_n9604_; 
wire u2__abc_52138_new_n9605_; 
wire u2__abc_52138_new_n9606_; 
wire u2__abc_52138_new_n9607_; 
wire u2__abc_52138_new_n9608_; 
wire u2__abc_52138_new_n9609_; 
wire u2__abc_52138_new_n9610_; 
wire u2__abc_52138_new_n9612_; 
wire u2__abc_52138_new_n9613_; 
wire u2__abc_52138_new_n9614_; 
wire u2__abc_52138_new_n9615_; 
wire u2__abc_52138_new_n9616_; 
wire u2__abc_52138_new_n9617_; 
wire u2__abc_52138_new_n9618_; 
wire u2__abc_52138_new_n9619_; 
wire u2__abc_52138_new_n9620_; 
wire u2__abc_52138_new_n9621_; 
wire u2__abc_52138_new_n9622_; 
wire u2__abc_52138_new_n9623_; 
wire u2__abc_52138_new_n9624_; 
wire u2__abc_52138_new_n9625_; 
wire u2__abc_52138_new_n9626_; 
wire u2__abc_52138_new_n9627_; 
wire u2__abc_52138_new_n9628_; 
wire u2__abc_52138_new_n9629_; 
wire u2__abc_52138_new_n9631_; 
wire u2__abc_52138_new_n9632_; 
wire u2__abc_52138_new_n9633_; 
wire u2__abc_52138_new_n9634_; 
wire u2__abc_52138_new_n9635_; 
wire u2__abc_52138_new_n9636_; 
wire u2__abc_52138_new_n9637_; 
wire u2__abc_52138_new_n9639_; 
wire u2__abc_52138_new_n9640_; 
wire u2__abc_52138_new_n9641_; 
wire u2__abc_52138_new_n9642_; 
wire u2__abc_52138_new_n9643_; 
wire u2__abc_52138_new_n9644_; 
wire u2__abc_52138_new_n9645_; 
wire u2__abc_52138_new_n9646_; 
wire u2__abc_52138_new_n9647_; 
wire u2__abc_52138_new_n9648_; 
wire u2__abc_52138_new_n9650_; 
wire u2__abc_52138_new_n9651_; 
wire u2__abc_52138_new_n9652_; 
wire u2__abc_52138_new_n9653_; 
wire u2__abc_52138_new_n9654_; 
wire u2__abc_52138_new_n9655_; 
wire u2__abc_52138_new_n9656_; 
wire u2__abc_52138_new_n9657_; 
wire u2__abc_52138_new_n9659_; 
wire u2__abc_52138_new_n9660_; 
wire u2__abc_52138_new_n9661_; 
wire u2__abc_52138_new_n9662_; 
wire u2__abc_52138_new_n9663_; 
wire u2__abc_52138_new_n9664_; 
wire u2__abc_52138_new_n9665_; 
wire u2__abc_52138_new_n9666_; 
wire u2__abc_52138_new_n9667_; 
wire u2__abc_52138_new_n9668_; 
wire u2__abc_52138_new_n9669_; 
wire u2__abc_52138_new_n9670_; 
wire u2__abc_52138_new_n9671_; 
wire u2__abc_52138_new_n9672_; 
wire u2__abc_52138_new_n9673_; 
wire u2__abc_52138_new_n9675_; 
wire u2__abc_52138_new_n9676_; 
wire u2__abc_52138_new_n9677_; 
wire u2__abc_52138_new_n9678_; 
wire u2__abc_52138_new_n9679_; 
wire u2__abc_52138_new_n9680_; 
wire u2__abc_52138_new_n9681_; 
wire u2__abc_52138_new_n9683_; 
wire u2__abc_52138_new_n9684_; 
wire u2__abc_52138_new_n9685_; 
wire u2__abc_52138_new_n9686_; 
wire u2__abc_52138_new_n9687_; 
wire u2__abc_52138_new_n9688_; 
wire u2__abc_52138_new_n9689_; 
wire u2__abc_52138_new_n9690_; 
wire u2__abc_52138_new_n9691_; 
wire u2__abc_52138_new_n9692_; 
wire u2__abc_52138_new_n9694_; 
wire u2__abc_52138_new_n9695_; 
wire u2__abc_52138_new_n9696_; 
wire u2__abc_52138_new_n9697_; 
wire u2__abc_52138_new_n9698_; 
wire u2__abc_52138_new_n9699_; 
wire u2__abc_52138_new_n9700_; 
wire u2__abc_52138_new_n9701_; 
wire u2__abc_52138_new_n9703_; 
wire u2__abc_52138_new_n9704_; 
wire u2__abc_52138_new_n9705_; 
wire u2__abc_52138_new_n9706_; 
wire u2__abc_52138_new_n9707_; 
wire u2__abc_52138_new_n9708_; 
wire u2__abc_52138_new_n9709_; 
wire u2__abc_52138_new_n9710_; 
wire u2__abc_52138_new_n9711_; 
wire u2__abc_52138_new_n9712_; 
wire u2__abc_52138_new_n9713_; 
wire u2__abc_52138_new_n9715_; 
wire u2__abc_52138_new_n9716_; 
wire u2__abc_52138_new_n9717_; 
wire u2__abc_52138_new_n9718_; 
wire u2__abc_52138_new_n9719_; 
wire u2__abc_52138_new_n9720_; 
wire u2__abc_52138_new_n9721_; 
wire u2__abc_52138_new_n9722_; 
wire u2__abc_52138_new_n9723_; 
wire u2__abc_52138_new_n9725_; 
wire u2__abc_52138_new_n9726_; 
wire u2__abc_52138_new_n9727_; 
wire u2__abc_52138_new_n9728_; 
wire u2__abc_52138_new_n9729_; 
wire u2__abc_52138_new_n9730_; 
wire u2__abc_52138_new_n9731_; 
wire u2__abc_52138_new_n9732_; 
wire u2__abc_52138_new_n9733_; 
wire u2__abc_52138_new_n9735_; 
wire u2__abc_52138_new_n9736_; 
wire u2__abc_52138_new_n9737_; 
wire u2__abc_52138_new_n9738_; 
wire u2__abc_52138_new_n9739_; 
wire u2__abc_52138_new_n9740_; 
wire u2__abc_52138_new_n9741_; 
wire u2__abc_52138_new_n9742_; 
wire u2__abc_52138_new_n9744_; 
wire u2__abc_52138_new_n9745_; 
wire u2__abc_52138_new_n9746_; 
wire u2__abc_52138_new_n9747_; 
wire u2__abc_52138_new_n9748_; 
wire u2__abc_52138_new_n9749_; 
wire u2__abc_52138_new_n9750_; 
wire u2__abc_52138_new_n9751_; 
wire u2__abc_52138_new_n9752_; 
wire u2__abc_52138_new_n9753_; 
wire u2__abc_52138_new_n9754_; 
wire u2__abc_52138_new_n9755_; 
wire u2__abc_52138_new_n9757_; 
wire u2__abc_52138_new_n9758_; 
wire u2__abc_52138_new_n9759_; 
wire u2__abc_52138_new_n9760_; 
wire u2__abc_52138_new_n9761_; 
wire u2__abc_52138_new_n9762_; 
wire u2__abc_52138_new_n9763_; 
wire u2__abc_52138_new_n9765_; 
wire u2__abc_52138_new_n9766_; 
wire u2__abc_52138_new_n9767_; 
wire u2__abc_52138_new_n9768_; 
wire u2__abc_52138_new_n9769_; 
wire u2__abc_52138_new_n9770_; 
wire u2__abc_52138_new_n9771_; 
wire u2__abc_52138_new_n9772_; 
wire u2__abc_52138_new_n9773_; 
wire u2__abc_52138_new_n9774_; 
wire u2__abc_52138_new_n9775_; 
wire u2__abc_52138_new_n9777_; 
wire u2__abc_52138_new_n9778_; 
wire u2__abc_52138_new_n9779_; 
wire u2__abc_52138_new_n9780_; 
wire u2__abc_52138_new_n9781_; 
wire u2__abc_52138_new_n9782_; 
wire u2__abc_52138_new_n9783_; 
wire u2__abc_52138_new_n9784_; 
wire u2__abc_52138_new_n9786_; 
wire u2__abc_52138_new_n9787_; 
wire u2__abc_52138_new_n9788_; 
wire u2__abc_52138_new_n9789_; 
wire u2__abc_52138_new_n9790_; 
wire u2__abc_52138_new_n9791_; 
wire u2__abc_52138_new_n9792_; 
wire u2__abc_52138_new_n9793_; 
wire u2__abc_52138_new_n9794_; 
wire u2__abc_52138_new_n9795_; 
wire u2__abc_52138_new_n9796_; 
wire u2__abc_52138_new_n9797_; 
wire u2__abc_52138_new_n9798_; 
wire u2__abc_52138_new_n9799_; 
wire u2__abc_52138_new_n9801_; 
wire u2__abc_52138_new_n9802_; 
wire u2__abc_52138_new_n9803_; 
wire u2__abc_52138_new_n9804_; 
wire u2__abc_52138_new_n9805_; 
wire u2__abc_52138_new_n9806_; 
wire u2__abc_52138_new_n9807_; 
wire u2__abc_52138_new_n9808_; 
wire u2__abc_52138_new_n9809_; 
wire u2__abc_52138_new_n9811_; 
wire u2__abc_52138_new_n9812_; 
wire u2__abc_52138_new_n9813_; 
wire u2__abc_52138_new_n9814_; 
wire u2__abc_52138_new_n9815_; 
wire u2__abc_52138_new_n9816_; 
wire u2__abc_52138_new_n9817_; 
wire u2__abc_52138_new_n9818_; 
wire u2__abc_52138_new_n9820_; 
wire u2__abc_52138_new_n9821_; 
wire u2__abc_52138_new_n9822_; 
wire u2__abc_52138_new_n9823_; 
wire u2__abc_52138_new_n9824_; 
wire u2__abc_52138_new_n9825_; 
wire u2__abc_52138_new_n9826_; 
wire u2__abc_52138_new_n9827_; 
wire u2__abc_52138_new_n9829_; 
wire u2__abc_52138_new_n9830_; 
wire u2__abc_52138_new_n9831_; 
wire u2__abc_52138_new_n9832_; 
wire u2__abc_52138_new_n9833_; 
wire u2__abc_52138_new_n9834_; 
wire u2__abc_52138_new_n9835_; 
wire u2__abc_52138_new_n9836_; 
wire u2__abc_52138_new_n9837_; 
wire u2__abc_52138_new_n9838_; 
wire u2__abc_52138_new_n9839_; 
wire u2__abc_52138_new_n9840_; 
wire u2__abc_52138_new_n9841_; 
wire u2__abc_52138_new_n9843_; 
wire u2__abc_52138_new_n9844_; 
wire u2__abc_52138_new_n9845_; 
wire u2__abc_52138_new_n9846_; 
wire u2__abc_52138_new_n9847_; 
wire u2__abc_52138_new_n9848_; 
wire u2__abc_52138_new_n9849_; 
wire u2__abc_52138_new_n9850_; 
wire u2__abc_52138_new_n9851_; 
wire u2__abc_52138_new_n9853_; 
wire u2__abc_52138_new_n9854_; 
wire u2__abc_52138_new_n9855_; 
wire u2__abc_52138_new_n9856_; 
wire u2__abc_52138_new_n9857_; 
wire u2__abc_52138_new_n9858_; 
wire u2__abc_52138_new_n9859_; 
wire u2__abc_52138_new_n9860_; 
wire u2__abc_52138_new_n9862_; 
wire u2__abc_52138_new_n9863_; 
wire u2__abc_52138_new_n9864_; 
wire u2__abc_52138_new_n9865_; 
wire u2__abc_52138_new_n9866_; 
wire u2__abc_52138_new_n9867_; 
wire u2__abc_52138_new_n9868_; 
wire u2__abc_52138_new_n9869_; 
wire u2__abc_52138_new_n9871_; 
wire u2__abc_52138_new_n9872_; 
wire u2__abc_52138_new_n9873_; 
wire u2__abc_52138_new_n9874_; 
wire u2__abc_52138_new_n9875_; 
wire u2__abc_52138_new_n9876_; 
wire u2__abc_52138_new_n9877_; 
wire u2__abc_52138_new_n9878_; 
wire u2__abc_52138_new_n9879_; 
wire u2__abc_52138_new_n9880_; 
wire u2__abc_52138_new_n9881_; 
wire u2__abc_52138_new_n9882_; 
wire u2__abc_52138_new_n9883_; 
wire u2__abc_52138_new_n9885_; 
wire u2__abc_52138_new_n9886_; 
wire u2__abc_52138_new_n9887_; 
wire u2__abc_52138_new_n9888_; 
wire u2__abc_52138_new_n9889_; 
wire u2__abc_52138_new_n9890_; 
wire u2__abc_52138_new_n9891_; 
wire u2__abc_52138_new_n9893_; 
wire u2__abc_52138_new_n9894_; 
wire u2__abc_52138_new_n9895_; 
wire u2__abc_52138_new_n9896_; 
wire u2__abc_52138_new_n9897_; 
wire u2__abc_52138_new_n9898_; 
wire u2__abc_52138_new_n9899_; 
wire u2__abc_52138_new_n9900_; 
wire u2__abc_52138_new_n9901_; 
wire u2__abc_52138_new_n9902_; 
wire u2__abc_52138_new_n9904_; 
wire u2__abc_52138_new_n9905_; 
wire u2__abc_52138_new_n9906_; 
wire u2__abc_52138_new_n9907_; 
wire u2__abc_52138_new_n9908_; 
wire u2__abc_52138_new_n9909_; 
wire u2__abc_52138_new_n9910_; 
wire u2__abc_52138_new_n9911_; 
wire u2__abc_52138_new_n9913_; 
wire u2__abc_52138_new_n9914_; 
wire u2__abc_52138_new_n9915_; 
wire u2__abc_52138_new_n9916_; 
wire u2__abc_52138_new_n9917_; 
wire u2__abc_52138_new_n9918_; 
wire u2__abc_52138_new_n9919_; 
wire u2__abc_52138_new_n9920_; 
wire u2__abc_52138_new_n9921_; 
wire u2__abc_52138_new_n9922_; 
wire u2__abc_52138_new_n9923_; 
wire u2__abc_52138_new_n9924_; 
wire u2__abc_52138_new_n9925_; 
wire u2__abc_52138_new_n9926_; 
wire u2__abc_52138_new_n9928_; 
wire u2__abc_52138_new_n9929_; 
wire u2__abc_52138_new_n9930_; 
wire u2__abc_52138_new_n9931_; 
wire u2__abc_52138_new_n9932_; 
wire u2__abc_52138_new_n9933_; 
wire u2__abc_52138_new_n9934_; 
wire u2__abc_52138_new_n9936_; 
wire u2__abc_52138_new_n9937_; 
wire u2__abc_52138_new_n9938_; 
wire u2__abc_52138_new_n9939_; 
wire u2__abc_52138_new_n9940_; 
wire u2__abc_52138_new_n9941_; 
wire u2__abc_52138_new_n9942_; 
wire u2__abc_52138_new_n9943_; 
wire u2__abc_52138_new_n9944_; 
wire u2__abc_52138_new_n9945_; 
wire u2__abc_52138_new_n9947_; 
wire u2__abc_52138_new_n9948_; 
wire u2__abc_52138_new_n9949_; 
wire u2__abc_52138_new_n9950_; 
wire u2__abc_52138_new_n9951_; 
wire u2__abc_52138_new_n9952_; 
wire u2__abc_52138_new_n9953_; 
wire u2__abc_52138_new_n9954_; 
wire u2__abc_52138_new_n9956_; 
wire u2__abc_52138_new_n9957_; 
wire u2__abc_52138_new_n9958_; 
wire u2__abc_52138_new_n9959_; 
wire u2__abc_52138_new_n9960_; 
wire u2__abc_52138_new_n9961_; 
wire u2__abc_52138_new_n9962_; 
wire u2__abc_52138_new_n9963_; 
wire u2__abc_52138_new_n9964_; 
wire u2__abc_52138_new_n9965_; 
wire u2__abc_52138_new_n9966_; 
wire u2__abc_52138_new_n9967_; 
wire u2__abc_52138_new_n9968_; 
wire u2__abc_52138_new_n9969_; 
wire u2__abc_52138_new_n9970_; 
wire u2__abc_52138_new_n9971_; 
wire u2__abc_52138_new_n9972_; 
wire u2__abc_52138_new_n9973_; 
wire u2__abc_52138_new_n9975_; 
wire u2__abc_52138_new_n9976_; 
wire u2__abc_52138_new_n9977_; 
wire u2__abc_52138_new_n9978_; 
wire u2__abc_52138_new_n9979_; 
wire u2__abc_52138_new_n9980_; 
wire u2__abc_52138_new_n9981_; 
wire u2__abc_52138_new_n9982_; 
wire u2__abc_52138_new_n9984_; 
wire u2__abc_52138_new_n9985_; 
wire u2__abc_52138_new_n9986_; 
wire u2__abc_52138_new_n9987_; 
wire u2__abc_52138_new_n9988_; 
wire u2__abc_52138_new_n9989_; 
wire u2__abc_52138_new_n9990_; 
wire u2__abc_52138_new_n9991_; 
wire u2__abc_52138_new_n9992_; 
wire u2__abc_52138_new_n9993_; 
wire u2__abc_52138_new_n9994_; 
wire u2__abc_52138_new_n9996_; 
wire u2__abc_52138_new_n9997_; 
wire u2__abc_52138_new_n9998_; 
wire u2__abc_52138_new_n9999_; 
wire u2_cnt_0_; 
wire u2_cnt_1_; 
wire u2_cnt_2_; 
wire u2_cnt_3_; 
wire u2_cnt_4_; 
wire u2_cnt_5_; 
wire u2_cnt_6_; 
wire u2_cnt_7_; 
wire u2_o_226_; 
wire u2_o_227_; 
wire u2_o_228_; 
wire u2_o_229_; 
wire u2_o_230_; 
wire u2_o_231_; 
wire u2_o_232_; 
wire u2_o_233_; 
wire u2_o_234_; 
wire u2_o_235_; 
wire u2_o_236_; 
wire u2_o_237_; 
wire u2_o_238_; 
wire u2_o_239_; 
wire u2_o_240_; 
wire u2_o_241_; 
wire u2_o_242_; 
wire u2_o_243_; 
wire u2_o_244_; 
wire u2_o_245_; 
wire u2_o_246_; 
wire u2_o_247_; 
wire u2_o_248_; 
wire u2_o_249_; 
wire u2_o_250_; 
wire u2_o_251_; 
wire u2_o_252_; 
wire u2_o_253_; 
wire u2_o_254_; 
wire u2_o_255_; 
wire u2_o_256_; 
wire u2_o_257_; 
wire u2_o_258_; 
wire u2_o_259_; 
wire u2_o_260_; 
wire u2_o_261_; 
wire u2_o_262_; 
wire u2_o_263_; 
wire u2_o_264_; 
wire u2_o_265_; 
wire u2_o_266_; 
wire u2_o_267_; 
wire u2_o_268_; 
wire u2_o_269_; 
wire u2_o_270_; 
wire u2_o_271_; 
wire u2_o_272_; 
wire u2_o_273_; 
wire u2_o_274_; 
wire u2_o_275_; 
wire u2_o_276_; 
wire u2_o_277_; 
wire u2_o_278_; 
wire u2_o_279_; 
wire u2_o_280_; 
wire u2_o_281_; 
wire u2_o_282_; 
wire u2_o_283_; 
wire u2_o_284_; 
wire u2_o_285_; 
wire u2_o_286_; 
wire u2_o_287_; 
wire u2_o_288_; 
wire u2_o_289_; 
wire u2_o_290_; 
wire u2_o_291_; 
wire u2_o_292_; 
wire u2_o_293_; 
wire u2_o_294_; 
wire u2_o_295_; 
wire u2_o_296_; 
wire u2_o_297_; 
wire u2_o_298_; 
wire u2_o_299_; 
wire u2_o_300_; 
wire u2_o_301_; 
wire u2_o_302_; 
wire u2_o_303_; 
wire u2_o_304_; 
wire u2_o_305_; 
wire u2_o_306_; 
wire u2_o_307_; 
wire u2_o_308_; 
wire u2_o_309_; 
wire u2_o_310_; 
wire u2_o_311_; 
wire u2_o_312_; 
wire u2_o_313_; 
wire u2_o_314_; 
wire u2_o_315_; 
wire u2_o_316_; 
wire u2_o_317_; 
wire u2_o_318_; 
wire u2_o_319_; 
wire u2_o_320_; 
wire u2_o_321_; 
wire u2_o_322_; 
wire u2_o_323_; 
wire u2_o_324_; 
wire u2_o_325_; 
wire u2_o_326_; 
wire u2_o_327_; 
wire u2_o_328_; 
wire u2_o_329_; 
wire u2_o_330_; 
wire u2_o_331_; 
wire u2_o_332_; 
wire u2_o_333_; 
wire u2_o_334_; 
wire u2_o_335_; 
wire u2_o_336_; 
wire u2_o_337_; 
wire u2_o_338_; 
wire u2_o_339_; 
wire u2_o_340_; 
wire u2_o_341_; 
wire u2_o_342_; 
wire u2_o_343_; 
wire u2_o_344_; 
wire u2_o_345_; 
wire u2_o_346_; 
wire u2_o_347_; 
wire u2_o_348_; 
wire u2_o_349_; 
wire u2_o_350_; 
wire u2_o_351_; 
wire u2_o_352_; 
wire u2_o_353_; 
wire u2_o_354_; 
wire u2_o_355_; 
wire u2_o_356_; 
wire u2_o_357_; 
wire u2_o_358_; 
wire u2_o_359_; 
wire u2_o_360_; 
wire u2_o_361_; 
wire u2_o_362_; 
wire u2_o_363_; 
wire u2_o_364_; 
wire u2_o_365_; 
wire u2_o_366_; 
wire u2_o_367_; 
wire u2_o_368_; 
wire u2_o_369_; 
wire u2_o_370_; 
wire u2_o_371_; 
wire u2_o_372_; 
wire u2_o_373_; 
wire u2_o_374_; 
wire u2_o_375_; 
wire u2_o_376_; 
wire u2_o_377_; 
wire u2_o_378_; 
wire u2_o_379_; 
wire u2_o_380_; 
wire u2_o_381_; 
wire u2_o_382_; 
wire u2_o_383_; 
wire u2_o_384_; 
wire u2_o_385_; 
wire u2_o_386_; 
wire u2_o_387_; 
wire u2_o_388_; 
wire u2_o_389_; 
wire u2_o_390_; 
wire u2_o_391_; 
wire u2_o_392_; 
wire u2_o_393_; 
wire u2_o_394_; 
wire u2_o_395_; 
wire u2_o_396_; 
wire u2_o_397_; 
wire u2_o_398_; 
wire u2_o_399_; 
wire u2_o_400_; 
wire u2_o_401_; 
wire u2_o_402_; 
wire u2_o_403_; 
wire u2_o_404_; 
wire u2_o_405_; 
wire u2_o_406_; 
wire u2_o_407_; 
wire u2_o_408_; 
wire u2_o_409_; 
wire u2_o_410_; 
wire u2_o_411_; 
wire u2_o_412_; 
wire u2_o_413_; 
wire u2_o_414_; 
wire u2_o_415_; 
wire u2_o_416_; 
wire u2_o_417_; 
wire u2_o_418_; 
wire u2_o_419_; 
wire u2_o_420_; 
wire u2_o_421_; 
wire u2_o_422_; 
wire u2_o_423_; 
wire u2_o_424_; 
wire u2_o_425_; 
wire u2_o_426_; 
wire u2_o_427_; 
wire u2_o_428_; 
wire u2_o_429_; 
wire u2_o_430_; 
wire u2_o_431_; 
wire u2_o_432_; 
wire u2_o_433_; 
wire u2_o_434_; 
wire u2_o_435_; 
wire u2_o_436_; 
wire u2_o_437_; 
wire u2_o_438_; 
wire u2_o_439_; 
wire u2_o_440_; 
wire u2_o_441_; 
wire u2_o_442_; 
wire u2_o_443_; 
wire u2_o_444_; 
wire u2_o_445_; 
wire u2_o_446_; 
wire u2_o_447_; 
wire u2_o_448_; 
wire u2_o_449_; 
wire u2_remHiShift_0_; 
wire u2_remHiShift_1_; 
wire u2_remHi_0_; 
wire u2_remHi_100_; 
wire u2_remHi_101_; 
wire u2_remHi_102_; 
wire u2_remHi_103_; 
wire u2_remHi_104_; 
wire u2_remHi_105_; 
wire u2_remHi_106_; 
wire u2_remHi_107_; 
wire u2_remHi_108_; 
wire u2_remHi_109_; 
wire u2_remHi_10_; 
wire u2_remHi_110_; 
wire u2_remHi_111_; 
wire u2_remHi_112_; 
wire u2_remHi_113_; 
wire u2_remHi_114_; 
wire u2_remHi_115_; 
wire u2_remHi_116_; 
wire u2_remHi_117_; 
wire u2_remHi_118_; 
wire u2_remHi_119_; 
wire u2_remHi_11_; 
wire u2_remHi_120_; 
wire u2_remHi_121_; 
wire u2_remHi_122_; 
wire u2_remHi_123_; 
wire u2_remHi_124_; 
wire u2_remHi_125_; 
wire u2_remHi_126_; 
wire u2_remHi_127_; 
wire u2_remHi_128_; 
wire u2_remHi_129_; 
wire u2_remHi_12_; 
wire u2_remHi_130_; 
wire u2_remHi_131_; 
wire u2_remHi_132_; 
wire u2_remHi_133_; 
wire u2_remHi_134_; 
wire u2_remHi_135_; 
wire u2_remHi_136_; 
wire u2_remHi_137_; 
wire u2_remHi_138_; 
wire u2_remHi_139_; 
wire u2_remHi_13_; 
wire u2_remHi_140_; 
wire u2_remHi_141_; 
wire u2_remHi_142_; 
wire u2_remHi_143_; 
wire u2_remHi_144_; 
wire u2_remHi_145_; 
wire u2_remHi_146_; 
wire u2_remHi_147_; 
wire u2_remHi_148_; 
wire u2_remHi_149_; 
wire u2_remHi_14_; 
wire u2_remHi_150_; 
wire u2_remHi_151_; 
wire u2_remHi_152_; 
wire u2_remHi_153_; 
wire u2_remHi_154_; 
wire u2_remHi_155_; 
wire u2_remHi_156_; 
wire u2_remHi_157_; 
wire u2_remHi_158_; 
wire u2_remHi_159_; 
wire u2_remHi_15_; 
wire u2_remHi_160_; 
wire u2_remHi_161_; 
wire u2_remHi_162_; 
wire u2_remHi_163_; 
wire u2_remHi_164_; 
wire u2_remHi_165_; 
wire u2_remHi_166_; 
wire u2_remHi_167_; 
wire u2_remHi_168_; 
wire u2_remHi_169_; 
wire u2_remHi_16_; 
wire u2_remHi_170_; 
wire u2_remHi_171_; 
wire u2_remHi_172_; 
wire u2_remHi_173_; 
wire u2_remHi_174_; 
wire u2_remHi_175_; 
wire u2_remHi_176_; 
wire u2_remHi_177_; 
wire u2_remHi_178_; 
wire u2_remHi_179_; 
wire u2_remHi_17_; 
wire u2_remHi_180_; 
wire u2_remHi_181_; 
wire u2_remHi_182_; 
wire u2_remHi_183_; 
wire u2_remHi_184_; 
wire u2_remHi_185_; 
wire u2_remHi_186_; 
wire u2_remHi_187_; 
wire u2_remHi_188_; 
wire u2_remHi_189_; 
wire u2_remHi_18_; 
wire u2_remHi_190_; 
wire u2_remHi_191_; 
wire u2_remHi_192_; 
wire u2_remHi_193_; 
wire u2_remHi_194_; 
wire u2_remHi_195_; 
wire u2_remHi_196_; 
wire u2_remHi_197_; 
wire u2_remHi_198_; 
wire u2_remHi_199_; 
wire u2_remHi_19_; 
wire u2_remHi_1_; 
wire u2_remHi_200_; 
wire u2_remHi_201_; 
wire u2_remHi_202_; 
wire u2_remHi_203_; 
wire u2_remHi_204_; 
wire u2_remHi_205_; 
wire u2_remHi_206_; 
wire u2_remHi_207_; 
wire u2_remHi_208_; 
wire u2_remHi_209_; 
wire u2_remHi_20_; 
wire u2_remHi_210_; 
wire u2_remHi_211_; 
wire u2_remHi_212_; 
wire u2_remHi_213_; 
wire u2_remHi_214_; 
wire u2_remHi_215_; 
wire u2_remHi_216_; 
wire u2_remHi_217_; 
wire u2_remHi_218_; 
wire u2_remHi_219_; 
wire u2_remHi_21_; 
wire u2_remHi_220_; 
wire u2_remHi_221_; 
wire u2_remHi_222_; 
wire u2_remHi_223_; 
wire u2_remHi_224_; 
wire u2_remHi_225_; 
wire u2_remHi_226_; 
wire u2_remHi_227_; 
wire u2_remHi_228_; 
wire u2_remHi_229_; 
wire u2_remHi_22_; 
wire u2_remHi_230_; 
wire u2_remHi_231_; 
wire u2_remHi_232_; 
wire u2_remHi_233_; 
wire u2_remHi_234_; 
wire u2_remHi_235_; 
wire u2_remHi_236_; 
wire u2_remHi_237_; 
wire u2_remHi_238_; 
wire u2_remHi_239_; 
wire u2_remHi_23_; 
wire u2_remHi_240_; 
wire u2_remHi_241_; 
wire u2_remHi_242_; 
wire u2_remHi_243_; 
wire u2_remHi_244_; 
wire u2_remHi_245_; 
wire u2_remHi_246_; 
wire u2_remHi_247_; 
wire u2_remHi_248_; 
wire u2_remHi_249_; 
wire u2_remHi_24_; 
wire u2_remHi_250_; 
wire u2_remHi_251_; 
wire u2_remHi_252_; 
wire u2_remHi_253_; 
wire u2_remHi_254_; 
wire u2_remHi_255_; 
wire u2_remHi_256_; 
wire u2_remHi_257_; 
wire u2_remHi_258_; 
wire u2_remHi_259_; 
wire u2_remHi_25_; 
wire u2_remHi_260_; 
wire u2_remHi_261_; 
wire u2_remHi_262_; 
wire u2_remHi_263_; 
wire u2_remHi_264_; 
wire u2_remHi_265_; 
wire u2_remHi_266_; 
wire u2_remHi_267_; 
wire u2_remHi_268_; 
wire u2_remHi_269_; 
wire u2_remHi_26_; 
wire u2_remHi_270_; 
wire u2_remHi_271_; 
wire u2_remHi_272_; 
wire u2_remHi_273_; 
wire u2_remHi_274_; 
wire u2_remHi_275_; 
wire u2_remHi_276_; 
wire u2_remHi_277_; 
wire u2_remHi_278_; 
wire u2_remHi_279_; 
wire u2_remHi_27_; 
wire u2_remHi_280_; 
wire u2_remHi_281_; 
wire u2_remHi_282_; 
wire u2_remHi_283_; 
wire u2_remHi_284_; 
wire u2_remHi_285_; 
wire u2_remHi_286_; 
wire u2_remHi_287_; 
wire u2_remHi_288_; 
wire u2_remHi_289_; 
wire u2_remHi_28_; 
wire u2_remHi_290_; 
wire u2_remHi_291_; 
wire u2_remHi_292_; 
wire u2_remHi_293_; 
wire u2_remHi_294_; 
wire u2_remHi_295_; 
wire u2_remHi_296_; 
wire u2_remHi_297_; 
wire u2_remHi_298_; 
wire u2_remHi_299_; 
wire u2_remHi_29_; 
wire u2_remHi_2_; 
wire u2_remHi_300_; 
wire u2_remHi_301_; 
wire u2_remHi_302_; 
wire u2_remHi_303_; 
wire u2_remHi_304_; 
wire u2_remHi_305_; 
wire u2_remHi_306_; 
wire u2_remHi_307_; 
wire u2_remHi_308_; 
wire u2_remHi_309_; 
wire u2_remHi_30_; 
wire u2_remHi_310_; 
wire u2_remHi_311_; 
wire u2_remHi_312_; 
wire u2_remHi_313_; 
wire u2_remHi_314_; 
wire u2_remHi_315_; 
wire u2_remHi_316_; 
wire u2_remHi_317_; 
wire u2_remHi_318_; 
wire u2_remHi_319_; 
wire u2_remHi_31_; 
wire u2_remHi_320_; 
wire u2_remHi_321_; 
wire u2_remHi_322_; 
wire u2_remHi_323_; 
wire u2_remHi_324_; 
wire u2_remHi_325_; 
wire u2_remHi_326_; 
wire u2_remHi_327_; 
wire u2_remHi_328_; 
wire u2_remHi_329_; 
wire u2_remHi_32_; 
wire u2_remHi_330_; 
wire u2_remHi_331_; 
wire u2_remHi_332_; 
wire u2_remHi_333_; 
wire u2_remHi_334_; 
wire u2_remHi_335_; 
wire u2_remHi_336_; 
wire u2_remHi_337_; 
wire u2_remHi_338_; 
wire u2_remHi_339_; 
wire u2_remHi_33_; 
wire u2_remHi_340_; 
wire u2_remHi_341_; 
wire u2_remHi_342_; 
wire u2_remHi_343_; 
wire u2_remHi_344_; 
wire u2_remHi_345_; 
wire u2_remHi_346_; 
wire u2_remHi_347_; 
wire u2_remHi_348_; 
wire u2_remHi_349_; 
wire u2_remHi_34_; 
wire u2_remHi_350_; 
wire u2_remHi_351_; 
wire u2_remHi_352_; 
wire u2_remHi_353_; 
wire u2_remHi_354_; 
wire u2_remHi_355_; 
wire u2_remHi_356_; 
wire u2_remHi_357_; 
wire u2_remHi_358_; 
wire u2_remHi_359_; 
wire u2_remHi_35_; 
wire u2_remHi_360_; 
wire u2_remHi_361_; 
wire u2_remHi_362_; 
wire u2_remHi_363_; 
wire u2_remHi_364_; 
wire u2_remHi_365_; 
wire u2_remHi_366_; 
wire u2_remHi_367_; 
wire u2_remHi_368_; 
wire u2_remHi_369_; 
wire u2_remHi_36_; 
wire u2_remHi_370_; 
wire u2_remHi_371_; 
wire u2_remHi_372_; 
wire u2_remHi_373_; 
wire u2_remHi_374_; 
wire u2_remHi_375_; 
wire u2_remHi_376_; 
wire u2_remHi_377_; 
wire u2_remHi_378_; 
wire u2_remHi_379_; 
wire u2_remHi_37_; 
wire u2_remHi_380_; 
wire u2_remHi_381_; 
wire u2_remHi_382_; 
wire u2_remHi_383_; 
wire u2_remHi_384_; 
wire u2_remHi_385_; 
wire u2_remHi_386_; 
wire u2_remHi_387_; 
wire u2_remHi_388_; 
wire u2_remHi_389_; 
wire u2_remHi_38_; 
wire u2_remHi_390_; 
wire u2_remHi_391_; 
wire u2_remHi_392_; 
wire u2_remHi_393_; 
wire u2_remHi_394_; 
wire u2_remHi_395_; 
wire u2_remHi_396_; 
wire u2_remHi_397_; 
wire u2_remHi_398_; 
wire u2_remHi_399_; 
wire u2_remHi_39_; 
wire u2_remHi_3_; 
wire u2_remHi_400_; 
wire u2_remHi_401_; 
wire u2_remHi_402_; 
wire u2_remHi_403_; 
wire u2_remHi_404_; 
wire u2_remHi_405_; 
wire u2_remHi_406_; 
wire u2_remHi_407_; 
wire u2_remHi_408_; 
wire u2_remHi_409_; 
wire u2_remHi_40_; 
wire u2_remHi_410_; 
wire u2_remHi_411_; 
wire u2_remHi_412_; 
wire u2_remHi_413_; 
wire u2_remHi_414_; 
wire u2_remHi_415_; 
wire u2_remHi_416_; 
wire u2_remHi_417_; 
wire u2_remHi_418_; 
wire u2_remHi_419_; 
wire u2_remHi_41_; 
wire u2_remHi_420_; 
wire u2_remHi_421_; 
wire u2_remHi_422_; 
wire u2_remHi_423_; 
wire u2_remHi_424_; 
wire u2_remHi_425_; 
wire u2_remHi_426_; 
wire u2_remHi_427_; 
wire u2_remHi_428_; 
wire u2_remHi_429_; 
wire u2_remHi_42_; 
wire u2_remHi_430_; 
wire u2_remHi_431_; 
wire u2_remHi_432_; 
wire u2_remHi_433_; 
wire u2_remHi_434_; 
wire u2_remHi_435_; 
wire u2_remHi_436_; 
wire u2_remHi_437_; 
wire u2_remHi_438_; 
wire u2_remHi_439_; 
wire u2_remHi_43_; 
wire u2_remHi_440_; 
wire u2_remHi_441_; 
wire u2_remHi_442_; 
wire u2_remHi_443_; 
wire u2_remHi_444_; 
wire u2_remHi_445_; 
wire u2_remHi_446_; 
wire u2_remHi_447_; 
wire u2_remHi_448_; 
wire u2_remHi_449_; 
wire u2_remHi_44_; 
wire u2_remHi_45_; 
wire u2_remHi_46_; 
wire u2_remHi_47_; 
wire u2_remHi_48_; 
wire u2_remHi_49_; 
wire u2_remHi_4_; 
wire u2_remHi_50_; 
wire u2_remHi_51_; 
wire u2_remHi_52_; 
wire u2_remHi_53_; 
wire u2_remHi_54_; 
wire u2_remHi_55_; 
wire u2_remHi_56_; 
wire u2_remHi_57_; 
wire u2_remHi_58_; 
wire u2_remHi_59_; 
wire u2_remHi_5_; 
wire u2_remHi_60_; 
wire u2_remHi_61_; 
wire u2_remHi_62_; 
wire u2_remHi_63_; 
wire u2_remHi_64_; 
wire u2_remHi_65_; 
wire u2_remHi_66_; 
wire u2_remHi_67_; 
wire u2_remHi_68_; 
wire u2_remHi_69_; 
wire u2_remHi_6_; 
wire u2_remHi_70_; 
wire u2_remHi_71_; 
wire u2_remHi_72_; 
wire u2_remHi_73_; 
wire u2_remHi_74_; 
wire u2_remHi_75_; 
wire u2_remHi_76_; 
wire u2_remHi_77_; 
wire u2_remHi_78_; 
wire u2_remHi_79_; 
wire u2_remHi_7_; 
wire u2_remHi_80_; 
wire u2_remHi_81_; 
wire u2_remHi_82_; 
wire u2_remHi_83_; 
wire u2_remHi_84_; 
wire u2_remHi_85_; 
wire u2_remHi_86_; 
wire u2_remHi_87_; 
wire u2_remHi_88_; 
wire u2_remHi_89_; 
wire u2_remHi_8_; 
wire u2_remHi_90_; 
wire u2_remHi_91_; 
wire u2_remHi_92_; 
wire u2_remHi_93_; 
wire u2_remHi_94_; 
wire u2_remHi_95_; 
wire u2_remHi_96_; 
wire u2_remHi_97_; 
wire u2_remHi_98_; 
wire u2_remHi_99_; 
wire u2_remHi_9_; 
wire u2_remLo_0_; 
wire u2_remLo_100_; 
wire u2_remLo_101_; 
wire u2_remLo_102_; 
wire u2_remLo_103_; 
wire u2_remLo_104_; 
wire u2_remLo_105_; 
wire u2_remLo_106_; 
wire u2_remLo_107_; 
wire u2_remLo_108_; 
wire u2_remLo_109_; 
wire u2_remLo_10_; 
wire u2_remLo_110_; 
wire u2_remLo_111_; 
wire u2_remLo_112_; 
wire u2_remLo_113_; 
wire u2_remLo_114_; 
wire u2_remLo_115_; 
wire u2_remLo_116_; 
wire u2_remLo_117_; 
wire u2_remLo_118_; 
wire u2_remLo_119_; 
wire u2_remLo_11_; 
wire u2_remLo_120_; 
wire u2_remLo_121_; 
wire u2_remLo_122_; 
wire u2_remLo_123_; 
wire u2_remLo_124_; 
wire u2_remLo_125_; 
wire u2_remLo_126_; 
wire u2_remLo_127_; 
wire u2_remLo_128_; 
wire u2_remLo_129_; 
wire u2_remLo_12_; 
wire u2_remLo_130_; 
wire u2_remLo_131_; 
wire u2_remLo_132_; 
wire u2_remLo_133_; 
wire u2_remLo_134_; 
wire u2_remLo_135_; 
wire u2_remLo_136_; 
wire u2_remLo_137_; 
wire u2_remLo_138_; 
wire u2_remLo_139_; 
wire u2_remLo_13_; 
wire u2_remLo_140_; 
wire u2_remLo_141_; 
wire u2_remLo_142_; 
wire u2_remLo_143_; 
wire u2_remLo_144_; 
wire u2_remLo_145_; 
wire u2_remLo_146_; 
wire u2_remLo_147_; 
wire u2_remLo_148_; 
wire u2_remLo_149_; 
wire u2_remLo_14_; 
wire u2_remLo_150_; 
wire u2_remLo_151_; 
wire u2_remLo_152_; 
wire u2_remLo_153_; 
wire u2_remLo_154_; 
wire u2_remLo_155_; 
wire u2_remLo_156_; 
wire u2_remLo_157_; 
wire u2_remLo_158_; 
wire u2_remLo_159_; 
wire u2_remLo_15_; 
wire u2_remLo_160_; 
wire u2_remLo_161_; 
wire u2_remLo_162_; 
wire u2_remLo_163_; 
wire u2_remLo_164_; 
wire u2_remLo_165_; 
wire u2_remLo_166_; 
wire u2_remLo_167_; 
wire u2_remLo_168_; 
wire u2_remLo_169_; 
wire u2_remLo_16_; 
wire u2_remLo_170_; 
wire u2_remLo_171_; 
wire u2_remLo_172_; 
wire u2_remLo_173_; 
wire u2_remLo_174_; 
wire u2_remLo_175_; 
wire u2_remLo_176_; 
wire u2_remLo_177_; 
wire u2_remLo_178_; 
wire u2_remLo_179_; 
wire u2_remLo_17_; 
wire u2_remLo_180_; 
wire u2_remLo_181_; 
wire u2_remLo_182_; 
wire u2_remLo_183_; 
wire u2_remLo_184_; 
wire u2_remLo_185_; 
wire u2_remLo_186_; 
wire u2_remLo_187_; 
wire u2_remLo_188_; 
wire u2_remLo_189_; 
wire u2_remLo_18_; 
wire u2_remLo_190_; 
wire u2_remLo_191_; 
wire u2_remLo_192_; 
wire u2_remLo_193_; 
wire u2_remLo_194_; 
wire u2_remLo_195_; 
wire u2_remLo_196_; 
wire u2_remLo_197_; 
wire u2_remLo_198_; 
wire u2_remLo_199_; 
wire u2_remLo_19_; 
wire u2_remLo_1_; 
wire u2_remLo_200_; 
wire u2_remLo_201_; 
wire u2_remLo_202_; 
wire u2_remLo_203_; 
wire u2_remLo_204_; 
wire u2_remLo_205_; 
wire u2_remLo_206_; 
wire u2_remLo_207_; 
wire u2_remLo_208_; 
wire u2_remLo_209_; 
wire u2_remLo_20_; 
wire u2_remLo_210_; 
wire u2_remLo_211_; 
wire u2_remLo_212_; 
wire u2_remLo_213_; 
wire u2_remLo_214_; 
wire u2_remLo_215_; 
wire u2_remLo_216_; 
wire u2_remLo_217_; 
wire u2_remLo_218_; 
wire u2_remLo_219_; 
wire u2_remLo_21_; 
wire u2_remLo_220_; 
wire u2_remLo_221_; 
wire u2_remLo_222_; 
wire u2_remLo_223_; 
wire u2_remLo_224_; 
wire u2_remLo_225_; 
wire u2_remLo_226_; 
wire u2_remLo_227_; 
wire u2_remLo_228_; 
wire u2_remLo_229_; 
wire u2_remLo_22_; 
wire u2_remLo_230_; 
wire u2_remLo_231_; 
wire u2_remLo_232_; 
wire u2_remLo_233_; 
wire u2_remLo_234_; 
wire u2_remLo_235_; 
wire u2_remLo_236_; 
wire u2_remLo_237_; 
wire u2_remLo_238_; 
wire u2_remLo_239_; 
wire u2_remLo_23_; 
wire u2_remLo_240_; 
wire u2_remLo_241_; 
wire u2_remLo_242_; 
wire u2_remLo_243_; 
wire u2_remLo_244_; 
wire u2_remLo_245_; 
wire u2_remLo_246_; 
wire u2_remLo_247_; 
wire u2_remLo_248_; 
wire u2_remLo_249_; 
wire u2_remLo_24_; 
wire u2_remLo_250_; 
wire u2_remLo_251_; 
wire u2_remLo_252_; 
wire u2_remLo_253_; 
wire u2_remLo_254_; 
wire u2_remLo_255_; 
wire u2_remLo_256_; 
wire u2_remLo_257_; 
wire u2_remLo_258_; 
wire u2_remLo_259_; 
wire u2_remLo_25_; 
wire u2_remLo_260_; 
wire u2_remLo_261_; 
wire u2_remLo_262_; 
wire u2_remLo_263_; 
wire u2_remLo_264_; 
wire u2_remLo_265_; 
wire u2_remLo_266_; 
wire u2_remLo_267_; 
wire u2_remLo_268_; 
wire u2_remLo_269_; 
wire u2_remLo_26_; 
wire u2_remLo_270_; 
wire u2_remLo_271_; 
wire u2_remLo_272_; 
wire u2_remLo_273_; 
wire u2_remLo_274_; 
wire u2_remLo_275_; 
wire u2_remLo_276_; 
wire u2_remLo_277_; 
wire u2_remLo_278_; 
wire u2_remLo_279_; 
wire u2_remLo_27_; 
wire u2_remLo_280_; 
wire u2_remLo_281_; 
wire u2_remLo_282_; 
wire u2_remLo_283_; 
wire u2_remLo_284_; 
wire u2_remLo_285_; 
wire u2_remLo_286_; 
wire u2_remLo_287_; 
wire u2_remLo_288_; 
wire u2_remLo_289_; 
wire u2_remLo_28_; 
wire u2_remLo_290_; 
wire u2_remLo_291_; 
wire u2_remLo_292_; 
wire u2_remLo_293_; 
wire u2_remLo_294_; 
wire u2_remLo_295_; 
wire u2_remLo_296_; 
wire u2_remLo_297_; 
wire u2_remLo_298_; 
wire u2_remLo_299_; 
wire u2_remLo_29_; 
wire u2_remLo_2_; 
wire u2_remLo_300_; 
wire u2_remLo_301_; 
wire u2_remLo_302_; 
wire u2_remLo_303_; 
wire u2_remLo_304_; 
wire u2_remLo_305_; 
wire u2_remLo_306_; 
wire u2_remLo_307_; 
wire u2_remLo_308_; 
wire u2_remLo_309_; 
wire u2_remLo_30_; 
wire u2_remLo_310_; 
wire u2_remLo_311_; 
wire u2_remLo_312_; 
wire u2_remLo_313_; 
wire u2_remLo_314_; 
wire u2_remLo_315_; 
wire u2_remLo_316_; 
wire u2_remLo_317_; 
wire u2_remLo_318_; 
wire u2_remLo_319_; 
wire u2_remLo_31_; 
wire u2_remLo_320_; 
wire u2_remLo_321_; 
wire u2_remLo_322_; 
wire u2_remLo_323_; 
wire u2_remLo_324_; 
wire u2_remLo_325_; 
wire u2_remLo_326_; 
wire u2_remLo_327_; 
wire u2_remLo_328_; 
wire u2_remLo_329_; 
wire u2_remLo_32_; 
wire u2_remLo_330_; 
wire u2_remLo_331_; 
wire u2_remLo_332_; 
wire u2_remLo_333_; 
wire u2_remLo_334_; 
wire u2_remLo_335_; 
wire u2_remLo_336_; 
wire u2_remLo_337_; 
wire u2_remLo_338_; 
wire u2_remLo_339_; 
wire u2_remLo_33_; 
wire u2_remLo_340_; 
wire u2_remLo_341_; 
wire u2_remLo_342_; 
wire u2_remLo_343_; 
wire u2_remLo_344_; 
wire u2_remLo_345_; 
wire u2_remLo_346_; 
wire u2_remLo_347_; 
wire u2_remLo_348_; 
wire u2_remLo_349_; 
wire u2_remLo_34_; 
wire u2_remLo_350_; 
wire u2_remLo_351_; 
wire u2_remLo_352_; 
wire u2_remLo_353_; 
wire u2_remLo_354_; 
wire u2_remLo_355_; 
wire u2_remLo_356_; 
wire u2_remLo_357_; 
wire u2_remLo_358_; 
wire u2_remLo_359_; 
wire u2_remLo_35_; 
wire u2_remLo_360_; 
wire u2_remLo_361_; 
wire u2_remLo_362_; 
wire u2_remLo_363_; 
wire u2_remLo_364_; 
wire u2_remLo_365_; 
wire u2_remLo_366_; 
wire u2_remLo_367_; 
wire u2_remLo_368_; 
wire u2_remLo_369_; 
wire u2_remLo_36_; 
wire u2_remLo_370_; 
wire u2_remLo_371_; 
wire u2_remLo_372_; 
wire u2_remLo_373_; 
wire u2_remLo_374_; 
wire u2_remLo_375_; 
wire u2_remLo_376_; 
wire u2_remLo_377_; 
wire u2_remLo_378_; 
wire u2_remLo_379_; 
wire u2_remLo_37_; 
wire u2_remLo_380_; 
wire u2_remLo_381_; 
wire u2_remLo_382_; 
wire u2_remLo_383_; 
wire u2_remLo_384_; 
wire u2_remLo_385_; 
wire u2_remLo_386_; 
wire u2_remLo_387_; 
wire u2_remLo_388_; 
wire u2_remLo_389_; 
wire u2_remLo_38_; 
wire u2_remLo_390_; 
wire u2_remLo_391_; 
wire u2_remLo_392_; 
wire u2_remLo_393_; 
wire u2_remLo_394_; 
wire u2_remLo_395_; 
wire u2_remLo_396_; 
wire u2_remLo_397_; 
wire u2_remLo_398_; 
wire u2_remLo_399_; 
wire u2_remLo_39_; 
wire u2_remLo_3_; 
wire u2_remLo_400_; 
wire u2_remLo_401_; 
wire u2_remLo_402_; 
wire u2_remLo_403_; 
wire u2_remLo_404_; 
wire u2_remLo_405_; 
wire u2_remLo_406_; 
wire u2_remLo_407_; 
wire u2_remLo_408_; 
wire u2_remLo_409_; 
wire u2_remLo_40_; 
wire u2_remLo_410_; 
wire u2_remLo_411_; 
wire u2_remLo_412_; 
wire u2_remLo_413_; 
wire u2_remLo_414_; 
wire u2_remLo_415_; 
wire u2_remLo_416_; 
wire u2_remLo_417_; 
wire u2_remLo_418_; 
wire u2_remLo_419_; 
wire u2_remLo_41_; 
wire u2_remLo_420_; 
wire u2_remLo_421_; 
wire u2_remLo_422_; 
wire u2_remLo_423_; 
wire u2_remLo_424_; 
wire u2_remLo_425_; 
wire u2_remLo_426_; 
wire u2_remLo_427_; 
wire u2_remLo_428_; 
wire u2_remLo_429_; 
wire u2_remLo_42_; 
wire u2_remLo_430_; 
wire u2_remLo_431_; 
wire u2_remLo_432_; 
wire u2_remLo_433_; 
wire u2_remLo_434_; 
wire u2_remLo_435_; 
wire u2_remLo_436_; 
wire u2_remLo_437_; 
wire u2_remLo_438_; 
wire u2_remLo_439_; 
wire u2_remLo_43_; 
wire u2_remLo_440_; 
wire u2_remLo_441_; 
wire u2_remLo_442_; 
wire u2_remLo_443_; 
wire u2_remLo_444_; 
wire u2_remLo_445_; 
wire u2_remLo_446_; 
wire u2_remLo_447_; 
wire u2_remLo_448_; 
wire u2_remLo_449_; 
wire u2_remLo_44_; 
wire u2_remLo_45_; 
wire u2_remLo_46_; 
wire u2_remLo_47_; 
wire u2_remLo_48_; 
wire u2_remLo_49_; 
wire u2_remLo_4_; 
wire u2_remLo_50_; 
wire u2_remLo_51_; 
wire u2_remLo_52_; 
wire u2_remLo_53_; 
wire u2_remLo_54_; 
wire u2_remLo_55_; 
wire u2_remLo_56_; 
wire u2_remLo_57_; 
wire u2_remLo_58_; 
wire u2_remLo_59_; 
wire u2_remLo_5_; 
wire u2_remLo_60_; 
wire u2_remLo_61_; 
wire u2_remLo_62_; 
wire u2_remLo_63_; 
wire u2_remLo_64_; 
wire u2_remLo_65_; 
wire u2_remLo_66_; 
wire u2_remLo_67_; 
wire u2_remLo_68_; 
wire u2_remLo_69_; 
wire u2_remLo_6_; 
wire u2_remLo_70_; 
wire u2_remLo_71_; 
wire u2_remLo_72_; 
wire u2_remLo_73_; 
wire u2_remLo_74_; 
wire u2_remLo_75_; 
wire u2_remLo_76_; 
wire u2_remLo_77_; 
wire u2_remLo_78_; 
wire u2_remLo_79_; 
wire u2_remLo_7_; 
wire u2_remLo_80_; 
wire u2_remLo_81_; 
wire u2_remLo_82_; 
wire u2_remLo_83_; 
wire u2_remLo_84_; 
wire u2_remLo_85_; 
wire u2_remLo_86_; 
wire u2_remLo_87_; 
wire u2_remLo_88_; 
wire u2_remLo_89_; 
wire u2_remLo_8_; 
wire u2_remLo_90_; 
wire u2_remLo_91_; 
wire u2_remLo_92_; 
wire u2_remLo_93_; 
wire u2_remLo_94_; 
wire u2_remLo_95_; 
wire u2_remLo_96_; 
wire u2_remLo_97_; 
wire u2_remLo_98_; 
wire u2_remLo_99_; 
wire u2_remLo_9_; 
wire u2_root_0_; 
wire u2_state_0_; 
wire u2_state_2_; 
AND2X2 AND2X2_1 ( .A(_abc_65734_new_n753_), .B(sqrto_0_), .Y(\o[36] ));
AND2X2 AND2X2_10 ( .A(_abc_65734_new_n753_), .B(sqrto_9_), .Y(\o[45] ));
AND2X2 AND2X2_100 ( .A(u2__abc_52138_new_n3345_), .B(u2__abc_52138_new_n3356_), .Y(u2__abc_52138_new_n3425_));
AND2X2 AND2X2_101 ( .A(u2__abc_52138_new_n3368_), .B(u2__abc_52138_new_n3379_), .Y(u2__abc_52138_new_n3426_));
AND2X2 AND2X2_102 ( .A(u2__abc_52138_new_n3560_), .B(u2__abc_52138_new_n3571_), .Y(u2__abc_52138_new_n3572_));
AND2X2 AND2X2_103 ( .A(u2__abc_52138_new_n3675_), .B(u2__abc_52138_new_n3686_), .Y(u2__abc_52138_new_n3687_));
AND2X2 AND2X2_104 ( .A(u2__abc_52138_new_n3750_), .B(u2__abc_52138_new_n3752_), .Y(u2__abc_52138_new_n3753_));
AND2X2 AND2X2_105 ( .A(u2__abc_52138_new_n3755_), .B(u2__abc_52138_new_n3757_), .Y(u2__abc_52138_new_n3758_));
AND2X2 AND2X2_106 ( .A(u2__abc_52138_new_n3771_), .B(u2__abc_52138_new_n3782_), .Y(u2__abc_52138_new_n3783_));
AND2X2 AND2X2_107 ( .A(u2__abc_52138_new_n3798_), .B(u2__abc_52138_new_n3800_), .Y(u2__abc_52138_new_n3801_));
AND2X2 AND2X2_108 ( .A(u2__abc_52138_new_n3842_), .B(u2__abc_52138_new_n3853_), .Y(u2__abc_52138_new_n3854_));
AND2X2 AND2X2_109 ( .A(u2__abc_52138_new_n3916_), .B(u2__abc_52138_new_n3775_), .Y(u2__abc_52138_new_n3917_));
AND2X2 AND2X2_11 ( .A(_abc_65734_new_n753_), .B(sqrto_10_), .Y(\o[46] ));
AND2X2 AND2X2_110 ( .A(u2__abc_52138_new_n3956_), .B(u2__abc_52138_new_n3611_), .Y(u2__abc_52138_new_n3957_));
AND2X2 AND2X2_111 ( .A(u2__abc_52138_new_n4091_), .B(u2__abc_52138_new_n4093_), .Y(u2__abc_52138_new_n4094_));
AND2X2 AND2X2_112 ( .A(u2__abc_52138_new_n4089_), .B(u2__abc_52138_new_n4094_), .Y(u2__abc_52138_new_n4095_));
AND2X2 AND2X2_113 ( .A(u2__abc_52138_new_n4095_), .B(u2__abc_52138_new_n4084_), .Y(u2__abc_52138_new_n4096_));
AND2X2 AND2X2_114 ( .A(u2__abc_52138_new_n4234_), .B(u2__abc_52138_new_n4236_), .Y(u2__abc_52138_new_n4237_));
AND2X2 AND2X2_115 ( .A(u2__abc_52138_new_n4341_), .B(u2__abc_52138_new_n4352_), .Y(u2__abc_52138_new_n4353_));
AND2X2 AND2X2_116 ( .A(u2__abc_52138_new_n4376_), .B(u2__abc_52138_new_n4363_), .Y(u2__abc_52138_new_n4377_));
AND2X2 AND2X2_117 ( .A(u2__abc_52138_new_n4546_), .B(u2__abc_52138_new_n4535_), .Y(u2__abc_52138_new_n4547_));
AND2X2 AND2X2_118 ( .A(u2__abc_52138_new_n4558_), .B(u2__abc_52138_new_n4569_), .Y(u2__abc_52138_new_n4570_));
AND2X2 AND2X2_119 ( .A(u2__abc_52138_new_n4629_), .B(u2__abc_52138_new_n4640_), .Y(u2__abc_52138_new_n4641_));
AND2X2 AND2X2_12 ( .A(_abc_65734_new_n753_), .B(sqrto_11_), .Y(\o[47] ));
AND2X2 AND2X2_120 ( .A(u2__abc_52138_new_n4643_), .B(u2__abc_52138_new_n4645_), .Y(u2__abc_52138_new_n4646_));
AND2X2 AND2X2_121 ( .A(u2__abc_52138_new_n4676_), .B(u2__abc_52138_new_n4687_), .Y(u2__abc_52138_new_n4688_));
AND2X2 AND2X2_122 ( .A(u2__abc_52138_new_n4699_), .B(u2__abc_52138_new_n4710_), .Y(u2__abc_52138_new_n4711_));
AND2X2 AND2X2_123 ( .A(u2__abc_52138_new_n4745_), .B(u2__abc_52138_new_n4747_), .Y(u2__abc_52138_new_n4748_));
AND2X2 AND2X2_124 ( .A(u2__abc_52138_new_n4803_), .B(u2__abc_52138_new_n4650_), .Y(u2__abc_52138_new_n4804_));
AND2X2 AND2X2_125 ( .A(u2__abc_52138_new_n4924_), .B(u2__abc_52138_new_n4923_), .Y(u2__abc_52138_new_n4925_));
AND2X2 AND2X2_126 ( .A(u2__abc_52138_new_n4036_), .B(u2__abc_52138_new_n4047_), .Y(u2__abc_52138_new_n4971_));
AND2X2 AND2X2_127 ( .A(u2__abc_52138_new_n5054_), .B(u2__abc_52138_new_n5055_), .Y(u2__abc_52138_new_n5056_));
AND2X2 AND2X2_128 ( .A(u2__abc_52138_new_n5083_), .B(u2__abc_52138_new_n5085_), .Y(u2__abc_52138_new_n5086_));
AND2X2 AND2X2_129 ( .A(u2__abc_52138_new_n5097_), .B(u2__abc_52138_new_n5099_), .Y(u2__abc_52138_new_n5100_));
AND2X2 AND2X2_13 ( .A(_abc_65734_new_n753_), .B(sqrto_12_), .Y(\o[48] ));
AND2X2 AND2X2_130 ( .A(u2__abc_52138_new_n5108_), .B(u2__abc_52138_new_n5110_), .Y(u2__abc_52138_new_n5111_));
AND2X2 AND2X2_131 ( .A(u2__abc_52138_new_n5181_), .B(u2__abc_52138_new_n5090_), .Y(u2__abc_52138_new_n5182_));
AND2X2 AND2X2_132 ( .A(u2__abc_52138_new_n5184_), .B(u2__abc_52138_new_n5186_), .Y(u2__abc_52138_new_n5187_));
AND2X2 AND2X2_133 ( .A(u2__abc_52138_new_n5250_), .B(u2__abc_52138_new_n5252_), .Y(u2__abc_52138_new_n5253_));
AND2X2 AND2X2_134 ( .A(u2__abc_52138_new_n5263_), .B(u2__abc_52138_new_n5264_), .Y(u2__abc_52138_new_n5265_));
AND2X2 AND2X2_135 ( .A(u2__abc_52138_new_n5280_), .B(u2__abc_52138_new_n5282_), .Y(u2__abc_52138_new_n5283_));
AND2X2 AND2X2_136 ( .A(u2__abc_52138_new_n5319_), .B(u2__abc_52138_new_n5296_), .Y(u2__abc_52138_new_n5320_));
AND2X2 AND2X2_137 ( .A(u2__abc_52138_new_n5334_), .B(u2__abc_52138_new_n5336_), .Y(u2__abc_52138_new_n5337_));
AND2X2 AND2X2_138 ( .A(u2__abc_52138_new_n5347_), .B(u2__abc_52138_new_n5349_), .Y(u2__abc_52138_new_n5350_));
AND2X2 AND2X2_139 ( .A(u2__abc_52138_new_n5461_), .B(u2__abc_52138_new_n5463_), .Y(u2__abc_52138_new_n5464_));
AND2X2 AND2X2_14 ( .A(_abc_65734_new_n753_), .B(sqrto_13_), .Y(\o[49] ));
AND2X2 AND2X2_140 ( .A(u2__abc_52138_new_n5591_), .B(u2__abc_52138_new_n5585_), .Y(u2__abc_52138_new_n5775_));
AND2X2 AND2X2_141 ( .A(u2__abc_52138_new_n5317_), .B(u2__abc_52138_new_n5311_), .Y(u2__abc_52138_new_n5855_));
AND2X2 AND2X2_142 ( .A(u2__abc_52138_new_n6322_), .B(u2__abc_52138_new_n6323_), .Y(u2__abc_52138_new_n6324_));
AND2X2 AND2X2_143 ( .A(u2__abc_52138_new_n6330_), .B(u2__abc_52138_new_n6184_), .Y(u2__abc_52138_new_n6331_));
AND2X2 AND2X2_144 ( .A(u2__abc_52138_new_n6398_), .B(u2__abc_52138_new_n6083_), .Y(u2__abc_52138_new_n6399_));
AND2X2 AND2X2_145 ( .A(u2__abc_52138_new_n6413_), .B(u2__abc_52138_new_n6417_), .Y(u2__abc_52138_new_n6418_));
AND2X2 AND2X2_146 ( .A(u2__abc_52138_new_n3689_), .B(u2__abc_52138_new_n3869_), .Y(u2__abc_52138_new_n6451_));
AND2X2 AND2X2_147 ( .A(u2__abc_52138_new_n6478_), .B(u2__abc_52138_new_n6472_), .Y(u2__abc_52138_new_n6479_));
AND2X2 AND2X2_148 ( .A(u2__abc_52138_new_n3594_), .B(u2__abc_52138_new_n3572_), .Y(u2__abc_52138_new_n6483_));
AND2X2 AND2X2_149 ( .A(u2__abc_52138_new_n3712_), .B(u2__abc_52138_new_n3736_), .Y(u2__abc_52138_new_n6484_));
AND2X2 AND2X2_15 ( .A(_abc_65734_new_n753_), .B(sqrto_14_), .Y(\o[50] ));
AND2X2 AND2X2_150 ( .A(u2__abc_52138_new_n6493_), .B(u2__abc_52138_new_n6494_), .Y(u2__abc_52138_new_n6495_));
AND2X2 AND2X2_151 ( .A(u2__abc_52138_new_n6666_), .B(u2__abc_52138_new_n6671_), .Y(u2__abc_52138_new_n6672_));
AND2X2 AND2X2_152 ( .A(u2__abc_52138_new_n6872_), .B(u2__abc_52138_new_n3387_), .Y(u2__abc_52138_new_n6874_));
AND2X2 AND2X2_153 ( .A(u2__abc_52138_new_n3370_), .B(u2__abc_52138_new_n3375_), .Y(u2__abc_52138_new_n6989_));
AND2X2 AND2X2_154 ( .A(u2__abc_52138_new_n7161_), .B(u2__abc_52138_new_n7162_), .Y(u2__abc_52138_new_n7163_));
AND2X2 AND2X2_155 ( .A(u2__abc_52138_new_n7098_), .B(u2__abc_52138_new_n3286_), .Y(u2__abc_52138_new_n7177_));
AND2X2 AND2X2_156 ( .A(u2__abc_52138_new_n7188_), .B(u2__abc_52138_new_n3833_), .Y(u2__abc_52138_new_n7195_));
AND2X2 AND2X2_157 ( .A(u2__abc_52138_new_n7288_), .B(u2__abc_52138_new_n3895_), .Y(u2__abc_52138_new_n7289_));
AND2X2 AND2X2_158 ( .A(u2__abc_52138_new_n7631_), .B(u2__abc_52138_new_n3618_), .Y(u2__abc_52138_new_n7674_));
AND2X2 AND2X2_159 ( .A(u2__abc_52138_new_n3631_), .B(u2__abc_52138_new_n3633_), .Y(u2__abc_52138_new_n7684_));
AND2X2 AND2X2_16 ( .A(_abc_65734_new_n753_), .B(sqrto_15_), .Y(\o[51] ));
AND2X2 AND2X2_160 ( .A(u2__abc_52138_new_n7789_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__118_));
AND2X2 AND2X2_161 ( .A(u2__abc_52138_new_n7806_), .B(u2__abc_52138_new_n3579_), .Y(u2__abc_52138_new_n7807_));
AND2X2 AND2X2_162 ( .A(u2__abc_52138_new_n7811_), .B(u2__abc_52138_new_n7812_), .Y(u2__abc_52138_new_n7813_));
AND2X2 AND2X2_163 ( .A(u2__abc_52138_new_n7859_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__124_));
AND2X2 AND2X2_164 ( .A(u2__abc_52138_new_n3596_), .B(u2__abc_52138_new_n3689_), .Y(u2__abc_52138_new_n7892_));
AND2X2 AND2X2_165 ( .A(u2__abc_52138_new_n8151_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__150_));
AND2X2 AND2X2_166 ( .A(u2__abc_52138_new_n8218_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__156_));
AND2X2 AND2X2_167 ( .A(u2__abc_52138_new_n8230_), .B(u2__abc_52138_new_n8229_), .Y(u2__abc_52138_new_n8249_));
AND2X2 AND2X2_168 ( .A(u2__abc_52138_new_n8347_), .B(u2__abc_52138_new_n8348_), .Y(u2__abc_52138_new_n8349_));
AND2X2 AND2X2_169 ( .A(u2__abc_52138_new_n8390_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__172_));
AND2X2 AND2X2_17 ( .A(_abc_65734_new_n753_), .B(sqrto_16_), .Y(\o[52] ));
AND2X2 AND2X2_170 ( .A(u2__abc_52138_new_n8433_), .B(u2__abc_52138_new_n8431_), .Y(u2__abc_52138_new_n8434_));
AND2X2 AND2X2_171 ( .A(u2__abc_52138_new_n8460_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__178_));
AND2X2 AND2X2_172 ( .A(u2__abc_52138_new_n8481_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__180_));
AND2X2 AND2X2_173 ( .A(u2__abc_52138_new_n8520_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__184_));
AND2X2 AND2X2_174 ( .A(u2__abc_52138_new_n8674_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__198_));
AND2X2 AND2X2_175 ( .A(u2__abc_52138_new_n8738_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__204_));
AND2X2 AND2X2_176 ( .A(u2__abc_52138_new_n8750_), .B(u2__abc_52138_new_n4904_), .Y(u2__abc_52138_new_n8770_));
AND2X2 AND2X2_177 ( .A(u2__abc_52138_new_n8769_), .B(u2__abc_52138_new_n8772_), .Y(u2__abc_52138_new_n8773_));
AND2X2 AND2X2_178 ( .A(u2__abc_52138_new_n8603_), .B(u2__abc_52138_new_n4379_), .Y(u2__abc_52138_new_n8775_));
AND2X2 AND2X2_179 ( .A(u2__abc_52138_new_n8782_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__208_));
AND2X2 AND2X2_18 ( .A(_abc_65734_new_n753_), .B(sqrto_17_), .Y(\o[53] ));
AND2X2 AND2X2_180 ( .A(u2__abc_52138_new_n8823_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__212_));
AND2X2 AND2X2_181 ( .A(u2__abc_52138_new_n4268_), .B(u2__abc_52138_new_n4273_), .Y(u2__abc_52138_new_n8851_));
AND2X2 AND2X2_182 ( .A(u2__abc_52138_new_n8863_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__216_));
AND2X2 AND2X2_183 ( .A(u2__abc_52138_new_n8990_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__228_));
AND2X2 AND2X2_184 ( .A(u2__abc_52138_new_n4179_), .B(u2__abc_52138_new_n9001_), .Y(u2__abc_52138_new_n9019_));
AND2X2 AND2X2_185 ( .A(u2__abc_52138_new_n9031_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__232_));
AND2X2 AND2X2_186 ( .A(u2__abc_52138_new_n9190_), .B(u2__abc_52138_new_n9189_), .Y(u2__abc_52138_new_n9191_));
AND2X2 AND2X2_187 ( .A(u2__abc_52138_new_n9253_), .B(u2__abc_52138_new_n7779_), .Y(u2__0remHi_451_0__254_));
AND2X2 AND2X2_188 ( .A(u2__abc_52138_new_n4098_), .B(u2__abc_52138_new_n4192_), .Y(u2__abc_52138_new_n9267_));
AND2X2 AND2X2_189 ( .A(u2__abc_52138_new_n9270_), .B(u2__abc_52138_new_n9272_), .Y(u2__abc_52138_new_n9273_));
AND2X2 AND2X2_19 ( .A(_abc_65734_new_n753_), .B(sqrto_18_), .Y(\o[54] ));
AND2X2 AND2X2_190 ( .A(u2__abc_52138_new_n5689_), .B(u2__abc_52138_new_n5693_), .Y(u2__abc_52138_new_n9286_));
AND2X2 AND2X2_191 ( .A(u2__abc_52138_new_n9342_), .B(u2__abc_52138_new_n5713_), .Y(u2__abc_52138_new_n9343_));
AND2X2 AND2X2_192 ( .A(u2__abc_52138_new_n9401_), .B(u2__abc_52138_new_n5655_), .Y(u2__abc_52138_new_n9402_));
AND2X2 AND2X2_193 ( .A(u2__abc_52138_new_n9444_), .B(u2__abc_52138_new_n5638_), .Y(u2__abc_52138_new_n9613_));
AND2X2 AND2X2_194 ( .A(u2__abc_52138_new_n9278_), .B(u2__abc_52138_new_n5734_), .Y(u2__abc_52138_new_n9620_));
AND2X2 AND2X2_195 ( .A(u2__abc_52138_new_n10313_), .B(u2__abc_52138_new_n5181_), .Y(u2__abc_52138_new_n10485_));
AND2X2 AND2X2_196 ( .A(u2__abc_52138_new_n10589_), .B(u2__abc_52138_new_n10590_), .Y(u2__abc_52138_new_n10591_));
AND2X2 AND2X2_197 ( .A(u2__abc_52138_new_n11248_), .B(u2__abc_52138_new_n11245_), .Y(u2__abc_52138_new_n11249_));
AND2X2 AND2X2_198 ( .A(u2__abc_52138_new_n11379_), .B(u2__abc_52138_new_n11380_), .Y(u2__0cnt_7_0__0_));
AND2X2 AND2X2_199 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_31_), .Y(u2__abc_52138_new_n11513_));
AND2X2 AND2X2_2 ( .A(_abc_65734_new_n753_), .B(sqrto_1_), .Y(\o[37] ));
AND2X2 AND2X2_20 ( .A(_abc_65734_new_n753_), .B(sqrto_19_), .Y(\o[55] ));
AND2X2 AND2X2_200 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_34_), .Y(u2__abc_52138_new_n11525_));
AND2X2 AND2X2_201 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_46_), .Y(u2__abc_52138_new_n11564_));
AND2X2 AND2X2_202 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_65_), .Y(u2__abc_52138_new_n11624_));
AND2X2 AND2X2_203 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_74_), .Y(u2__abc_52138_new_n11654_));
AND2X2 AND2X2_204 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_97_), .Y(u2__abc_52138_new_n11729_));
AND2X2 AND2X2_205 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_114_), .Y(u2__abc_52138_new_n11783_));
AND2X2 AND2X2_206 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_129_), .Y(u2__abc_52138_new_n11831_));
AND2X2 AND2X2_207 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_161_), .Y(u2__abc_52138_new_n11931_));
AND2X2 AND2X2_208 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_193_), .Y(u2__abc_52138_new_n12031_));
AND2X2 AND2X2_209 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_202_), .Y(u2__abc_52138_new_n12061_));
AND2X2 AND2X2_21 ( .A(_abc_65734_new_n753_), .B(sqrto_20_), .Y(\o[56] ));
AND2X2 AND2X2_210 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_225_), .Y(u2__abc_52138_new_n12134_));
AND2X2 AND2X2_211 ( .A(u2__abc_52138_new_n11509_), .B(u2_remLo_226_), .Y(u2__abc_52138_new_n12140_));
AND2X2 AND2X2_212 ( .A(u2__abc_52138_new_n12823_), .B(u2__abc_52138_new_n3077_), .Y(u2__abc_52138_new_n12824_));
AND2X2 AND2X2_213 ( .A(u2__abc_52138_new_n4122_), .B(u2__abc_52138_new_n4144_), .Y(u2__abc_52138_new_n13019_));
AND2X2 AND2X2_214 ( .A(u2__abc_52138_new_n4972_), .B(u2__abc_52138_new_n4024_), .Y(u2__abc_52138_new_n13024_));
AND2X2 AND2X2_215 ( .A(u2__abc_52138_new_n5755_), .B(u2__abc_52138_new_n5780_), .Y(u2__abc_52138_new_n13032_));
AND2X2 AND2X2_216 ( .A(u2__abc_52138_new_n5807_), .B(u2__abc_52138_new_n5833_), .Y(u2__abc_52138_new_n13033_));
AND2X2 AND2X2_217 ( .A(u2__abc_52138_new_n5901_), .B(u2__abc_52138_new_n5939_), .Y(u2__abc_52138_new_n13036_));
AND2X2 AND2X2_22 ( .A(_abc_65734_new_n753_), .B(sqrto_21_), .Y(\o[57] ));
AND2X2 AND2X2_23 ( .A(_abc_65734_new_n753_), .B(sqrto_22_), .Y(\o[58] ));
AND2X2 AND2X2_24 ( .A(_abc_65734_new_n753_), .B(sqrto_23_), .Y(\o[59] ));
AND2X2 AND2X2_25 ( .A(_abc_65734_new_n753_), .B(sqrto_24_), .Y(\o[60] ));
AND2X2 AND2X2_26 ( .A(_abc_65734_new_n753_), .B(sqrto_25_), .Y(\o[61] ));
AND2X2 AND2X2_27 ( .A(_abc_65734_new_n753_), .B(sqrto_26_), .Y(\o[62] ));
AND2X2 AND2X2_28 ( .A(_abc_65734_new_n753_), .B(sqrto_27_), .Y(\o[63] ));
AND2X2 AND2X2_29 ( .A(_abc_65734_new_n753_), .B(sqrto_28_), .Y(\o[64] ));
AND2X2 AND2X2_3 ( .A(_abc_65734_new_n753_), .B(sqrto_2_), .Y(\o[38] ));
AND2X2 AND2X2_30 ( .A(_abc_65734_new_n753_), .B(sqrto_29_), .Y(\o[65] ));
AND2X2 AND2X2_31 ( .A(_abc_65734_new_n753_), .B(sqrto_30_), .Y(\o[66] ));
AND2X2 AND2X2_32 ( .A(_abc_65734_new_n753_), .B(sqrto_31_), .Y(\o[67] ));
AND2X2 AND2X2_33 ( .A(_abc_65734_new_n753_), .B(sqrto_32_), .Y(\o[68] ));
AND2X2 AND2X2_34 ( .A(_abc_65734_new_n753_), .B(sqrto_33_), .Y(\o[69] ));
AND2X2 AND2X2_35 ( .A(_abc_65734_new_n753_), .B(sqrto_34_), .Y(\o[70] ));
AND2X2 AND2X2_36 ( .A(_abc_65734_new_n753_), .B(sqrto_35_), .Y(\o[71] ));
AND2X2 AND2X2_37 ( .A(_abc_65734_new_n753_), .B(sqrto_36_), .Y(\o[72] ));
AND2X2 AND2X2_38 ( .A(_abc_65734_new_n753_), .B(sqrto_37_), .Y(\o[73] ));
AND2X2 AND2X2_39 ( .A(_abc_65734_new_n753_), .B(sqrto_38_), .Y(\o[74] ));
AND2X2 AND2X2_4 ( .A(_abc_65734_new_n753_), .B(sqrto_3_), .Y(\o[39] ));
AND2X2 AND2X2_40 ( .A(_abc_65734_new_n753_), .B(sqrto_39_), .Y(\o[75] ));
AND2X2 AND2X2_41 ( .A(_abc_65734_new_n753_), .B(sqrto_40_), .Y(\o[76] ));
AND2X2 AND2X2_42 ( .A(_abc_65734_new_n753_), .B(sqrto_41_), .Y(\o[77] ));
AND2X2 AND2X2_43 ( .A(_abc_65734_new_n753_), .B(sqrto_42_), .Y(\o[78] ));
AND2X2 AND2X2_44 ( .A(_abc_65734_new_n753_), .B(sqrto_43_), .Y(\o[79] ));
AND2X2 AND2X2_45 ( .A(_abc_65734_new_n753_), .B(sqrto_44_), .Y(\o[80] ));
AND2X2 AND2X2_46 ( .A(_abc_65734_new_n753_), .B(sqrto_45_), .Y(\o[81] ));
AND2X2 AND2X2_47 ( .A(_abc_65734_new_n753_), .B(sqrto_46_), .Y(\o[82] ));
AND2X2 AND2X2_48 ( .A(_abc_65734_new_n753_), .B(sqrto_47_), .Y(\o[83] ));
AND2X2 AND2X2_49 ( .A(_abc_65734_new_n753_), .B(sqrto_48_), .Y(\o[84] ));
AND2X2 AND2X2_5 ( .A(_abc_65734_new_n753_), .B(sqrto_4_), .Y(\o[40] ));
AND2X2 AND2X2_50 ( .A(_abc_65734_new_n753_), .B(sqrto_49_), .Y(\o[85] ));
AND2X2 AND2X2_51 ( .A(_abc_65734_new_n753_), .B(sqrto_50_), .Y(\o[86] ));
AND2X2 AND2X2_52 ( .A(_abc_65734_new_n753_), .B(sqrto_51_), .Y(\o[87] ));
AND2X2 AND2X2_53 ( .A(_abc_65734_new_n753_), .B(sqrto_52_), .Y(\o[88] ));
AND2X2 AND2X2_54 ( .A(_abc_65734_new_n753_), .B(sqrto_53_), .Y(\o[89] ));
AND2X2 AND2X2_55 ( .A(_abc_65734_new_n753_), .B(sqrto_54_), .Y(\o[90] ));
AND2X2 AND2X2_56 ( .A(_abc_65734_new_n753_), .B(sqrto_55_), .Y(\o[91] ));
AND2X2 AND2X2_57 ( .A(_abc_65734_new_n753_), .B(sqrto_56_), .Y(\o[92] ));
AND2X2 AND2X2_58 ( .A(_abc_65734_new_n753_), .B(sqrto_57_), .Y(\o[93] ));
AND2X2 AND2X2_59 ( .A(_abc_65734_new_n753_), .B(sqrto_58_), .Y(\o[94] ));
AND2X2 AND2X2_6 ( .A(_abc_65734_new_n753_), .B(sqrto_5_), .Y(\o[41] ));
AND2X2 AND2X2_60 ( .A(_abc_65734_new_n753_), .B(sqrto_59_), .Y(\o[95] ));
AND2X2 AND2X2_61 ( .A(_abc_65734_new_n753_), .B(sqrto_60_), .Y(\o[96] ));
AND2X2 AND2X2_62 ( .A(_abc_65734_new_n753_), .B(sqrto_61_), .Y(\o[97] ));
AND2X2 AND2X2_63 ( .A(_abc_65734_new_n753_), .B(sqrto_62_), .Y(\o[98] ));
AND2X2 AND2X2_64 ( .A(_abc_65734_new_n753_), .B(sqrto_63_), .Y(\o[99] ));
AND2X2 AND2X2_65 ( .A(_abc_65734_new_n753_), .B(sqrto_64_), .Y(\o[100] ));
AND2X2 AND2X2_66 ( .A(_abc_65734_new_n753_), .B(sqrto_65_), .Y(\o[101] ));
AND2X2 AND2X2_67 ( .A(_abc_65734_new_n753_), .B(sqrto_66_), .Y(\o[102] ));
AND2X2 AND2X2_68 ( .A(_abc_65734_new_n753_), .B(sqrto_67_), .Y(\o[103] ));
AND2X2 AND2X2_69 ( .A(_abc_65734_new_n753_), .B(sqrto_68_), .Y(\o[104] ));
AND2X2 AND2X2_7 ( .A(_abc_65734_new_n753_), .B(sqrto_6_), .Y(\o[42] ));
AND2X2 AND2X2_70 ( .A(_abc_65734_new_n753_), .B(sqrto_69_), .Y(\o[105] ));
AND2X2 AND2X2_71 ( .A(_abc_65734_new_n753_), .B(sqrto_70_), .Y(\o[106] ));
AND2X2 AND2X2_72 ( .A(_abc_65734_new_n753_), .B(sqrto_71_), .Y(\o[107] ));
AND2X2 AND2X2_73 ( .A(_abc_65734_new_n753_), .B(sqrto_72_), .Y(\o[108] ));
AND2X2 AND2X2_74 ( .A(_abc_65734_new_n753_), .B(sqrto_73_), .Y(\o[109] ));
AND2X2 AND2X2_75 ( .A(_abc_65734_new_n753_), .B(sqrto_74_), .Y(\o[110] ));
AND2X2 AND2X2_76 ( .A(_abc_65734_new_n753_), .B(sqrto_75_), .Y(\o[111] ));
AND2X2 AND2X2_77 ( .A(_abc_65734_new_n753_), .B(sqrto_189_), .Y(\o[225] ));
AND2X2 AND2X2_78 ( .A(\a[112] ), .B(\a[113] ), .Y(_abc_65734_new_n1452_));
AND2X2 AND2X2_79 ( .A(\a[114] ), .B(\a[115] ), .Y(_abc_65734_new_n1470_));
AND2X2 AND2X2_8 ( .A(_abc_65734_new_n753_), .B(sqrto_7_), .Y(\o[43] ));
AND2X2 AND2X2_80 ( .A(_abc_65734_new_n1526_), .B(_abc_65734_new_n1525_), .Y(_abc_65734_new_n1529_));
AND2X2 AND2X2_81 ( .A(_abc_65734_new_n1537_), .B(_abc_65734_new_n1536_), .Y(_abc_65734_new_n1540_));
AND2X2 AND2X2_82 ( .A(_abc_65734_new_n1560_), .B(_abc_65734_new_n1557_), .Y(_abc_65734_new_n1561_));
AND2X2 AND2X2_83 ( .A(_abc_65734_new_n1580_), .B(\a[122] ), .Y(_abc_65734_new_n1581_));
AND2X2 AND2X2_84 ( .A(aNan), .B(\a[127] ), .Y(\o[241] ));
AND2X2 AND2X2_85 ( .A(\a[113] ), .B(\a[114] ), .Y(u1__abc_51895_new_n160_));
AND2X2 AND2X2_86 ( .A(u1__abc_51895_new_n297_), .B(u1__abc_51895_new_n328_), .Y(u1__abc_51895_new_n329_));
AND2X2 AND2X2_87 ( .A(u2_cnt_5_), .B(u2_cnt_6_), .Y(u2__abc_52138_new_n2969_));
AND2X2 AND2X2_88 ( .A(u2__abc_52138_new_n3007_), .B(u2__abc_52138_new_n3012_), .Y(u2__abc_52138_new_n3013_));
AND2X2 AND2X2_89 ( .A(u2__abc_52138_new_n3023_), .B(u2__abc_52138_new_n3025_), .Y(u2__abc_52138_new_n3026_));
AND2X2 AND2X2_9 ( .A(_abc_65734_new_n753_), .B(sqrto_8_), .Y(\o[44] ));
AND2X2 AND2X2_90 ( .A(u2__abc_52138_new_n3028_), .B(u2__abc_52138_new_n3030_), .Y(u2__abc_52138_new_n3031_));
AND2X2 AND2X2_91 ( .A(u2__abc_52138_new_n3041_), .B(u2__abc_52138_new_n3043_), .Y(u2__abc_52138_new_n3044_));
AND2X2 AND2X2_92 ( .A(u2__abc_52138_new_n3046_), .B(u2__abc_52138_new_n3048_), .Y(u2__abc_52138_new_n3049_));
AND2X2 AND2X2_93 ( .A(u2__abc_52138_new_n3098_), .B(u2__abc_52138_new_n3038_), .Y(u2__abc_52138_new_n3099_));
AND2X2 AND2X2_94 ( .A(u2__abc_52138_new_n3169_), .B(u2__abc_52138_new_n3180_), .Y(u2__abc_52138_new_n3181_));
AND2X2 AND2X2_95 ( .A(u2__abc_52138_new_n3145_), .B(u2__abc_52138_new_n3156_), .Y(u2__abc_52138_new_n3218_));
AND2X2 AND2X2_96 ( .A(u2__abc_52138_new_n3113_), .B(u2__abc_52138_new_n3115_), .Y(u2__abc_52138_new_n3219_));
AND2X2 AND2X2_97 ( .A(u2__abc_52138_new_n3118_), .B(u2__abc_52138_new_n3120_), .Y(u2__abc_52138_new_n3220_));
AND2X2 AND2X2_98 ( .A(u2__abc_52138_new_n3321_), .B(u2__abc_52138_new_n3332_), .Y(u2__abc_52138_new_n3333_));
AND2X2 AND2X2_99 ( .A(u2__abc_52138_new_n3413_), .B(u2__abc_52138_new_n3415_), .Y(u2__abc_52138_new_n3416_));
AOI21X1 AOI21X1_1 ( .A(\a[114] ), .B(_abc_65734_new_n1461_), .C(_abc_65734_new_n1457_), .Y(_abc_65734_new_n1466_));
AOI21X1 AOI21X1_10 ( .A(u2__abc_52138_new_n3094_), .B(u2__abc_52138_new_n3041_), .C(u2__abc_52138_new_n3093_), .Y(u2__abc_52138_new_n3095_));
AOI21X1 AOI21X1_100 ( .A(u2__abc_52138_new_n5738_), .B(u2__abc_52138_new_n5700_), .C(u2__abc_52138_new_n5705_), .Y(u2__abc_52138_new_n5739_));
AOI21X1 AOI21X1_1000 ( .A(u2__abc_52138_new_n9982_), .B(u2__abc_52138_new_n9975_), .C(rst), .Y(u2__0remHi_451_0__321_));
AOI21X1 AOI21X1_1001 ( .A(u2__abc_52138_new_n5356_), .B(u2__abc_52138_new_n9988_), .C(u2__abc_52138_new_n9989_), .Y(u2__abc_52138_new_n9990_));
AOI21X1 AOI21X1_1002 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n9992_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9993_));
AOI21X1 AOI21X1_1003 ( .A(u2__abc_52138_new_n9994_), .B(u2__abc_52138_new_n9984_), .C(rst), .Y(u2__0remHi_451_0__322_));
AOI21X1 AOI21X1_1004 ( .A(u2__abc_52138_new_n5361_), .B(u2__abc_52138_new_n9998_), .C(u2__abc_52138_new_n9999_), .Y(u2__abc_52138_new_n10000_));
AOI21X1 AOI21X1_1005 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5335_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10002_));
AOI21X1 AOI21X1_1006 ( .A(u2__abc_52138_new_n10003_), .B(u2__abc_52138_new_n9996_), .C(rst), .Y(u2__0remHi_451_0__323_));
AOI21X1 AOI21X1_1007 ( .A(u2__abc_52138_new_n5361_), .B(u2__abc_52138_new_n5353_), .C(u2__abc_52138_new_n5358_), .Y(u2__abc_52138_new_n10006_));
AOI21X1 AOI21X1_1008 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5323_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10015_));
AOI21X1 AOI21X1_1009 ( .A(u2__abc_52138_new_n10016_), .B(u2__abc_52138_new_n10005_), .C(rst), .Y(u2__0remHi_451_0__324_));
AOI21X1 AOI21X1_101 ( .A(u2__abc_52138_new_n5718_), .B(u2__abc_52138_new_n5712_), .C(u2__abc_52138_new_n5717_), .Y(u2__abc_52138_new_n5743_));
AOI21X1 AOI21X1_1010 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5328_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10023_));
AOI21X1 AOI21X1_1011 ( .A(u2__abc_52138_new_n10024_), .B(u2__abc_52138_new_n10018_), .C(rst), .Y(u2__0remHi_451_0__325_));
AOI21X1 AOI21X1_1012 ( .A(u2__abc_52138_new_n5325_), .B(u2__abc_52138_new_n10029_), .C(u2__abc_52138_new_n10030_), .Y(u2__abc_52138_new_n10031_));
AOI21X1 AOI21X1_1013 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5276_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10033_));
AOI21X1 AOI21X1_1014 ( .A(u2__abc_52138_new_n10034_), .B(u2__abc_52138_new_n10026_), .C(rst), .Y(u2__0remHi_451_0__326_));
AOI21X1 AOI21X1_1015 ( .A(u2__abc_52138_new_n5330_), .B(u2__abc_52138_new_n10038_), .C(u2__abc_52138_new_n10039_), .Y(u2__abc_52138_new_n10040_));
AOI21X1 AOI21X1_1016 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5279_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10042_));
AOI21X1 AOI21X1_1017 ( .A(u2__abc_52138_new_n10043_), .B(u2__abc_52138_new_n10036_), .C(rst), .Y(u2__0remHi_451_0__327_));
AOI21X1 AOI21X1_1018 ( .A(u2__abc_52138_new_n5330_), .B(u2__abc_52138_new_n5324_), .C(u2__abc_52138_new_n5329_), .Y(u2__abc_52138_new_n10048_));
AOI21X1 AOI21X1_1019 ( .A(u2__abc_52138_new_n5278_), .B(u2__abc_52138_new_n10052_), .C(u2__abc_52138_new_n10053_), .Y(u2__abc_52138_new_n10054_));
AOI21X1 AOI21X1_102 ( .A(u2__abc_52138_new_n5740_), .B(u2__abc_52138_new_n5731_), .C(u2__abc_52138_new_n5744_), .Y(u2__abc_52138_new_n5745_));
AOI21X1 AOI21X1_1020 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5285_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10056_));
AOI21X1 AOI21X1_1021 ( .A(u2__abc_52138_new_n10057_), .B(u2__abc_52138_new_n10045_), .C(rst), .Y(u2__0remHi_451_0__328_));
AOI21X1 AOI21X1_1022 ( .A(u2__abc_52138_new_n5283_), .B(u2__abc_52138_new_n10062_), .C(u2__abc_52138_new_n10063_), .Y(u2__abc_52138_new_n10064_));
AOI21X1 AOI21X1_1023 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5290_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10066_));
AOI21X1 AOI21X1_1024 ( .A(u2__abc_52138_new_n10067_), .B(u2__abc_52138_new_n10059_), .C(rst), .Y(u2__0remHi_451_0__329_));
AOI21X1 AOI21X1_1025 ( .A(u2__abc_52138_new_n5289_), .B(u2__abc_52138_new_n10072_), .C(u2__abc_52138_new_n10073_), .Y(u2__abc_52138_new_n10074_));
AOI21X1 AOI21X1_1026 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5308_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10076_));
AOI21X1 AOI21X1_1027 ( .A(u2__abc_52138_new_n10077_), .B(u2__abc_52138_new_n10069_), .C(rst), .Y(u2__0remHi_451_0__330_));
AOI21X1 AOI21X1_1028 ( .A(u2__abc_52138_new_n5294_), .B(u2__abc_52138_new_n10081_), .C(u2__abc_52138_new_n10082_), .Y(u2__abc_52138_new_n10083_));
AOI21X1 AOI21X1_1029 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5313_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10085_));
AOI21X1 AOI21X1_103 ( .A(u2__abc_52138_new_n5683_), .B(u2__abc_52138_new_n5675_), .C(u2__abc_52138_new_n5680_), .Y(u2__abc_52138_new_n5747_));
AOI21X1 AOI21X1_1030 ( .A(u2__abc_52138_new_n10086_), .B(u2__abc_52138_new_n10079_), .C(rst), .Y(u2__0remHi_451_0__331_));
AOI21X1 AOI21X1_1031 ( .A(u2__abc_52138_new_n5294_), .B(u2__abc_52138_new_n5286_), .C(u2__abc_52138_new_n5291_), .Y(u2__abc_52138_new_n10089_));
AOI21X1 AOI21X1_1032 ( .A(u2__abc_52138_new_n10052_), .B(u2__abc_52138_new_n5296_), .C(u2__abc_52138_new_n10090_), .Y(u2__abc_52138_new_n10091_));
AOI21X1 AOI21X1_1033 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5297_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10098_));
AOI21X1 AOI21X1_1034 ( .A(u2__abc_52138_new_n10099_), .B(u2__abc_52138_new_n10088_), .C(rst), .Y(u2__0remHi_451_0__332_));
AOI21X1 AOI21X1_1035 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5302_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10107_));
AOI21X1 AOI21X1_1036 ( .A(u2__abc_52138_new_n10108_), .B(u2__abc_52138_new_n10101_), .C(rst), .Y(u2__0remHi_451_0__333_));
AOI21X1 AOI21X1_1037 ( .A(u2__abc_52138_new_n5301_), .B(u2__abc_52138_new_n10114_), .C(u2__abc_52138_new_n10115_), .Y(u2__abc_52138_new_n10116_));
AOI21X1 AOI21X1_1038 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5874_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10118_));
AOI21X1 AOI21X1_1039 ( .A(u2__abc_52138_new_n10119_), .B(u2__abc_52138_new_n10110_), .C(rst), .Y(u2__0remHi_451_0__334_));
AOI21X1 AOI21X1_104 ( .A(u2__abc_52138_new_n5672_), .B(u2__abc_52138_new_n5666_), .C(u2__abc_52138_new_n5671_), .Y(u2__abc_52138_new_n5748_));
AOI21X1 AOI21X1_1040 ( .A(u2__abc_52138_new_n5306_), .B(u2__abc_52138_new_n10123_), .C(u2__abc_52138_new_n10124_), .Y(u2__abc_52138_new_n10125_));
AOI21X1 AOI21X1_1041 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5244_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10127_));
AOI21X1 AOI21X1_1042 ( .A(u2__abc_52138_new_n10128_), .B(u2__abc_52138_new_n10121_), .C(rst), .Y(u2__0remHi_451_0__335_));
AOI21X1 AOI21X1_1043 ( .A(u2__abc_52138_new_n10090_), .B(u2__abc_52138_new_n5319_), .C(u2__abc_52138_new_n5303_), .Y(u2__abc_52138_new_n10134_));
AOI21X1 AOI21X1_1044 ( .A(u2__abc_52138_new_n10131_), .B(u2__abc_52138_new_n5320_), .C(u2__abc_52138_new_n10135_), .Y(u2__abc_52138_new_n10136_));
AOI21X1 AOI21X1_1045 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5229_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10143_));
AOI21X1 AOI21X1_1046 ( .A(u2__abc_52138_new_n10144_), .B(u2__abc_52138_new_n10130_), .C(rst), .Y(u2__0remHi_451_0__336_));
AOI21X1 AOI21X1_1047 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5234_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10151_));
AOI21X1 AOI21X1_1048 ( .A(u2__abc_52138_new_n10152_), .B(u2__abc_52138_new_n10146_), .C(rst), .Y(u2__0remHi_451_0__337_));
AOI21X1 AOI21X1_1049 ( .A(u2__abc_52138_new_n5233_), .B(u2__abc_52138_new_n10157_), .C(u2__abc_52138_new_n10158_), .Y(u2__abc_52138_new_n10159_));
AOI21X1 AOI21X1_105 ( .A(u2__abc_52138_new_n5649_), .B(u2__abc_52138_new_n5641_), .C(u2__abc_52138_new_n5646_), .Y(u2__abc_52138_new_n5751_));
AOI21X1 AOI21X1_1050 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5261_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10161_));
AOI21X1 AOI21X1_1051 ( .A(u2__abc_52138_new_n10162_), .B(u2__abc_52138_new_n10154_), .C(rst), .Y(u2__0remHi_451_0__338_));
AOI21X1 AOI21X1_1052 ( .A(u2__abc_52138_new_n5238_), .B(u2__abc_52138_new_n10166_), .C(u2__abc_52138_new_n10167_), .Y(u2__abc_52138_new_n10168_));
AOI21X1 AOI21X1_1053 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5266_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10170_));
AOI21X1 AOI21X1_1054 ( .A(u2__abc_52138_new_n10171_), .B(u2__abc_52138_new_n10164_), .C(rst), .Y(u2__0remHi_451_0__339_));
AOI21X1 AOI21X1_1055 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5251_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10186_));
AOI21X1 AOI21X1_1056 ( .A(u2__abc_52138_new_n10187_), .B(u2__abc_52138_new_n10173_), .C(rst), .Y(u2__0remHi_451_0__340_));
AOI21X1 AOI21X1_1057 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5254_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10194_));
AOI21X1 AOI21X1_1058 ( .A(u2__abc_52138_new_n10195_), .B(u2__abc_52138_new_n10189_), .C(rst), .Y(u2__0remHi_451_0__341_));
AOI21X1 AOI21X1_1059 ( .A(u2__abc_52138_new_n5253_), .B(u2__abc_52138_new_n10200_), .C(u2__abc_52138_new_n10201_), .Y(u2__abc_52138_new_n10202_));
AOI21X1 AOI21X1_106 ( .A(u2__abc_52138_new_n5660_), .B(u2__abc_52138_new_n5654_), .C(u2__abc_52138_new_n5659_), .Y(u2__abc_52138_new_n5752_));
AOI21X1 AOI21X1_1060 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5195_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10204_));
AOI21X1 AOI21X1_1061 ( .A(u2__abc_52138_new_n10205_), .B(u2__abc_52138_new_n10197_), .C(rst), .Y(u2__0remHi_451_0__342_));
AOI21X1 AOI21X1_1062 ( .A(u2__abc_52138_new_n5258_), .B(u2__abc_52138_new_n10209_), .C(u2__abc_52138_new_n10210_), .Y(u2__abc_52138_new_n10211_));
AOI21X1 AOI21X1_1063 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5200_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10213_));
AOI21X1 AOI21X1_1064 ( .A(u2__abc_52138_new_n10214_), .B(u2__abc_52138_new_n10207_), .C(rst), .Y(u2__0remHi_451_0__343_));
AOI21X1 AOI21X1_1065 ( .A(u2__abc_52138_new_n10217_), .B(u2__abc_52138_new_n10198_), .C(u2__abc_52138_new_n10219_), .Y(u2__abc_52138_new_n10220_));
AOI21X1 AOI21X1_1066 ( .A(u2__abc_52138_new_n10137_), .B(u2__abc_52138_new_n5272_), .C(u2__abc_52138_new_n10221_), .Y(u2__abc_52138_new_n10222_));
AOI21X1 AOI21X1_1067 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5185_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10229_));
AOI21X1 AOI21X1_1068 ( .A(u2__abc_52138_new_n10230_), .B(u2__abc_52138_new_n10216_), .C(rst), .Y(u2__0remHi_451_0__344_));
AOI21X1 AOI21X1_1069 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5188_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10238_));
AOI21X1 AOI21X1_107 ( .A(u2__abc_52138_new_n5604_), .B(u2__abc_52138_new_n5598_), .C(u2__abc_52138_new_n5603_), .Y(u2__abc_52138_new_n5758_));
AOI21X1 AOI21X1_1070 ( .A(u2__abc_52138_new_n10239_), .B(u2__abc_52138_new_n10232_), .C(rst), .Y(u2__0remHi_451_0__345_));
AOI21X1 AOI21X1_1071 ( .A(u2__abc_52138_new_n5187_), .B(u2__abc_52138_new_n10245_), .C(u2__abc_52138_new_n10246_), .Y(u2__abc_52138_new_n10247_));
AOI21X1 AOI21X1_1072 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5216_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10249_));
AOI21X1 AOI21X1_1073 ( .A(u2__abc_52138_new_n10250_), .B(u2__abc_52138_new_n10241_), .C(rst), .Y(u2__0remHi_451_0__346_));
AOI21X1 AOI21X1_1074 ( .A(u2__abc_52138_new_n5192_), .B(u2__abc_52138_new_n10254_), .C(u2__abc_52138_new_n10255_), .Y(u2__abc_52138_new_n10256_));
AOI21X1 AOI21X1_1075 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5221_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10258_));
AOI21X1 AOI21X1_1076 ( .A(u2__abc_52138_new_n10259_), .B(u2__abc_52138_new_n10252_), .C(rst), .Y(u2__0remHi_451_0__347_));
AOI21X1 AOI21X1_1077 ( .A(u2__abc_52138_new_n5862_), .B(u2__abc_52138_new_n10263_), .C(u2__abc_52138_new_n5189_), .Y(u2__abc_52138_new_n10264_));
AOI21X1 AOI21X1_1078 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5208_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10273_));
AOI21X1 AOI21X1_1079 ( .A(u2__abc_52138_new_n10274_), .B(u2__abc_52138_new_n10261_), .C(rst), .Y(u2__0remHi_451_0__348_));
AOI21X1 AOI21X1_108 ( .A(u2__abc_52138_new_n5627_), .B(u2__abc_52138_new_n5621_), .C(u2__abc_52138_new_n5626_), .Y(u2__abc_52138_new_n5760_));
AOI21X1 AOI21X1_1080 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5210_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10281_));
AOI21X1 AOI21X1_1081 ( .A(u2__abc_52138_new_n10282_), .B(u2__abc_52138_new_n10276_), .C(rst), .Y(u2__0remHi_451_0__349_));
AOI21X1 AOI21X1_1082 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5145_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10293_));
AOI21X1 AOI21X1_1083 ( .A(u2__abc_52138_new_n10294_), .B(u2__abc_52138_new_n10284_), .C(rst), .Y(u2__0remHi_451_0__350_));
AOI21X1 AOI21X1_1084 ( .A(u2__abc_52138_new_n5214_), .B(u2__abc_52138_new_n10297_), .C(u2__abc_52138_new_n10298_), .Y(u2__abc_52138_new_n10299_));
AOI21X1 AOI21X1_1085 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5150_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10301_));
AOI21X1 AOI21X1_1086 ( .A(u2__abc_52138_new_n10302_), .B(u2__abc_52138_new_n10296_), .C(rst), .Y(u2__0remHi_451_0__351_));
AOI21X1 AOI21X1_1087 ( .A(u2__abc_52138_new_n10221_), .B(u2__abc_52138_new_n5228_), .C(u2__abc_52138_new_n10308_), .Y(u2__abc_52138_new_n10309_));
AOI21X1 AOI21X1_1088 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5134_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10319_));
AOI21X1 AOI21X1_1089 ( .A(u2__abc_52138_new_n10320_), .B(u2__abc_52138_new_n10304_), .C(rst), .Y(u2__0remHi_451_0__352_));
AOI21X1 AOI21X1_109 ( .A(u2__abc_52138_new_n5759_), .B(u2__abc_52138_new_n5636_), .C(u2__abc_52138_new_n5765_), .Y(u2__abc_52138_new_n5766_));
AOI21X1 AOI21X1_1090 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5139_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10327_));
AOI21X1 AOI21X1_1091 ( .A(u2__abc_52138_new_n10328_), .B(u2__abc_52138_new_n10322_), .C(rst), .Y(u2__0remHi_451_0__353_));
AOI21X1 AOI21X1_1092 ( .A(u2__abc_52138_new_n5138_), .B(u2__abc_52138_new_n10333_), .C(u2__abc_52138_new_n10334_), .Y(u2__abc_52138_new_n10335_));
AOI21X1 AOI21X1_1093 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5168_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10337_));
AOI21X1 AOI21X1_1094 ( .A(u2__abc_52138_new_n10338_), .B(u2__abc_52138_new_n10330_), .C(rst), .Y(u2__0remHi_451_0__354_));
AOI21X1 AOI21X1_1095 ( .A(u2__abc_52138_new_n5143_), .B(u2__abc_52138_new_n10342_), .C(u2__abc_52138_new_n10343_), .Y(u2__abc_52138_new_n10344_));
AOI21X1 AOI21X1_1096 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5173_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10346_));
AOI21X1 AOI21X1_1097 ( .A(u2__abc_52138_new_n10347_), .B(u2__abc_52138_new_n10340_), .C(rst), .Y(u2__0remHi_451_0__355_));
AOI21X1 AOI21X1_1098 ( .A(u2__abc_52138_new_n10313_), .B(u2__abc_52138_new_n5156_), .C(u2__abc_52138_new_n10353_), .Y(u2__abc_52138_new_n10354_));
AOI21X1 AOI21X1_1099 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5157_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10361_));
AOI21X1 AOI21X1_11 ( .A(u2__abc_52138_new_n3103_), .B(u2__abc_52138_new_n3020_), .C(u2__abc_52138_new_n3104_), .Y(u2__abc_52138_new_n3105_));
AOI21X1 AOI21X1_110 ( .A(u2__abc_52138_new_n5770_), .B(u2__abc_52138_new_n5551_), .C(u2__abc_52138_new_n5556_), .Y(u2__abc_52138_new_n5771_));
AOI21X1 AOI21X1_1100 ( .A(u2__abc_52138_new_n10362_), .B(u2__abc_52138_new_n10349_), .C(rst), .Y(u2__0remHi_451_0__356_));
AOI21X1 AOI21X1_1101 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5162_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10370_));
AOI21X1 AOI21X1_1102 ( .A(u2__abc_52138_new_n10371_), .B(u2__abc_52138_new_n10364_), .C(rst), .Y(u2__0remHi_451_0__357_));
AOI21X1 AOI21X1_1103 ( .A(u2__abc_52138_new_n5161_), .B(u2__abc_52138_new_n10377_), .C(u2__abc_52138_new_n10378_), .Y(u2__abc_52138_new_n10379_));
AOI21X1 AOI21X1_1104 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5093_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10381_));
AOI21X1 AOI21X1_1105 ( .A(u2__abc_52138_new_n10382_), .B(u2__abc_52138_new_n10373_), .C(rst), .Y(u2__0remHi_451_0__358_));
AOI21X1 AOI21X1_1106 ( .A(u2__abc_52138_new_n5166_), .B(u2__abc_52138_new_n10386_), .C(u2__abc_52138_new_n10387_), .Y(u2__abc_52138_new_n10388_));
AOI21X1 AOI21X1_1107 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5096_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10390_));
AOI21X1 AOI21X1_1108 ( .A(u2__abc_52138_new_n10391_), .B(u2__abc_52138_new_n10384_), .C(rst), .Y(u2__0remHi_451_0__359_));
AOI21X1 AOI21X1_1109 ( .A(u2__abc_52138_new_n5166_), .B(u2__abc_52138_new_n5158_), .C(u2__abc_52138_new_n5163_), .Y(u2__abc_52138_new_n10395_));
AOI21X1 AOI21X1_111 ( .A(u2__abc_52138_new_n5534_), .B(u2__abc_52138_new_n5528_), .C(u2__abc_52138_new_n5533_), .Y(u2__abc_52138_new_n5791_));
AOI21X1 AOI21X1_1110 ( .A(u2__abc_52138_new_n10353_), .B(u2__abc_52138_new_n5179_), .C(u2__abc_52138_new_n10396_), .Y(u2__abc_52138_new_n10397_));
AOI21X1 AOI21X1_1111 ( .A(u2__abc_52138_new_n10312_), .B(u2__abc_52138_new_n10311_), .C(u2__abc_52138_new_n5180_), .Y(u2__abc_52138_new_n10399_));
AOI21X1 AOI21X1_1112 ( .A(u2__abc_52138_new_n5095_), .B(u2__abc_52138_new_n10401_), .C(u2__abc_52138_new_n10402_), .Y(u2__abc_52138_new_n10403_));
AOI21X1 AOI21X1_1113 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5102_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10405_));
AOI21X1 AOI21X1_1114 ( .A(u2__abc_52138_new_n10406_), .B(u2__abc_52138_new_n10393_), .C(rst), .Y(u2__0remHi_451_0__360_));
AOI21X1 AOI21X1_1115 ( .A(u2__abc_52138_new_n5100_), .B(u2__abc_52138_new_n10410_), .C(u2__abc_52138_new_n10411_), .Y(u2__abc_52138_new_n10412_));
AOI21X1 AOI21X1_1116 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5109_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10414_));
AOI21X1 AOI21X1_1117 ( .A(u2__abc_52138_new_n10415_), .B(u2__abc_52138_new_n10408_), .C(rst), .Y(u2__0remHi_451_0__361_));
AOI21X1 AOI21X1_1118 ( .A(u2__abc_52138_new_n5106_), .B(u2__abc_52138_new_n10421_), .C(u2__abc_52138_new_n10422_), .Y(u2__abc_52138_new_n10423_));
AOI21X1 AOI21X1_1119 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n10425_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10426_));
AOI21X1 AOI21X1_112 ( .A(u2__abc_52138_new_n5786_), .B(u2__abc_52138_new_n5543_), .C(u2__abc_52138_new_n5792_), .Y(u2__abc_52138_new_n5793_));
AOI21X1 AOI21X1_1120 ( .A(u2__abc_52138_new_n10427_), .B(u2__abc_52138_new_n10417_), .C(rst), .Y(u2__0remHi_451_0__362_));
AOI21X1 AOI21X1_1121 ( .A(u2__abc_52138_new_n5111_), .B(u2__abc_52138_new_n10431_), .C(u2__abc_52138_new_n10432_), .Y(u2__abc_52138_new_n10433_));
AOI21X1 AOI21X1_1122 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5126_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10435_));
AOI21X1 AOI21X1_1123 ( .A(u2__abc_52138_new_n10436_), .B(u2__abc_52138_new_n10429_), .C(rst), .Y(u2__0remHi_451_0__363_));
AOI21X1 AOI21X1_1124 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5114_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10449_));
AOI21X1 AOI21X1_1125 ( .A(u2__abc_52138_new_n10450_), .B(u2__abc_52138_new_n10438_), .C(rst), .Y(u2__0remHi_451_0__364_));
AOI21X1 AOI21X1_1126 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5119_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10457_));
AOI21X1 AOI21X1_1127 ( .A(u2__abc_52138_new_n10458_), .B(u2__abc_52138_new_n10452_), .C(rst), .Y(u2__0remHi_451_0__365_));
AOI21X1 AOI21X1_1128 ( .A(u2__abc_52138_new_n5118_), .B(u2__abc_52138_new_n10463_), .C(u2__abc_52138_new_n10464_), .Y(u2__abc_52138_new_n10465_));
AOI21X1 AOI21X1_1129 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5052_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10467_));
AOI21X1 AOI21X1_113 ( .A(u2__abc_52138_new_n5797_), .B(u2__abc_52138_new_n5469_), .C(u2__abc_52138_new_n5474_), .Y(u2__abc_52138_new_n5798_));
AOI21X1 AOI21X1_1130 ( .A(u2__abc_52138_new_n10468_), .B(u2__abc_52138_new_n10460_), .C(rst), .Y(u2__0remHi_451_0__366_));
AOI21X1 AOI21X1_1131 ( .A(u2__abc_52138_new_n5123_), .B(u2__abc_52138_new_n10472_), .C(u2__abc_52138_new_n10473_), .Y(u2__abc_52138_new_n10474_));
AOI21X1 AOI21X1_1132 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5059_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10476_));
AOI21X1 AOI21X1_1133 ( .A(u2__abc_52138_new_n10477_), .B(u2__abc_52138_new_n10470_), .C(rst), .Y(u2__0remHi_451_0__367_));
AOI21X1 AOI21X1_1134 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5045_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10493_));
AOI21X1 AOI21X1_1135 ( .A(u2__abc_52138_new_n10494_), .B(u2__abc_52138_new_n10479_), .C(rst), .Y(u2__0remHi_451_0__368_));
AOI21X1 AOI21X1_1136 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5886_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10501_));
AOI21X1 AOI21X1_1137 ( .A(u2__abc_52138_new_n10502_), .B(u2__abc_52138_new_n10496_), .C(rst), .Y(u2__0remHi_451_0__369_));
AOI21X1 AOI21X1_1138 ( .A(u2__abc_52138_new_n5049_), .B(u2__abc_52138_new_n10507_), .C(u2__abc_52138_new_n10508_), .Y(u2__abc_52138_new_n10509_));
AOI21X1 AOI21X1_1139 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5084_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10511_));
AOI21X1 AOI21X1_114 ( .A(u2__abc_52138_new_n5487_), .B(u2__abc_52138_new_n5481_), .C(u2__abc_52138_new_n5486_), .Y(u2__abc_52138_new_n5805_));
AOI21X1 AOI21X1_1140 ( .A(u2__abc_52138_new_n10512_), .B(u2__abc_52138_new_n10504_), .C(rst), .Y(u2__0remHi_451_0__370_));
AOI21X1 AOI21X1_1141 ( .A(u2__abc_52138_new_n5050_), .B(u2__abc_52138_new_n10516_), .C(u2__abc_52138_new_n10517_), .Y(u2__abc_52138_new_n10518_));
AOI21X1 AOI21X1_1142 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5078_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10520_));
AOI21X1 AOI21X1_1143 ( .A(u2__abc_52138_new_n10521_), .B(u2__abc_52138_new_n10514_), .C(rst), .Y(u2__0remHi_451_0__371_));
AOI21X1 AOI21X1_1144 ( .A(u2__abc_52138_new_n5059_), .B(u2_o_367_), .C(u2__abc_52138_new_n5051_), .Y(u2__abc_52138_new_n10525_));
AOI21X1 AOI21X1_1145 ( .A(u2__abc_52138_new_n5086_), .B(u2__abc_52138_new_n10528_), .C(u2__abc_52138_new_n10529_), .Y(u2__abc_52138_new_n10530_));
AOI21X1 AOI21X1_1146 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5065_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10532_));
AOI21X1 AOI21X1_1147 ( .A(u2__abc_52138_new_n10533_), .B(u2__abc_52138_new_n10523_), .C(rst), .Y(u2__0remHi_451_0__372_));
AOI21X1 AOI21X1_1148 ( .A(u2__abc_52138_new_n5081_), .B(u2__abc_52138_new_n10537_), .C(u2__abc_52138_new_n10538_), .Y(u2__abc_52138_new_n10539_));
AOI21X1 AOI21X1_1149 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5070_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10541_));
AOI21X1 AOI21X1_115 ( .A(u2__abc_52138_new_n5808_), .B(u2__abc_52138_new_n5390_), .C(u2__abc_52138_new_n5395_), .Y(u2__abc_52138_new_n5809_));
AOI21X1 AOI21X1_1150 ( .A(u2__abc_52138_new_n10542_), .B(u2__abc_52138_new_n10535_), .C(rst), .Y(u2__0remHi_451_0__373_));
AOI21X1 AOI21X1_1151 ( .A(u2__abc_52138_new_n5069_), .B(u2__abc_52138_new_n10546_), .C(u2__abc_52138_new_n10547_), .Y(u2__abc_52138_new_n10548_));
AOI21X1 AOI21X1_1152 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5020_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10550_));
AOI21X1 AOI21X1_1153 ( .A(u2__abc_52138_new_n10551_), .B(u2__abc_52138_new_n10544_), .C(rst), .Y(u2__0remHi_451_0__374_));
AOI21X1 AOI21X1_1154 ( .A(u2__abc_52138_new_n5074_), .B(u2__abc_52138_new_n10555_), .C(u2__abc_52138_new_n10556_), .Y(u2__abc_52138_new_n10557_));
AOI21X1 AOI21X1_1155 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5023_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10559_));
AOI21X1 AOI21X1_1156 ( .A(u2__abc_52138_new_n10560_), .B(u2__abc_52138_new_n10553_), .C(rst), .Y(u2__0remHi_451_0__375_));
AOI21X1 AOI21X1_1157 ( .A(u2__abc_52138_new_n5894_), .B(u2__abc_52138_new_n5066_), .C(u2__abc_52138_new_n5071_), .Y(u2__abc_52138_new_n10565_));
AOI21X1 AOI21X1_1158 ( .A(u2__abc_52138_new_n5895_), .B(u2__abc_52138_new_n10563_), .C(u2__abc_52138_new_n10566_), .Y(u2__abc_52138_new_n10567_));
AOI21X1 AOI21X1_1159 ( .A(u2__abc_52138_new_n5022_), .B(u2__abc_52138_new_n10568_), .C(u2__abc_52138_new_n10569_), .Y(u2__abc_52138_new_n10570_));
AOI21X1 AOI21X1_116 ( .A(u2__abc_52138_new_n5819_), .B(u2__abc_52138_new_n5820_), .C(u2__abc_52138_new_n5397_), .Y(u2__abc_52138_new_n5821_));
AOI21X1 AOI21X1_1160 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5030_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10572_));
AOI21X1 AOI21X1_1161 ( .A(u2__abc_52138_new_n10573_), .B(u2__abc_52138_new_n10562_), .C(rst), .Y(u2__0remHi_451_0__376_));
AOI21X1 AOI21X1_1162 ( .A(u2__abc_52138_new_n5028_), .B(u2__abc_52138_new_n10577_), .C(u2__abc_52138_new_n10578_), .Y(u2__abc_52138_new_n10579_));
AOI21X1 AOI21X1_1163 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5035_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10581_));
AOI21X1 AOI21X1_1164 ( .A(u2__abc_52138_new_n10582_), .B(u2__abc_52138_new_n10575_), .C(rst), .Y(u2__0remHi_451_0__377_));
AOI21X1 AOI21X1_1165 ( .A(u2__abc_52138_new_n10568_), .B(u2__abc_52138_new_n10585_), .C(u2__abc_52138_new_n10587_), .Y(u2__abc_52138_new_n10588_));
AOI21X1 AOI21X1_1166 ( .A(u2__abc_52138_new_n10588_), .B(u2__abc_52138_new_n5034_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n10590_));
AOI21X1 AOI21X1_1167 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n10593_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10594_));
AOI21X1 AOI21X1_1168 ( .A(u2__abc_52138_new_n10595_), .B(u2__abc_52138_new_n10584_), .C(rst), .Y(u2__0remHi_451_0__378_));
AOI21X1 AOI21X1_1169 ( .A(u2__abc_52138_new_n10598_), .B(u2__abc_52138_new_n10599_), .C(u2__abc_52138_new_n10600_), .Y(u2__abc_52138_new_n10601_));
AOI21X1 AOI21X1_117 ( .A(u2__abc_52138_new_n5416_), .B(u2__abc_52138_new_n5408_), .C(u2__abc_52138_new_n5413_), .Y(u2__abc_52138_new_n5824_));
AOI21X1 AOI21X1_1170 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5011_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10603_));
AOI21X1 AOI21X1_1171 ( .A(u2__abc_52138_new_n10604_), .B(u2__abc_52138_new_n10597_), .C(rst), .Y(u2__0remHi_451_0__379_));
AOI21X1 AOI21X1_1172 ( .A(u2__abc_52138_new_n5040_), .B(u2__abc_52138_new_n5031_), .C(u2__abc_52138_new_n5036_), .Y(u2__abc_52138_new_n10607_));
AOI21X1 AOI21X1_1173 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4999_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10614_));
AOI21X1 AOI21X1_1174 ( .A(u2__abc_52138_new_n10615_), .B(u2__abc_52138_new_n10606_), .C(rst), .Y(u2__0remHi_451_0__380_));
AOI21X1 AOI21X1_1175 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5006_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10622_));
AOI21X1 AOI21X1_1176 ( .A(u2__abc_52138_new_n10623_), .B(u2__abc_52138_new_n10617_), .C(rst), .Y(u2__0remHi_451_0__381_));
AOI21X1 AOI21X1_1177 ( .A(u2__abc_52138_new_n5003_), .B(u2__abc_52138_new_n10629_), .C(u2__abc_52138_new_n10630_), .Y(u2__abc_52138_new_n10631_));
AOI21X1 AOI21X1_1178 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6176_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10633_));
AOI21X1 AOI21X1_1179 ( .A(u2__abc_52138_new_n10634_), .B(u2__abc_52138_new_n10625_), .C(rst), .Y(u2__0remHi_451_0__382_));
AOI21X1 AOI21X1_118 ( .A(u2__abc_52138_new_n5825_), .B(u2__abc_52138_new_n5421_), .C(u2__abc_52138_new_n5426_), .Y(u2__abc_52138_new_n5826_));
AOI21X1 AOI21X1_1180 ( .A(u2__abc_52138_new_n5008_), .B(u2__abc_52138_new_n10638_), .C(u2__abc_52138_new_n10639_), .Y(u2__abc_52138_new_n10640_));
AOI21X1 AOI21X1_1181 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6173_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10642_));
AOI21X1 AOI21X1_1182 ( .A(u2__abc_52138_new_n10643_), .B(u2__abc_52138_new_n10636_), .C(rst), .Y(u2__0remHi_451_0__383_));
AOI21X1 AOI21X1_1183 ( .A(u2__abc_52138_new_n5008_), .B(u2__abc_52138_new_n5000_), .C(u2__abc_52138_new_n5007_), .Y(u2__abc_52138_new_n10654_));
AOI21X1 AOI21X1_1184 ( .A(u2__abc_52138_new_n10652_), .B(u2__abc_52138_new_n5017_), .C(u2__abc_52138_new_n10655_), .Y(u2__abc_52138_new_n10656_));
AOI21X1 AOI21X1_1185 ( .A(u2__abc_52138_new_n10484_), .B(u2__abc_52138_new_n5090_), .C(u2__abc_52138_new_n10657_), .Y(u2__abc_52138_new_n10658_));
AOI21X1 AOI21X1_1186 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6160_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10667_));
AOI21X1 AOI21X1_1187 ( .A(u2__abc_52138_new_n10668_), .B(u2__abc_52138_new_n10645_), .C(rst), .Y(u2__0remHi_451_0__384_));
AOI21X1 AOI21X1_1188 ( .A(u2__abc_52138_new_n6175_), .B(u2__abc_52138_new_n10671_), .C(u2__abc_52138_new_n10672_), .Y(u2__abc_52138_new_n10673_));
AOI21X1 AOI21X1_1189 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6167_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10675_));
AOI21X1 AOI21X1_119 ( .A(u2__abc_52138_new_n5445_), .B(u2__abc_52138_new_n5449_), .C(u2__abc_52138_new_n5444_), .Y(u2__abc_52138_new_n5828_));
AOI21X1 AOI21X1_1190 ( .A(u2__abc_52138_new_n10676_), .B(u2__abc_52138_new_n10670_), .C(rst), .Y(u2__0remHi_451_0__385_));
AOI21X1 AOI21X1_1191 ( .A(u2__abc_52138_new_n6164_), .B(u2__abc_52138_new_n10682_), .C(u2__abc_52138_new_n10683_), .Y(u2__abc_52138_new_n10684_));
AOI21X1 AOI21X1_1192 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6152_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10686_));
AOI21X1 AOI21X1_1193 ( .A(u2__abc_52138_new_n10687_), .B(u2__abc_52138_new_n10678_), .C(rst), .Y(u2__0remHi_451_0__386_));
AOI21X1 AOI21X1_1194 ( .A(u2__abc_52138_new_n6169_), .B(u2__abc_52138_new_n10691_), .C(u2__abc_52138_new_n10692_), .Y(u2__abc_52138_new_n10693_));
AOI21X1 AOI21X1_1195 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6149_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10695_));
AOI21X1 AOI21X1_1196 ( .A(u2__abc_52138_new_n10696_), .B(u2__abc_52138_new_n10689_), .C(rst), .Y(u2__0remHi_451_0__387_));
AOI21X1 AOI21X1_1197 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6136_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10710_));
AOI21X1 AOI21X1_1198 ( .A(u2__abc_52138_new_n10711_), .B(u2__abc_52138_new_n10698_), .C(rst), .Y(u2__0remHi_451_0__388_));
AOI21X1 AOI21X1_1199 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6141_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10718_));
AOI21X1 AOI21X1_12 ( .A(u2__abc_52138_new_n3107_), .B(u2__abc_52138_new_n3023_), .C(u2__abc_52138_new_n3106_), .Y(u2__abc_52138_new_n3108_));
AOI21X1 AOI21X1_120 ( .A(u2__abc_52138_new_n5439_), .B(u2__abc_52138_new_n5433_), .C(u2__abc_52138_new_n5438_), .Y(u2__abc_52138_new_n5829_));
AOI21X1 AOI21X1_1200 ( .A(u2__abc_52138_new_n10719_), .B(u2__abc_52138_new_n10713_), .C(rst), .Y(u2__0remHi_451_0__389_));
AOI21X1 AOI21X1_1201 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6292_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10731_));
AOI21X1 AOI21X1_1202 ( .A(u2__abc_52138_new_n10732_), .B(u2__abc_52138_new_n10721_), .C(rst), .Y(u2__0remHi_451_0__390_));
AOI21X1 AOI21X1_1203 ( .A(u2__abc_52138_new_n6145_), .B(u2__abc_52138_new_n10736_), .C(u2__abc_52138_new_n10737_), .Y(u2__abc_52138_new_n10738_));
AOI21X1 AOI21X1_1204 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6297_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10740_));
AOI21X1 AOI21X1_1205 ( .A(u2__abc_52138_new_n10741_), .B(u2__abc_52138_new_n10734_), .C(rst), .Y(u2__0remHi_451_0__391_));
AOI21X1 AOI21X1_1206 ( .A(u2__abc_52138_new_n10744_), .B(u2__abc_52138_new_n10724_), .C(u2__abc_52138_new_n10746_), .Y(u2__abc_52138_new_n10747_));
AOI21X1 AOI21X1_1207 ( .A(u2__abc_52138_new_n6296_), .B(u2__abc_52138_new_n10751_), .C(u2__abc_52138_new_n10752_), .Y(u2__abc_52138_new_n10753_));
AOI21X1 AOI21X1_1208 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6280_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10755_));
AOI21X1 AOI21X1_1209 ( .A(u2__abc_52138_new_n10756_), .B(u2__abc_52138_new_n10743_), .C(rst), .Y(u2__0remHi_451_0__392_));
AOI21X1 AOI21X1_121 ( .A(u2__abc_52138_new_n5827_), .B(u2__abc_52138_new_n5452_), .C(u2__abc_52138_new_n5830_), .Y(u2__abc_52138_new_n5831_));
AOI21X1 AOI21X1_1210 ( .A(u2__abc_52138_new_n10763_), .B(u2__abc_52138_new_n10761_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n10764_));
AOI21X1 AOI21X1_1211 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6352_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10766_));
AOI21X1 AOI21X1_1212 ( .A(u2__abc_52138_new_n10767_), .B(u2__abc_52138_new_n10758_), .C(rst), .Y(u2__0remHi_451_0__393_));
AOI21X1 AOI21X1_1213 ( .A(u2__abc_52138_new_n6284_), .B(u2__abc_52138_new_n10770_), .C(u2__abc_52138_new_n10771_), .Y(u2__abc_52138_new_n10772_));
AOI21X1 AOI21X1_1214 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6320_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10774_));
AOI21X1 AOI21X1_1215 ( .A(u2__abc_52138_new_n10775_), .B(u2__abc_52138_new_n10769_), .C(rst), .Y(u2__0remHi_451_0__394_));
AOI21X1 AOI21X1_1216 ( .A(u2__abc_52138_new_n6290_), .B(u2__abc_52138_new_n10779_), .C(u2__abc_52138_new_n10780_), .Y(u2__abc_52138_new_n10781_));
AOI21X1 AOI21X1_1217 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6317_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10783_));
AOI21X1 AOI21X1_1218 ( .A(u2__abc_52138_new_n10784_), .B(u2__abc_52138_new_n10777_), .C(rst), .Y(u2__0remHi_451_0__395_));
AOI21X1 AOI21X1_1219 ( .A(u2__abc_52138_new_n10751_), .B(u2__abc_52138_new_n6303_), .C(u2__abc_52138_new_n10791_), .Y(u2__abc_52138_new_n10792_));
AOI21X1 AOI21X1_122 ( .A(u2__abc_52138_new_n5781_), .B(u2__abc_52138_new_n5547_), .C(u2__abc_52138_new_n5834_), .Y(u2__abc_52138_new_n5835_));
AOI21X1 AOI21X1_1220 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6304_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10799_));
AOI21X1 AOI21X1_1221 ( .A(u2__abc_52138_new_n10800_), .B(u2__abc_52138_new_n10786_), .C(rst), .Y(u2__0remHi_451_0__396_));
AOI21X1 AOI21X1_1222 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6309_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10807_));
AOI21X1 AOI21X1_1223 ( .A(u2__abc_52138_new_n10808_), .B(u2__abc_52138_new_n10802_), .C(rst), .Y(u2__0remHi_451_0__397_));
AOI21X1 AOI21X1_1224 ( .A(u2__abc_52138_new_n6308_), .B(u2__abc_52138_new_n10813_), .C(u2__abc_52138_new_n10814_), .Y(u2__abc_52138_new_n10815_));
AOI21X1 AOI21X1_1225 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6232_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10817_));
AOI21X1 AOI21X1_1226 ( .A(u2__abc_52138_new_n10818_), .B(u2__abc_52138_new_n10810_), .C(rst), .Y(u2__0remHi_451_0__398_));
AOI21X1 AOI21X1_1227 ( .A(u2__abc_52138_new_n6313_), .B(u2__abc_52138_new_n10822_), .C(u2__abc_52138_new_n10823_), .Y(u2__abc_52138_new_n10824_));
AOI21X1 AOI21X1_1228 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6239_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10826_));
AOI21X1 AOI21X1_1229 ( .A(u2__abc_52138_new_n10827_), .B(u2__abc_52138_new_n10820_), .C(rst), .Y(u2__0remHi_451_0__399_));
AOI21X1 AOI21X1_123 ( .A(u2__abc_52138_new_n5838_), .B(u2__abc_52138_new_n5355_), .C(u2__abc_52138_new_n5360_), .Y(u2__abc_52138_new_n5839_));
AOI21X1 AOI21X1_1230 ( .A(u2__abc_52138_new_n10791_), .B(u2__abc_52138_new_n6326_), .C(u2__abc_52138_new_n6310_), .Y(u2__abc_52138_new_n10832_));
AOI21X1 AOI21X1_1231 ( .A(u2__abc_52138_new_n10750_), .B(u2__abc_52138_new_n10749_), .C(u2__abc_52138_new_n6327_), .Y(u2__abc_52138_new_n10834_));
AOI21X1 AOI21X1_1232 ( .A(u2__abc_52138_new_n6236_), .B(u2__abc_52138_new_n10836_), .C(u2__abc_52138_new_n10837_), .Y(u2__abc_52138_new_n10838_));
AOI21X1 AOI21X1_1233 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6243_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10840_));
AOI21X1 AOI21X1_1234 ( .A(u2__abc_52138_new_n10841_), .B(u2__abc_52138_new_n10829_), .C(rst), .Y(u2__0remHi_451_0__400_));
AOI21X1 AOI21X1_1235 ( .A(u2__abc_52138_new_n6241_), .B(u2__abc_52138_new_n10845_), .C(u2__abc_52138_new_n10846_), .Y(u2__abc_52138_new_n10847_));
AOI21X1 AOI21X1_1236 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6250_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10849_));
AOI21X1 AOI21X1_1237 ( .A(u2__abc_52138_new_n10850_), .B(u2__abc_52138_new_n10843_), .C(rst), .Y(u2__0remHi_451_0__401_));
AOI21X1 AOI21X1_1238 ( .A(u2__abc_52138_new_n6247_), .B(u2__abc_52138_new_n10855_), .C(u2__abc_52138_new_n10856_), .Y(u2__abc_52138_new_n10857_));
AOI21X1 AOI21X1_1239 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6271_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10859_));
AOI21X1 AOI21X1_124 ( .A(u2__abc_52138_new_n5330_), .B(u2__abc_52138_new_n5322_), .C(u2__abc_52138_new_n5327_), .Y(u2__abc_52138_new_n5842_));
AOI21X1 AOI21X1_1240 ( .A(u2__abc_52138_new_n10860_), .B(u2__abc_52138_new_n10852_), .C(rst), .Y(u2__0remHi_451_0__402_));
AOI21X1 AOI21X1_1241 ( .A(u2__abc_52138_new_n6252_), .B(u2__abc_52138_new_n10864_), .C(u2__abc_52138_new_n10865_), .Y(u2__abc_52138_new_n10866_));
AOI21X1 AOI21X1_1242 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6268_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10868_));
AOI21X1 AOI21X1_1243 ( .A(u2__abc_52138_new_n10869_), .B(u2__abc_52138_new_n10862_), .C(rst), .Y(u2__0remHi_451_0__403_));
AOI21X1 AOI21X1_1244 ( .A(u2__abc_52138_new_n10873_), .B(u2__abc_52138_new_n10853_), .C(u2__abc_52138_new_n10875_), .Y(u2__abc_52138_new_n10876_));
AOI21X1 AOI21X1_1245 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6255_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10883_));
AOI21X1 AOI21X1_1246 ( .A(u2__abc_52138_new_n10884_), .B(u2__abc_52138_new_n10871_), .C(rst), .Y(u2__0remHi_451_0__404_));
AOI21X1 AOI21X1_1247 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6260_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10891_));
AOI21X1 AOI21X1_1248 ( .A(u2__abc_52138_new_n10892_), .B(u2__abc_52138_new_n10886_), .C(rst), .Y(u2__0remHi_451_0__405_));
AOI21X1 AOI21X1_1249 ( .A(u2__abc_52138_new_n6259_), .B(u2__abc_52138_new_n10898_), .C(u2__abc_52138_new_n10899_), .Y(u2__abc_52138_new_n10900_));
AOI21X1 AOI21X1_125 ( .A(u2__abc_52138_new_n5850_), .B(u2__abc_52138_new_n5288_), .C(u2__abc_52138_new_n5293_), .Y(u2__abc_52138_new_n5851_));
AOI21X1 AOI21X1_1250 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6201_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10902_));
AOI21X1 AOI21X1_1251 ( .A(u2__abc_52138_new_n10903_), .B(u2__abc_52138_new_n10894_), .C(rst), .Y(u2__0remHi_451_0__406_));
AOI21X1 AOI21X1_1252 ( .A(u2__abc_52138_new_n6264_), .B(u2__abc_52138_new_n10907_), .C(u2__abc_52138_new_n10908_), .Y(u2__abc_52138_new_n10909_));
AOI21X1 AOI21X1_1253 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6198_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10911_));
AOI21X1 AOI21X1_1254 ( .A(u2__abc_52138_new_n10912_), .B(u2__abc_52138_new_n10905_), .C(rst), .Y(u2__0remHi_451_0__407_));
AOI21X1 AOI21X1_1255 ( .A(u2__abc_52138_new_n6264_), .B(u2__abc_52138_new_n6256_), .C(u2__abc_52138_new_n6261_), .Y(u2__abc_52138_new_n10918_));
AOI21X1 AOI21X1_1256 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6185_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10927_));
AOI21X1 AOI21X1_1257 ( .A(u2__abc_52138_new_n10928_), .B(u2__abc_52138_new_n10914_), .C(rst), .Y(u2__0remHi_451_0__408_));
AOI21X1 AOI21X1_1258 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6192_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10935_));
AOI21X1 AOI21X1_1259 ( .A(u2__abc_52138_new_n10936_), .B(u2__abc_52138_new_n10930_), .C(rst), .Y(u2__0remHi_451_0__409_));
AOI21X1 AOI21X1_126 ( .A(u2__abc_52138_new_n5306_), .B(u2__abc_52138_new_n5300_), .C(u2__abc_52138_new_n5305_), .Y(u2__abc_52138_new_n5857_));
AOI21X1 AOI21X1_1260 ( .A(u2__abc_52138_new_n6189_), .B(u2__abc_52138_new_n10942_), .C(u2__abc_52138_new_n10943_), .Y(u2__abc_52138_new_n10944_));
AOI21X1 AOI21X1_1261 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6224_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10946_));
AOI21X1 AOI21X1_1262 ( .A(u2__abc_52138_new_n10947_), .B(u2__abc_52138_new_n10938_), .C(rst), .Y(u2__0remHi_451_0__410_));
AOI21X1 AOI21X1_1263 ( .A(u2__abc_52138_new_n6194_), .B(u2__abc_52138_new_n10951_), .C(u2__abc_52138_new_n10952_), .Y(u2__abc_52138_new_n10953_));
AOI21X1 AOI21X1_1264 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6221_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10955_));
AOI21X1 AOI21X1_1265 ( .A(u2__abc_52138_new_n10956_), .B(u2__abc_52138_new_n10949_), .C(rst), .Y(u2__0remHi_451_0__411_));
AOI21X1 AOI21X1_1266 ( .A(u2__abc_52138_new_n10921_), .B(u2__abc_52138_new_n6207_), .C(u2__abc_52138_new_n10962_), .Y(u2__abc_52138_new_n10963_));
AOI21X1 AOI21X1_1267 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6208_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10970_));
AOI21X1 AOI21X1_1268 ( .A(u2__abc_52138_new_n10971_), .B(u2__abc_52138_new_n10958_), .C(rst), .Y(u2__0remHi_451_0__412_));
AOI21X1 AOI21X1_1269 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6213_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10979_));
AOI21X1 AOI21X1_127 ( .A(u2__abc_52138_new_n5847_), .B(u2__abc_52138_new_n5320_), .C(u2__abc_52138_new_n5858_), .Y(u2__abc_52138_new_n5859_));
AOI21X1 AOI21X1_1270 ( .A(u2__abc_52138_new_n10980_), .B(u2__abc_52138_new_n10973_), .C(rst), .Y(u2__0remHi_451_0__413_));
AOI21X1 AOI21X1_1271 ( .A(u2__abc_52138_new_n6212_), .B(u2__abc_52138_new_n10985_), .C(u2__abc_52138_new_n10986_), .Y(u2__abc_52138_new_n10987_));
AOI21X1 AOI21X1_1272 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6125_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10989_));
AOI21X1 AOI21X1_1273 ( .A(u2__abc_52138_new_n10990_), .B(u2__abc_52138_new_n10982_), .C(rst), .Y(u2__0remHi_451_0__414_));
AOI21X1 AOI21X1_1274 ( .A(u2__abc_52138_new_n6217_), .B(u2__abc_52138_new_n10994_), .C(u2__abc_52138_new_n10995_), .Y(u2__abc_52138_new_n10996_));
AOI21X1 AOI21X1_1275 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6122_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n10998_));
AOI21X1 AOI21X1_1276 ( .A(u2__abc_52138_new_n10999_), .B(u2__abc_52138_new_n10992_), .C(rst), .Y(u2__0remHi_451_0__415_));
AOI21X1 AOI21X1_1277 ( .A(u2__abc_52138_new_n6230_), .B(u2__abc_52138_new_n10962_), .C(u2__abc_52138_new_n11005_), .Y(u2__abc_52138_new_n11006_));
AOI21X1 AOI21X1_1278 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6110_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11017_));
AOI21X1 AOI21X1_1279 ( .A(u2__abc_52138_new_n11018_), .B(u2__abc_52138_new_n11001_), .C(rst), .Y(u2__0remHi_451_0__416_));
AOI21X1 AOI21X1_128 ( .A(u2__abc_52138_new_n5861_), .B(u2__abc_52138_new_n5194_), .C(u2__abc_52138_new_n5863_), .Y(u2__abc_52138_new_n5864_));
AOI21X1 AOI21X1_1280 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6113_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11025_));
AOI21X1 AOI21X1_1281 ( .A(u2__abc_52138_new_n11026_), .B(u2__abc_52138_new_n11020_), .C(rst), .Y(u2__0remHi_451_0__417_));
AOI21X1 AOI21X1_1282 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6101_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11037_));
AOI21X1 AOI21X1_1283 ( .A(u2__abc_52138_new_n11038_), .B(u2__abc_52138_new_n11028_), .C(rst), .Y(u2__0remHi_451_0__418_));
AOI21X1 AOI21X1_1284 ( .A(u2__abc_52138_new_n11041_), .B(u2__abc_52138_new_n11042_), .C(u2__abc_52138_new_n11043_), .Y(u2__abc_52138_new_n11044_));
AOI21X1 AOI21X1_1285 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6098_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11046_));
AOI21X1 AOI21X1_1286 ( .A(u2__abc_52138_new_n11047_), .B(u2__abc_52138_new_n11040_), .C(rst), .Y(u2__0remHi_451_0__419_));
AOI21X1 AOI21X1_1287 ( .A(u2__abc_52138_new_n11011_), .B(u2__abc_52138_new_n6131_), .C(u2__abc_52138_new_n11053_), .Y(u2__abc_52138_new_n11054_));
AOI21X1 AOI21X1_1288 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6086_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11061_));
AOI21X1 AOI21X1_1289 ( .A(u2__abc_52138_new_n11062_), .B(u2__abc_52138_new_n11049_), .C(rst), .Y(u2__0remHi_451_0__420_));
AOI21X1 AOI21X1_129 ( .A(u2__abc_52138_new_n5866_), .B(u2__abc_52138_new_n5865_), .C(u2__abc_52138_new_n5215_), .Y(u2__abc_52138_new_n5867_));
AOI21X1 AOI21X1_1290 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6091_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11070_));
AOI21X1 AOI21X1_1291 ( .A(u2__abc_52138_new_n11071_), .B(u2__abc_52138_new_n11064_), .C(rst), .Y(u2__0remHi_451_0__421_));
AOI21X1 AOI21X1_1292 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6047_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11081_));
AOI21X1 AOI21X1_1293 ( .A(u2__abc_52138_new_n11082_), .B(u2__abc_52138_new_n11073_), .C(rst), .Y(u2__0remHi_451_0__422_));
AOI21X1 AOI21X1_1294 ( .A(u2__abc_52138_new_n11085_), .B(u2__abc_52138_new_n11086_), .C(u2__abc_52138_new_n11087_), .Y(u2__abc_52138_new_n11088_));
AOI21X1 AOI21X1_1295 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6054_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11090_));
AOI21X1 AOI21X1_1296 ( .A(u2__abc_52138_new_n11091_), .B(u2__abc_52138_new_n11084_), .C(rst), .Y(u2__0remHi_451_0__423_));
AOI21X1 AOI21X1_1297 ( .A(u2__abc_52138_new_n11095_), .B(u2__abc_52138_new_n11074_), .C(u2__abc_52138_new_n11096_), .Y(u2__abc_52138_new_n11097_));
AOI21X1 AOI21X1_1298 ( .A(u2__abc_52138_new_n11011_), .B(u2__abc_52138_new_n6133_), .C(u2__abc_52138_new_n11098_), .Y(u2__abc_52138_new_n11099_));
AOI21X1 AOI21X1_1299 ( .A(u2__abc_52138_new_n6051_), .B(u2__abc_52138_new_n11100_), .C(u2__abc_52138_new_n11101_), .Y(u2__abc_52138_new_n11102_));
AOI21X1 AOI21X1_13 ( .A(u2__abc_52138_new_n3100_), .B(u2__abc_52138_new_n3033_), .C(u2__abc_52138_new_n3109_), .Y(u2__abc_52138_new_n3110_));
AOI21X1 AOI21X1_130 ( .A(u2__abc_52138_new_n5260_), .B(u2__abc_52138_new_n5881_), .C(u2__abc_52138_new_n5879_), .Y(u2__abc_52138_new_n5882_));
AOI21X1 AOI21X1_1300 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6038_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11104_));
AOI21X1 AOI21X1_1301 ( .A(u2__abc_52138_new_n11105_), .B(u2__abc_52138_new_n11093_), .C(rst), .Y(u2__0remHi_451_0__424_));
AOI21X1 AOI21X1_1302 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6041_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11113_));
AOI21X1 AOI21X1_1303 ( .A(u2__abc_52138_new_n11114_), .B(u2__abc_52138_new_n11107_), .C(rst), .Y(u2__0remHi_451_0__425_));
AOI21X1 AOI21X1_1304 ( .A(u2__abc_52138_new_n11109_), .B(u2__abc_52138_new_n11117_), .C(u2__abc_52138_new_n6055_), .Y(u2__abc_52138_new_n11118_));
AOI21X1 AOI21X1_1305 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6075_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11124_));
AOI21X1 AOI21X1_1306 ( .A(u2__abc_52138_new_n11125_), .B(u2__abc_52138_new_n11116_), .C(rst), .Y(u2__0remHi_451_0__426_));
AOI21X1 AOI21X1_1307 ( .A(u2__abc_52138_new_n11128_), .B(u2__abc_52138_new_n11129_), .C(u2__abc_52138_new_n11130_), .Y(u2__abc_52138_new_n11131_));
AOI21X1 AOI21X1_1308 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6072_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11133_));
AOI21X1 AOI21X1_1309 ( .A(u2__abc_52138_new_n11134_), .B(u2__abc_52138_new_n11127_), .C(rst), .Y(u2__0remHi_451_0__427_));
AOI21X1 AOI21X1_131 ( .A(u2__abc_52138_new_n5883_), .B(u2__abc_52138_new_n5228_), .C(u2__abc_52138_new_n5871_), .Y(u2__abc_52138_new_n5884_));
AOI21X1 AOI21X1_1310 ( .A(u2__abc_52138_new_n11108_), .B(u2__abc_52138_new_n6401_), .C(u2__abc_52138_new_n6053_), .Y(u2__abc_52138_new_n11137_));
AOI21X1 AOI21X1_1311 ( .A(u2__abc_52138_new_n11137_), .B(u2__abc_52138_new_n6046_), .C(u2__abc_52138_new_n11138_), .Y(u2__abc_52138_new_n11139_));
AOI21X1 AOI21X1_1312 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6060_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11146_));
AOI21X1 AOI21X1_1313 ( .A(u2__abc_52138_new_n11147_), .B(u2__abc_52138_new_n11136_), .C(rst), .Y(u2__0remHi_451_0__428_));
AOI21X1 AOI21X1_1314 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6065_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11154_));
AOI21X1 AOI21X1_1315 ( .A(u2__abc_52138_new_n11155_), .B(u2__abc_52138_new_n11149_), .C(rst), .Y(u2__0remHi_451_0__429_));
AOI21X1 AOI21X1_1316 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6010_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11166_));
AOI21X1 AOI21X1_1317 ( .A(u2__abc_52138_new_n11167_), .B(u2__abc_52138_new_n11157_), .C(rst), .Y(u2__0remHi_451_0__430_));
AOI21X1 AOI21X1_1318 ( .A(u2__abc_52138_new_n11170_), .B(u2__abc_52138_new_n11171_), .C(u2__abc_52138_new_n11172_), .Y(u2__abc_52138_new_n11173_));
AOI21X1 AOI21X1_1319 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6017_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11175_));
AOI21X1 AOI21X1_132 ( .A(u2__abc_52138_new_n5893_), .B(u2__abc_52138_new_n5088_), .C(u2__abc_52138_new_n5899_), .Y(u2__abc_52138_new_n5900_));
AOI21X1 AOI21X1_1320 ( .A(u2__abc_52138_new_n11176_), .B(u2__abc_52138_new_n11169_), .C(rst), .Y(u2__0remHi_451_0__431_));
AOI21X1 AOI21X1_1321 ( .A(u2__abc_52138_new_n11180_), .B(u2__abc_52138_new_n6068_), .C(u2__abc_52138_new_n11181_), .Y(u2__abc_52138_new_n11182_));
AOI21X1 AOI21X1_1322 ( .A(u2__abc_52138_new_n11098_), .B(u2__abc_52138_new_n6083_), .C(u2__abc_52138_new_n11183_), .Y(u2__abc_52138_new_n11184_));
AOI21X1 AOI21X1_1323 ( .A(u2__abc_52138_new_n6014_), .B(u2__abc_52138_new_n11185_), .C(u2__abc_52138_new_n11186_), .Y(u2__abc_52138_new_n11187_));
AOI21X1 AOI21X1_1324 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6021_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11189_));
AOI21X1 AOI21X1_1325 ( .A(u2__abc_52138_new_n11190_), .B(u2__abc_52138_new_n11178_), .C(rst), .Y(u2__0remHi_451_0__432_));
AOI21X1 AOI21X1_1326 ( .A(u2__abc_52138_new_n6019_), .B(u2__abc_52138_new_n11195_), .C(u2__abc_52138_new_n11196_), .Y(u2__abc_52138_new_n11197_));
AOI21X1 AOI21X1_1327 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6028_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11199_));
AOI21X1 AOI21X1_1328 ( .A(u2__abc_52138_new_n11200_), .B(u2__abc_52138_new_n11192_), .C(rst), .Y(u2__0remHi_451_0__433_));
AOI21X1 AOI21X1_1329 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6003_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11211_));
AOI21X1 AOI21X1_133 ( .A(u2__abc_52138_new_n5915_), .B(u2__abc_52138_new_n5117_), .C(u2__abc_52138_new_n5122_), .Y(u2__abc_52138_new_n5916_));
AOI21X1 AOI21X1_1330 ( .A(u2__abc_52138_new_n11212_), .B(u2__abc_52138_new_n11202_), .C(rst), .Y(u2__0remHi_451_0__434_));
AOI21X1 AOI21X1_1331 ( .A(u2__abc_52138_new_n6030_), .B(u2__abc_52138_new_n11215_), .C(u2__abc_52138_new_n11216_), .Y(u2__abc_52138_new_n11217_));
AOI21X1 AOI21X1_1332 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6000_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11219_));
AOI21X1 AOI21X1_1333 ( .A(u2__abc_52138_new_n11220_), .B(u2__abc_52138_new_n11214_), .C(rst), .Y(u2__0remHi_451_0__435_));
AOI21X1 AOI21X1_1334 ( .A(u2__abc_52138_new_n6007_), .B(u2__abc_52138_new_n11226_), .C(u2__abc_52138_new_n11227_), .Y(u2__abc_52138_new_n11228_));
AOI21X1 AOI21X1_1335 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5987_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11230_));
AOI21X1 AOI21X1_1336 ( .A(u2__abc_52138_new_n11231_), .B(u2__abc_52138_new_n11222_), .C(rst), .Y(u2__0remHi_451_0__436_));
AOI21X1 AOI21X1_1337 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5992_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11241_));
AOI21X1 AOI21X1_1338 ( .A(u2__abc_52138_new_n11242_), .B(u2__abc_52138_new_n11233_), .C(rst), .Y(u2__0remHi_451_0__437_));
AOI21X1 AOI21X1_1339 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5967_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11251_));
AOI21X1 AOI21X1_134 ( .A(u2__abc_52138_new_n5166_), .B(u2__abc_52138_new_n5160_), .C(u2__abc_52138_new_n5165_), .Y(u2__abc_52138_new_n5923_));
AOI21X1 AOI21X1_1340 ( .A(u2__abc_52138_new_n11252_), .B(u2__abc_52138_new_n11244_), .C(rst), .Y(u2__0remHi_451_0__438_));
AOI21X1 AOI21X1_1341 ( .A(u2__abc_52138_new_n5996_), .B(u2__abc_52138_new_n11255_), .C(u2__abc_52138_new_n11256_), .Y(u2__abc_52138_new_n11257_));
AOI21X1 AOI21X1_1342 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6415_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11259_));
AOI21X1 AOI21X1_1343 ( .A(u2__abc_52138_new_n11260_), .B(u2__abc_52138_new_n11254_), .C(rst), .Y(u2__0remHi_451_0__439_));
AOI21X1 AOI21X1_1344 ( .A(u2__abc_52138_new_n6002_), .B(u2__abc_52138_new_n6004_), .C(u2__abc_52138_new_n6001_), .Y(u2__abc_52138_new_n11265_));
AOI21X1 AOI21X1_1345 ( .A(u2__abc_52138_new_n5996_), .B(u2__abc_52138_new_n5988_), .C(u2__abc_52138_new_n5993_), .Y(u2__abc_52138_new_n11266_));
AOI21X1 AOI21X1_1346 ( .A(u2__abc_52138_new_n11264_), .B(u2__abc_52138_new_n6009_), .C(u2__abc_52138_new_n11267_), .Y(u2__abc_52138_new_n11268_));
AOI21X1 AOI21X1_1347 ( .A(u2__abc_52138_new_n5971_), .B(u2__abc_52138_new_n11269_), .C(u2__abc_52138_new_n11270_), .Y(u2__abc_52138_new_n11271_));
AOI21X1 AOI21X1_1348 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5974_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11273_));
AOI21X1 AOI21X1_1349 ( .A(u2__abc_52138_new_n11274_), .B(u2__abc_52138_new_n11262_), .C(rst), .Y(u2__0remHi_451_0__440_));
AOI21X1 AOI21X1_135 ( .A(u2__abc_52138_new_n5177_), .B(u2__abc_52138_new_n5171_), .C(u2__abc_52138_new_n5176_), .Y(u2__abc_52138_new_n5924_));
AOI21X1 AOI21X1_1350 ( .A(u2__abc_52138_new_n5972_), .B(u2__abc_52138_new_n11278_), .C(u2__abc_52138_new_n11279_), .Y(u2__abc_52138_new_n11280_));
AOI21X1 AOI21X1_1351 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5981_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11282_));
AOI21X1 AOI21X1_1352 ( .A(u2__abc_52138_new_n11283_), .B(u2__abc_52138_new_n11276_), .C(rst), .Y(u2__0remHi_451_0__441_));
AOI21X1 AOI21X1_1353 ( .A(u2__abc_52138_new_n11269_), .B(u2__abc_52138_new_n11287_), .C(u2__abc_52138_new_n11289_), .Y(u2__abc_52138_new_n11290_));
AOI21X1 AOI21X1_1354 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5960_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11296_));
AOI21X1 AOI21X1_1355 ( .A(u2__abc_52138_new_n11297_), .B(u2__abc_52138_new_n11285_), .C(rst), .Y(u2__0remHi_451_0__442_));
AOI21X1 AOI21X1_1356 ( .A(u2__abc_52138_new_n5983_), .B(u2__abc_52138_new_n11301_), .C(u2__abc_52138_new_n11302_), .Y(u2__abc_52138_new_n11303_));
AOI21X1 AOI21X1_1357 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5957_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11305_));
AOI21X1 AOI21X1_1358 ( .A(u2__abc_52138_new_n11306_), .B(u2__abc_52138_new_n11299_), .C(rst), .Y(u2__0remHi_451_0__443_));
AOI21X1 AOI21X1_1359 ( .A(u2__abc_52138_new_n6413_), .B(u2__abc_52138_new_n11289_), .C(u2__abc_52138_new_n11310_), .Y(u2__abc_52138_new_n11311_));
AOI21X1 AOI21X1_136 ( .A(u2__abc_52138_new_n5922_), .B(u2__abc_52138_new_n5179_), .C(u2__abc_52138_new_n5925_), .Y(u2__abc_52138_new_n5926_));
AOI21X1 AOI21X1_1360 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5944_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11319_));
AOI21X1 AOI21X1_1361 ( .A(u2__abc_52138_new_n11320_), .B(u2__abc_52138_new_n11308_), .C(rst), .Y(u2__0remHi_451_0__444_));
AOI21X1 AOI21X1_1362 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5951_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11327_));
AOI21X1 AOI21X1_1363 ( .A(u2__abc_52138_new_n11328_), .B(u2__abc_52138_new_n11322_), .C(rst), .Y(u2__0remHi_451_0__445_));
AOI21X1 AOI21X1_1364 ( .A(u2__abc_52138_new_n5948_), .B(u2__abc_52138_new_n11335_), .C(u2__abc_52138_new_n11336_), .Y(u2__abc_52138_new_n11337_));
AOI21X1 AOI21X1_1365 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3008_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11339_));
AOI21X1 AOI21X1_1366 ( .A(u2__abc_52138_new_n11340_), .B(u2__abc_52138_new_n11330_), .C(rst), .Y(u2__0remHi_451_0__446_));
AOI21X1 AOI21X1_1367 ( .A(u2__abc_52138_new_n5953_), .B(u2__abc_52138_new_n11344_), .C(u2__abc_52138_new_n11345_), .Y(u2__abc_52138_new_n11346_));
AOI21X1 AOI21X1_1368 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3003_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11348_));
AOI21X1 AOI21X1_1369 ( .A(u2__abc_52138_new_n11349_), .B(u2__abc_52138_new_n11342_), .C(rst), .Y(u2__0remHi_451_0__447_));
AOI21X1 AOI21X1_137 ( .A(u2__abc_52138_new_n5008_), .B(u2__abc_52138_new_n5002_), .C(u2__abc_52138_new_n5005_), .Y(u2__abc_52138_new_n5937_));
AOI21X1 AOI21X1_1370 ( .A(u2__abc_52138_new_n11355_), .B(u2__abc_52138_new_n11333_), .C(u2__abc_52138_new_n11354_), .Y(u2__abc_52138_new_n11356_));
AOI21X1 AOI21X1_1371 ( .A(u2__abc_52138_new_n11011_), .B(u2__abc_52138_new_n6135_), .C(u2__abc_52138_new_n11359_), .Y(u2__abc_52138_new_n11360_));
AOI21X1 AOI21X1_1372 ( .A(u2__abc_52138_new_n3012_), .B(u2__abc_52138_new_n11361_), .C(u2__abc_52138_new_n11362_), .Y(u2__abc_52138_new_n11363_));
AOI21X1 AOI21X1_1373 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n2999_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11365_));
AOI21X1 AOI21X1_1374 ( .A(u2__abc_52138_new_n11366_), .B(u2__abc_52138_new_n11351_), .C(rst), .Y(u2__0remHi_451_0__448_));
AOI21X1 AOI21X1_1375 ( .A(u2__abc_52138_new_n3007_), .B(u2__abc_52138_new_n11370_), .C(u2__abc_52138_new_n11371_), .Y(u2__abc_52138_new_n11372_));
AOI21X1 AOI21X1_1376 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6447_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n11374_));
AOI21X1 AOI21X1_1377 ( .A(u2__abc_52138_new_n11375_), .B(u2__abc_52138_new_n11368_), .C(rst), .Y(u2__0remHi_451_0__449_));
AOI21X1 AOI21X1_1378 ( .A(u2_cnt_1_), .B(u2__abc_52138_new_n2982_), .C(u2__abc_52138_new_n11383_), .Y(u2__abc_52138_new_n11384_));
AOI21X1 AOI21X1_1379 ( .A(u2__abc_52138_new_n11377_), .B(u2__abc_52138_new_n2974_), .C(u2__abc_52138_new_n11384_), .Y(u2__0cnt_7_0__1_));
AOI21X1 AOI21X1_138 ( .A(u2__abc_52138_new_n5017_), .B(u2__abc_52138_new_n5932_), .C(u2__abc_52138_new_n5938_), .Y(u2__abc_52138_new_n5939_));
AOI21X1 AOI21X1_1380 ( .A(u2__abc_52138_new_n11382_), .B(ce), .C(rst), .Y(u2__abc_52138_new_n11387_));
AOI21X1 AOI21X1_1381 ( .A(u2__abc_52138_new_n11417_), .B(u2__abc_52138_new_n11418_), .C(rst), .Y(u2__0remLo_451_0__2_));
AOI21X1 AOI21X1_1382 ( .A(u2__abc_52138_new_n11420_), .B(u2__abc_52138_new_n11421_), .C(rst), .Y(u2__0remLo_451_0__3_));
AOI21X1 AOI21X1_1383 ( .A(u2__abc_52138_new_n11423_), .B(u2__abc_52138_new_n11424_), .C(rst), .Y(u2__0remLo_451_0__4_));
AOI21X1 AOI21X1_1384 ( .A(u2__abc_52138_new_n11426_), .B(u2__abc_52138_new_n11427_), .C(rst), .Y(u2__0remLo_451_0__5_));
AOI21X1 AOI21X1_1385 ( .A(u2__abc_52138_new_n11429_), .B(u2__abc_52138_new_n11430_), .C(rst), .Y(u2__0remLo_451_0__6_));
AOI21X1 AOI21X1_1386 ( .A(u2__abc_52138_new_n11432_), .B(u2__abc_52138_new_n11433_), .C(rst), .Y(u2__0remLo_451_0__7_));
AOI21X1 AOI21X1_1387 ( .A(u2__abc_52138_new_n11435_), .B(u2__abc_52138_new_n11436_), .C(rst), .Y(u2__0remLo_451_0__8_));
AOI21X1 AOI21X1_1388 ( .A(u2__abc_52138_new_n11438_), .B(u2__abc_52138_new_n11439_), .C(rst), .Y(u2__0remLo_451_0__9_));
AOI21X1 AOI21X1_1389 ( .A(u2__abc_52138_new_n11441_), .B(u2__abc_52138_new_n11442_), .C(rst), .Y(u2__0remLo_451_0__10_));
AOI21X1 AOI21X1_139 ( .A(u2__abc_52138_new_n5182_), .B(u2__abc_52138_new_n5885_), .C(u2__abc_52138_new_n5940_), .Y(u2__abc_52138_new_n5941_));
AOI21X1 AOI21X1_1390 ( .A(u2__abc_52138_new_n11444_), .B(u2__abc_52138_new_n11445_), .C(rst), .Y(u2__0remLo_451_0__11_));
AOI21X1 AOI21X1_1391 ( .A(u2__abc_52138_new_n11447_), .B(u2__abc_52138_new_n11448_), .C(rst), .Y(u2__0remLo_451_0__12_));
AOI21X1 AOI21X1_1392 ( .A(u2__abc_52138_new_n11450_), .B(u2__abc_52138_new_n11451_), .C(rst), .Y(u2__0remLo_451_0__13_));
AOI21X1 AOI21X1_1393 ( .A(u2__abc_52138_new_n11453_), .B(u2__abc_52138_new_n11454_), .C(rst), .Y(u2__0remLo_451_0__14_));
AOI21X1 AOI21X1_1394 ( .A(u2__abc_52138_new_n11456_), .B(u2__abc_52138_new_n11457_), .C(rst), .Y(u2__0remLo_451_0__15_));
AOI21X1 AOI21X1_1395 ( .A(u2__abc_52138_new_n11459_), .B(u2__abc_52138_new_n11460_), .C(rst), .Y(u2__0remLo_451_0__16_));
AOI21X1 AOI21X1_1396 ( .A(u2__abc_52138_new_n11462_), .B(u2__abc_52138_new_n11463_), .C(rst), .Y(u2__0remLo_451_0__17_));
AOI21X1 AOI21X1_1397 ( .A(u2__abc_52138_new_n11465_), .B(u2__abc_52138_new_n11466_), .C(rst), .Y(u2__0remLo_451_0__18_));
AOI21X1 AOI21X1_1398 ( .A(u2__abc_52138_new_n11468_), .B(u2__abc_52138_new_n11469_), .C(rst), .Y(u2__0remLo_451_0__19_));
AOI21X1 AOI21X1_1399 ( .A(u2__abc_52138_new_n11471_), .B(u2__abc_52138_new_n11472_), .C(rst), .Y(u2__0remLo_451_0__20_));
AOI21X1 AOI21X1_14 ( .A(u2__abc_52138_new_n3199_), .B(u2__abc_52138_new_n3176_), .C(u2__abc_52138_new_n3200_), .Y(u2__abc_52138_new_n3201_));
AOI21X1 AOI21X1_140 ( .A(u2__abc_52138_new_n4998_), .B(u2__abc_52138_new_n5736_), .C(u2__abc_52138_new_n5942_), .Y(u2__abc_52138_new_n5943_));
AOI21X1 AOI21X1_1400 ( .A(u2__abc_52138_new_n11474_), .B(u2__abc_52138_new_n11475_), .C(rst), .Y(u2__0remLo_451_0__21_));
AOI21X1 AOI21X1_1401 ( .A(u2__abc_52138_new_n11477_), .B(u2__abc_52138_new_n11478_), .C(rst), .Y(u2__0remLo_451_0__22_));
AOI21X1 AOI21X1_1402 ( .A(u2__abc_52138_new_n11480_), .B(u2__abc_52138_new_n11481_), .C(rst), .Y(u2__0remLo_451_0__23_));
AOI21X1 AOI21X1_1403 ( .A(u2__abc_52138_new_n11483_), .B(u2__abc_52138_new_n11484_), .C(rst), .Y(u2__0remLo_451_0__24_));
AOI21X1 AOI21X1_1404 ( .A(u2__abc_52138_new_n11486_), .B(u2__abc_52138_new_n11487_), .C(rst), .Y(u2__0remLo_451_0__25_));
AOI21X1 AOI21X1_1405 ( .A(u2__abc_52138_new_n11489_), .B(u2__abc_52138_new_n11490_), .C(rst), .Y(u2__0remLo_451_0__26_));
AOI21X1 AOI21X1_1406 ( .A(u2__abc_52138_new_n11492_), .B(u2__abc_52138_new_n11493_), .C(rst), .Y(u2__0remLo_451_0__27_));
AOI21X1 AOI21X1_1407 ( .A(u2__abc_52138_new_n11495_), .B(u2__abc_52138_new_n11496_), .C(rst), .Y(u2__0remLo_451_0__28_));
AOI21X1 AOI21X1_1408 ( .A(u2__abc_52138_new_n11498_), .B(u2__abc_52138_new_n11499_), .C(rst), .Y(u2__0remLo_451_0__29_));
AOI21X1 AOI21X1_1409 ( .A(u2__abc_52138_new_n11501_), .B(u2__abc_52138_new_n11502_), .C(rst), .Y(u2__0remLo_451_0__30_));
AOI21X1 AOI21X1_141 ( .A(u2__abc_52138_new_n6334_), .B(u2__abc_52138_new_n6179_), .C(u2__abc_52138_new_n6172_), .Y(u2__abc_52138_new_n6335_));
AOI21X1 AOI21X1_1410 ( .A(u2__abc_52138_new_n11504_), .B(u2__abc_52138_new_n11505_), .C(rst), .Y(u2__0remLo_451_0__31_));
AOI21X1 AOI21X1_1411 ( .A(u2__abc_52138_new_n12234_), .B(u2__abc_52138_new_n12235_), .C(rst), .Y(u2__0remLo_451_0__258_));
AOI21X1 AOI21X1_1412 ( .A(u2__abc_52138_new_n12237_), .B(u2__abc_52138_new_n12238_), .C(rst), .Y(u2__0remLo_451_0__259_));
AOI21X1 AOI21X1_1413 ( .A(u2__abc_52138_new_n12240_), .B(u2__abc_52138_new_n12241_), .C(rst), .Y(u2__0remLo_451_0__260_));
AOI21X1 AOI21X1_1414 ( .A(u2__abc_52138_new_n12243_), .B(u2__abc_52138_new_n12244_), .C(rst), .Y(u2__0remLo_451_0__261_));
AOI21X1 AOI21X1_1415 ( .A(u2__abc_52138_new_n12246_), .B(u2__abc_52138_new_n12247_), .C(rst), .Y(u2__0remLo_451_0__262_));
AOI21X1 AOI21X1_1416 ( .A(u2__abc_52138_new_n12249_), .B(u2__abc_52138_new_n12250_), .C(rst), .Y(u2__0remLo_451_0__263_));
AOI21X1 AOI21X1_1417 ( .A(u2__abc_52138_new_n12252_), .B(u2__abc_52138_new_n12253_), .C(rst), .Y(u2__0remLo_451_0__264_));
AOI21X1 AOI21X1_1418 ( .A(u2__abc_52138_new_n12255_), .B(u2__abc_52138_new_n12256_), .C(rst), .Y(u2__0remLo_451_0__265_));
AOI21X1 AOI21X1_1419 ( .A(u2__abc_52138_new_n12258_), .B(u2__abc_52138_new_n12259_), .C(rst), .Y(u2__0remLo_451_0__266_));
AOI21X1 AOI21X1_142 ( .A(u2__abc_52138_new_n6336_), .B(u2__abc_52138_new_n6163_), .C(u2__abc_52138_new_n6166_), .Y(u2__abc_52138_new_n6337_));
AOI21X1 AOI21X1_1420 ( .A(u2__abc_52138_new_n12261_), .B(u2__abc_52138_new_n12262_), .C(rst), .Y(u2__0remLo_451_0__267_));
AOI21X1 AOI21X1_1421 ( .A(u2__abc_52138_new_n12264_), .B(u2__abc_52138_new_n12265_), .C(rst), .Y(u2__0remLo_451_0__268_));
AOI21X1 AOI21X1_1422 ( .A(u2__abc_52138_new_n12267_), .B(u2__abc_52138_new_n12268_), .C(rst), .Y(u2__0remLo_451_0__269_));
AOI21X1 AOI21X1_1423 ( .A(u2__abc_52138_new_n12270_), .B(u2__abc_52138_new_n12271_), .C(rst), .Y(u2__0remLo_451_0__270_));
AOI21X1 AOI21X1_1424 ( .A(u2__abc_52138_new_n12273_), .B(u2__abc_52138_new_n12274_), .C(rst), .Y(u2__0remLo_451_0__271_));
AOI21X1 AOI21X1_1425 ( .A(u2__abc_52138_new_n12276_), .B(u2__abc_52138_new_n12277_), .C(rst), .Y(u2__0remLo_451_0__272_));
AOI21X1 AOI21X1_1426 ( .A(u2__abc_52138_new_n12279_), .B(u2__abc_52138_new_n12280_), .C(rst), .Y(u2__0remLo_451_0__273_));
AOI21X1 AOI21X1_1427 ( .A(u2__abc_52138_new_n12282_), .B(u2__abc_52138_new_n12283_), .C(rst), .Y(u2__0remLo_451_0__274_));
AOI21X1 AOI21X1_1428 ( .A(u2__abc_52138_new_n12285_), .B(u2__abc_52138_new_n12286_), .C(rst), .Y(u2__0remLo_451_0__275_));
AOI21X1 AOI21X1_1429 ( .A(u2__abc_52138_new_n12288_), .B(u2__abc_52138_new_n12289_), .C(rst), .Y(u2__0remLo_451_0__276_));
AOI21X1 AOI21X1_143 ( .A(u2__abc_52138_new_n6339_), .B(u2__abc_52138_new_n6155_), .C(u2__abc_52138_new_n6148_), .Y(u2__abc_52138_new_n6340_));
AOI21X1 AOI21X1_1430 ( .A(u2__abc_52138_new_n12291_), .B(u2__abc_52138_new_n12292_), .C(rst), .Y(u2__0remLo_451_0__277_));
AOI21X1 AOI21X1_1431 ( .A(u2__abc_52138_new_n12294_), .B(u2__abc_52138_new_n12295_), .C(rst), .Y(u2__0remLo_451_0__278_));
AOI21X1 AOI21X1_1432 ( .A(u2__abc_52138_new_n12297_), .B(u2__abc_52138_new_n12298_), .C(rst), .Y(u2__0remLo_451_0__279_));
AOI21X1 AOI21X1_1433 ( .A(u2__abc_52138_new_n12300_), .B(u2__abc_52138_new_n12301_), .C(rst), .Y(u2__0remLo_451_0__280_));
AOI21X1 AOI21X1_1434 ( .A(u2__abc_52138_new_n12303_), .B(u2__abc_52138_new_n12304_), .C(rst), .Y(u2__0remLo_451_0__281_));
AOI21X1 AOI21X1_1435 ( .A(u2__abc_52138_new_n12306_), .B(u2__abc_52138_new_n12307_), .C(rst), .Y(u2__0remLo_451_0__282_));
AOI21X1 AOI21X1_1436 ( .A(u2__abc_52138_new_n12309_), .B(u2__abc_52138_new_n12310_), .C(rst), .Y(u2__0remLo_451_0__283_));
AOI21X1 AOI21X1_1437 ( .A(u2__abc_52138_new_n12312_), .B(u2__abc_52138_new_n12313_), .C(rst), .Y(u2__0remLo_451_0__284_));
AOI21X1 AOI21X1_1438 ( .A(u2__abc_52138_new_n12315_), .B(u2__abc_52138_new_n12316_), .C(rst), .Y(u2__0remLo_451_0__285_));
AOI21X1 AOI21X1_1439 ( .A(u2__abc_52138_new_n12318_), .B(u2__abc_52138_new_n12319_), .C(rst), .Y(u2__0remLo_451_0__286_));
AOI21X1 AOI21X1_144 ( .A(u2__abc_52138_new_n6145_), .B(u2__abc_52138_new_n6139_), .C(u2__abc_52138_new_n6144_), .Y(u2__abc_52138_new_n6341_));
AOI21X1 AOI21X1_1440 ( .A(u2__abc_52138_new_n12321_), .B(u2__abc_52138_new_n12322_), .C(rst), .Y(u2__0remLo_451_0__287_));
AOI21X1 AOI21X1_1441 ( .A(u2__abc_52138_new_n12324_), .B(u2__abc_52138_new_n12325_), .C(rst), .Y(u2__0remLo_451_0__288_));
AOI21X1 AOI21X1_1442 ( .A(u2__abc_52138_new_n12327_), .B(u2__abc_52138_new_n12328_), .C(rst), .Y(u2__0remLo_451_0__289_));
AOI21X1 AOI21X1_1443 ( .A(u2__abc_52138_new_n12330_), .B(u2__abc_52138_new_n12331_), .C(rst), .Y(u2__0remLo_451_0__290_));
AOI21X1 AOI21X1_1444 ( .A(u2__abc_52138_new_n12333_), .B(u2__abc_52138_new_n12334_), .C(rst), .Y(u2__0remLo_451_0__291_));
AOI21X1 AOI21X1_1445 ( .A(u2__abc_52138_new_n12336_), .B(u2__abc_52138_new_n12337_), .C(rst), .Y(u2__0remLo_451_0__292_));
AOI21X1 AOI21X1_1446 ( .A(u2__abc_52138_new_n12339_), .B(u2__abc_52138_new_n12340_), .C(rst), .Y(u2__0remLo_451_0__293_));
AOI21X1 AOI21X1_1447 ( .A(u2__abc_52138_new_n12342_), .B(u2__abc_52138_new_n12343_), .C(rst), .Y(u2__0remLo_451_0__294_));
AOI21X1 AOI21X1_1448 ( .A(u2__abc_52138_new_n12345_), .B(u2__abc_52138_new_n12346_), .C(rst), .Y(u2__0remLo_451_0__295_));
AOI21X1 AOI21X1_1449 ( .A(u2__abc_52138_new_n12348_), .B(u2__abc_52138_new_n12349_), .C(rst), .Y(u2__0remLo_451_0__296_));
AOI21X1 AOI21X1_145 ( .A(u2__abc_52138_new_n6338_), .B(u2__abc_52138_new_n6158_), .C(u2__abc_52138_new_n6342_), .Y(u2__abc_52138_new_n6343_));
AOI21X1 AOI21X1_1450 ( .A(u2__abc_52138_new_n12351_), .B(u2__abc_52138_new_n12352_), .C(rst), .Y(u2__0remLo_451_0__297_));
AOI21X1 AOI21X1_1451 ( .A(u2__abc_52138_new_n12354_), .B(u2__abc_52138_new_n12355_), .C(rst), .Y(u2__0remLo_451_0__298_));
AOI21X1 AOI21X1_1452 ( .A(u2__abc_52138_new_n12357_), .B(u2__abc_52138_new_n12358_), .C(rst), .Y(u2__0remLo_451_0__299_));
AOI21X1 AOI21X1_1453 ( .A(u2__abc_52138_new_n12360_), .B(u2__abc_52138_new_n12361_), .C(rst), .Y(u2__0remLo_451_0__300_));
AOI21X1 AOI21X1_1454 ( .A(u2__abc_52138_new_n12363_), .B(u2__abc_52138_new_n12364_), .C(rst), .Y(u2__0remLo_451_0__301_));
AOI21X1 AOI21X1_1455 ( .A(u2__abc_52138_new_n12366_), .B(u2__abc_52138_new_n12367_), .C(rst), .Y(u2__0remLo_451_0__302_));
AOI21X1 AOI21X1_1456 ( .A(u2__abc_52138_new_n12369_), .B(u2__abc_52138_new_n12370_), .C(rst), .Y(u2__0remLo_451_0__303_));
AOI21X1 AOI21X1_1457 ( .A(u2__abc_52138_new_n12372_), .B(u2__abc_52138_new_n12373_), .C(rst), .Y(u2__0remLo_451_0__304_));
AOI21X1 AOI21X1_1458 ( .A(u2__abc_52138_new_n12375_), .B(u2__abc_52138_new_n12376_), .C(rst), .Y(u2__0remLo_451_0__305_));
AOI21X1 AOI21X1_1459 ( .A(u2__abc_52138_new_n12378_), .B(u2__abc_52138_new_n12379_), .C(rst), .Y(u2__0remLo_451_0__306_));
AOI21X1 AOI21X1_146 ( .A(u2__abc_52138_new_n6313_), .B(u2__abc_52138_new_n6307_), .C(u2__abc_52138_new_n6312_), .Y(u2__abc_52138_new_n6349_));
AOI21X1 AOI21X1_1460 ( .A(u2__abc_52138_new_n12381_), .B(u2__abc_52138_new_n12382_), .C(rst), .Y(u2__0remLo_451_0__307_));
AOI21X1 AOI21X1_1461 ( .A(u2__abc_52138_new_n12384_), .B(u2__abc_52138_new_n12385_), .C(rst), .Y(u2__0remLo_451_0__308_));
AOI21X1 AOI21X1_1462 ( .A(u2__abc_52138_new_n12387_), .B(u2__abc_52138_new_n12388_), .C(rst), .Y(u2__0remLo_451_0__309_));
AOI21X1 AOI21X1_1463 ( .A(u2__abc_52138_new_n12390_), .B(u2__abc_52138_new_n12391_), .C(rst), .Y(u2__0remLo_451_0__310_));
AOI21X1 AOI21X1_1464 ( .A(u2__abc_52138_new_n12393_), .B(u2__abc_52138_new_n12394_), .C(rst), .Y(u2__0remLo_451_0__311_));
AOI21X1 AOI21X1_1465 ( .A(u2__abc_52138_new_n12396_), .B(u2__abc_52138_new_n12397_), .C(rst), .Y(u2__0remLo_451_0__312_));
AOI21X1 AOI21X1_1466 ( .A(u2__abc_52138_new_n12399_), .B(u2__abc_52138_new_n12400_), .C(rst), .Y(u2__0remLo_451_0__313_));
AOI21X1 AOI21X1_1467 ( .A(u2__abc_52138_new_n12402_), .B(u2__abc_52138_new_n12403_), .C(rst), .Y(u2__0remLo_451_0__314_));
AOI21X1 AOI21X1_1468 ( .A(u2__abc_52138_new_n12405_), .B(u2__abc_52138_new_n12406_), .C(rst), .Y(u2__0remLo_451_0__315_));
AOI21X1 AOI21X1_1469 ( .A(u2__abc_52138_new_n12408_), .B(u2__abc_52138_new_n12409_), .C(rst), .Y(u2__0remLo_451_0__316_));
AOI21X1 AOI21X1_147 ( .A(u2__abc_52138_new_n6350_), .B(u2__abc_52138_new_n6295_), .C(u2__abc_52138_new_n6299_), .Y(u2__abc_52138_new_n6351_));
AOI21X1 AOI21X1_1470 ( .A(u2__abc_52138_new_n12411_), .B(u2__abc_52138_new_n12412_), .C(rst), .Y(u2__0remLo_451_0__317_));
AOI21X1 AOI21X1_1471 ( .A(u2__abc_52138_new_n12414_), .B(u2__abc_52138_new_n12415_), .C(rst), .Y(u2__0remLo_451_0__318_));
AOI21X1 AOI21X1_1472 ( .A(u2__abc_52138_new_n12417_), .B(u2__abc_52138_new_n12418_), .C(rst), .Y(u2__0remLo_451_0__319_));
AOI21X1 AOI21X1_1473 ( .A(u2__abc_52138_new_n12420_), .B(u2__abc_52138_new_n12421_), .C(rst), .Y(u2__0remLo_451_0__320_));
AOI21X1 AOI21X1_1474 ( .A(u2__abc_52138_new_n12423_), .B(u2__abc_52138_new_n12424_), .C(rst), .Y(u2__0remLo_451_0__321_));
AOI21X1 AOI21X1_1475 ( .A(u2__abc_52138_new_n12426_), .B(u2__abc_52138_new_n12427_), .C(rst), .Y(u2__0remLo_451_0__322_));
AOI21X1 AOI21X1_1476 ( .A(u2__abc_52138_new_n12429_), .B(u2__abc_52138_new_n12430_), .C(rst), .Y(u2__0remLo_451_0__323_));
AOI21X1 AOI21X1_1477 ( .A(u2__abc_52138_new_n12432_), .B(u2__abc_52138_new_n12433_), .C(rst), .Y(u2__0remLo_451_0__324_));
AOI21X1 AOI21X1_1478 ( .A(u2__abc_52138_new_n12435_), .B(u2__abc_52138_new_n12436_), .C(rst), .Y(u2__0remLo_451_0__325_));
AOI21X1 AOI21X1_1479 ( .A(u2__abc_52138_new_n12438_), .B(u2__abc_52138_new_n12439_), .C(rst), .Y(u2__0remLo_451_0__326_));
AOI21X1 AOI21X1_148 ( .A(u2__abc_52138_new_n6358_), .B(u2__abc_52138_new_n6204_), .C(u2__abc_52138_new_n6197_), .Y(u2__abc_52138_new_n6359_));
AOI21X1 AOI21X1_1480 ( .A(u2__abc_52138_new_n12441_), .B(u2__abc_52138_new_n12442_), .C(rst), .Y(u2__0remLo_451_0__327_));
AOI21X1 AOI21X1_1481 ( .A(u2__abc_52138_new_n12444_), .B(u2__abc_52138_new_n12445_), .C(rst), .Y(u2__0remLo_451_0__328_));
AOI21X1 AOI21X1_1482 ( .A(u2__abc_52138_new_n12447_), .B(u2__abc_52138_new_n12448_), .C(rst), .Y(u2__0remLo_451_0__329_));
AOI21X1 AOI21X1_1483 ( .A(u2__abc_52138_new_n12450_), .B(u2__abc_52138_new_n12451_), .C(rst), .Y(u2__0remLo_451_0__330_));
AOI21X1 AOI21X1_1484 ( .A(u2__abc_52138_new_n12453_), .B(u2__abc_52138_new_n12454_), .C(rst), .Y(u2__0remLo_451_0__331_));
AOI21X1 AOI21X1_1485 ( .A(u2__abc_52138_new_n12456_), .B(u2__abc_52138_new_n12457_), .C(rst), .Y(u2__0remLo_451_0__332_));
AOI21X1 AOI21X1_1486 ( .A(u2__abc_52138_new_n12459_), .B(u2__abc_52138_new_n12460_), .C(rst), .Y(u2__0remLo_451_0__333_));
AOI21X1 AOI21X1_1487 ( .A(u2__abc_52138_new_n12462_), .B(u2__abc_52138_new_n12463_), .C(rst), .Y(u2__0remLo_451_0__334_));
AOI21X1 AOI21X1_1488 ( .A(u2__abc_52138_new_n12465_), .B(u2__abc_52138_new_n12466_), .C(rst), .Y(u2__0remLo_451_0__335_));
AOI21X1 AOI21X1_1489 ( .A(u2__abc_52138_new_n12468_), .B(u2__abc_52138_new_n12469_), .C(rst), .Y(u2__0remLo_451_0__336_));
AOI21X1 AOI21X1_149 ( .A(u2__abc_52138_new_n6360_), .B(u2__abc_52138_new_n6188_), .C(u2__abc_52138_new_n6191_), .Y(u2__abc_52138_new_n6361_));
AOI21X1 AOI21X1_1490 ( .A(u2__abc_52138_new_n12471_), .B(u2__abc_52138_new_n12472_), .C(rst), .Y(u2__0remLo_451_0__337_));
AOI21X1 AOI21X1_1491 ( .A(u2__abc_52138_new_n12474_), .B(u2__abc_52138_new_n12475_), .C(rst), .Y(u2__0remLo_451_0__338_));
AOI21X1 AOI21X1_1492 ( .A(u2__abc_52138_new_n12477_), .B(u2__abc_52138_new_n12478_), .C(rst), .Y(u2__0remLo_451_0__339_));
AOI21X1 AOI21X1_1493 ( .A(u2__abc_52138_new_n12480_), .B(u2__abc_52138_new_n12481_), .C(rst), .Y(u2__0remLo_451_0__340_));
AOI21X1 AOI21X1_1494 ( .A(u2__abc_52138_new_n12483_), .B(u2__abc_52138_new_n12484_), .C(rst), .Y(u2__0remLo_451_0__341_));
AOI21X1 AOI21X1_1495 ( .A(u2__abc_52138_new_n12486_), .B(u2__abc_52138_new_n12487_), .C(rst), .Y(u2__0remLo_451_0__342_));
AOI21X1 AOI21X1_1496 ( .A(u2__abc_52138_new_n12489_), .B(u2__abc_52138_new_n12490_), .C(rst), .Y(u2__0remLo_451_0__343_));
AOI21X1 AOI21X1_1497 ( .A(u2__abc_52138_new_n12492_), .B(u2__abc_52138_new_n12493_), .C(rst), .Y(u2__0remLo_451_0__344_));
AOI21X1 AOI21X1_1498 ( .A(u2__abc_52138_new_n12495_), .B(u2__abc_52138_new_n12496_), .C(rst), .Y(u2__0remLo_451_0__345_));
AOI21X1 AOI21X1_1499 ( .A(u2__abc_52138_new_n12498_), .B(u2__abc_52138_new_n12499_), .C(rst), .Y(u2__0remLo_451_0__346_));
AOI21X1 AOI21X1_15 ( .A(u2__abc_52138_new_n3202_), .B(u2__abc_52138_new_n3165_), .C(u2__abc_52138_new_n3203_), .Y(u2__abc_52138_new_n3204_));
AOI21X1 AOI21X1_150 ( .A(u2__abc_52138_new_n6368_), .B(u2__abc_52138_new_n6211_), .C(u2__abc_52138_new_n6216_), .Y(u2__abc_52138_new_n6369_));
AOI21X1 AOI21X1_1500 ( .A(u2__abc_52138_new_n12501_), .B(u2__abc_52138_new_n12502_), .C(rst), .Y(u2__0remLo_451_0__347_));
AOI21X1 AOI21X1_1501 ( .A(u2__abc_52138_new_n12504_), .B(u2__abc_52138_new_n12505_), .C(rst), .Y(u2__0remLo_451_0__348_));
AOI21X1 AOI21X1_1502 ( .A(u2__abc_52138_new_n12507_), .B(u2__abc_52138_new_n12508_), .C(rst), .Y(u2__0remLo_451_0__349_));
AOI21X1 AOI21X1_1503 ( .A(u2__abc_52138_new_n12510_), .B(u2__abc_52138_new_n12511_), .C(rst), .Y(u2__0remLo_451_0__350_));
AOI21X1 AOI21X1_1504 ( .A(u2__abc_52138_new_n12513_), .B(u2__abc_52138_new_n12514_), .C(rst), .Y(u2__0remLo_451_0__351_));
AOI21X1 AOI21X1_1505 ( .A(u2__abc_52138_new_n12516_), .B(u2__abc_52138_new_n12517_), .C(rst), .Y(u2__0remLo_451_0__352_));
AOI21X1 AOI21X1_1506 ( .A(u2__abc_52138_new_n12519_), .B(u2__abc_52138_new_n12520_), .C(rst), .Y(u2__0remLo_451_0__353_));
AOI21X1 AOI21X1_1507 ( .A(u2__abc_52138_new_n12522_), .B(u2__abc_52138_new_n12523_), .C(rst), .Y(u2__0remLo_451_0__354_));
AOI21X1 AOI21X1_1508 ( .A(u2__abc_52138_new_n12525_), .B(u2__abc_52138_new_n12526_), .C(rst), .Y(u2__0remLo_451_0__355_));
AOI21X1 AOI21X1_1509 ( .A(u2__abc_52138_new_n12528_), .B(u2__abc_52138_new_n12529_), .C(rst), .Y(u2__0remLo_451_0__356_));
AOI21X1 AOI21X1_151 ( .A(u2__abc_52138_new_n6364_), .B(u2__abc_52138_new_n6367_), .C(u2__abc_52138_new_n6370_), .Y(u2__abc_52138_new_n6371_));
AOI21X1 AOI21X1_1510 ( .A(u2__abc_52138_new_n12531_), .B(u2__abc_52138_new_n12532_), .C(rst), .Y(u2__0remLo_451_0__357_));
AOI21X1 AOI21X1_1511 ( .A(u2__abc_52138_new_n12534_), .B(u2__abc_52138_new_n12535_), .C(rst), .Y(u2__0remLo_451_0__358_));
AOI21X1 AOI21X1_1512 ( .A(u2__abc_52138_new_n12537_), .B(u2__abc_52138_new_n12538_), .C(rst), .Y(u2__0remLo_451_0__359_));
AOI21X1 AOI21X1_1513 ( .A(u2__abc_52138_new_n12540_), .B(u2__abc_52138_new_n12541_), .C(rst), .Y(u2__0remLo_451_0__360_));
AOI21X1 AOI21X1_1514 ( .A(u2__abc_52138_new_n12543_), .B(u2__abc_52138_new_n12544_), .C(rst), .Y(u2__0remLo_451_0__361_));
AOI21X1 AOI21X1_1515 ( .A(u2__abc_52138_new_n12546_), .B(u2__abc_52138_new_n12547_), .C(rst), .Y(u2__0remLo_451_0__362_));
AOI21X1 AOI21X1_1516 ( .A(u2__abc_52138_new_n12549_), .B(u2__abc_52138_new_n12550_), .C(rst), .Y(u2__0remLo_451_0__363_));
AOI21X1 AOI21X1_1517 ( .A(u2__abc_52138_new_n12552_), .B(u2__abc_52138_new_n12553_), .C(rst), .Y(u2__0remLo_451_0__364_));
AOI21X1 AOI21X1_1518 ( .A(u2__abc_52138_new_n12555_), .B(u2__abc_52138_new_n12556_), .C(rst), .Y(u2__0remLo_451_0__365_));
AOI21X1 AOI21X1_1519 ( .A(u2__abc_52138_new_n12558_), .B(u2__abc_52138_new_n12559_), .C(rst), .Y(u2__0remLo_451_0__366_));
AOI21X1 AOI21X1_152 ( .A(u2__abc_52138_new_n6373_), .B(u2__abc_52138_new_n6235_), .C(u2__abc_52138_new_n6238_), .Y(u2__abc_52138_new_n6374_));
AOI21X1 AOI21X1_1520 ( .A(u2__abc_52138_new_n12561_), .B(u2__abc_52138_new_n12562_), .C(rst), .Y(u2__0remLo_451_0__367_));
AOI21X1 AOI21X1_1521 ( .A(u2__abc_52138_new_n12564_), .B(u2__abc_52138_new_n12565_), .C(rst), .Y(u2__0remLo_451_0__368_));
AOI21X1 AOI21X1_1522 ( .A(u2__abc_52138_new_n12567_), .B(u2__abc_52138_new_n12568_), .C(rst), .Y(u2__0remLo_451_0__369_));
AOI21X1 AOI21X1_1523 ( .A(u2__abc_52138_new_n12570_), .B(u2__abc_52138_new_n12571_), .C(rst), .Y(u2__0remLo_451_0__370_));
AOI21X1 AOI21X1_1524 ( .A(u2__abc_52138_new_n12573_), .B(u2__abc_52138_new_n12574_), .C(rst), .Y(u2__0remLo_451_0__371_));
AOI21X1 AOI21X1_1525 ( .A(u2__abc_52138_new_n12576_), .B(u2__abc_52138_new_n12577_), .C(rst), .Y(u2__0remLo_451_0__372_));
AOI21X1 AOI21X1_1526 ( .A(u2__abc_52138_new_n12579_), .B(u2__abc_52138_new_n12580_), .C(rst), .Y(u2__0remLo_451_0__373_));
AOI21X1 AOI21X1_1527 ( .A(u2__abc_52138_new_n12582_), .B(u2__abc_52138_new_n12583_), .C(rst), .Y(u2__0remLo_451_0__374_));
AOI21X1 AOI21X1_1528 ( .A(u2__abc_52138_new_n12585_), .B(u2__abc_52138_new_n12586_), .C(rst), .Y(u2__0remLo_451_0__375_));
AOI21X1 AOI21X1_1529 ( .A(u2__abc_52138_new_n12588_), .B(u2__abc_52138_new_n12589_), .C(rst), .Y(u2__0remLo_451_0__376_));
AOI21X1 AOI21X1_153 ( .A(u2__abc_52138_new_n6375_), .B(u2__abc_52138_new_n6246_), .C(u2__abc_52138_new_n6249_), .Y(u2__abc_52138_new_n6376_));
AOI21X1 AOI21X1_1530 ( .A(u2__abc_52138_new_n12591_), .B(u2__abc_52138_new_n12592_), .C(rst), .Y(u2__0remLo_451_0__377_));
AOI21X1 AOI21X1_1531 ( .A(u2__abc_52138_new_n12594_), .B(u2__abc_52138_new_n12595_), .C(rst), .Y(u2__0remLo_451_0__378_));
AOI21X1 AOI21X1_1532 ( .A(u2__abc_52138_new_n12597_), .B(u2__abc_52138_new_n12598_), .C(rst), .Y(u2__0remLo_451_0__379_));
AOI21X1 AOI21X1_1533 ( .A(u2__abc_52138_new_n12600_), .B(u2__abc_52138_new_n12601_), .C(rst), .Y(u2__0remLo_451_0__380_));
AOI21X1 AOI21X1_1534 ( .A(u2__abc_52138_new_n12603_), .B(u2__abc_52138_new_n12604_), .C(rst), .Y(u2__0remLo_451_0__381_));
AOI21X1 AOI21X1_1535 ( .A(u2__abc_52138_new_n12606_), .B(u2__abc_52138_new_n12607_), .C(rst), .Y(u2__0remLo_451_0__382_));
AOI21X1 AOI21X1_1536 ( .A(u2__abc_52138_new_n12609_), .B(u2__abc_52138_new_n12610_), .C(rst), .Y(u2__0remLo_451_0__383_));
AOI21X1 AOI21X1_1537 ( .A(u2__abc_52138_new_n12612_), .B(u2__abc_52138_new_n12613_), .C(rst), .Y(u2__0remLo_451_0__384_));
AOI21X1 AOI21X1_1538 ( .A(u2__abc_52138_new_n12615_), .B(u2__abc_52138_new_n12616_), .C(rst), .Y(u2__0remLo_451_0__385_));
AOI21X1 AOI21X1_1539 ( .A(u2__abc_52138_new_n12618_), .B(u2__abc_52138_new_n12619_), .C(rst), .Y(u2__0remLo_451_0__386_));
AOI21X1 AOI21X1_154 ( .A(u2__abc_52138_new_n6378_), .B(u2__abc_52138_new_n6274_), .C(u2__abc_52138_new_n6267_), .Y(u2__abc_52138_new_n6379_));
AOI21X1 AOI21X1_1540 ( .A(u2__abc_52138_new_n12621_), .B(u2__abc_52138_new_n12622_), .C(rst), .Y(u2__0remLo_451_0__387_));
AOI21X1 AOI21X1_1541 ( .A(u2__abc_52138_new_n12624_), .B(u2__abc_52138_new_n12625_), .C(rst), .Y(u2__0remLo_451_0__388_));
AOI21X1 AOI21X1_1542 ( .A(u2__abc_52138_new_n12627_), .B(u2__abc_52138_new_n12628_), .C(rst), .Y(u2__0remLo_451_0__389_));
AOI21X1 AOI21X1_1543 ( .A(u2__abc_52138_new_n12630_), .B(u2__abc_52138_new_n12631_), .C(rst), .Y(u2__0remLo_451_0__390_));
AOI21X1 AOI21X1_1544 ( .A(u2__abc_52138_new_n12633_), .B(u2__abc_52138_new_n12634_), .C(rst), .Y(u2__0remLo_451_0__391_));
AOI21X1 AOI21X1_1545 ( .A(u2__abc_52138_new_n12636_), .B(u2__abc_52138_new_n12637_), .C(rst), .Y(u2__0remLo_451_0__392_));
AOI21X1 AOI21X1_1546 ( .A(u2__abc_52138_new_n12639_), .B(u2__abc_52138_new_n12640_), .C(rst), .Y(u2__0remLo_451_0__393_));
AOI21X1 AOI21X1_1547 ( .A(u2__abc_52138_new_n12642_), .B(u2__abc_52138_new_n12643_), .C(rst), .Y(u2__0remLo_451_0__394_));
AOI21X1 AOI21X1_1548 ( .A(u2__abc_52138_new_n12645_), .B(u2__abc_52138_new_n12646_), .C(rst), .Y(u2__0remLo_451_0__395_));
AOI21X1 AOI21X1_1549 ( .A(u2__abc_52138_new_n12648_), .B(u2__abc_52138_new_n12649_), .C(rst), .Y(u2__0remLo_451_0__396_));
AOI21X1 AOI21X1_155 ( .A(u2__abc_52138_new_n6380_), .B(u2__abc_52138_new_n6258_), .C(u2__abc_52138_new_n6263_), .Y(u2__abc_52138_new_n6381_));
AOI21X1 AOI21X1_1550 ( .A(u2__abc_52138_new_n12651_), .B(u2__abc_52138_new_n12652_), .C(rst), .Y(u2__0remLo_451_0__397_));
AOI21X1 AOI21X1_1551 ( .A(u2__abc_52138_new_n12654_), .B(u2__abc_52138_new_n12655_), .C(rst), .Y(u2__0remLo_451_0__398_));
AOI21X1 AOI21X1_1552 ( .A(u2__abc_52138_new_n12657_), .B(u2__abc_52138_new_n12658_), .C(rst), .Y(u2__0remLo_451_0__399_));
AOI21X1 AOI21X1_1553 ( .A(u2__abc_52138_new_n12660_), .B(u2__abc_52138_new_n12661_), .C(rst), .Y(u2__0remLo_451_0__400_));
AOI21X1 AOI21X1_1554 ( .A(u2__abc_52138_new_n12663_), .B(u2__abc_52138_new_n12664_), .C(rst), .Y(u2__0remLo_451_0__401_));
AOI21X1 AOI21X1_1555 ( .A(u2__abc_52138_new_n12666_), .B(u2__abc_52138_new_n12667_), .C(rst), .Y(u2__0remLo_451_0__402_));
AOI21X1 AOI21X1_1556 ( .A(u2__abc_52138_new_n12669_), .B(u2__abc_52138_new_n12670_), .C(rst), .Y(u2__0remLo_451_0__403_));
AOI21X1 AOI21X1_1557 ( .A(u2__abc_52138_new_n12672_), .B(u2__abc_52138_new_n12673_), .C(rst), .Y(u2__0remLo_451_0__404_));
AOI21X1 AOI21X1_1558 ( .A(u2__abc_52138_new_n12675_), .B(u2__abc_52138_new_n12676_), .C(rst), .Y(u2__0remLo_451_0__405_));
AOI21X1 AOI21X1_1559 ( .A(u2__abc_52138_new_n12678_), .B(u2__abc_52138_new_n12679_), .C(rst), .Y(u2__0remLo_451_0__406_));
AOI21X1 AOI21X1_156 ( .A(u2__abc_52138_new_n6377_), .B(u2__abc_52138_new_n6277_), .C(u2__abc_52138_new_n6382_), .Y(u2__abc_52138_new_n6383_));
AOI21X1 AOI21X1_1560 ( .A(u2__abc_52138_new_n12681_), .B(u2__abc_52138_new_n12682_), .C(rst), .Y(u2__0remLo_451_0__407_));
AOI21X1 AOI21X1_1561 ( .A(u2__abc_52138_new_n12684_), .B(u2__abc_52138_new_n12685_), .C(rst), .Y(u2__0remLo_451_0__408_));
AOI21X1 AOI21X1_1562 ( .A(u2__abc_52138_new_n12687_), .B(u2__abc_52138_new_n12688_), .C(rst), .Y(u2__0remLo_451_0__409_));
AOI21X1 AOI21X1_1563 ( .A(u2__abc_52138_new_n12690_), .B(u2__abc_52138_new_n12691_), .C(rst), .Y(u2__0remLo_451_0__410_));
AOI21X1 AOI21X1_1564 ( .A(u2__abc_52138_new_n12693_), .B(u2__abc_52138_new_n12694_), .C(rst), .Y(u2__0remLo_451_0__411_));
AOI21X1 AOI21X1_1565 ( .A(u2__abc_52138_new_n12696_), .B(u2__abc_52138_new_n12697_), .C(rst), .Y(u2__0remLo_451_0__412_));
AOI21X1 AOI21X1_1566 ( .A(u2__abc_52138_new_n12699_), .B(u2__abc_52138_new_n12700_), .C(rst), .Y(u2__0remLo_451_0__413_));
AOI21X1 AOI21X1_1567 ( .A(u2__abc_52138_new_n12702_), .B(u2__abc_52138_new_n12703_), .C(rst), .Y(u2__0remLo_451_0__414_));
AOI21X1 AOI21X1_1568 ( .A(u2__abc_52138_new_n12705_), .B(u2__abc_52138_new_n12706_), .C(rst), .Y(u2__0remLo_451_0__415_));
AOI21X1 AOI21X1_1569 ( .A(u2__abc_52138_new_n12708_), .B(u2__abc_52138_new_n12709_), .C(rst), .Y(u2__0remLo_451_0__416_));
AOI21X1 AOI21X1_157 ( .A(u2__abc_52138_new_n6385_), .B(u2__abc_52138_new_n6357_), .C(u2__abc_52138_new_n6333_), .Y(u2__abc_52138_new_n6386_));
AOI21X1 AOI21X1_1570 ( .A(u2__abc_52138_new_n12711_), .B(u2__abc_52138_new_n12712_), .C(rst), .Y(u2__0remLo_451_0__417_));
AOI21X1 AOI21X1_1571 ( .A(u2__abc_52138_new_n12714_), .B(u2__abc_52138_new_n12715_), .C(rst), .Y(u2__0remLo_451_0__418_));
AOI21X1 AOI21X1_1572 ( .A(u2__abc_52138_new_n12717_), .B(u2__abc_52138_new_n12718_), .C(rst), .Y(u2__0remLo_451_0__419_));
AOI21X1 AOI21X1_1573 ( .A(u2__abc_52138_new_n12720_), .B(u2__abc_52138_new_n12721_), .C(rst), .Y(u2__0remLo_451_0__420_));
AOI21X1 AOI21X1_1574 ( .A(u2__abc_52138_new_n12723_), .B(u2__abc_52138_new_n12724_), .C(rst), .Y(u2__0remLo_451_0__421_));
AOI21X1 AOI21X1_1575 ( .A(u2__abc_52138_new_n12726_), .B(u2__abc_52138_new_n12727_), .C(rst), .Y(u2__0remLo_451_0__422_));
AOI21X1 AOI21X1_1576 ( .A(u2__abc_52138_new_n12729_), .B(u2__abc_52138_new_n12730_), .C(rst), .Y(u2__0remLo_451_0__423_));
AOI21X1 AOI21X1_1577 ( .A(u2__abc_52138_new_n12732_), .B(u2__abc_52138_new_n12733_), .C(rst), .Y(u2__0remLo_451_0__424_));
AOI21X1 AOI21X1_1578 ( .A(u2__abc_52138_new_n12735_), .B(u2__abc_52138_new_n12736_), .C(rst), .Y(u2__0remLo_451_0__425_));
AOI21X1 AOI21X1_1579 ( .A(u2__abc_52138_new_n12738_), .B(u2__abc_52138_new_n12739_), .C(rst), .Y(u2__0remLo_451_0__426_));
AOI21X1 AOI21X1_158 ( .A(u2__abc_52138_new_n6390_), .B(u2__abc_52138_new_n6118_), .C(u2__abc_52138_new_n6391_), .Y(u2__abc_52138_new_n6392_));
AOI21X1 AOI21X1_1580 ( .A(u2__abc_52138_new_n12741_), .B(u2__abc_52138_new_n12742_), .C(rst), .Y(u2__0remLo_451_0__427_));
AOI21X1 AOI21X1_1581 ( .A(u2__abc_52138_new_n12744_), .B(u2__abc_52138_new_n12745_), .C(rst), .Y(u2__0remLo_451_0__428_));
AOI21X1 AOI21X1_1582 ( .A(u2__abc_52138_new_n12747_), .B(u2__abc_52138_new_n12748_), .C(rst), .Y(u2__0remLo_451_0__429_));
AOI21X1 AOI21X1_1583 ( .A(u2__abc_52138_new_n12750_), .B(u2__abc_52138_new_n12751_), .C(rst), .Y(u2__0remLo_451_0__430_));
AOI21X1 AOI21X1_1584 ( .A(u2__abc_52138_new_n12753_), .B(u2__abc_52138_new_n12754_), .C(rst), .Y(u2__0remLo_451_0__431_));
AOI21X1 AOI21X1_1585 ( .A(u2__abc_52138_new_n12756_), .B(u2__abc_52138_new_n12757_), .C(rst), .Y(u2__0remLo_451_0__432_));
AOI21X1 AOI21X1_1586 ( .A(u2__abc_52138_new_n12759_), .B(u2__abc_52138_new_n12760_), .C(rst), .Y(u2__0remLo_451_0__433_));
AOI21X1 AOI21X1_1587 ( .A(u2__abc_52138_new_n12762_), .B(u2__abc_52138_new_n12763_), .C(rst), .Y(u2__0remLo_451_0__434_));
AOI21X1 AOI21X1_1588 ( .A(u2__abc_52138_new_n12765_), .B(u2__abc_52138_new_n12766_), .C(rst), .Y(u2__0remLo_451_0__435_));
AOI21X1 AOI21X1_1589 ( .A(u2__abc_52138_new_n12768_), .B(u2__abc_52138_new_n12769_), .C(rst), .Y(u2__0remLo_451_0__436_));
AOI21X1 AOI21X1_159 ( .A(u2__abc_52138_new_n6395_), .B(u2__abc_52138_new_n6094_), .C(u2__abc_52138_new_n6396_), .Y(u2__abc_52138_new_n6397_));
AOI21X1 AOI21X1_1590 ( .A(u2__abc_52138_new_n12771_), .B(u2__abc_52138_new_n12772_), .C(rst), .Y(u2__0remLo_451_0__437_));
AOI21X1 AOI21X1_1591 ( .A(u2__abc_52138_new_n12774_), .B(u2__abc_52138_new_n12775_), .C(rst), .Y(u2__0remLo_451_0__438_));
AOI21X1 AOI21X1_1592 ( .A(u2__abc_52138_new_n12777_), .B(u2__abc_52138_new_n12778_), .C(rst), .Y(u2__0remLo_451_0__439_));
AOI21X1 AOI21X1_1593 ( .A(u2__abc_52138_new_n12780_), .B(u2__abc_52138_new_n12781_), .C(rst), .Y(u2__0remLo_451_0__440_));
AOI21X1 AOI21X1_1594 ( .A(u2__abc_52138_new_n12783_), .B(u2__abc_52138_new_n12784_), .C(rst), .Y(u2__0remLo_451_0__441_));
AOI21X1 AOI21X1_1595 ( .A(u2__abc_52138_new_n12786_), .B(u2__abc_52138_new_n12787_), .C(rst), .Y(u2__0remLo_451_0__442_));
AOI21X1 AOI21X1_1596 ( .A(u2__abc_52138_new_n12789_), .B(u2__abc_52138_new_n12790_), .C(rst), .Y(u2__0remLo_451_0__443_));
AOI21X1 AOI21X1_1597 ( .A(u2__abc_52138_new_n12792_), .B(u2__abc_52138_new_n12793_), .C(rst), .Y(u2__0remLo_451_0__444_));
AOI21X1 AOI21X1_1598 ( .A(u2__abc_52138_new_n12795_), .B(u2__abc_52138_new_n12796_), .C(rst), .Y(u2__0remLo_451_0__445_));
AOI21X1 AOI21X1_1599 ( .A(u2__abc_52138_new_n12798_), .B(u2__abc_52138_new_n12799_), .C(rst), .Y(u2__0remLo_451_0__446_));
AOI21X1 AOI21X1_16 ( .A(u2__abc_52138_new_n3209_), .B(u2__abc_52138_new_n3207_), .C(u2__abc_52138_new_n3208_), .Y(u2__abc_52138_new_n3210_));
AOI21X1 AOI21X1_160 ( .A(u2__abc_52138_new_n6401_), .B(u2__abc_52138_new_n6050_), .C(u2__abc_52138_new_n6053_), .Y(u2__abc_52138_new_n6402_));
AOI21X1 AOI21X1_1600 ( .A(u2__abc_52138_new_n12801_), .B(u2__abc_52138_new_n12802_), .C(rst), .Y(u2__0remLo_451_0__447_));
AOI21X1 AOI21X1_1601 ( .A(u2__abc_52138_new_n12804_), .B(u2__abc_52138_new_n12805_), .C(rst), .Y(u2__0remLo_451_0__448_));
AOI21X1 AOI21X1_1602 ( .A(u2__abc_52138_new_n12807_), .B(u2__abc_52138_new_n12808_), .C(rst), .Y(u2__0remLo_451_0__449_));
AOI21X1 AOI21X1_1603 ( .A(u2__abc_52138_new_n12810_), .B(u2__abc_52138_new_n12811_), .C(rst), .Y(u2__0remLo_451_0__450_));
AOI21X1 AOI21X1_1604 ( .A(u2__abc_52138_new_n12813_), .B(u2__abc_52138_new_n12814_), .C(rst), .Y(u2__0remLo_451_0__451_));
AOI21X1 AOI21X1_1605 ( .A(u2__abc_52138_new_n12825_), .B(u2__abc_52138_new_n6462_), .C(u2__abc_52138_new_n12826_), .Y(u2__abc_52138_new_n12827_));
AOI21X1 AOI21X1_1606 ( .A(u2__abc_52138_new_n12820_), .B(u2__abc_52138_new_n12829_), .C(u2__abc_52138_new_n12830_), .Y(u2__abc_52138_new_n12831_));
AOI21X1 AOI21X1_1607 ( .A(u2__abc_52138_new_n12834_), .B(u2__abc_52138_new_n6668_), .C(u2__abc_52138_new_n12832_), .Y(u2__abc_52138_new_n12835_));
AOI21X1 AOI21X1_1608 ( .A(u2__abc_52138_new_n12828_), .B(u2__abc_52138_new_n12822_), .C(u2__abc_52138_new_n12836_), .Y(u2__abc_52138_new_n12837_));
AOI21X1 AOI21X1_1609 ( .A(u2__abc_52138_new_n3169_), .B(u2__abc_52138_new_n12841_), .C(u2__abc_52138_new_n12842_), .Y(u2__abc_52138_new_n12843_));
AOI21X1 AOI21X1_161 ( .A(u2__abc_52138_new_n6408_), .B(u2__abc_52138_new_n6068_), .C(u2__abc_52138_new_n6409_), .Y(u2__abc_52138_new_n6410_));
AOI21X1 AOI21X1_1610 ( .A(u2__abc_52138_new_n6758_), .B(u2__abc_52138_new_n12846_), .C(u2__abc_52138_new_n3214_), .Y(u2__abc_52138_new_n12847_));
AOI21X1 AOI21X1_1611 ( .A(u2__abc_52138_new_n12849_), .B(u2__abc_52138_new_n3122_), .C(u2__abc_52138_new_n3226_), .Y(u2__abc_52138_new_n12850_));
AOI21X1 AOI21X1_1612 ( .A(u2__abc_52138_new_n12852_), .B(u2__abc_52138_new_n3145_), .C(u2__abc_52138_new_n12851_), .Y(u2__abc_52138_new_n12853_));
AOI21X1 AOI21X1_1613 ( .A(u2__abc_52138_new_n12848_), .B(u2__abc_52138_new_n12838_), .C(u2__abc_52138_new_n12854_), .Y(u2__abc_52138_new_n12855_));
AOI21X1 AOI21X1_1614 ( .A(u2__abc_52138_new_n3388_), .B(u2__abc_52138_new_n12859_), .C(u2__abc_52138_new_n12861_), .Y(u2__abc_52138_new_n12862_));
AOI21X1 AOI21X1_1615 ( .A(u2__abc_52138_new_n12863_), .B(u2__abc_52138_new_n3411_), .C(u2__abc_52138_new_n12864_), .Y(u2__abc_52138_new_n12865_));
AOI21X1 AOI21X1_1616 ( .A(u2__abc_52138_new_n3345_), .B(u2__abc_52138_new_n12867_), .C(u2__abc_52138_new_n3457_), .Y(u2__abc_52138_new_n12868_));
AOI21X1 AOI21X1_1617 ( .A(u2__abc_52138_new_n3368_), .B(u2__abc_52138_new_n3461_), .C(u2__abc_52138_new_n3464_), .Y(u2__abc_52138_new_n12869_));
AOI21X1 AOI21X1_1618 ( .A(u2__abc_52138_new_n12866_), .B(u2__abc_52138_new_n3381_), .C(u2__abc_52138_new_n12870_), .Y(u2__abc_52138_new_n12871_));
AOI21X1 AOI21X1_1619 ( .A(u2__abc_52138_new_n12873_), .B(u2__abc_52138_new_n12874_), .C(u2__abc_52138_new_n3474_), .Y(u2__abc_52138_new_n12875_));
AOI21X1 AOI21X1_162 ( .A(u2__abc_52138_new_n5959_), .B(u2__abc_52138_new_n5963_), .C(u2__abc_52138_new_n5956_), .Y(u2__abc_52138_new_n6422_));
AOI21X1 AOI21X1_1620 ( .A(u2__abc_52138_new_n3321_), .B(u2__abc_52138_new_n3479_), .C(u2__abc_52138_new_n12876_), .Y(u2__abc_52138_new_n12877_));
AOI21X1 AOI21X1_1621 ( .A(u2__abc_52138_new_n12879_), .B(u2__abc_52138_new_n3250_), .C(u2__abc_52138_new_n3491_), .Y(u2__abc_52138_new_n12880_));
AOI21X1 AOI21X1_1622 ( .A(u2__abc_52138_new_n3273_), .B(u2__abc_52138_new_n3495_), .C(u2__abc_52138_new_n12881_), .Y(u2__abc_52138_new_n12882_));
AOI21X1 AOI21X1_1623 ( .A(u2__abc_52138_new_n12878_), .B(u2__abc_52138_new_n3286_), .C(u2__abc_52138_new_n12883_), .Y(u2__abc_52138_new_n12884_));
AOI21X1 AOI21X1_1624 ( .A(u2__abc_52138_new_n12856_), .B(u2__abc_52138_new_n12857_), .C(u2__abc_52138_new_n12885_), .Y(u2__abc_52138_new_n12886_));
AOI21X1 AOI21X1_1625 ( .A(u2__abc_52138_new_n12891_), .B(u2__abc_52138_new_n3853_), .C(u2__abc_52138_new_n12892_), .Y(u2__abc_52138_new_n12893_));
AOI21X1 AOI21X1_1626 ( .A(u2__abc_52138_new_n12897_), .B(u2__abc_52138_new_n12895_), .C(u2__abc_52138_new_n3891_), .Y(u2__abc_52138_new_n12898_));
AOI21X1 AOI21X1_1627 ( .A(u2__abc_52138_new_n12901_), .B(u2__abc_52138_new_n7309_), .C(u2__abc_52138_new_n12902_), .Y(u2__abc_52138_new_n12903_));
AOI21X1 AOI21X1_1628 ( .A(u2__abc_52138_new_n7354_), .B(u2__abc_52138_new_n12905_), .C(u2__abc_52138_new_n12906_), .Y(u2__abc_52138_new_n12907_));
AOI21X1 AOI21X1_1629 ( .A(u2__abc_52138_new_n12899_), .B(u2__abc_52138_new_n12889_), .C(u2__abc_52138_new_n12908_), .Y(u2__abc_52138_new_n12909_));
AOI21X1 AOI21X1_163 ( .A(u2__abc_52138_new_n6424_), .B(u2__abc_52138_new_n5947_), .C(u2__abc_52138_new_n5950_), .Y(u2__abc_52138_new_n6425_));
AOI21X1 AOI21X1_1630 ( .A(u2__abc_52138_new_n12910_), .B(u2__abc_52138_new_n7403_), .C(u2__abc_52138_new_n12911_), .Y(u2__abc_52138_new_n12912_));
AOI21X1 AOI21X1_1631 ( .A(u2__abc_52138_new_n3771_), .B(u2__abc_52138_new_n12913_), .C(u2__abc_52138_new_n3919_), .Y(u2__abc_52138_new_n12914_));
AOI21X1 AOI21X1_1632 ( .A(u2__abc_52138_new_n12920_), .B(u2__abc_52138_new_n12918_), .C(u2__abc_52138_new_n3925_), .Y(u2__abc_52138_new_n12921_));
AOI21X1 AOI21X1_1633 ( .A(u2__abc_52138_new_n3930_), .B(u2__abc_52138_new_n3928_), .C(u2__abc_52138_new_n3933_), .Y(u2__abc_52138_new_n12922_));
AOI21X1 AOI21X1_1634 ( .A(u2__abc_52138_new_n6484_), .B(u2__abc_52138_new_n12915_), .C(u2__abc_52138_new_n12923_), .Y(u2__abc_52138_new_n12924_));
AOI21X1 AOI21X1_1635 ( .A(u2__abc_52138_new_n12928_), .B(u2__abc_52138_new_n12927_), .C(u2__abc_52138_new_n3944_), .Y(u2__abc_52138_new_n12929_));
AOI21X1 AOI21X1_1636 ( .A(u2__abc_52138_new_n12930_), .B(u2__abc_52138_new_n3675_), .C(u2__abc_52138_new_n12931_), .Y(u2__abc_52138_new_n12932_));
AOI21X1 AOI21X1_1637 ( .A(u2__abc_52138_new_n12935_), .B(u2__abc_52138_new_n12934_), .C(u2__abc_52138_new_n3959_), .Y(u2__abc_52138_new_n12936_));
AOI21X1 AOI21X1_1638 ( .A(u2__abc_52138_new_n3964_), .B(u2__abc_52138_new_n3962_), .C(u2__abc_52138_new_n12937_), .Y(u2__abc_52138_new_n12938_));
AOI21X1 AOI21X1_1639 ( .A(u2__abc_52138_new_n12933_), .B(u2__abc_52138_new_n7715_), .C(u2__abc_52138_new_n12939_), .Y(u2__abc_52138_new_n12940_));
AOI21X1 AOI21X1_164 ( .A(u2__abc_52138_new_n6427_), .B(u2__abc_52138_new_n6013_), .C(u2__abc_52138_new_n6016_), .Y(u2__abc_52138_new_n6428_));
AOI21X1 AOI21X1_1640 ( .A(u2__abc_52138_new_n12943_), .B(u2__abc_52138_new_n3571_), .C(u2__abc_52138_new_n3976_), .Y(u2__abc_52138_new_n12944_));
AOI21X1 AOI21X1_1641 ( .A(u2__abc_52138_new_n7803_), .B(u2__abc_52138_new_n3983_), .C(u2__abc_52138_new_n3980_), .Y(u2__abc_52138_new_n12945_));
AOI21X1 AOI21X1_1642 ( .A(u2__abc_52138_new_n3526_), .B(u2__abc_52138_new_n3987_), .C(u2__abc_52138_new_n12947_), .Y(u2__abc_52138_new_n12948_));
AOI21X1 AOI21X1_1643 ( .A(u2__abc_52138_new_n6489_), .B(u2__abc_52138_new_n12946_), .C(u2__abc_52138_new_n12949_), .Y(u2__abc_52138_new_n12950_));
AOI21X1 AOI21X1_1644 ( .A(u2__abc_52138_new_n12925_), .B(u2__abc_52138_new_n7892_), .C(u2__abc_52138_new_n12951_), .Y(u2__abc_52138_new_n12952_));
AOI21X1 AOI21X1_1645 ( .A(u2__abc_52138_new_n7939_), .B(u2__abc_52138_new_n12956_), .C(u2__abc_52138_new_n12958_), .Y(u2__abc_52138_new_n12959_));
AOI21X1 AOI21X1_1646 ( .A(u2__abc_52138_new_n4743_), .B(u2__abc_52138_new_n4778_), .C(u2__abc_52138_new_n4781_), .Y(u2__abc_52138_new_n12960_));
AOI21X1 AOI21X1_1647 ( .A(u2__abc_52138_new_n4676_), .B(u2__abc_52138_new_n12962_), .C(u2__abc_52138_new_n4790_), .Y(u2__abc_52138_new_n12963_));
AOI21X1 AOI21X1_1648 ( .A(u2__abc_52138_new_n4699_), .B(u2__abc_52138_new_n4794_), .C(u2__abc_52138_new_n4796_), .Y(u2__abc_52138_new_n12964_));
AOI21X1 AOI21X1_1649 ( .A(u2__abc_52138_new_n12961_), .B(u2__abc_52138_new_n8071_), .C(u2__abc_52138_new_n12965_), .Y(u2__abc_52138_new_n12966_));
AOI21X1 AOI21X1_165 ( .A(u2__abc_52138_new_n6030_), .B(u2__abc_52138_new_n6024_), .C(u2__abc_52138_new_n6027_), .Y(u2__abc_52138_new_n6429_));
AOI21X1 AOI21X1_1650 ( .A(u2__abc_52138_new_n12970_), .B(u2__abc_52138_new_n12968_), .C(u2__abc_52138_new_n12971_), .Y(u2__abc_52138_new_n12972_));
AOI21X1 AOI21X1_1651 ( .A(u2__abc_52138_new_n4629_), .B(u2__abc_52138_new_n4808_), .C(u2__abc_52138_new_n12973_), .Y(u2__abc_52138_new_n12974_));
AOI21X1 AOI21X1_1652 ( .A(u2__abc_52138_new_n4583_), .B(u2__abc_52138_new_n4817_), .C(u2__abc_52138_new_n4819_), .Y(u2__abc_52138_new_n12976_));
AOI21X1 AOI21X1_1653 ( .A(u2__abc_52138_new_n4823_), .B(u2__abc_52138_new_n4606_), .C(u2__abc_52138_new_n4825_), .Y(u2__abc_52138_new_n12977_));
AOI21X1 AOI21X1_1654 ( .A(u2__abc_52138_new_n12975_), .B(u2__abc_52138_new_n4618_), .C(u2__abc_52138_new_n12978_), .Y(u2__abc_52138_new_n12979_));
AOI21X1 AOI21X1_1655 ( .A(u2__abc_52138_new_n12982_), .B(u2__abc_52138_new_n4535_), .C(u2__abc_52138_new_n4834_), .Y(u2__abc_52138_new_n12983_));
AOI21X1 AOI21X1_1656 ( .A(u2__abc_52138_new_n4558_), .B(u2__abc_52138_new_n4839_), .C(u2__abc_52138_new_n4841_), .Y(u2__abc_52138_new_n12984_));
AOI21X1 AOI21X1_1657 ( .A(u2__abc_52138_new_n4846_), .B(u2__abc_52138_new_n4511_), .C(u2__abc_52138_new_n4848_), .Y(u2__abc_52138_new_n12986_));
AOI21X1 AOI21X1_1658 ( .A(u2__abc_52138_new_n4851_), .B(u2__abc_52138_new_n4488_), .C(u2__abc_52138_new_n12987_), .Y(u2__abc_52138_new_n12988_));
AOI21X1 AOI21X1_1659 ( .A(u2__abc_52138_new_n4524_), .B(u2__abc_52138_new_n12985_), .C(u2__abc_52138_new_n12989_), .Y(u2__abc_52138_new_n12990_));
AOI21X1 AOI21X1_166 ( .A(u2__abc_52138_new_n6431_), .B(u2__abc_52138_new_n6006_), .C(u2__abc_52138_new_n5999_), .Y(u2__abc_52138_new_n6432_));
AOI21X1 AOI21X1_1660 ( .A(u2__abc_52138_new_n4866_), .B(u2__abc_52138_new_n4428_), .C(u2__abc_52138_new_n4875_), .Y(u2__abc_52138_new_n12991_));
AOI21X1 AOI21X1_1661 ( .A(u2__abc_52138_new_n12980_), .B(u2__abc_52138_new_n4572_), .C(u2__abc_52138_new_n12992_), .Y(u2__abc_52138_new_n12993_));
AOI21X1 AOI21X1_1662 ( .A(u2__abc_52138_new_n4363_), .B(u2__abc_52138_new_n12996_), .C(u2__abc_52138_new_n12997_), .Y(u2__abc_52138_new_n12998_));
AOI21X1 AOI21X1_1663 ( .A(u2__abc_52138_new_n4341_), .B(u2__abc_52138_new_n4890_), .C(u2__abc_52138_new_n4893_), .Y(u2__abc_52138_new_n12999_));
AOI21X1 AOI21X1_1664 ( .A(u2__abc_52138_new_n4299_), .B(u2__abc_52138_new_n4899_), .C(u2__abc_52138_new_n4901_), .Y(u2__abc_52138_new_n13001_));
AOI21X1 AOI21X1_1665 ( .A(u2__abc_52138_new_n4322_), .B(u2__abc_52138_new_n4907_), .C(u2__abc_52138_new_n13002_), .Y(u2__abc_52138_new_n13003_));
AOI21X1 AOI21X1_1666 ( .A(u2__abc_52138_new_n13000_), .B(u2__abc_52138_new_n8768_), .C(u2__abc_52138_new_n13004_), .Y(u2__abc_52138_new_n13005_));
AOI21X1 AOI21X1_1667 ( .A(u2__abc_52138_new_n13007_), .B(u2__abc_52138_new_n8811_), .C(u2__abc_52138_new_n13008_), .Y(u2__abc_52138_new_n13009_));
AOI21X1 AOI21X1_1668 ( .A(u2__abc_52138_new_n8851_), .B(u2__abc_52138_new_n13011_), .C(u2__abc_52138_new_n13012_), .Y(u2__abc_52138_new_n13013_));
AOI21X1 AOI21X1_1669 ( .A(u2__abc_52138_new_n4929_), .B(u2__abc_52138_new_n4928_), .C(u2__abc_52138_new_n4931_), .Y(u2__abc_52138_new_n13015_));
AOI21X1 AOI21X1_167 ( .A(u2__abc_52138_new_n6433_), .B(u2__abc_52138_new_n5990_), .C(u2__abc_52138_new_n5995_), .Y(u2__abc_52138_new_n6434_));
AOI21X1 AOI21X1_1670 ( .A(u2__abc_52138_new_n13014_), .B(u2__abc_52138_new_n13006_), .C(u2__abc_52138_new_n13016_), .Y(u2__abc_52138_new_n13017_));
AOI21X1 AOI21X1_1671 ( .A(u2__abc_52138_new_n4156_), .B(u2__abc_52138_new_n4946_), .C(u2__abc_52138_new_n4948_), .Y(u2__abc_52138_new_n13020_));
AOI21X1 AOI21X1_1672 ( .A(u2__abc_52138_new_n4952_), .B(u2__abc_52138_new_n4179_), .C(u2__abc_52138_new_n4955_), .Y(u2__abc_52138_new_n13021_));
AOI21X1 AOI21X1_1673 ( .A(u2__abc_52138_new_n13019_), .B(u2__abc_52138_new_n13022_), .C(u2__abc_52138_new_n4968_), .Y(u2__abc_52138_new_n13023_));
AOI21X1 AOI21X1_1674 ( .A(u2__abc_52138_new_n4992_), .B(u2__abc_52138_new_n4982_), .C(u2__abc_52138_new_n13026_), .Y(u2__abc_52138_new_n13027_));
AOI21X1 AOI21X1_1675 ( .A(u2__abc_52138_new_n13018_), .B(u2__abc_52138_new_n9267_), .C(u2__abc_52138_new_n13028_), .Y(u2__abc_52138_new_n13029_));
AOI21X1 AOI21X1_1676 ( .A(u2__abc_52138_new_n12953_), .B(u2__abc_52138_new_n12954_), .C(u2__abc_52138_new_n13030_), .Y(u2__abc_52138_new_n13031_));
AOI21X1 AOI21X1_1677 ( .A(u2__abc_52138_new_n10648_), .B(u2__abc_52138_new_n13034_), .C(u2__abc_52138_new_n13037_), .Y(u2__abc_52138_new_n13038_));
AOI21X1 AOI21X1_1678 ( .A(u2__abc_52138_new_n13039_), .B(u2__abc_52138_new_n13040_), .C(u2__abc_52138_new_n13041_), .Y(u2__abc_52138_new_n13042_));
AOI21X1 AOI21X1_1679 ( .A(u2__abc_52138_new_n13043_), .B(u2__abc_52138_new_n6540_), .C(u2__abc_52138_new_n3069_), .Y(u2__abc_52138_new_n13044_));
AOI21X1 AOI21X1_168 ( .A(u2__abc_52138_new_n6430_), .B(u2__abc_52138_new_n6009_), .C(u2__abc_52138_new_n6435_), .Y(u2__abc_52138_new_n6436_));
AOI21X1 AOI21X1_1680 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3072_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13047_));
AOI21X1 AOI21X1_1681 ( .A(u2__abc_52138_new_n13048_), .B(u2__abc_52138_new_n12818_), .C(rst), .Y(u2__0root_452_0__1_));
AOI21X1 AOI21X1_1682 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3074_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13054_));
AOI21X1 AOI21X1_1683 ( .A(u2__abc_52138_new_n13055_), .B(u2__abc_52138_new_n13050_), .C(rst), .Y(u2__0root_452_0__2_));
AOI21X1 AOI21X1_1684 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3060_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13062_));
AOI21X1 AOI21X1_1685 ( .A(u2__abc_52138_new_n13063_), .B(u2__abc_52138_new_n13057_), .C(rst), .Y(u2__0root_452_0__3_));
AOI21X1 AOI21X1_1686 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3079_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13070_));
AOI21X1 AOI21X1_1687 ( .A(u2__abc_52138_new_n13071_), .B(u2__abc_52138_new_n13065_), .C(rst), .Y(u2__0root_452_0__4_));
AOI21X1 AOI21X1_1688 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6458_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13078_));
AOI21X1 AOI21X1_1689 ( .A(u2__abc_52138_new_n13079_), .B(u2__abc_52138_new_n13073_), .C(rst), .Y(u2__0root_452_0__5_));
AOI21X1 AOI21X1_169 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n6502_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6506_));
AOI21X1 AOI21X1_1690 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3056_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13085_));
AOI21X1 AOI21X1_1691 ( .A(u2__abc_52138_new_n13086_), .B(u2__abc_52138_new_n13081_), .C(rst), .Y(u2__0root_452_0__6_));
AOI21X1 AOI21X1_1692 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3045_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13093_));
AOI21X1 AOI21X1_1693 ( .A(u2__abc_52138_new_n13094_), .B(u2__abc_52138_new_n13088_), .C(rst), .Y(u2__0root_452_0__7_));
AOI21X1 AOI21X1_1694 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3040_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13101_));
AOI21X1 AOI21X1_1695 ( .A(u2__abc_52138_new_n13102_), .B(u2__abc_52138_new_n13096_), .C(rst), .Y(u2__0root_452_0__8_));
AOI21X1 AOI21X1_1696 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3096_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13109_));
AOI21X1 AOI21X1_1697 ( .A(u2__abc_52138_new_n13110_), .B(u2__abc_52138_new_n13104_), .C(rst), .Y(u2__0root_452_0__9_));
AOI21X1 AOI21X1_1698 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3035_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13116_));
AOI21X1 AOI21X1_1699 ( .A(u2__abc_52138_new_n13117_), .B(u2__abc_52138_new_n13112_), .C(rst), .Y(u2__0root_452_0__10_));
AOI21X1 AOI21X1_17 ( .A(u2__abc_52138_new_n3205_), .B(u2__abc_52138_new_n3194_), .C(u2__abc_52138_new_n3216_), .Y(u2__abc_52138_new_n3217_));
AOI21X1 AOI21X1_170 ( .A(u2__abc_52138_new_n6507_), .B(u2__abc_52138_new_n2995_), .C(rst), .Y(u2__0remHi_451_0__0_));
AOI21X1 AOI21X1_1700 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3027_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13124_));
AOI21X1 AOI21X1_1701 ( .A(u2__abc_52138_new_n13125_), .B(u2__abc_52138_new_n13119_), .C(rst), .Y(u2__0root_452_0__11_));
AOI21X1 AOI21X1_1702 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3022_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13132_));
AOI21X1 AOI21X1_1703 ( .A(u2__abc_52138_new_n13133_), .B(u2__abc_52138_new_n13127_), .C(rst), .Y(u2__0root_452_0__12_));
AOI21X1 AOI21X1_1704 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6654_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13140_));
AOI21X1 AOI21X1_1705 ( .A(u2__abc_52138_new_n13141_), .B(u2__abc_52138_new_n13135_), .C(rst), .Y(u2__0root_452_0__13_));
AOI21X1 AOI21X1_1706 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3019_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13147_));
AOI21X1 AOI21X1_1707 ( .A(u2__abc_52138_new_n13148_), .B(u2__abc_52138_new_n13143_), .C(rst), .Y(u2__0root_452_0__14_));
AOI21X1 AOI21X1_1708 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3170_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13155_));
AOI21X1 AOI21X1_1709 ( .A(u2__abc_52138_new_n13156_), .B(u2__abc_52138_new_n13150_), .C(rst), .Y(u2__0root_452_0__15_));
AOI21X1 AOI21X1_171 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n6515_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6516_));
AOI21X1 AOI21X1_1710 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3175_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13163_));
AOI21X1 AOI21X1_1711 ( .A(u2__abc_52138_new_n13164_), .B(u2__abc_52138_new_n13158_), .C(rst), .Y(u2__0root_452_0__16_));
AOI21X1 AOI21X1_1712 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3159_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13171_));
AOI21X1 AOI21X1_1713 ( .A(u2__abc_52138_new_n13172_), .B(u2__abc_52138_new_n13166_), .C(rst), .Y(u2__0root_452_0__17_));
AOI21X1 AOI21X1_1714 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3164_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13178_));
AOI21X1 AOI21X1_1715 ( .A(u2__abc_52138_new_n13179_), .B(u2__abc_52138_new_n13174_), .C(rst), .Y(u2__0root_452_0__18_));
AOI21X1 AOI21X1_1716 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3189_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13186_));
AOI21X1 AOI21X1_1717 ( .A(u2__abc_52138_new_n13187_), .B(u2__abc_52138_new_n13181_), .C(rst), .Y(u2__0root_452_0__19_));
AOI21X1 AOI21X1_1718 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3206_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13194_));
AOI21X1 AOI21X1_1719 ( .A(u2__abc_52138_new_n13195_), .B(u2__abc_52138_new_n13189_), .C(rst), .Y(u2__0root_452_0__20_));
AOI21X1 AOI21X1_172 ( .A(u2__abc_52138_new_n6517_), .B(u2__abc_52138_new_n6509_), .C(rst), .Y(u2__0remHi_451_0__1_));
AOI21X1 AOI21X1_1720 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6733_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13202_));
AOI21X1 AOI21X1_1721 ( .A(u2__abc_52138_new_n13203_), .B(u2__abc_52138_new_n13197_), .C(rst), .Y(u2__0root_452_0__21_));
AOI21X1 AOI21X1_1722 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3183_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13209_));
AOI21X1 AOI21X1_1723 ( .A(u2__abc_52138_new_n13210_), .B(u2__abc_52138_new_n13205_), .C(rst), .Y(u2__0root_452_0__22_));
AOI21X1 AOI21X1_1724 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3128_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13217_));
AOI21X1 AOI21X1_1725 ( .A(u2__abc_52138_new_n13218_), .B(u2__abc_52138_new_n13212_), .C(rst), .Y(u2__0root_452_0__23_));
AOI21X1 AOI21X1_1726 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3123_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13225_));
AOI21X1 AOI21X1_1727 ( .A(u2__abc_52138_new_n13226_), .B(u2__abc_52138_new_n13220_), .C(rst), .Y(u2__0root_452_0__24_));
AOI21X1 AOI21X1_1728 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3112_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13233_));
AOI21X1 AOI21X1_1729 ( .A(u2__abc_52138_new_n13234_), .B(u2__abc_52138_new_n13228_), .C(rst), .Y(u2__0root_452_0__25_));
AOI21X1 AOI21X1_173 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3062_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6525_));
AOI21X1 AOI21X1_1730 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3117_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13240_));
AOI21X1 AOI21X1_1731 ( .A(u2__abc_52138_new_n13241_), .B(u2__abc_52138_new_n13236_), .C(rst), .Y(u2__0root_452_0__26_));
AOI21X1 AOI21X1_1732 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3151_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13248_));
AOI21X1 AOI21X1_1733 ( .A(u2__abc_52138_new_n13249_), .B(u2__abc_52138_new_n13243_), .C(rst), .Y(u2__0root_452_0__27_));
AOI21X1 AOI21X1_1734 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3146_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13256_));
AOI21X1 AOI21X1_1735 ( .A(u2__abc_52138_new_n13257_), .B(u2__abc_52138_new_n13251_), .C(rst), .Y(u2__0root_452_0__28_));
AOI21X1 AOI21X1_1736 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3135_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13264_));
AOI21X1 AOI21X1_1737 ( .A(u2__abc_52138_new_n13265_), .B(u2__abc_52138_new_n13259_), .C(rst), .Y(u2__0root_452_0__29_));
AOI21X1 AOI21X1_1738 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3142_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13271_));
AOI21X1 AOI21X1_1739 ( .A(u2__abc_52138_new_n13272_), .B(u2__abc_52138_new_n13267_), .C(rst), .Y(u2__0root_452_0__30_));
AOI21X1 AOI21X1_174 ( .A(u2__abc_52138_new_n6526_), .B(u2__abc_52138_new_n6519_), .C(rst), .Y(u2__0remHi_451_0__2_));
AOI21X1 AOI21X1_1740 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3389_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13279_));
AOI21X1 AOI21X1_1741 ( .A(u2__abc_52138_new_n13280_), .B(u2__abc_52138_new_n13274_), .C(rst), .Y(u2__0root_452_0__31_));
AOI21X1 AOI21X1_1742 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3394_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13287_));
AOI21X1 AOI21X1_1743 ( .A(u2__abc_52138_new_n13288_), .B(u2__abc_52138_new_n13282_), .C(rst), .Y(u2__0root_452_0__32_));
AOI21X1 AOI21X1_1744 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3437_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13295_));
AOI21X1 AOI21X1_1745 ( .A(u2__abc_52138_new_n13296_), .B(u2__abc_52138_new_n13290_), .C(rst), .Y(u2__0root_452_0__33_));
AOI21X1 AOI21X1_1746 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3383_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13302_));
AOI21X1 AOI21X1_1747 ( .A(u2__abc_52138_new_n13303_), .B(u2__abc_52138_new_n13298_), .C(rst), .Y(u2__0root_452_0__34_));
AOI21X1 AOI21X1_1748 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n13310_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13311_));
AOI21X1 AOI21X1_1749 ( .A(u2__abc_52138_new_n13312_), .B(u2__abc_52138_new_n13305_), .C(rst), .Y(u2__0root_452_0__35_));
AOI21X1 AOI21X1_175 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3081_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6534_));
AOI21X1 AOI21X1_1750 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3412_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13319_));
AOI21X1 AOI21X1_1751 ( .A(u2__abc_52138_new_n13320_), .B(u2__abc_52138_new_n13314_), .C(rst), .Y(u2__0root_452_0__36_));
AOI21X1 AOI21X1_1752 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3401_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13327_));
AOI21X1 AOI21X1_1753 ( .A(u2__abc_52138_new_n13328_), .B(u2__abc_52138_new_n13322_), .C(rst), .Y(u2__0root_452_0__37_));
AOI21X1 AOI21X1_1754 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3406_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13334_));
AOI21X1 AOI21X1_1755 ( .A(u2__abc_52138_new_n13335_), .B(u2__abc_52138_new_n13330_), .C(rst), .Y(u2__0root_452_0__38_));
AOI21X1 AOI21X1_1756 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3346_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13342_));
AOI21X1 AOI21X1_1757 ( .A(u2__abc_52138_new_n13343_), .B(u2__abc_52138_new_n13337_), .C(rst), .Y(u2__0root_452_0__39_));
AOI21X1 AOI21X1_1758 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3351_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13350_));
AOI21X1 AOI21X1_1759 ( .A(u2__abc_52138_new_n13351_), .B(u2__abc_52138_new_n13345_), .C(rst), .Y(u2__0root_452_0__40_));
AOI21X1 AOI21X1_176 ( .A(u2__abc_52138_new_n6535_), .B(u2__abc_52138_new_n6528_), .C(rst), .Y(u2__0remHi_451_0__3_));
AOI21X1 AOI21X1_1760 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3335_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13358_));
AOI21X1 AOI21X1_1761 ( .A(u2__abc_52138_new_n13359_), .B(u2__abc_52138_new_n13353_), .C(rst), .Y(u2__0root_452_0__41_));
AOI21X1 AOI21X1_1762 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3340_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13365_));
AOI21X1 AOI21X1_1763 ( .A(u2__abc_52138_new_n13366_), .B(u2__abc_52138_new_n13361_), .C(rst), .Y(u2__0root_452_0__42_));
AOI21X1 AOI21X1_1764 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3374_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13373_));
AOI21X1 AOI21X1_1765 ( .A(u2__abc_52138_new_n13374_), .B(u2__abc_52138_new_n13368_), .C(rst), .Y(u2__0root_452_0__43_));
AOI21X1 AOI21X1_1766 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3369_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13381_));
AOI21X1 AOI21X1_1767 ( .A(u2__abc_52138_new_n13382_), .B(u2__abc_52138_new_n13376_), .C(rst), .Y(u2__0root_452_0__44_));
AOI21X1 AOI21X1_1768 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3358_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13389_));
AOI21X1 AOI21X1_1769 ( .A(u2__abc_52138_new_n13390_), .B(u2__abc_52138_new_n13384_), .C(rst), .Y(u2__0root_452_0__45_));
AOI21X1 AOI21X1_177 ( .A(u2__abc_52138_new_n6441_), .B(u2__abc_52138_new_n3015_), .C(u2__abc_52138_new_n6538_), .Y(u2__abc_52138_new_n6539_));
AOI21X1 AOI21X1_1770 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3363_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13396_));
AOI21X1 AOI21X1_1771 ( .A(u2__abc_52138_new_n13397_), .B(u2__abc_52138_new_n13392_), .C(rst), .Y(u2__0root_452_0__46_));
AOI21X1 AOI21X1_1772 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3303_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13404_));
AOI21X1 AOI21X1_1773 ( .A(u2__abc_52138_new_n13405_), .B(u2__abc_52138_new_n13399_), .C(rst), .Y(u2__0root_452_0__47_));
AOI21X1 AOI21X1_1774 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3300_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13412_));
AOI21X1 AOI21X1_1775 ( .A(u2__abc_52138_new_n13413_), .B(u2__abc_52138_new_n13407_), .C(rst), .Y(u2__0root_452_0__48_));
AOI21X1 AOI21X1_1776 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3289_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13420_));
AOI21X1 AOI21X1_1777 ( .A(u2__abc_52138_new_n13421_), .B(u2__abc_52138_new_n13415_), .C(rst), .Y(u2__0root_452_0__49_));
AOI21X1 AOI21X1_1778 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3294_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13427_));
AOI21X1 AOI21X1_1779 ( .A(u2__abc_52138_new_n13428_), .B(u2__abc_52138_new_n13423_), .C(rst), .Y(u2__0root_452_0__50_));
AOI21X1 AOI21X1_178 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3086_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6546_));
AOI21X1 AOI21X1_1780 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3327_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13435_));
AOI21X1 AOI21X1_1781 ( .A(u2__abc_52138_new_n13436_), .B(u2__abc_52138_new_n13430_), .C(rst), .Y(u2__0root_452_0__51_));
AOI21X1 AOI21X1_1782 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3322_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13443_));
AOI21X1 AOI21X1_1783 ( .A(u2__abc_52138_new_n13444_), .B(u2__abc_52138_new_n13438_), .C(rst), .Y(u2__0root_452_0__52_));
AOI21X1 AOI21X1_1784 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3311_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13451_));
AOI21X1 AOI21X1_1785 ( .A(u2__abc_52138_new_n13452_), .B(u2__abc_52138_new_n13446_), .C(rst), .Y(u2__0root_452_0__53_));
AOI21X1 AOI21X1_1786 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3316_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13458_));
AOI21X1 AOI21X1_1787 ( .A(u2__abc_52138_new_n13459_), .B(u2__abc_52138_new_n13454_), .C(rst), .Y(u2__0root_452_0__54_));
AOI21X1 AOI21X1_1788 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3251_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13466_));
AOI21X1 AOI21X1_1789 ( .A(u2__abc_52138_new_n13467_), .B(u2__abc_52138_new_n13461_), .C(rst), .Y(u2__0root_452_0__55_));
AOI21X1 AOI21X1_179 ( .A(u2__abc_52138_new_n6547_), .B(u2__abc_52138_new_n6537_), .C(rst), .Y(u2__0remHi_451_0__4_));
AOI21X1 AOI21X1_1790 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3256_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13474_));
AOI21X1 AOI21X1_1791 ( .A(u2__abc_52138_new_n13475_), .B(u2__abc_52138_new_n13469_), .C(rst), .Y(u2__0root_452_0__56_));
AOI21X1 AOI21X1_1792 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3240_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13482_));
AOI21X1 AOI21X1_1793 ( .A(u2__abc_52138_new_n13483_), .B(u2__abc_52138_new_n13477_), .C(rst), .Y(u2__0root_452_0__57_));
AOI21X1 AOI21X1_1794 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3245_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13489_));
AOI21X1 AOI21X1_1795 ( .A(u2__abc_52138_new_n13490_), .B(u2__abc_52138_new_n13485_), .C(rst), .Y(u2__0root_452_0__58_));
AOI21X1 AOI21X1_1796 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3279_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13497_));
AOI21X1 AOI21X1_1797 ( .A(u2__abc_52138_new_n13498_), .B(u2__abc_52138_new_n13492_), .C(rst), .Y(u2__0root_452_0__59_));
AOI21X1 AOI21X1_1798 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3274_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13505_));
AOI21X1 AOI21X1_1799 ( .A(u2__abc_52138_new_n13506_), .B(u2__abc_52138_new_n13500_), .C(rst), .Y(u2__0root_452_0__60_));
AOI21X1 AOI21X1_18 ( .A(u2__abc_52138_new_n3223_), .B(u2__abc_52138_new_n3124_), .C(u2__abc_52138_new_n3222_), .Y(u2__abc_52138_new_n3224_));
AOI21X1 AOI21X1_180 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3054_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6555_));
AOI21X1 AOI21X1_1800 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3263_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13513_));
AOI21X1 AOI21X1_1801 ( .A(u2__abc_52138_new_n13514_), .B(u2__abc_52138_new_n13508_), .C(rst), .Y(u2__0root_452_0__61_));
AOI21X1 AOI21X1_1802 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3270_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13520_));
AOI21X1 AOI21X1_1803 ( .A(u2__abc_52138_new_n13521_), .B(u2__abc_52138_new_n13516_), .C(rst), .Y(u2__0root_452_0__62_));
AOI21X1 AOI21X1_1804 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3832_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13528_));
AOI21X1 AOI21X1_1805 ( .A(u2__abc_52138_new_n13529_), .B(u2__abc_52138_new_n13523_), .C(rst), .Y(u2__0root_452_0__63_));
AOI21X1 AOI21X1_1806 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3837_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13536_));
AOI21X1 AOI21X1_1807 ( .A(u2__abc_52138_new_n13537_), .B(u2__abc_52138_new_n13531_), .C(rst), .Y(u2__0root_452_0__64_));
AOI21X1 AOI21X1_1808 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3843_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13544_));
AOI21X1 AOI21X1_1809 ( .A(u2__abc_52138_new_n13545_), .B(u2__abc_52138_new_n13539_), .C(rst), .Y(u2__0root_452_0__65_));
AOI21X1 AOI21X1_181 ( .A(u2__abc_52138_new_n6556_), .B(u2__abc_52138_new_n6549_), .C(rst), .Y(u2__0remHi_451_0__5_));
AOI21X1 AOI21X1_1810 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3848_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13551_));
AOI21X1 AOI21X1_1811 ( .A(u2__abc_52138_new_n13552_), .B(u2__abc_52138_new_n13547_), .C(rst), .Y(u2__0root_452_0__66_));
AOI21X1 AOI21X1_1812 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3862_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13559_));
AOI21X1 AOI21X1_1813 ( .A(u2__abc_52138_new_n13560_), .B(u2__abc_52138_new_n13554_), .C(rst), .Y(u2__0root_452_0__67_));
AOI21X1 AOI21X1_1814 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3881_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13567_));
AOI21X1 AOI21X1_1815 ( .A(u2__abc_52138_new_n13568_), .B(u2__abc_52138_new_n13562_), .C(rst), .Y(u2__0root_452_0__68_));
AOI21X1 AOI21X1_1816 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7264_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13575_));
AOI21X1 AOI21X1_1817 ( .A(u2__abc_52138_new_n13576_), .B(u2__abc_52138_new_n13570_), .C(rst), .Y(u2__0root_452_0__69_));
AOI21X1 AOI21X1_1818 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3856_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13582_));
AOI21X1 AOI21X1_1819 ( .A(u2__abc_52138_new_n13583_), .B(u2__abc_52138_new_n13578_), .C(rst), .Y(u2__0root_452_0__70_));
AOI21X1 AOI21X1_182 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3047_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6564_));
AOI21X1 AOI21X1_1820 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3788_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13590_));
AOI21X1 AOI21X1_1821 ( .A(u2__abc_52138_new_n13591_), .B(u2__abc_52138_new_n13585_), .C(rst), .Y(u2__0root_452_0__71_));
AOI21X1 AOI21X1_1822 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3793_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13598_));
AOI21X1 AOI21X1_1823 ( .A(u2__abc_52138_new_n13599_), .B(u2__abc_52138_new_n13593_), .C(rst), .Y(u2__0root_452_0__72_));
AOI21X1 AOI21X1_1824 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3797_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13606_));
AOI21X1 AOI21X1_1825 ( .A(u2__abc_52138_new_n13607_), .B(u2__abc_52138_new_n13601_), .C(rst), .Y(u2__0root_452_0__73_));
AOI21X1 AOI21X1_1826 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3802_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13613_));
AOI21X1 AOI21X1_1827 ( .A(u2__abc_52138_new_n13614_), .B(u2__abc_52138_new_n13609_), .C(rst), .Y(u2__0root_452_0__74_));
AOI21X1 AOI21X1_1828 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3826_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13621_));
AOI21X1 AOI21X1_1829 ( .A(u2__abc_52138_new_n13622_), .B(u2__abc_52138_new_n13616_), .C(rst), .Y(u2__0root_452_0__75_));
AOI21X1 AOI21X1_183 ( .A(u2__abc_52138_new_n6565_), .B(u2__abc_52138_new_n6558_), .C(rst), .Y(u2__0remHi_451_0__6_));
AOI21X1 AOI21X1_1830 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3821_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13629_));
AOI21X1 AOI21X1_1831 ( .A(u2__abc_52138_new_n13630_), .B(u2__abc_52138_new_n13624_), .C(rst), .Y(u2__0root_452_0__76_));
AOI21X1 AOI21X1_1832 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3810_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13637_));
AOI21X1 AOI21X1_1833 ( .A(u2__abc_52138_new_n13638_), .B(u2__abc_52138_new_n13632_), .C(rst), .Y(u2__0root_452_0__77_));
AOI21X1 AOI21X1_1834 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3815_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13644_));
AOI21X1 AOI21X1_1835 ( .A(u2__abc_52138_new_n13645_), .B(u2__abc_52138_new_n13640_), .C(rst), .Y(u2__0root_452_0__78_));
AOI21X1 AOI21X1_1836 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3738_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13652_));
AOI21X1 AOI21X1_1837 ( .A(u2__abc_52138_new_n13653_), .B(u2__abc_52138_new_n13647_), .C(rst), .Y(u2__0root_452_0__79_));
AOI21X1 AOI21X1_1838 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3743_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13660_));
AOI21X1 AOI21X1_1839 ( .A(u2__abc_52138_new_n13661_), .B(u2__abc_52138_new_n13655_), .C(rst), .Y(u2__0root_452_0__80_));
AOI21X1 AOI21X1_184 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3042_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6572_));
AOI21X1 AOI21X1_1840 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3749_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13668_));
AOI21X1 AOI21X1_1841 ( .A(u2__abc_52138_new_n13669_), .B(u2__abc_52138_new_n13663_), .C(rst), .Y(u2__0root_452_0__81_));
AOI21X1 AOI21X1_1842 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3754_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13675_));
AOI21X1 AOI21X1_1843 ( .A(u2__abc_52138_new_n13676_), .B(u2__abc_52138_new_n13671_), .C(rst), .Y(u2__0root_452_0__82_));
AOI21X1 AOI21X1_1844 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3777_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13683_));
AOI21X1 AOI21X1_1845 ( .A(u2__abc_52138_new_n13684_), .B(u2__abc_52138_new_n13678_), .C(rst), .Y(u2__0root_452_0__83_));
AOI21X1 AOI21X1_1846 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3772_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13691_));
AOI21X1 AOI21X1_1847 ( .A(u2__abc_52138_new_n13692_), .B(u2__abc_52138_new_n13686_), .C(rst), .Y(u2__0root_452_0__84_));
AOI21X1 AOI21X1_1848 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3761_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13699_));
AOI21X1 AOI21X1_1849 ( .A(u2__abc_52138_new_n13700_), .B(u2__abc_52138_new_n13694_), .C(rst), .Y(u2__0root_452_0__85_));
AOI21X1 AOI21X1_185 ( .A(u2__abc_52138_new_n6573_), .B(u2__abc_52138_new_n6567_), .C(rst), .Y(u2__0remHi_451_0__7_));
AOI21X1 AOI21X1_1850 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3766_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13706_));
AOI21X1 AOI21X1_1851 ( .A(u2__abc_52138_new_n13707_), .B(u2__abc_52138_new_n13702_), .C(rst), .Y(u2__0root_452_0__86_));
AOI21X1 AOI21X1_1852 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3732_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13714_));
AOI21X1 AOI21X1_1853 ( .A(u2__abc_52138_new_n13715_), .B(u2__abc_52138_new_n13709_), .C(rst), .Y(u2__0root_452_0__87_));
AOI21X1 AOI21X1_1854 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3727_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13722_));
AOI21X1 AOI21X1_1855 ( .A(u2__abc_52138_new_n13723_), .B(u2__abc_52138_new_n13717_), .C(rst), .Y(u2__0root_452_0__88_));
AOI21X1 AOI21X1_1856 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3713_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13730_));
AOI21X1 AOI21X1_1857 ( .A(u2__abc_52138_new_n13731_), .B(u2__abc_52138_new_n13725_), .C(rst), .Y(u2__0root_452_0__89_));
AOI21X1 AOI21X1_1858 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3718_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13737_));
AOI21X1 AOI21X1_1859 ( .A(u2__abc_52138_new_n13738_), .B(u2__abc_52138_new_n13733_), .C(rst), .Y(u2__0root_452_0__90_));
AOI21X1 AOI21X1_186 ( .A(u2__abc_52138_new_n6578_), .B(u2__abc_52138_new_n3055_), .C(u2__abc_52138_new_n6579_), .Y(u2__abc_52138_new_n6580_));
AOI21X1 AOI21X1_1860 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3708_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13745_));
AOI21X1 AOI21X1_1861 ( .A(u2__abc_52138_new_n13746_), .B(u2__abc_52138_new_n13740_), .C(rst), .Y(u2__0root_452_0__91_));
AOI21X1 AOI21X1_1862 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3702_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13753_));
AOI21X1 AOI21X1_1863 ( .A(u2__abc_52138_new_n13754_), .B(u2__abc_52138_new_n13748_), .C(rst), .Y(u2__0root_452_0__92_));
AOI21X1 AOI21X1_1864 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3691_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13761_));
AOI21X1 AOI21X1_1865 ( .A(u2__abc_52138_new_n13762_), .B(u2__abc_52138_new_n13756_), .C(rst), .Y(u2__0root_452_0__93_));
AOI21X1 AOI21X1_1866 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3696_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13768_));
AOI21X1 AOI21X1_1867 ( .A(u2__abc_52138_new_n13769_), .B(u2__abc_52138_new_n13764_), .C(rst), .Y(u2__0root_452_0__94_));
AOI21X1 AOI21X1_1868 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3658_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13776_));
AOI21X1 AOI21X1_1869 ( .A(u2__abc_52138_new_n13777_), .B(u2__abc_52138_new_n13771_), .C(rst), .Y(u2__0root_452_0__95_));
AOI21X1 AOI21X1_187 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n6586_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6587_));
AOI21X1 AOI21X1_1870 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3653_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13784_));
AOI21X1 AOI21X1_1871 ( .A(u2__abc_52138_new_n13785_), .B(u2__abc_52138_new_n13779_), .C(rst), .Y(u2__0root_452_0__96_));
AOI21X1 AOI21X1_1872 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3644_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13792_));
AOI21X1 AOI21X1_1873 ( .A(u2__abc_52138_new_n13793_), .B(u2__abc_52138_new_n13787_), .C(rst), .Y(u2__0root_452_0__97_));
AOI21X1 AOI21X1_1874 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3649_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13799_));
AOI21X1 AOI21X1_1875 ( .A(u2__abc_52138_new_n13800_), .B(u2__abc_52138_new_n13795_), .C(rst), .Y(u2__0root_452_0__98_));
AOI21X1 AOI21X1_1876 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3681_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13807_));
AOI21X1 AOI21X1_1877 ( .A(u2__abc_52138_new_n13808_), .B(u2__abc_52138_new_n13802_), .C(rst), .Y(u2__0root_452_0__99_));
AOI21X1 AOI21X1_1878 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3676_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13815_));
AOI21X1 AOI21X1_1879 ( .A(u2__abc_52138_new_n13816_), .B(u2__abc_52138_new_n13810_), .C(rst), .Y(u2__0root_452_0__100_));
AOI21X1 AOI21X1_188 ( .A(u2__abc_52138_new_n6588_), .B(u2__abc_52138_new_n6575_), .C(rst), .Y(u2__0remHi_451_0__8_));
AOI21X1 AOI21X1_1880 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3665_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13823_));
AOI21X1 AOI21X1_1881 ( .A(u2__abc_52138_new_n13824_), .B(u2__abc_52138_new_n13818_), .C(rst), .Y(u2__0root_452_0__101_));
AOI21X1 AOI21X1_1882 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3670_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13830_));
AOI21X1 AOI21X1_1883 ( .A(u2__abc_52138_new_n13831_), .B(u2__abc_52138_new_n13826_), .C(rst), .Y(u2__0root_452_0__102_));
AOI21X1 AOI21X1_1884 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3614_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13838_));
AOI21X1 AOI21X1_1885 ( .A(u2__abc_52138_new_n13839_), .B(u2__abc_52138_new_n13833_), .C(rst), .Y(u2__0root_452_0__103_));
AOI21X1 AOI21X1_1886 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3608_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13846_));
AOI21X1 AOI21X1_1887 ( .A(u2__abc_52138_new_n13847_), .B(u2__abc_52138_new_n13841_), .C(rst), .Y(u2__0root_452_0__104_));
AOI21X1 AOI21X1_1888 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3597_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13854_));
AOI21X1 AOI21X1_1889 ( .A(u2__abc_52138_new_n13855_), .B(u2__abc_52138_new_n13849_), .C(rst), .Y(u2__0root_452_0__105_));
AOI21X1 AOI21X1_189 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3037_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6595_));
AOI21X1 AOI21X1_1890 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3602_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13861_));
AOI21X1 AOI21X1_1891 ( .A(u2__abc_52138_new_n13862_), .B(u2__abc_52138_new_n13857_), .C(rst), .Y(u2__0root_452_0__106_));
AOI21X1 AOI21X1_1892 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3636_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13869_));
AOI21X1 AOI21X1_1893 ( .A(u2__abc_52138_new_n13870_), .B(u2__abc_52138_new_n13864_), .C(rst), .Y(u2__0root_452_0__107_));
AOI21X1 AOI21X1_1894 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3630_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13877_));
AOI21X1 AOI21X1_1895 ( .A(u2__abc_52138_new_n13878_), .B(u2__abc_52138_new_n13872_), .C(rst), .Y(u2__0root_452_0__108_));
AOI21X1 AOI21X1_1896 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3619_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13885_));
AOI21X1 AOI21X1_1897 ( .A(u2__abc_52138_new_n13886_), .B(u2__abc_52138_new_n13880_), .C(rst), .Y(u2__0root_452_0__109_));
AOI21X1 AOI21X1_1898 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3624_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13892_));
AOI21X1 AOI21X1_1899 ( .A(u2__abc_52138_new_n13893_), .B(u2__abc_52138_new_n13888_), .C(rst), .Y(u2__0root_452_0__110_));
AOI21X1 AOI21X1_19 ( .A(u2__abc_52138_new_n3230_), .B(u2__abc_52138_new_n3143_), .C(u2__abc_52138_new_n3231_), .Y(u2__abc_52138_new_n3232_));
AOI21X1 AOI21X1_190 ( .A(u2__abc_52138_new_n6596_), .B(u2__abc_52138_new_n6590_), .C(rst), .Y(u2__0remHi_451_0__9_));
AOI21X1 AOI21X1_1900 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3550_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13900_));
AOI21X1 AOI21X1_1901 ( .A(u2__abc_52138_new_n13901_), .B(u2__abc_52138_new_n13895_), .C(rst), .Y(u2__0root_452_0__111_));
AOI21X1 AOI21X1_1902 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3555_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13908_));
AOI21X1 AOI21X1_1903 ( .A(u2__abc_52138_new_n13909_), .B(u2__abc_52138_new_n13903_), .C(rst), .Y(u2__0root_452_0__112_));
AOI21X1 AOI21X1_1904 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3561_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13916_));
AOI21X1 AOI21X1_1905 ( .A(u2__abc_52138_new_n13917_), .B(u2__abc_52138_new_n13911_), .C(rst), .Y(u2__0root_452_0__113_));
AOI21X1 AOI21X1_1906 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3566_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13923_));
AOI21X1 AOI21X1_1907 ( .A(u2__abc_52138_new_n13924_), .B(u2__abc_52138_new_n13919_), .C(rst), .Y(u2__0root_452_0__114_));
AOI21X1 AOI21X1_1908 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3588_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13931_));
AOI21X1 AOI21X1_1909 ( .A(u2__abc_52138_new_n13932_), .B(u2__abc_52138_new_n13926_), .C(rst), .Y(u2__0root_452_0__115_));
AOI21X1 AOI21X1_191 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3029_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6610_));
AOI21X1 AOI21X1_1910 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3583_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13939_));
AOI21X1 AOI21X1_1911 ( .A(u2__abc_52138_new_n13940_), .B(u2__abc_52138_new_n13934_), .C(rst), .Y(u2__0root_452_0__116_));
AOI21X1 AOI21X1_1912 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3575_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13947_));
AOI21X1 AOI21X1_1913 ( .A(u2__abc_52138_new_n13948_), .B(u2__abc_52138_new_n13942_), .C(rst), .Y(u2__0root_452_0__117_));
AOI21X1 AOI21X1_1914 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3578_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13954_));
AOI21X1 AOI21X1_1915 ( .A(u2__abc_52138_new_n13955_), .B(u2__abc_52138_new_n13950_), .C(rst), .Y(u2__0root_452_0__118_));
AOI21X1 AOI21X1_1916 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n13962_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13963_));
AOI21X1 AOI21X1_1917 ( .A(u2__abc_52138_new_n13964_), .B(u2__abc_52138_new_n13957_), .C(rst), .Y(u2__0root_452_0__119_));
AOI21X1 AOI21X1_1918 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3511_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13971_));
AOI21X1 AOI21X1_1919 ( .A(u2__abc_52138_new_n13972_), .B(u2__abc_52138_new_n13966_), .C(rst), .Y(u2__0root_452_0__120_));
AOI21X1 AOI21X1_192 ( .A(u2__abc_52138_new_n6611_), .B(u2__abc_52138_new_n6598_), .C(rst), .Y(u2__0remHi_451_0__10_));
AOI21X1 AOI21X1_1920 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3516_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13979_));
AOI21X1 AOI21X1_1921 ( .A(u2__abc_52138_new_n13980_), .B(u2__abc_52138_new_n13974_), .C(rst), .Y(u2__0root_452_0__121_));
AOI21X1 AOI21X1_1922 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3521_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13986_));
AOI21X1 AOI21X1_1923 ( .A(u2__abc_52138_new_n13987_), .B(u2__abc_52138_new_n13982_), .C(rst), .Y(u2__0root_452_0__122_));
AOI21X1 AOI21X1_1924 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3544_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n13994_));
AOI21X1 AOI21X1_1925 ( .A(u2__abc_52138_new_n13995_), .B(u2__abc_52138_new_n13989_), .C(rst), .Y(u2__0root_452_0__123_));
AOI21X1 AOI21X1_1926 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3538_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14002_));
AOI21X1 AOI21X1_1927 ( .A(u2__abc_52138_new_n14003_), .B(u2__abc_52138_new_n13997_), .C(rst), .Y(u2__0root_452_0__124_));
AOI21X1 AOI21X1_1928 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3527_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14010_));
AOI21X1 AOI21X1_1929 ( .A(u2__abc_52138_new_n14011_), .B(u2__abc_52138_new_n14005_), .C(rst), .Y(u2__0root_452_0__125_));
AOI21X1 AOI21X1_193 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3024_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6620_));
AOI21X1 AOI21X1_1930 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3534_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14017_));
AOI21X1 AOI21X1_1931 ( .A(u2__abc_52138_new_n14018_), .B(u2__abc_52138_new_n14013_), .C(rst), .Y(u2__0root_452_0__126_));
AOI21X1 AOI21X1_1932 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4713_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14025_));
AOI21X1 AOI21X1_1933 ( .A(u2__abc_52138_new_n14026_), .B(u2__abc_52138_new_n14020_), .C(rst), .Y(u2__0root_452_0__127_));
AOI21X1 AOI21X1_1934 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4719_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14033_));
AOI21X1 AOI21X1_1935 ( .A(u2__abc_52138_new_n14034_), .B(u2__abc_52138_new_n14028_), .C(rst), .Y(u2__0root_452_0__128_));
AOI21X1 AOI21X1_1936 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4770_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14041_));
AOI21X1 AOI21X1_1937 ( .A(u2__abc_52138_new_n14042_), .B(u2__abc_52138_new_n14036_), .C(rst), .Y(u2__0root_452_0__129_));
AOI21X1 AOI21X1_1938 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4727_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14048_));
AOI21X1 AOI21X1_1939 ( .A(u2__abc_52138_new_n14049_), .B(u2__abc_52138_new_n14044_), .C(rst), .Y(u2__0root_452_0__130_));
AOI21X1 AOI21X1_194 ( .A(u2__abc_52138_new_n6621_), .B(u2__abc_52138_new_n6613_), .C(rst), .Y(u2__0remHi_451_0__11_));
AOI21X1 AOI21X1_1940 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n14056_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14057_));
AOI21X1 AOI21X1_1941 ( .A(u2__abc_52138_new_n14058_), .B(u2__abc_52138_new_n14051_), .C(rst), .Y(u2__0root_452_0__131_));
AOI21X1 AOI21X1_1942 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4744_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14065_));
AOI21X1 AOI21X1_1943 ( .A(u2__abc_52138_new_n14066_), .B(u2__abc_52138_new_n14060_), .C(rst), .Y(u2__0root_452_0__132_));
AOI21X1 AOI21X1_1944 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4733_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14073_));
AOI21X1 AOI21X1_1945 ( .A(u2__abc_52138_new_n14074_), .B(u2__abc_52138_new_n14068_), .C(rst), .Y(u2__0root_452_0__133_));
AOI21X1 AOI21X1_1946 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4738_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14080_));
AOI21X1 AOI21X1_1947 ( .A(u2__abc_52138_new_n14081_), .B(u2__abc_52138_new_n14076_), .C(rst), .Y(u2__0root_452_0__134_));
AOI21X1 AOI21X1_1948 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4677_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14088_));
AOI21X1 AOI21X1_1949 ( .A(u2__abc_52138_new_n14089_), .B(u2__abc_52138_new_n14083_), .C(rst), .Y(u2__0root_452_0__135_));
AOI21X1 AOI21X1_195 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3101_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6631_));
AOI21X1 AOI21X1_1950 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4682_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14096_));
AOI21X1 AOI21X1_1951 ( .A(u2__abc_52138_new_n14097_), .B(u2__abc_52138_new_n14091_), .C(rst), .Y(u2__0root_452_0__136_));
AOI21X1 AOI21X1_1952 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4666_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14104_));
AOI21X1 AOI21X1_1953 ( .A(u2__abc_52138_new_n14105_), .B(u2__abc_52138_new_n14099_), .C(rst), .Y(u2__0root_452_0__137_));
AOI21X1 AOI21X1_1954 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4671_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14111_));
AOI21X1 AOI21X1_1955 ( .A(u2__abc_52138_new_n14112_), .B(u2__abc_52138_new_n14107_), .C(rst), .Y(u2__0root_452_0__138_));
AOI21X1 AOI21X1_1956 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4705_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14119_));
AOI21X1 AOI21X1_1957 ( .A(u2__abc_52138_new_n14120_), .B(u2__abc_52138_new_n14114_), .C(rst), .Y(u2__0root_452_0__139_));
AOI21X1 AOI21X1_1958 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4700_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14127_));
AOI21X1 AOI21X1_1959 ( .A(u2__abc_52138_new_n14128_), .B(u2__abc_52138_new_n14122_), .C(rst), .Y(u2__0root_452_0__140_));
AOI21X1 AOI21X1_196 ( .A(u2__abc_52138_new_n6632_), .B(u2__abc_52138_new_n6623_), .C(rst), .Y(u2__0remHi_451_0__12_));
AOI21X1 AOI21X1_1960 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4689_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14135_));
AOI21X1 AOI21X1_1961 ( .A(u2__abc_52138_new_n14136_), .B(u2__abc_52138_new_n14130_), .C(rst), .Y(u2__0root_452_0__141_));
AOI21X1 AOI21X1_1962 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4694_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14142_));
AOI21X1 AOI21X1_1963 ( .A(u2__abc_52138_new_n14143_), .B(u2__abc_52138_new_n14138_), .C(rst), .Y(u2__0root_452_0__142_));
AOI21X1 AOI21X1_1964 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4660_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14150_));
AOI21X1 AOI21X1_1965 ( .A(u2__abc_52138_new_n14151_), .B(u2__abc_52138_new_n14145_), .C(rst), .Y(u2__0root_452_0__143_));
AOI21X1 AOI21X1_1966 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4655_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14158_));
AOI21X1 AOI21X1_1967 ( .A(u2__abc_52138_new_n14159_), .B(u2__abc_52138_new_n14153_), .C(rst), .Y(u2__0root_452_0__144_));
AOI21X1 AOI21X1_1968 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4642_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14166_));
AOI21X1 AOI21X1_1969 ( .A(u2__abc_52138_new_n14167_), .B(u2__abc_52138_new_n14161_), .C(rst), .Y(u2__0root_452_0__145_));
AOI21X1 AOI21X1_197 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3017_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6639_));
AOI21X1 AOI21X1_1970 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4647_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14173_));
AOI21X1 AOI21X1_1971 ( .A(u2__abc_52138_new_n14174_), .B(u2__abc_52138_new_n14169_), .C(rst), .Y(u2__0root_452_0__146_));
AOI21X1 AOI21X1_1972 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4635_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14181_));
AOI21X1 AOI21X1_1973 ( .A(u2__abc_52138_new_n14182_), .B(u2__abc_52138_new_n14176_), .C(rst), .Y(u2__0root_452_0__147_));
AOI21X1 AOI21X1_1974 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4630_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14189_));
AOI21X1 AOI21X1_1975 ( .A(u2__abc_52138_new_n14190_), .B(u2__abc_52138_new_n14184_), .C(rst), .Y(u2__0root_452_0__148_));
AOI21X1 AOI21X1_1976 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4619_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14197_));
AOI21X1 AOI21X1_1977 ( .A(u2__abc_52138_new_n14198_), .B(u2__abc_52138_new_n14192_), .C(rst), .Y(u2__0root_452_0__149_));
AOI21X1 AOI21X1_1978 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4624_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14204_));
AOI21X1 AOI21X1_1979 ( .A(u2__abc_52138_new_n14205_), .B(u2__abc_52138_new_n14200_), .C(rst), .Y(u2__0root_452_0__150_));
AOI21X1 AOI21X1_198 ( .A(u2__abc_52138_new_n6640_), .B(u2__abc_52138_new_n6634_), .C(rst), .Y(u2__0remHi_451_0__13_));
AOI21X1 AOI21X1_1980 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4589_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14212_));
AOI21X1 AOI21X1_1981 ( .A(u2__abc_52138_new_n14213_), .B(u2__abc_52138_new_n14207_), .C(rst), .Y(u2__0root_452_0__151_));
AOI21X1 AOI21X1_1982 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4584_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14220_));
AOI21X1 AOI21X1_1983 ( .A(u2__abc_52138_new_n14221_), .B(u2__abc_52138_new_n14215_), .C(rst), .Y(u2__0root_452_0__152_));
AOI21X1 AOI21X1_1984 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4573_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14228_));
AOI21X1 AOI21X1_1985 ( .A(u2__abc_52138_new_n14229_), .B(u2__abc_52138_new_n14223_), .C(rst), .Y(u2__0root_452_0__153_));
AOI21X1 AOI21X1_1986 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4578_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14235_));
AOI21X1 AOI21X1_1987 ( .A(u2__abc_52138_new_n14236_), .B(u2__abc_52138_new_n14231_), .C(rst), .Y(u2__0root_452_0__154_));
AOI21X1 AOI21X1_1988 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4614_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14243_));
AOI21X1 AOI21X1_1989 ( .A(u2__abc_52138_new_n14244_), .B(u2__abc_52138_new_n14238_), .C(rst), .Y(u2__0root_452_0__155_));
AOI21X1 AOI21X1_199 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3172_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6649_));
AOI21X1 AOI21X1_1990 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4609_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14251_));
AOI21X1 AOI21X1_1991 ( .A(u2__abc_52138_new_n14252_), .B(u2__abc_52138_new_n14246_), .C(rst), .Y(u2__0root_452_0__156_));
AOI21X1 AOI21X1_1992 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4596_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14259_));
AOI21X1 AOI21X1_1993 ( .A(u2__abc_52138_new_n14260_), .B(u2__abc_52138_new_n14254_), .C(rst), .Y(u2__0root_452_0__157_));
AOI21X1 AOI21X1_1994 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4601_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14266_));
AOI21X1 AOI21X1_1995 ( .A(u2__abc_52138_new_n14267_), .B(u2__abc_52138_new_n14262_), .C(rst), .Y(u2__0root_452_0__158_));
AOI21X1 AOI21X1_1996 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4543_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14274_));
AOI21X1 AOI21X1_1997 ( .A(u2__abc_52138_new_n14275_), .B(u2__abc_52138_new_n14269_), .C(rst), .Y(u2__0root_452_0__159_));
AOI21X1 AOI21X1_1998 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4536_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14282_));
AOI21X1 AOI21X1_1999 ( .A(u2__abc_52138_new_n14283_), .B(u2__abc_52138_new_n14277_), .C(rst), .Y(u2__0root_452_0__160_));
AOI21X1 AOI21X1_2 ( .A(_abc_65734_new_n1479_), .B(\a[116] ), .C(\a[117] ), .Y(_abc_65734_new_n1480_));
AOI21X1 AOI21X1_20 ( .A(u2__abc_52138_new_n3234_), .B(u2__abc_52138_new_n3147_), .C(u2__abc_52138_new_n3233_), .Y(u2__abc_52138_new_n3235_));
AOI21X1 AOI21X1_200 ( .A(u2__abc_52138_new_n6650_), .B(u2__abc_52138_new_n6642_), .C(rst), .Y(u2__0remHi_451_0__14_));
AOI21X1 AOI21X1_2000 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4525_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14290_));
AOI21X1 AOI21X1_2001 ( .A(u2__abc_52138_new_n14291_), .B(u2__abc_52138_new_n14285_), .C(rst), .Y(u2__0root_452_0__161_));
AOI21X1 AOI21X1_2002 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4530_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14297_));
AOI21X1 AOI21X1_2003 ( .A(u2__abc_52138_new_n14298_), .B(u2__abc_52138_new_n14293_), .C(rst), .Y(u2__0root_452_0__162_));
AOI21X1 AOI21X1_2004 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4564_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14305_));
AOI21X1 AOI21X1_2005 ( .A(u2__abc_52138_new_n14306_), .B(u2__abc_52138_new_n14300_), .C(rst), .Y(u2__0root_452_0__163_));
AOI21X1 AOI21X1_2006 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4559_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14313_));
AOI21X1 AOI21X1_2007 ( .A(u2__abc_52138_new_n14314_), .B(u2__abc_52138_new_n14308_), .C(rst), .Y(u2__0root_452_0__164_));
AOI21X1 AOI21X1_2008 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4548_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14321_));
AOI21X1 AOI21X1_2009 ( .A(u2__abc_52138_new_n14322_), .B(u2__abc_52138_new_n14316_), .C(rst), .Y(u2__0root_452_0__165_));
AOI21X1 AOI21X1_201 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3177_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6660_));
AOI21X1 AOI21X1_2010 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4553_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14328_));
AOI21X1 AOI21X1_2011 ( .A(u2__abc_52138_new_n14329_), .B(u2__abc_52138_new_n14324_), .C(rst), .Y(u2__0root_452_0__166_));
AOI21X1 AOI21X1_2012 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4519_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14336_));
AOI21X1 AOI21X1_2013 ( .A(u2__abc_52138_new_n14337_), .B(u2__abc_52138_new_n14331_), .C(rst), .Y(u2__0root_452_0__167_));
AOI21X1 AOI21X1_2014 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4512_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14344_));
AOI21X1 AOI21X1_2015 ( .A(u2__abc_52138_new_n14345_), .B(u2__abc_52138_new_n14339_), .C(rst), .Y(u2__0root_452_0__168_));
AOI21X1 AOI21X1_2016 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4501_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14352_));
AOI21X1 AOI21X1_2017 ( .A(u2__abc_52138_new_n14353_), .B(u2__abc_52138_new_n14347_), .C(rst), .Y(u2__0root_452_0__169_));
AOI21X1 AOI21X1_2018 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4506_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14359_));
AOI21X1 AOI21X1_2019 ( .A(u2__abc_52138_new_n14360_), .B(u2__abc_52138_new_n14355_), .C(rst), .Y(u2__0root_452_0__170_));
AOI21X1 AOI21X1_202 ( .A(u2__abc_52138_new_n6661_), .B(u2__abc_52138_new_n6652_), .C(rst), .Y(u2__0remHi_451_0__15_));
AOI21X1 AOI21X1_2020 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4494_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14367_));
AOI21X1 AOI21X1_2021 ( .A(u2__abc_52138_new_n14368_), .B(u2__abc_52138_new_n14362_), .C(rst), .Y(u2__0root_452_0__171_));
AOI21X1 AOI21X1_2022 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4489_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14375_));
AOI21X1 AOI21X1_2023 ( .A(u2__abc_52138_new_n14376_), .B(u2__abc_52138_new_n14370_), .C(rst), .Y(u2__0root_452_0__172_));
AOI21X1 AOI21X1_2024 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4478_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14383_));
AOI21X1 AOI21X1_2025 ( .A(u2__abc_52138_new_n14384_), .B(u2__abc_52138_new_n14378_), .C(rst), .Y(u2__0root_452_0__173_));
AOI21X1 AOI21X1_2026 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4483_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14390_));
AOI21X1 AOI21X1_2027 ( .A(u2__abc_52138_new_n14391_), .B(u2__abc_52138_new_n14386_), .C(rst), .Y(u2__0root_452_0__174_));
AOI21X1 AOI21X1_2028 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4463_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14398_));
AOI21X1 AOI21X1_2029 ( .A(u2__abc_52138_new_n14399_), .B(u2__abc_52138_new_n14393_), .C(rst), .Y(u2__0root_452_0__175_));
AOI21X1 AOI21X1_203 ( .A(u2__abc_52138_new_n6668_), .B(u2__abc_52138_new_n6669_), .C(u2__abc_52138_new_n6670_), .Y(u2__abc_52138_new_n6671_));
AOI21X1 AOI21X1_2030 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4469_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14406_));
AOI21X1 AOI21X1_2031 ( .A(u2__abc_52138_new_n14407_), .B(u2__abc_52138_new_n14401_), .C(rst), .Y(u2__0root_452_0__176_));
AOI21X1 AOI21X1_2032 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4452_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14414_));
AOI21X1 AOI21X1_2033 ( .A(u2__abc_52138_new_n14415_), .B(u2__abc_52138_new_n14409_), .C(rst), .Y(u2__0root_452_0__177_));
AOI21X1 AOI21X1_2034 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4457_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14421_));
AOI21X1 AOI21X1_2035 ( .A(u2__abc_52138_new_n14422_), .B(u2__abc_52138_new_n14417_), .C(rst), .Y(u2__0root_452_0__178_));
AOI21X1 AOI21X1_2036 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4445_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14429_));
AOI21X1 AOI21X1_2037 ( .A(u2__abc_52138_new_n14430_), .B(u2__abc_52138_new_n14424_), .C(rst), .Y(u2__0root_452_0__179_));
AOI21X1 AOI21X1_2038 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4440_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14437_));
AOI21X1 AOI21X1_2039 ( .A(u2__abc_52138_new_n14438_), .B(u2__abc_52138_new_n14432_), .C(rst), .Y(u2__0root_452_0__180_));
AOI21X1 AOI21X1_204 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3161_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6679_));
AOI21X1 AOI21X1_2040 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4429_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14445_));
AOI21X1 AOI21X1_2041 ( .A(u2__abc_52138_new_n14446_), .B(u2__abc_52138_new_n14440_), .C(rst), .Y(u2__0root_452_0__181_));
AOI21X1 AOI21X1_2042 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4434_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14452_));
AOI21X1 AOI21X1_2043 ( .A(u2__abc_52138_new_n14453_), .B(u2__abc_52138_new_n14448_), .C(rst), .Y(u2__0root_452_0__182_));
AOI21X1 AOI21X1_2044 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4382_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14460_));
AOI21X1 AOI21X1_2045 ( .A(u2__abc_52138_new_n14461_), .B(u2__abc_52138_new_n14455_), .C(rst), .Y(u2__0root_452_0__183_));
AOI21X1 AOI21X1_2046 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4387_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14468_));
AOI21X1 AOI21X1_2047 ( .A(u2__abc_52138_new_n14469_), .B(u2__abc_52138_new_n14463_), .C(rst), .Y(u2__0root_452_0__184_));
AOI21X1 AOI21X1_2048 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4393_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14476_));
AOI21X1 AOI21X1_2049 ( .A(u2__abc_52138_new_n14477_), .B(u2__abc_52138_new_n14471_), .C(rst), .Y(u2__0root_452_0__185_));
AOI21X1 AOI21X1_205 ( .A(u2__abc_52138_new_n6680_), .B(u2__abc_52138_new_n6663_), .C(rst), .Y(u2__0remHi_451_0__16_));
AOI21X1 AOI21X1_2050 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4398_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14483_));
AOI21X1 AOI21X1_2051 ( .A(u2__abc_52138_new_n14484_), .B(u2__abc_52138_new_n14479_), .C(rst), .Y(u2__0root_452_0__186_));
AOI21X1 AOI21X1_2052 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4421_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14491_));
AOI21X1 AOI21X1_2053 ( .A(u2__abc_52138_new_n14492_), .B(u2__abc_52138_new_n14486_), .C(rst), .Y(u2__0root_452_0__187_));
AOI21X1 AOI21X1_2054 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4416_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14499_));
AOI21X1 AOI21X1_2055 ( .A(u2__abc_52138_new_n14500_), .B(u2__abc_52138_new_n14494_), .C(rst), .Y(u2__0root_452_0__188_));
AOI21X1 AOI21X1_2056 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4405_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14507_));
AOI21X1 AOI21X1_2057 ( .A(u2__abc_52138_new_n14508_), .B(u2__abc_52138_new_n14502_), .C(rst), .Y(u2__0root_452_0__189_));
AOI21X1 AOI21X1_2058 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4410_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14514_));
AOI21X1 AOI21X1_2059 ( .A(u2__abc_52138_new_n14515_), .B(u2__abc_52138_new_n14510_), .C(rst), .Y(u2__0root_452_0__190_));
AOI21X1 AOI21X1_206 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3166_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6687_));
AOI21X1 AOI21X1_2060 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4366_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14522_));
AOI21X1 AOI21X1_2061 ( .A(u2__abc_52138_new_n14523_), .B(u2__abc_52138_new_n14517_), .C(rst), .Y(u2__0root_452_0__191_));
AOI21X1 AOI21X1_2062 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4372_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14530_));
AOI21X1 AOI21X1_2063 ( .A(u2__abc_52138_new_n14531_), .B(u2__abc_52138_new_n14525_), .C(rst), .Y(u2__0root_452_0__192_));
AOI21X1 AOI21X1_2064 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4356_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14538_));
AOI21X1 AOI21X1_2065 ( .A(u2__abc_52138_new_n14539_), .B(u2__abc_52138_new_n14533_), .C(rst), .Y(u2__0root_452_0__193_));
AOI21X1 AOI21X1_2066 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4358_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14545_));
AOI21X1 AOI21X1_2067 ( .A(u2__abc_52138_new_n14546_), .B(u2__abc_52138_new_n14541_), .C(rst), .Y(u2__0root_452_0__194_));
AOI21X1 AOI21X1_2068 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4347_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14553_));
AOI21X1 AOI21X1_2069 ( .A(u2__abc_52138_new_n14554_), .B(u2__abc_52138_new_n14548_), .C(rst), .Y(u2__0root_452_0__195_));
AOI21X1 AOI21X1_207 ( .A(u2__abc_52138_new_n6688_), .B(u2__abc_52138_new_n6682_), .C(rst), .Y(u2__0remHi_451_0__17_));
AOI21X1 AOI21X1_2070 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4342_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14561_));
AOI21X1 AOI21X1_2071 ( .A(u2__abc_52138_new_n14562_), .B(u2__abc_52138_new_n14556_), .C(rst), .Y(u2__0root_452_0__196_));
AOI21X1 AOI21X1_2072 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4331_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14569_));
AOI21X1 AOI21X1_2073 ( .A(u2__abc_52138_new_n14570_), .B(u2__abc_52138_new_n14564_), .C(rst), .Y(u2__0root_452_0__197_));
AOI21X1 AOI21X1_2074 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4336_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14576_));
AOI21X1 AOI21X1_2075 ( .A(u2__abc_52138_new_n14577_), .B(u2__abc_52138_new_n14572_), .C(rst), .Y(u2__0root_452_0__198_));
AOI21X1 AOI21X1_2076 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4305_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14584_));
AOI21X1 AOI21X1_2077 ( .A(u2__abc_52138_new_n14585_), .B(u2__abc_52138_new_n14579_), .C(rst), .Y(u2__0root_452_0__199_));
AOI21X1 AOI21X1_2078 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4300_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14592_));
AOI21X1 AOI21X1_2079 ( .A(u2__abc_52138_new_n14593_), .B(u2__abc_52138_new_n14587_), .C(rst), .Y(u2__0root_452_0__200_));
AOI21X1 AOI21X1_208 ( .A(u2__abc_52138_new_n6683_), .B(u2__abc_52138_new_n3178_), .C(u2__abc_52138_new_n6692_), .Y(u2__abc_52138_new_n6693_));
AOI21X1 AOI21X1_2080 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4289_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14600_));
AOI21X1 AOI21X1_2081 ( .A(u2__abc_52138_new_n14601_), .B(u2__abc_52138_new_n14595_), .C(rst), .Y(u2__0root_452_0__201_));
AOI21X1 AOI21X1_2082 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4294_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14607_));
AOI21X1 AOI21X1_2083 ( .A(u2__abc_52138_new_n14608_), .B(u2__abc_52138_new_n14603_), .C(rst), .Y(u2__0root_452_0__202_));
AOI21X1 AOI21X1_2084 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n14615_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14616_));
AOI21X1 AOI21X1_2085 ( .A(u2__abc_52138_new_n14617_), .B(u2__abc_52138_new_n14610_), .C(rst), .Y(u2__0root_452_0__203_));
AOI21X1 AOI21X1_2086 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4325_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14624_));
AOI21X1 AOI21X1_2087 ( .A(u2__abc_52138_new_n14625_), .B(u2__abc_52138_new_n14619_), .C(rst), .Y(u2__0root_452_0__204_));
AOI21X1 AOI21X1_2088 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4312_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14632_));
AOI21X1 AOI21X1_2089 ( .A(u2__abc_52138_new_n14633_), .B(u2__abc_52138_new_n14627_), .C(rst), .Y(u2__0root_452_0__205_));
AOI21X1 AOI21X1_209 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3191_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6698_));
AOI21X1 AOI21X1_2090 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4317_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14639_));
AOI21X1 AOI21X1_2091 ( .A(u2__abc_52138_new_n14640_), .B(u2__abc_52138_new_n14635_), .C(rst), .Y(u2__0root_452_0__206_));
AOI21X1 AOI21X1_2092 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4252_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14647_));
AOI21X1 AOI21X1_2093 ( .A(u2__abc_52138_new_n14648_), .B(u2__abc_52138_new_n14642_), .C(rst), .Y(u2__0root_452_0__207_));
AOI21X1 AOI21X1_2094 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4257_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14655_));
AOI21X1 AOI21X1_2095 ( .A(u2__abc_52138_new_n14656_), .B(u2__abc_52138_new_n14650_), .C(rst), .Y(u2__0root_452_0__208_));
AOI21X1 AOI21X1_2096 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4241_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14663_));
AOI21X1 AOI21X1_2097 ( .A(u2__abc_52138_new_n14664_), .B(u2__abc_52138_new_n14658_), .C(rst), .Y(u2__0root_452_0__209_));
AOI21X1 AOI21X1_2098 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4246_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14670_));
AOI21X1 AOI21X1_2099 ( .A(u2__abc_52138_new_n14671_), .B(u2__abc_52138_new_n14666_), .C(rst), .Y(u2__0root_452_0__210_));
AOI21X1 AOI21X1_21 ( .A(u2__abc_52138_new_n3228_), .B(u2__abc_52138_new_n3218_), .C(u2__abc_52138_new_n3236_), .Y(u2__abc_52138_new_n3237_));
AOI21X1 AOI21X1_210 ( .A(u2__abc_52138_new_n6699_), .B(u2__abc_52138_new_n6690_), .C(rst), .Y(u2__0remHi_451_0__18_));
AOI21X1 AOI21X1_2100 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4282_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14678_));
AOI21X1 AOI21X1_2101 ( .A(u2__abc_52138_new_n14679_), .B(u2__abc_52138_new_n14673_), .C(rst), .Y(u2__0root_452_0__211_));
AOI21X1 AOI21X1_2102 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4277_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14686_));
AOI21X1 AOI21X1_2103 ( .A(u2__abc_52138_new_n14687_), .B(u2__abc_52138_new_n14681_), .C(rst), .Y(u2__0root_452_0__212_));
AOI21X1 AOI21X1_2104 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4266_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14694_));
AOI21X1 AOI21X1_2105 ( .A(u2__abc_52138_new_n14695_), .B(u2__abc_52138_new_n14689_), .C(rst), .Y(u2__0root_452_0__213_));
AOI21X1 AOI21X1_2106 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4271_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14701_));
AOI21X1 AOI21X1_2107 ( .A(u2__abc_52138_new_n14702_), .B(u2__abc_52138_new_n14697_), .C(rst), .Y(u2__0root_452_0__214_));
AOI21X1 AOI21X1_2108 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4205_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14709_));
AOI21X1 AOI21X1_2109 ( .A(u2__abc_52138_new_n14710_), .B(u2__abc_52138_new_n14704_), .C(rst), .Y(u2__0root_452_0__215_));
AOI21X1 AOI21X1_211 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n6706_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6707_));
AOI21X1 AOI21X1_2110 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4210_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14717_));
AOI21X1 AOI21X1_2111 ( .A(u2__abc_52138_new_n14718_), .B(u2__abc_52138_new_n14712_), .C(rst), .Y(u2__0root_452_0__216_));
AOI21X1 AOI21X1_2112 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4194_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14725_));
AOI21X1 AOI21X1_2113 ( .A(u2__abc_52138_new_n14726_), .B(u2__abc_52138_new_n14720_), .C(rst), .Y(u2__0root_452_0__217_));
AOI21X1 AOI21X1_2114 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4199_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14732_));
AOI21X1 AOI21X1_2115 ( .A(u2__abc_52138_new_n14733_), .B(u2__abc_52138_new_n14728_), .C(rst), .Y(u2__0root_452_0__218_));
AOI21X1 AOI21X1_2116 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4233_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14740_));
AOI21X1 AOI21X1_2117 ( .A(u2__abc_52138_new_n14741_), .B(u2__abc_52138_new_n14735_), .C(rst), .Y(u2__0root_452_0__219_));
AOI21X1 AOI21X1_2118 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4230_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14748_));
AOI21X1 AOI21X1_2119 ( .A(u2__abc_52138_new_n14749_), .B(u2__abc_52138_new_n14743_), .C(rst), .Y(u2__0root_452_0__220_));
AOI21X1 AOI21X1_212 ( .A(u2__abc_52138_new_n6708_), .B(u2__abc_52138_new_n6701_), .C(rst), .Y(u2__0remHi_451_0__19_));
AOI21X1 AOI21X1_2120 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4217_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14756_));
AOI21X1 AOI21X1_2121 ( .A(u2__abc_52138_new_n14757_), .B(u2__abc_52138_new_n14751_), .C(rst), .Y(u2__0root_452_0__221_));
AOI21X1 AOI21X1_2122 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4222_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14763_));
AOI21X1 AOI21X1_2123 ( .A(u2__abc_52138_new_n14764_), .B(u2__abc_52138_new_n14759_), .C(rst), .Y(u2__0root_452_0__222_));
AOI21X1 AOI21X1_2124 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4162_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14771_));
AOI21X1 AOI21X1_2125 ( .A(u2__abc_52138_new_n14772_), .B(u2__abc_52138_new_n14766_), .C(rst), .Y(u2__0root_452_0__223_));
AOI21X1 AOI21X1_2126 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4157_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14779_));
AOI21X1 AOI21X1_2127 ( .A(u2__abc_52138_new_n14780_), .B(u2__abc_52138_new_n14774_), .C(rst), .Y(u2__0root_452_0__224_));
AOI21X1 AOI21X1_2128 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4146_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14787_));
AOI21X1 AOI21X1_2129 ( .A(u2__abc_52138_new_n14788_), .B(u2__abc_52138_new_n14782_), .C(rst), .Y(u2__0root_452_0__225_));
AOI21X1 AOI21X1_213 ( .A(u2__abc_52138_new_n6691_), .B(u2__abc_52138_new_n3167_), .C(u2__abc_52138_new_n6713_), .Y(u2__abc_52138_new_n6714_));
AOI21X1 AOI21X1_2130 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4151_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14794_));
AOI21X1 AOI21X1_2131 ( .A(u2__abc_52138_new_n14795_), .B(u2__abc_52138_new_n14790_), .C(rst), .Y(u2__0root_452_0__226_));
AOI21X1 AOI21X1_2132 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4187_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14802_));
AOI21X1 AOI21X1_2133 ( .A(u2__abc_52138_new_n14803_), .B(u2__abc_52138_new_n14797_), .C(rst), .Y(u2__0root_452_0__227_));
AOI21X1 AOI21X1_2134 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4182_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14810_));
AOI21X1 AOI21X1_2135 ( .A(u2__abc_52138_new_n14811_), .B(u2__abc_52138_new_n14805_), .C(rst), .Y(u2__0root_452_0__228_));
AOI21X1 AOI21X1_2136 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4169_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14818_));
AOI21X1 AOI21X1_2137 ( .A(u2__abc_52138_new_n14819_), .B(u2__abc_52138_new_n14813_), .C(rst), .Y(u2__0root_452_0__229_));
AOI21X1 AOI21X1_2138 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4174_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14825_));
AOI21X1 AOI21X1_2139 ( .A(u2__abc_52138_new_n14826_), .B(u2__abc_52138_new_n14821_), .C(rst), .Y(u2__0root_452_0__230_));
AOI21X1 AOI21X1_214 ( .A(u2__abc_52138_new_n6673_), .B(u2__abc_52138_new_n3181_), .C(u2__abc_52138_new_n6715_), .Y(u2__abc_52138_new_n6716_));
AOI21X1 AOI21X1_2140 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4140_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14833_));
AOI21X1 AOI21X1_2141 ( .A(u2__abc_52138_new_n14834_), .B(u2__abc_52138_new_n14828_), .C(rst), .Y(u2__0root_452_0__231_));
AOI21X1 AOI21X1_2142 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4960_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14841_));
AOI21X1 AOI21X1_2143 ( .A(u2__abc_52138_new_n14842_), .B(u2__abc_52138_new_n14836_), .C(rst), .Y(u2__0root_452_0__232_));
AOI21X1 AOI21X1_2144 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4123_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14849_));
AOI21X1 AOI21X1_2145 ( .A(u2__abc_52138_new_n14850_), .B(u2__abc_52138_new_n14844_), .C(rst), .Y(u2__0root_452_0__233_));
AOI21X1 AOI21X1_2146 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4128_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14856_));
AOI21X1 AOI21X1_2147 ( .A(u2__abc_52138_new_n14857_), .B(u2__abc_52138_new_n14852_), .C(rst), .Y(u2__0root_452_0__234_));
AOI21X1 AOI21X1_2148 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4115_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14864_));
AOI21X1 AOI21X1_2149 ( .A(u2__abc_52138_new_n14865_), .B(u2__abc_52138_new_n14859_), .C(rst), .Y(u2__0root_452_0__235_));
AOI21X1 AOI21X1_215 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3211_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6721_));
AOI21X1 AOI21X1_2150 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4110_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14872_));
AOI21X1 AOI21X1_2151 ( .A(u2__abc_52138_new_n14873_), .B(u2__abc_52138_new_n14867_), .C(rst), .Y(u2__0root_452_0__236_));
AOI21X1 AOI21X1_2152 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4099_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14880_));
AOI21X1 AOI21X1_2153 ( .A(u2__abc_52138_new_n14881_), .B(u2__abc_52138_new_n14875_), .C(rst), .Y(u2__0root_452_0__237_));
AOI21X1 AOI21X1_2154 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4104_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14887_));
AOI21X1 AOI21X1_2155 ( .A(u2__abc_52138_new_n14888_), .B(u2__abc_52138_new_n14883_), .C(rst), .Y(u2__0root_452_0__238_));
AOI21X1 AOI21X1_2156 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4050_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14895_));
AOI21X1 AOI21X1_2157 ( .A(u2__abc_52138_new_n14896_), .B(u2__abc_52138_new_n14890_), .C(rst), .Y(u2__0root_452_0__239_));
AOI21X1 AOI21X1_2158 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4055_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14903_));
AOI21X1 AOI21X1_2159 ( .A(u2__abc_52138_new_n14904_), .B(u2__abc_52138_new_n14898_), .C(rst), .Y(u2__0root_452_0__240_));
AOI21X1 AOI21X1_216 ( .A(u2__abc_52138_new_n6722_), .B(u2__abc_52138_new_n6710_), .C(rst), .Y(u2__0remHi_451_0__20_));
AOI21X1 AOI21X1_2160 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4061_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14911_));
AOI21X1 AOI21X1_2161 ( .A(u2__abc_52138_new_n14912_), .B(u2__abc_52138_new_n14906_), .C(rst), .Y(u2__0root_452_0__241_));
AOI21X1 AOI21X1_2162 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4066_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14918_));
AOI21X1 AOI21X1_2163 ( .A(u2__abc_52138_new_n14919_), .B(u2__abc_52138_new_n14914_), .C(rst), .Y(u2__0root_452_0__242_));
AOI21X1 AOI21X1_2164 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4090_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14926_));
AOI21X1 AOI21X1_2165 ( .A(u2__abc_52138_new_n14927_), .B(u2__abc_52138_new_n14921_), .C(rst), .Y(u2__0root_452_0__243_));
AOI21X1 AOI21X1_2166 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4087_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14934_));
AOI21X1 AOI21X1_2167 ( .A(u2__abc_52138_new_n14935_), .B(u2__abc_52138_new_n14929_), .C(rst), .Y(u2__0root_452_0__244_));
AOI21X1 AOI21X1_2168 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4074_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14942_));
AOI21X1 AOI21X1_2169 ( .A(u2__abc_52138_new_n14943_), .B(u2__abc_52138_new_n14937_), .C(rst), .Y(u2__0root_452_0__245_));
AOI21X1 AOI21X1_217 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3185_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6729_));
AOI21X1 AOI21X1_2170 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4079_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14949_));
AOI21X1 AOI21X1_2171 ( .A(u2__abc_52138_new_n14950_), .B(u2__abc_52138_new_n14945_), .C(rst), .Y(u2__0root_452_0__246_));
AOI21X1 AOI21X1_2172 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4003_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14957_));
AOI21X1 AOI21X1_2173 ( .A(u2__abc_52138_new_n14958_), .B(u2__abc_52138_new_n14952_), .C(rst), .Y(u2__0root_452_0__247_));
AOI21X1 AOI21X1_2174 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4008_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14965_));
AOI21X1 AOI21X1_2175 ( .A(u2__abc_52138_new_n14966_), .B(u2__abc_52138_new_n14960_), .C(rst), .Y(u2__0root_452_0__248_));
AOI21X1 AOI21X1_2176 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4014_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14973_));
AOI21X1 AOI21X1_2177 ( .A(u2__abc_52138_new_n14974_), .B(u2__abc_52138_new_n14968_), .C(rst), .Y(u2__0root_452_0__249_));
AOI21X1 AOI21X1_2178 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4019_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14980_));
AOI21X1 AOI21X1_2179 ( .A(u2__abc_52138_new_n14981_), .B(u2__abc_52138_new_n14976_), .C(rst), .Y(u2__0root_452_0__250_));
AOI21X1 AOI21X1_218 ( .A(u2__abc_52138_new_n6730_), .B(u2__abc_52138_new_n6724_), .C(rst), .Y(u2__0remHi_451_0__21_));
AOI21X1 AOI21X1_2180 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4042_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14988_));
AOI21X1 AOI21X1_2181 ( .A(u2__abc_52138_new_n14989_), .B(u2__abc_52138_new_n14983_), .C(rst), .Y(u2__0root_452_0__251_));
AOI21X1 AOI21X1_2182 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4037_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n14996_));
AOI21X1 AOI21X1_2183 ( .A(u2__abc_52138_new_n14997_), .B(u2__abc_52138_new_n14991_), .C(rst), .Y(u2__0root_452_0__252_));
AOI21X1 AOI21X1_2184 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4026_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15004_));
AOI21X1 AOI21X1_2185 ( .A(u2__abc_52138_new_n15005_), .B(u2__abc_52138_new_n14999_), .C(rst), .Y(u2__0root_452_0__253_));
AOI21X1 AOI21X1_2186 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4033_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15011_));
AOI21X1 AOI21X1_2187 ( .A(u2__abc_52138_new_n15012_), .B(u2__abc_52138_new_n15007_), .C(rst), .Y(u2__0root_452_0__254_));
AOI21X1 AOI21X1_2188 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5687_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15019_));
AOI21X1 AOI21X1_2189 ( .A(u2__abc_52138_new_n15020_), .B(u2__abc_52138_new_n15014_), .C(rst), .Y(u2__0root_452_0__255_));
AOI21X1 AOI21X1_219 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3130_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6743_));
AOI21X1 AOI21X1_2190 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5692_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15027_));
AOI21X1 AOI21X1_2191 ( .A(u2__abc_52138_new_n15028_), .B(u2__abc_52138_new_n15022_), .C(rst), .Y(u2__0root_452_0__256_));
AOI21X1 AOI21X1_2192 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5699_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15035_));
AOI21X1 AOI21X1_2193 ( .A(u2__abc_52138_new_n15036_), .B(u2__abc_52138_new_n15030_), .C(rst), .Y(u2__0root_452_0__257_));
AOI21X1 AOI21X1_2194 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5704_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15042_));
AOI21X1 AOI21X1_2195 ( .A(u2__abc_52138_new_n15043_), .B(u2__abc_52138_new_n15038_), .C(rst), .Y(u2__0root_452_0__258_));
AOI21X1 AOI21X1_2196 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5722_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15050_));
AOI21X1 AOI21X1_2197 ( .A(u2__abc_52138_new_n15051_), .B(u2__abc_52138_new_n15045_), .C(rst), .Y(u2__0root_452_0__259_));
AOI21X1 AOI21X1_2198 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5727_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15058_));
AOI21X1 AOI21X1_2199 ( .A(u2__abc_52138_new_n15059_), .B(u2__abc_52138_new_n15053_), .C(rst), .Y(u2__0root_452_0__260_));
AOI21X1 AOI21X1_22 ( .A(u2__abc_52138_new_n3196_), .B(u2__abc_52138_new_n3111_), .C(u2__abc_52138_new_n3238_), .Y(u2__abc_52138_new_n3239_));
AOI21X1 AOI21X1_220 ( .A(u2__abc_52138_new_n6744_), .B(u2__abc_52138_new_n6732_), .C(rst), .Y(u2__0remHi_451_0__22_));
AOI21X1 AOI21X1_2200 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5711_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15066_));
AOI21X1 AOI21X1_2201 ( .A(u2__abc_52138_new_n15067_), .B(u2__abc_52138_new_n15061_), .C(rst), .Y(u2__0root_452_0__261_));
AOI21X1 AOI21X1_2202 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5716_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15073_));
AOI21X1 AOI21X1_2203 ( .A(u2__abc_52138_new_n15074_), .B(u2__abc_52138_new_n15069_), .C(rst), .Y(u2__0root_452_0__262_));
AOI21X1 AOI21X1_2204 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5674_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15081_));
AOI21X1 AOI21X1_2205 ( .A(u2__abc_52138_new_n15082_), .B(u2__abc_52138_new_n15076_), .C(rst), .Y(u2__0root_452_0__263_));
AOI21X1 AOI21X1_2206 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5679_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15089_));
AOI21X1 AOI21X1_2207 ( .A(u2__abc_52138_new_n15090_), .B(u2__abc_52138_new_n15084_), .C(rst), .Y(u2__0root_452_0__264_));
AOI21X1 AOI21X1_2208 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5665_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15097_));
AOI21X1 AOI21X1_2209 ( .A(u2__abc_52138_new_n15098_), .B(u2__abc_52138_new_n15092_), .C(rst), .Y(u2__0root_452_0__265_));
AOI21X1 AOI21X1_221 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3125_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6752_));
AOI21X1 AOI21X1_2210 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5670_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15104_));
AOI21X1 AOI21X1_2211 ( .A(u2__abc_52138_new_n15105_), .B(u2__abc_52138_new_n15100_), .C(rst), .Y(u2__0root_452_0__266_));
AOI21X1 AOI21X1_2212 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5653_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15112_));
AOI21X1 AOI21X1_2213 ( .A(u2__abc_52138_new_n15113_), .B(u2__abc_52138_new_n15107_), .C(rst), .Y(u2__0root_452_0__267_));
AOI21X1 AOI21X1_2214 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5658_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15120_));
AOI21X1 AOI21X1_2215 ( .A(u2__abc_52138_new_n15121_), .B(u2__abc_52138_new_n15115_), .C(rst), .Y(u2__0root_452_0__268_));
AOI21X1 AOI21X1_2216 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5640_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15128_));
AOI21X1 AOI21X1_2217 ( .A(u2__abc_52138_new_n15129_), .B(u2__abc_52138_new_n15123_), .C(rst), .Y(u2__0root_452_0__269_));
AOI21X1 AOI21X1_2218 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5645_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15135_));
AOI21X1 AOI21X1_2219 ( .A(u2__abc_52138_new_n15136_), .B(u2__abc_52138_new_n15131_), .C(rst), .Y(u2__0root_452_0__270_));
AOI21X1 AOI21X1_222 ( .A(u2__abc_52138_new_n6753_), .B(u2__abc_52138_new_n6746_), .C(rst), .Y(u2__0remHi_451_0__23_));
AOI21X1 AOI21X1_2220 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5608_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15143_));
AOI21X1 AOI21X1_2221 ( .A(u2__abc_52138_new_n15144_), .B(u2__abc_52138_new_n15138_), .C(rst), .Y(u2__0root_452_0__271_));
AOI21X1 AOI21X1_2222 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5613_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15151_));
AOI21X1 AOI21X1_2223 ( .A(u2__abc_52138_new_n15152_), .B(u2__abc_52138_new_n15146_), .C(rst), .Y(u2__0root_452_0__272_));
AOI21X1 AOI21X1_2224 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5597_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15159_));
AOI21X1 AOI21X1_2225 ( .A(u2__abc_52138_new_n15160_), .B(u2__abc_52138_new_n15154_), .C(rst), .Y(u2__0root_452_0__273_));
AOI21X1 AOI21X1_2226 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5602_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15166_));
AOI21X1 AOI21X1_2227 ( .A(u2__abc_52138_new_n15167_), .B(u2__abc_52138_new_n15162_), .C(rst), .Y(u2__0root_452_0__274_));
AOI21X1 AOI21X1_2228 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5761_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15174_));
AOI21X1 AOI21X1_2229 ( .A(u2__abc_52138_new_n15175_), .B(u2__abc_52138_new_n15169_), .C(rst), .Y(u2__0root_452_0__275_));
AOI21X1 AOI21X1_223 ( .A(u2__abc_52138_new_n6760_), .B(u2__abc_52138_new_n3186_), .C(u2__abc_52138_new_n3213_), .Y(u2__abc_52138_new_n6761_));
AOI21X1 AOI21X1_2230 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5632_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15182_));
AOI21X1 AOI21X1_2231 ( .A(u2__abc_52138_new_n15183_), .B(u2__abc_52138_new_n15177_), .C(rst), .Y(u2__0root_452_0__276_));
AOI21X1 AOI21X1_2232 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5620_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15190_));
AOI21X1 AOI21X1_2233 ( .A(u2__abc_52138_new_n15191_), .B(u2__abc_52138_new_n15185_), .C(rst), .Y(u2__0root_452_0__277_));
AOI21X1 AOI21X1_2234 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5625_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15197_));
AOI21X1 AOI21X1_2235 ( .A(u2__abc_52138_new_n15198_), .B(u2__abc_52138_new_n15193_), .C(rst), .Y(u2__0root_452_0__278_));
AOI21X1 AOI21X1_2236 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5561_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15205_));
AOI21X1 AOI21X1_2237 ( .A(u2__abc_52138_new_n15206_), .B(u2__abc_52138_new_n15200_), .C(rst), .Y(u2__0root_452_0__279_));
AOI21X1 AOI21X1_2238 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5566_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15213_));
AOI21X1 AOI21X1_2239 ( .A(u2__abc_52138_new_n15214_), .B(u2__abc_52138_new_n15208_), .C(rst), .Y(u2__0root_452_0__280_));
AOI21X1 AOI21X1_224 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3114_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6769_));
AOI21X1 AOI21X1_2240 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5550_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15221_));
AOI21X1 AOI21X1_2241 ( .A(u2__abc_52138_new_n15222_), .B(u2__abc_52138_new_n15216_), .C(rst), .Y(u2__0root_452_0__281_));
AOI21X1 AOI21X1_2242 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5555_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15228_));
AOI21X1 AOI21X1_2243 ( .A(u2__abc_52138_new_n15229_), .B(u2__abc_52138_new_n15224_), .C(rst), .Y(u2__0root_452_0__282_));
AOI21X1 AOI21X1_2244 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5584_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15236_));
AOI21X1 AOI21X1_2245 ( .A(u2__abc_52138_new_n15237_), .B(u2__abc_52138_new_n15231_), .C(rst), .Y(u2__0root_452_0__283_));
AOI21X1 AOI21X1_2246 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5589_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15244_));
AOI21X1 AOI21X1_2247 ( .A(u2__abc_52138_new_n15245_), .B(u2__abc_52138_new_n15239_), .C(rst), .Y(u2__0root_452_0__284_));
AOI21X1 AOI21X1_2248 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5573_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15252_));
AOI21X1 AOI21X1_2249 ( .A(u2__abc_52138_new_n15253_), .B(u2__abc_52138_new_n15247_), .C(rst), .Y(u2__0root_452_0__285_));
AOI21X1 AOI21X1_225 ( .A(u2__abc_52138_new_n6770_), .B(u2__abc_52138_new_n6755_), .C(rst), .Y(u2__0remHi_451_0__24_));
AOI21X1 AOI21X1_2250 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5578_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15259_));
AOI21X1 AOI21X1_2251 ( .A(u2__abc_52138_new_n15260_), .B(u2__abc_52138_new_n15255_), .C(rst), .Y(u2__0root_452_0__286_));
AOI21X1 AOI21X1_2252 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5515_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15267_));
AOI21X1 AOI21X1_2253 ( .A(u2__abc_52138_new_n15268_), .B(u2__abc_52138_new_n15262_), .C(rst), .Y(u2__0root_452_0__287_));
AOI21X1 AOI21X1_2254 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5520_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15275_));
AOI21X1 AOI21X1_2255 ( .A(u2__abc_52138_new_n15276_), .B(u2__abc_52138_new_n15270_), .C(rst), .Y(u2__0root_452_0__288_));
AOI21X1 AOI21X1_2256 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5504_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15283_));
AOI21X1 AOI21X1_2257 ( .A(u2__abc_52138_new_n15284_), .B(u2__abc_52138_new_n15278_), .C(rst), .Y(u2__0root_452_0__289_));
AOI21X1 AOI21X1_2258 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5509_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15290_));
AOI21X1 AOI21X1_2259 ( .A(u2__abc_52138_new_n15291_), .B(u2__abc_52138_new_n15286_), .C(rst), .Y(u2__0root_452_0__290_));
AOI21X1 AOI21X1_226 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3119_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6777_));
AOI21X1 AOI21X1_2260 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5787_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15298_));
AOI21X1 AOI21X1_2261 ( .A(u2__abc_52138_new_n15299_), .B(u2__abc_52138_new_n15293_), .C(rst), .Y(u2__0root_452_0__291_));
AOI21X1 AOI21X1_2262 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5539_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15306_));
AOI21X1 AOI21X1_2263 ( .A(u2__abc_52138_new_n15307_), .B(u2__abc_52138_new_n15301_), .C(rst), .Y(u2__0root_452_0__292_));
AOI21X1 AOI21X1_2264 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5527_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15314_));
AOI21X1 AOI21X1_2265 ( .A(u2__abc_52138_new_n15315_), .B(u2__abc_52138_new_n15309_), .C(rst), .Y(u2__0root_452_0__293_));
AOI21X1 AOI21X1_2266 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5532_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15321_));
AOI21X1 AOI21X1_2267 ( .A(u2__abc_52138_new_n15322_), .B(u2__abc_52138_new_n15317_), .C(rst), .Y(u2__0root_452_0__294_));
AOI21X1 AOI21X1_2268 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5455_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15329_));
AOI21X1 AOI21X1_2269 ( .A(u2__abc_52138_new_n15330_), .B(u2__abc_52138_new_n15324_), .C(rst), .Y(u2__0root_452_0__295_));
AOI21X1 AOI21X1_227 ( .A(u2__abc_52138_new_n6778_), .B(u2__abc_52138_new_n6772_), .C(rst), .Y(u2__0remHi_451_0__25_));
AOI21X1 AOI21X1_2270 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5462_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15337_));
AOI21X1 AOI21X1_2271 ( .A(u2__abc_52138_new_n15338_), .B(u2__abc_52138_new_n15332_), .C(rst), .Y(u2__0root_452_0__296_));
AOI21X1 AOI21X1_2272 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5468_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15345_));
AOI21X1 AOI21X1_2273 ( .A(u2__abc_52138_new_n15346_), .B(u2__abc_52138_new_n15340_), .C(rst), .Y(u2__0root_452_0__297_));
AOI21X1 AOI21X1_2274 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5473_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15352_));
AOI21X1 AOI21X1_2275 ( .A(u2__abc_52138_new_n15353_), .B(u2__abc_52138_new_n15348_), .C(rst), .Y(u2__0root_452_0__298_));
AOI21X1 AOI21X1_2276 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5491_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15360_));
AOI21X1 AOI21X1_2277 ( .A(u2__abc_52138_new_n15361_), .B(u2__abc_52138_new_n15355_), .C(rst), .Y(u2__0root_452_0__299_));
AOI21X1 AOI21X1_2278 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5496_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15368_));
AOI21X1 AOI21X1_2279 ( .A(u2__abc_52138_new_n15369_), .B(u2__abc_52138_new_n15363_), .C(rst), .Y(u2__0root_452_0__300_));
AOI21X1 AOI21X1_228 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3153_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6789_));
AOI21X1 AOI21X1_2280 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5480_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15376_));
AOI21X1 AOI21X1_2281 ( .A(u2__abc_52138_new_n15377_), .B(u2__abc_52138_new_n15371_), .C(rst), .Y(u2__0root_452_0__301_));
AOI21X1 AOI21X1_2282 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5485_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15383_));
AOI21X1 AOI21X1_2283 ( .A(u2__abc_52138_new_n15384_), .B(u2__abc_52138_new_n15379_), .C(rst), .Y(u2__0root_452_0__302_));
AOI21X1 AOI21X1_2284 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5407_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15391_));
AOI21X1 AOI21X1_2285 ( .A(u2__abc_52138_new_n15392_), .B(u2__abc_52138_new_n15386_), .C(rst), .Y(u2__0root_452_0__303_));
AOI21X1 AOI21X1_2286 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5412_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15399_));
AOI21X1 AOI21X1_2287 ( .A(u2__abc_52138_new_n15400_), .B(u2__abc_52138_new_n15394_), .C(rst), .Y(u2__0root_452_0__304_));
AOI21X1 AOI21X1_2288 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5420_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15407_));
AOI21X1 AOI21X1_2289 ( .A(u2__abc_52138_new_n15408_), .B(u2__abc_52138_new_n15402_), .C(rst), .Y(u2__0root_452_0__305_));
AOI21X1 AOI21X1_229 ( .A(u2__abc_52138_new_n6790_), .B(u2__abc_52138_new_n6780_), .C(rst), .Y(u2__0remHi_451_0__26_));
AOI21X1 AOI21X1_2290 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5425_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15414_));
AOI21X1 AOI21X1_2291 ( .A(u2__abc_52138_new_n15415_), .B(u2__abc_52138_new_n15410_), .C(rst), .Y(u2__0root_452_0__306_));
AOI21X1 AOI21X1_2292 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5448_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15422_));
AOI21X1 AOI21X1_2293 ( .A(u2__abc_52138_new_n15423_), .B(u2__abc_52138_new_n15417_), .C(rst), .Y(u2__0root_452_0__307_));
AOI21X1 AOI21X1_2294 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5443_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15430_));
AOI21X1 AOI21X1_2295 ( .A(u2__abc_52138_new_n15431_), .B(u2__abc_52138_new_n15425_), .C(rst), .Y(u2__0root_452_0__308_));
AOI21X1 AOI21X1_2296 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5432_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15438_));
AOI21X1 AOI21X1_2297 ( .A(u2__abc_52138_new_n15439_), .B(u2__abc_52138_new_n15433_), .C(rst), .Y(u2__0root_452_0__309_));
AOI21X1 AOI21X1_2298 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5437_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15445_));
AOI21X1 AOI21X1_2299 ( .A(u2__abc_52138_new_n15446_), .B(u2__abc_52138_new_n15441_), .C(rst), .Y(u2__0root_452_0__310_));
AOI21X1 AOI21X1_23 ( .A(u2__abc_52138_new_n3434_), .B(u2__abc_52138_new_n3395_), .C(u2__abc_52138_new_n3435_), .Y(u2__abc_52138_new_n3436_));
AOI21X1 AOI21X1_230 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3148_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6797_));
AOI21X1 AOI21X1_2300 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5811_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15453_));
AOI21X1 AOI21X1_2301 ( .A(u2__abc_52138_new_n15454_), .B(u2__abc_52138_new_n15448_), .C(rst), .Y(u2__0root_452_0__311_));
AOI21X1 AOI21X1_2302 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5382_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15461_));
AOI21X1 AOI21X1_2303 ( .A(u2__abc_52138_new_n15462_), .B(u2__abc_52138_new_n15456_), .C(rst), .Y(u2__0root_452_0__312_));
AOI21X1 AOI21X1_2304 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5370_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15469_));
AOI21X1 AOI21X1_2305 ( .A(u2__abc_52138_new_n15470_), .B(u2__abc_52138_new_n15464_), .C(rst), .Y(u2__0root_452_0__313_));
AOI21X1 AOI21X1_2306 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5375_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15476_));
AOI21X1 AOI21X1_2307 ( .A(u2__abc_52138_new_n15477_), .B(u2__abc_52138_new_n15472_), .C(rst), .Y(u2__0root_452_0__314_));
AOI21X1 AOI21X1_2308 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n15484_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15485_));
AOI21X1 AOI21X1_2309 ( .A(u2__abc_52138_new_n15486_), .B(u2__abc_52138_new_n15479_), .C(rst), .Y(u2__0root_452_0__315_));
AOI21X1 AOI21X1_231 ( .A(u2__abc_52138_new_n6798_), .B(u2__abc_52138_new_n6792_), .C(rst), .Y(u2__0remHi_451_0__27_));
AOI21X1 AOI21X1_2310 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5401_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15493_));
AOI21X1 AOI21X1_2311 ( .A(u2__abc_52138_new_n15494_), .B(u2__abc_52138_new_n15488_), .C(rst), .Y(u2__0root_452_0__316_));
AOI21X1 AOI21X1_2312 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5389_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15501_));
AOI21X1 AOI21X1_2313 ( .A(u2__abc_52138_new_n15502_), .B(u2__abc_52138_new_n15496_), .C(rst), .Y(u2__0root_452_0__317_));
AOI21X1 AOI21X1_2314 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5394_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15508_));
AOI21X1 AOI21X1_2315 ( .A(u2__abc_52138_new_n15509_), .B(u2__abc_52138_new_n15504_), .C(rst), .Y(u2__0root_452_0__318_));
AOI21X1 AOI21X1_2316 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5341_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15516_));
AOI21X1 AOI21X1_2317 ( .A(u2__abc_52138_new_n15517_), .B(u2__abc_52138_new_n15511_), .C(rst), .Y(u2__0root_452_0__319_));
AOI21X1 AOI21X1_2318 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5348_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15524_));
AOI21X1 AOI21X1_2319 ( .A(u2__abc_52138_new_n15525_), .B(u2__abc_52138_new_n15519_), .C(rst), .Y(u2__0root_452_0__320_));
AOI21X1 AOI21X1_232 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3137_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6812_));
AOI21X1 AOI21X1_2320 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5354_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15532_));
AOI21X1 AOI21X1_2321 ( .A(u2__abc_52138_new_n15533_), .B(u2__abc_52138_new_n15527_), .C(rst), .Y(u2__0root_452_0__321_));
AOI21X1 AOI21X1_2322 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5359_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15539_));
AOI21X1 AOI21X1_2323 ( .A(u2__abc_52138_new_n15540_), .B(u2__abc_52138_new_n15535_), .C(rst), .Y(u2__0root_452_0__322_));
AOI21X1 AOI21X1_2324 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5844_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15547_));
AOI21X1 AOI21X1_2325 ( .A(u2__abc_52138_new_n15548_), .B(u2__abc_52138_new_n15542_), .C(rst), .Y(u2__0root_452_0__323_));
AOI21X1 AOI21X1_2326 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5333_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15555_));
AOI21X1 AOI21X1_2327 ( .A(u2__abc_52138_new_n15556_), .B(u2__abc_52138_new_n15550_), .C(rst), .Y(u2__0root_452_0__324_));
AOI21X1 AOI21X1_2328 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5321_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15563_));
AOI21X1 AOI21X1_2329 ( .A(u2__abc_52138_new_n15564_), .B(u2__abc_52138_new_n15558_), .C(rst), .Y(u2__0root_452_0__325_));
AOI21X1 AOI21X1_233 ( .A(u2__abc_52138_new_n6813_), .B(u2__abc_52138_new_n6800_), .C(rst), .Y(u2__0remHi_451_0__28_));
AOI21X1 AOI21X1_2330 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5326_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15570_));
AOI21X1 AOI21X1_2331 ( .A(u2__abc_52138_new_n15571_), .B(u2__abc_52138_new_n15566_), .C(rst), .Y(u2__0root_452_0__326_));
AOI21X1 AOI21X1_2332 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5274_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15578_));
AOI21X1 AOI21X1_2333 ( .A(u2__abc_52138_new_n15579_), .B(u2__abc_52138_new_n15573_), .C(rst), .Y(u2__0root_452_0__327_));
AOI21X1 AOI21X1_2334 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5281_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15586_));
AOI21X1 AOI21X1_2335 ( .A(u2__abc_52138_new_n15587_), .B(u2__abc_52138_new_n15581_), .C(rst), .Y(u2__0root_452_0__328_));
AOI21X1 AOI21X1_2336 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5287_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15594_));
AOI21X1 AOI21X1_2337 ( .A(u2__abc_52138_new_n15595_), .B(u2__abc_52138_new_n15589_), .C(rst), .Y(u2__0root_452_0__329_));
AOI21X1 AOI21X1_2338 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5292_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15601_));
AOI21X1 AOI21X1_2339 ( .A(u2__abc_52138_new_n15602_), .B(u2__abc_52138_new_n15597_), .C(rst), .Y(u2__0root_452_0__330_));
AOI21X1 AOI21X1_234 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3140_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6820_));
AOI21X1 AOI21X1_2340 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5310_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15609_));
AOI21X1 AOI21X1_2341 ( .A(u2__abc_52138_new_n15610_), .B(u2__abc_52138_new_n15604_), .C(rst), .Y(u2__0root_452_0__331_));
AOI21X1 AOI21X1_2342 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5315_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15617_));
AOI21X1 AOI21X1_2343 ( .A(u2__abc_52138_new_n15618_), .B(u2__abc_52138_new_n15612_), .C(rst), .Y(u2__0root_452_0__332_));
AOI21X1 AOI21X1_2344 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5299_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15625_));
AOI21X1 AOI21X1_2345 ( .A(u2__abc_52138_new_n15626_), .B(u2__abc_52138_new_n15620_), .C(rst), .Y(u2__0root_452_0__333_));
AOI21X1 AOI21X1_2346 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5304_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15632_));
AOI21X1 AOI21X1_2347 ( .A(u2__abc_52138_new_n15633_), .B(u2__abc_52138_new_n15628_), .C(rst), .Y(u2__0root_452_0__334_));
AOI21X1 AOI21X1_2348 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n15640_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15641_));
AOI21X1 AOI21X1_2349 ( .A(u2__abc_52138_new_n15642_), .B(u2__abc_52138_new_n15635_), .C(rst), .Y(u2__0root_452_0__335_));
AOI21X1 AOI21X1_235 ( .A(u2__abc_52138_new_n6821_), .B(u2__abc_52138_new_n6815_), .C(rst), .Y(u2__0remHi_451_0__29_));
AOI21X1 AOI21X1_2350 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5242_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15649_));
AOI21X1 AOI21X1_2351 ( .A(u2__abc_52138_new_n15650_), .B(u2__abc_52138_new_n15644_), .C(rst), .Y(u2__0root_452_0__336_));
AOI21X1 AOI21X1_2352 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5231_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15657_));
AOI21X1 AOI21X1_2353 ( .A(u2__abc_52138_new_n15658_), .B(u2__abc_52138_new_n15652_), .C(rst), .Y(u2__0root_452_0__337_));
AOI21X1 AOI21X1_2354 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5236_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15664_));
AOI21X1 AOI21X1_2355 ( .A(u2__abc_52138_new_n15665_), .B(u2__abc_52138_new_n15660_), .C(rst), .Y(u2__0root_452_0__338_));
AOI21X1 AOI21X1_2356 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n15672_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15673_));
AOI21X1 AOI21X1_2357 ( .A(u2__abc_52138_new_n15674_), .B(u2__abc_52138_new_n15667_), .C(rst), .Y(u2__0root_452_0__339_));
AOI21X1 AOI21X1_2358 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5268_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15681_));
AOI21X1 AOI21X1_2359 ( .A(u2__abc_52138_new_n15682_), .B(u2__abc_52138_new_n15676_), .C(rst), .Y(u2__0root_452_0__340_));
AOI21X1 AOI21X1_236 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3391_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6829_));
AOI21X1 AOI21X1_2360 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5249_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15689_));
AOI21X1 AOI21X1_2361 ( .A(u2__abc_52138_new_n15690_), .B(u2__abc_52138_new_n15684_), .C(rst), .Y(u2__0root_452_0__341_));
AOI21X1 AOI21X1_2362 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5256_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15696_));
AOI21X1 AOI21X1_2363 ( .A(u2__abc_52138_new_n15697_), .B(u2__abc_52138_new_n15692_), .C(rst), .Y(u2__0root_452_0__342_));
AOI21X1 AOI21X1_2364 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5197_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15704_));
AOI21X1 AOI21X1_2365 ( .A(u2__abc_52138_new_n15705_), .B(u2__abc_52138_new_n15699_), .C(rst), .Y(u2__0root_452_0__343_));
AOI21X1 AOI21X1_2366 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5202_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15712_));
AOI21X1 AOI21X1_2367 ( .A(u2__abc_52138_new_n15713_), .B(u2__abc_52138_new_n15707_), .C(rst), .Y(u2__0root_452_0__344_));
AOI21X1 AOI21X1_2368 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5183_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15720_));
AOI21X1 AOI21X1_2369 ( .A(u2__abc_52138_new_n15721_), .B(u2__abc_52138_new_n15715_), .C(rst), .Y(u2__0root_452_0__345_));
AOI21X1 AOI21X1_237 ( .A(u2__abc_52138_new_n6830_), .B(u2__abc_52138_new_n6823_), .C(rst), .Y(u2__0remHi_451_0__30_));
AOI21X1 AOI21X1_2370 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5190_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15727_));
AOI21X1 AOI21X1_2371 ( .A(u2__abc_52138_new_n15728_), .B(u2__abc_52138_new_n15723_), .C(rst), .Y(u2__0root_452_0__346_));
AOI21X1 AOI21X1_2372 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5218_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15735_));
AOI21X1 AOI21X1_2373 ( .A(u2__abc_52138_new_n15736_), .B(u2__abc_52138_new_n15730_), .C(rst), .Y(u2__0root_452_0__347_));
AOI21X1 AOI21X1_2374 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5223_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15743_));
AOI21X1 AOI21X1_2375 ( .A(u2__abc_52138_new_n15744_), .B(u2__abc_52138_new_n15738_), .C(rst), .Y(u2__0root_452_0__348_));
AOI21X1 AOI21X1_2376 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5206_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15751_));
AOI21X1 AOI21X1_2377 ( .A(u2__abc_52138_new_n15752_), .B(u2__abc_52138_new_n15746_), .C(rst), .Y(u2__0root_452_0__349_));
AOI21X1 AOI21X1_2378 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5212_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15758_));
AOI21X1 AOI21X1_2379 ( .A(u2__abc_52138_new_n15759_), .B(u2__abc_52138_new_n15754_), .C(rst), .Y(u2__0root_452_0__350_));
AOI21X1 AOI21X1_238 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3396_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6837_));
AOI21X1 AOI21X1_2380 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5147_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15766_));
AOI21X1 AOI21X1_2381 ( .A(u2__abc_52138_new_n15767_), .B(u2__abc_52138_new_n15761_), .C(rst), .Y(u2__0root_452_0__351_));
AOI21X1 AOI21X1_2382 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5152_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15774_));
AOI21X1 AOI21X1_2383 ( .A(u2__abc_52138_new_n15775_), .B(u2__abc_52138_new_n15769_), .C(rst), .Y(u2__0root_452_0__352_));
AOI21X1 AOI21X1_2384 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5136_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15782_));
AOI21X1 AOI21X1_2385 ( .A(u2__abc_52138_new_n15783_), .B(u2__abc_52138_new_n15777_), .C(rst), .Y(u2__0root_452_0__353_));
AOI21X1 AOI21X1_2386 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5141_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15789_));
AOI21X1 AOI21X1_2387 ( .A(u2__abc_52138_new_n15790_), .B(u2__abc_52138_new_n15785_), .C(rst), .Y(u2__0root_452_0__354_));
AOI21X1 AOI21X1_2388 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5170_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15797_));
AOI21X1 AOI21X1_2389 ( .A(u2__abc_52138_new_n15798_), .B(u2__abc_52138_new_n15792_), .C(rst), .Y(u2__0root_452_0__355_));
AOI21X1 AOI21X1_239 ( .A(u2__abc_52138_new_n6838_), .B(u2__abc_52138_new_n6832_), .C(rst), .Y(u2__0remHi_451_0__31_));
AOI21X1 AOI21X1_2390 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5175_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15805_));
AOI21X1 AOI21X1_2391 ( .A(u2__abc_52138_new_n15806_), .B(u2__abc_52138_new_n15800_), .C(rst), .Y(u2__0root_452_0__356_));
AOI21X1 AOI21X1_2392 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5159_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15813_));
AOI21X1 AOI21X1_2393 ( .A(u2__abc_52138_new_n15814_), .B(u2__abc_52138_new_n15808_), .C(rst), .Y(u2__0root_452_0__357_));
AOI21X1 AOI21X1_2394 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5164_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15820_));
AOI21X1 AOI21X1_2395 ( .A(u2__abc_52138_new_n15821_), .B(u2__abc_52138_new_n15816_), .C(rst), .Y(u2__0root_452_0__358_));
AOI21X1 AOI21X1_2396 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5091_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15828_));
AOI21X1 AOI21X1_2397 ( .A(u2__abc_52138_new_n15829_), .B(u2__abc_52138_new_n15823_), .C(rst), .Y(u2__0root_452_0__359_));
AOI21X1 AOI21X1_2398 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5098_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15836_));
AOI21X1 AOI21X1_2399 ( .A(u2__abc_52138_new_n15837_), .B(u2__abc_52138_new_n15831_), .C(rst), .Y(u2__0root_452_0__360_));
AOI21X1 AOI21X1_24 ( .A(u2__abc_52138_new_n3438_), .B(u2__abc_52138_new_n3384_), .C(u2__abc_52138_new_n3439_), .Y(u2__abc_52138_new_n3440_));
AOI21X1 AOI21X1_240 ( .A(u2__abc_52138_new_n6841_), .B(u2__abc_52138_new_n6824_), .C(u2__abc_52138_new_n6842_), .Y(u2__abc_52138_new_n6843_));
AOI21X1 AOI21X1_2400 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5104_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15844_));
AOI21X1 AOI21X1_2401 ( .A(u2__abc_52138_new_n15845_), .B(u2__abc_52138_new_n15839_), .C(rst), .Y(u2__0root_452_0__361_));
AOI21X1 AOI21X1_2402 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5107_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15851_));
AOI21X1 AOI21X1_2403 ( .A(u2__abc_52138_new_n15852_), .B(u2__abc_52138_new_n15847_), .C(rst), .Y(u2__0root_452_0__362_));
AOI21X1 AOI21X1_2404 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5911_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15859_));
AOI21X1 AOI21X1_2405 ( .A(u2__abc_52138_new_n15860_), .B(u2__abc_52138_new_n15854_), .C(rst), .Y(u2__0root_452_0__363_));
AOI21X1 AOI21X1_2406 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5128_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15867_));
AOI21X1 AOI21X1_2407 ( .A(u2__abc_52138_new_n15868_), .B(u2__abc_52138_new_n15862_), .C(rst), .Y(u2__0root_452_0__364_));
AOI21X1 AOI21X1_2408 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5116_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15875_));
AOI21X1 AOI21X1_2409 ( .A(u2__abc_52138_new_n15876_), .B(u2__abc_52138_new_n15870_), .C(rst), .Y(u2__0root_452_0__365_));
AOI21X1 AOI21X1_241 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n6848_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6849_));
AOI21X1 AOI21X1_2410 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5121_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15882_));
AOI21X1 AOI21X1_2411 ( .A(u2__abc_52138_new_n15883_), .B(u2__abc_52138_new_n15878_), .C(rst), .Y(u2__0root_452_0__366_));
AOI21X1 AOI21X1_2412 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5890_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15890_));
AOI21X1 AOI21X1_2413 ( .A(u2__abc_52138_new_n15891_), .B(u2__abc_52138_new_n15885_), .C(rst), .Y(u2__0root_452_0__367_));
AOI21X1 AOI21X1_2414 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5057_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15898_));
AOI21X1 AOI21X1_2415 ( .A(u2__abc_52138_new_n15899_), .B(u2__abc_52138_new_n15893_), .C(rst), .Y(u2__0root_452_0__368_));
AOI21X1 AOI21X1_2416 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5047_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15906_));
AOI21X1 AOI21X1_2417 ( .A(u2__abc_52138_new_n15907_), .B(u2__abc_52138_new_n15901_), .C(rst), .Y(u2__0root_452_0__369_));
AOI21X1 AOI21X1_2418 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n15913_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15914_));
AOI21X1 AOI21X1_2419 ( .A(u2__abc_52138_new_n15915_), .B(u2__abc_52138_new_n15909_), .C(rst), .Y(u2__0root_452_0__370_));
AOI21X1 AOI21X1_242 ( .A(u2__abc_52138_new_n6850_), .B(u2__abc_52138_new_n6840_), .C(rst), .Y(u2__0remHi_451_0__32_));
AOI21X1 AOI21X1_2420 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5082_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15922_));
AOI21X1 AOI21X1_2421 ( .A(u2__abc_52138_new_n15923_), .B(u2__abc_52138_new_n15917_), .C(rst), .Y(u2__0root_452_0__371_));
AOI21X1 AOI21X1_2422 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5076_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15930_));
AOI21X1 AOI21X1_2423 ( .A(u2__abc_52138_new_n15931_), .B(u2__abc_52138_new_n15925_), .C(rst), .Y(u2__0root_452_0__372_));
AOI21X1 AOI21X1_2424 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5067_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15938_));
AOI21X1 AOI21X1_2425 ( .A(u2__abc_52138_new_n15939_), .B(u2__abc_52138_new_n15933_), .C(rst), .Y(u2__0root_452_0__373_));
AOI21X1 AOI21X1_2426 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5072_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15945_));
AOI21X1 AOI21X1_2427 ( .A(u2__abc_52138_new_n15946_), .B(u2__abc_52138_new_n15941_), .C(rst), .Y(u2__0root_452_0__374_));
AOI21X1 AOI21X1_2428 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5018_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15953_));
AOI21X1 AOI21X1_2429 ( .A(u2__abc_52138_new_n15954_), .B(u2__abc_52138_new_n15948_), .C(rst), .Y(u2__0root_452_0__375_));
AOI21X1 AOI21X1_243 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3385_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6858_));
AOI21X1 AOI21X1_2430 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5025_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15961_));
AOI21X1 AOI21X1_2431 ( .A(u2__abc_52138_new_n15962_), .B(u2__abc_52138_new_n15956_), .C(rst), .Y(u2__0root_452_0__376_));
AOI21X1 AOI21X1_2432 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5032_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15969_));
AOI21X1 AOI21X1_2433 ( .A(u2__abc_52138_new_n15970_), .B(u2__abc_52138_new_n15964_), .C(rst), .Y(u2__0root_452_0__377_));
AOI21X1 AOI21X1_2434 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5038_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15976_));
AOI21X1 AOI21X1_2435 ( .A(u2__abc_52138_new_n15977_), .B(u2__abc_52138_new_n15972_), .C(rst), .Y(u2__0root_452_0__378_));
AOI21X1 AOI21X1_2436 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5933_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15984_));
AOI21X1 AOI21X1_2437 ( .A(u2__abc_52138_new_n15985_), .B(u2__abc_52138_new_n15979_), .C(rst), .Y(u2__0root_452_0__379_));
AOI21X1 AOI21X1_2438 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5013_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n15992_));
AOI21X1 AOI21X1_2439 ( .A(u2__abc_52138_new_n15993_), .B(u2__abc_52138_new_n15987_), .C(rst), .Y(u2__0root_452_0__380_));
AOI21X1 AOI21X1_244 ( .A(u2__abc_52138_new_n6859_), .B(u2__abc_52138_new_n6852_), .C(rst), .Y(u2__0remHi_451_0__33_));
AOI21X1 AOI21X1_2440 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5001_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16000_));
AOI21X1 AOI21X1_2441 ( .A(u2__abc_52138_new_n16001_), .B(u2__abc_52138_new_n15995_), .C(rst), .Y(u2__0root_452_0__381_));
AOI21X1 AOI21X1_2442 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5004_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16007_));
AOI21X1 AOI21X1_2443 ( .A(u2__abc_52138_new_n16008_), .B(u2__abc_52138_new_n16003_), .C(rst), .Y(u2__0root_452_0__382_));
AOI21X1 AOI21X1_2444 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6178_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16015_));
AOI21X1 AOI21X1_2445 ( .A(u2__abc_52138_new_n16016_), .B(u2__abc_52138_new_n16010_), .C(rst), .Y(u2__0root_452_0__383_));
AOI21X1 AOI21X1_2446 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6171_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16023_));
AOI21X1 AOI21X1_2447 ( .A(u2__abc_52138_new_n16024_), .B(u2__abc_52138_new_n16018_), .C(rst), .Y(u2__0root_452_0__384_));
AOI21X1 AOI21X1_2448 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6162_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16031_));
AOI21X1 AOI21X1_2449 ( .A(u2__abc_52138_new_n16032_), .B(u2__abc_52138_new_n16026_), .C(rst), .Y(u2__0root_452_0__385_));
AOI21X1 AOI21X1_245 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3443_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6868_));
AOI21X1 AOI21X1_2450 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6165_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16038_));
AOI21X1 AOI21X1_2451 ( .A(u2__abc_52138_new_n16039_), .B(u2__abc_52138_new_n16034_), .C(rst), .Y(u2__0root_452_0__386_));
AOI21X1 AOI21X1_2452 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6154_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16046_));
AOI21X1 AOI21X1_2453 ( .A(u2__abc_52138_new_n16047_), .B(u2__abc_52138_new_n16041_), .C(rst), .Y(u2__0root_452_0__387_));
AOI21X1 AOI21X1_2454 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6147_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16054_));
AOI21X1 AOI21X1_2455 ( .A(u2__abc_52138_new_n16055_), .B(u2__abc_52138_new_n16049_), .C(rst), .Y(u2__0root_452_0__388_));
AOI21X1 AOI21X1_2456 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6138_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16062_));
AOI21X1 AOI21X1_2457 ( .A(u2__abc_52138_new_n16063_), .B(u2__abc_52138_new_n16057_), .C(rst), .Y(u2__0root_452_0__389_));
AOI21X1 AOI21X1_2458 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6143_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16069_));
AOI21X1 AOI21X1_2459 ( .A(u2__abc_52138_new_n16070_), .B(u2__abc_52138_new_n16065_), .C(rst), .Y(u2__0root_452_0__390_));
AOI21X1 AOI21X1_246 ( .A(u2__abc_52138_new_n6869_), .B(u2__abc_52138_new_n6861_), .C(rst), .Y(u2__0remHi_451_0__34_));
AOI21X1 AOI21X1_2460 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n16077_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16078_));
AOI21X1 AOI21X1_2461 ( .A(u2__abc_52138_new_n16079_), .B(u2__abc_52138_new_n16072_), .C(rst), .Y(u2__0root_452_0__391_));
AOI21X1 AOI21X1_2462 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n16086_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16087_));
AOI21X1 AOI21X1_2463 ( .A(u2__abc_52138_new_n16088_), .B(u2__abc_52138_new_n16081_), .C(rst), .Y(u2__0root_452_0__392_));
AOI21X1 AOI21X1_2464 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6282_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16095_));
AOI21X1 AOI21X1_2465 ( .A(u2__abc_52138_new_n16096_), .B(u2__abc_52138_new_n16090_), .C(rst), .Y(u2__0root_452_0__393_));
AOI21X1 AOI21X1_2466 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6285_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16102_));
AOI21X1 AOI21X1_2467 ( .A(u2__abc_52138_new_n16103_), .B(u2__abc_52138_new_n16098_), .C(rst), .Y(u2__0root_452_0__394_));
AOI21X1 AOI21X1_2468 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n16110_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16111_));
AOI21X1 AOI21X1_2469 ( .A(u2__abc_52138_new_n16112_), .B(u2__abc_52138_new_n16105_), .C(rst), .Y(u2__0root_452_0__395_));
AOI21X1 AOI21X1_247 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3414_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6877_));
AOI21X1 AOI21X1_2470 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6315_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16119_));
AOI21X1 AOI21X1_2471 ( .A(u2__abc_52138_new_n16120_), .B(u2__abc_52138_new_n16114_), .C(rst), .Y(u2__0root_452_0__396_));
AOI21X1 AOI21X1_2472 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6306_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16127_));
AOI21X1 AOI21X1_2473 ( .A(u2__abc_52138_new_n16128_), .B(u2__abc_52138_new_n16122_), .C(rst), .Y(u2__0root_452_0__397_));
AOI21X1 AOI21X1_2474 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6311_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16134_));
AOI21X1 AOI21X1_2475 ( .A(u2__abc_52138_new_n16135_), .B(u2__abc_52138_new_n16130_), .C(rst), .Y(u2__0root_452_0__398_));
AOI21X1 AOI21X1_2476 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6234_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16142_));
AOI21X1 AOI21X1_2477 ( .A(u2__abc_52138_new_n16143_), .B(u2__abc_52138_new_n16137_), .C(rst), .Y(u2__0root_452_0__399_));
AOI21X1 AOI21X1_2478 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6237_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16150_));
AOI21X1 AOI21X1_2479 ( .A(u2__abc_52138_new_n16151_), .B(u2__abc_52138_new_n16145_), .C(rst), .Y(u2__0root_452_0__400_));
AOI21X1 AOI21X1_248 ( .A(u2__abc_52138_new_n6878_), .B(u2__abc_52138_new_n6871_), .C(rst), .Y(u2__0remHi_451_0__35_));
AOI21X1 AOI21X1_2480 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6245_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16158_));
AOI21X1 AOI21X1_2481 ( .A(u2__abc_52138_new_n16159_), .B(u2__abc_52138_new_n16153_), .C(rst), .Y(u2__0root_452_0__401_));
AOI21X1 AOI21X1_2482 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6248_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16165_));
AOI21X1 AOI21X1_2483 ( .A(u2__abc_52138_new_n16166_), .B(u2__abc_52138_new_n16161_), .C(rst), .Y(u2__0root_452_0__402_));
AOI21X1 AOI21X1_2484 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6273_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16173_));
AOI21X1 AOI21X1_2485 ( .A(u2__abc_52138_new_n16174_), .B(u2__abc_52138_new_n16168_), .C(rst), .Y(u2__0root_452_0__403_));
AOI21X1 AOI21X1_2486 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6266_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16181_));
AOI21X1 AOI21X1_2487 ( .A(u2__abc_52138_new_n16182_), .B(u2__abc_52138_new_n16176_), .C(rst), .Y(u2__0root_452_0__404_));
AOI21X1 AOI21X1_2488 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6257_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16189_));
AOI21X1 AOI21X1_2489 ( .A(u2__abc_52138_new_n16190_), .B(u2__abc_52138_new_n16184_), .C(rst), .Y(u2__0root_452_0__405_));
AOI21X1 AOI21X1_249 ( .A(u2__abc_52138_new_n6881_), .B(u2__abc_52138_new_n3388_), .C(u2__abc_52138_new_n6883_), .Y(u2__abc_52138_new_n6884_));
AOI21X1 AOI21X1_2490 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6262_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16196_));
AOI21X1 AOI21X1_2491 ( .A(u2__abc_52138_new_n16197_), .B(u2__abc_52138_new_n16192_), .C(rst), .Y(u2__0root_452_0__406_));
AOI21X1 AOI21X1_2492 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6203_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16204_));
AOI21X1 AOI21X1_2493 ( .A(u2__abc_52138_new_n16205_), .B(u2__abc_52138_new_n16199_), .C(rst), .Y(u2__0root_452_0__407_));
AOI21X1 AOI21X1_2494 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6196_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16212_));
AOI21X1 AOI21X1_2495 ( .A(u2__abc_52138_new_n16213_), .B(u2__abc_52138_new_n16207_), .C(rst), .Y(u2__0root_452_0__408_));
AOI21X1 AOI21X1_2496 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6187_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16220_));
AOI21X1 AOI21X1_2497 ( .A(u2__abc_52138_new_n16221_), .B(u2__abc_52138_new_n16215_), .C(rst), .Y(u2__0root_452_0__409_));
AOI21X1 AOI21X1_2498 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6190_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16227_));
AOI21X1 AOI21X1_2499 ( .A(u2__abc_52138_new_n16228_), .B(u2__abc_52138_new_n16223_), .C(rst), .Y(u2__0root_452_0__410_));
AOI21X1 AOI21X1_25 ( .A(u2__abc_52138_new_n3445_), .B(u2__abc_52138_new_n3413_), .C(u2__abc_52138_new_n3442_), .Y(u2__abc_52138_new_n3446_));
AOI21X1 AOI21X1_250 ( .A(u2__abc_52138_new_n6890_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6891_));
AOI21X1 AOI21X1_2500 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6226_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16235_));
AOI21X1 AOI21X1_2501 ( .A(u2__abc_52138_new_n16236_), .B(u2__abc_52138_new_n16230_), .C(rst), .Y(u2__0root_452_0__411_));
AOI21X1 AOI21X1_2502 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6219_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16243_));
AOI21X1 AOI21X1_2503 ( .A(u2__abc_52138_new_n16244_), .B(u2__abc_52138_new_n16238_), .C(rst), .Y(u2__0root_452_0__412_));
AOI21X1 AOI21X1_2504 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6210_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16251_));
AOI21X1 AOI21X1_2505 ( .A(u2__abc_52138_new_n16252_), .B(u2__abc_52138_new_n16246_), .C(rst), .Y(u2__0root_452_0__413_));
AOI21X1 AOI21X1_2506 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6215_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16258_));
AOI21X1 AOI21X1_2507 ( .A(u2__abc_52138_new_n16259_), .B(u2__abc_52138_new_n16254_), .C(rst), .Y(u2__0root_452_0__414_));
AOI21X1 AOI21X1_2508 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6127_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16266_));
AOI21X1 AOI21X1_2509 ( .A(u2__abc_52138_new_n16267_), .B(u2__abc_52138_new_n16261_), .C(rst), .Y(u2__0root_452_0__415_));
AOI21X1 AOI21X1_251 ( .A(u2__abc_52138_new_n6892_), .B(u2__abc_52138_new_n6880_), .C(rst), .Y(u2__0remHi_451_0__36_));
AOI21X1 AOI21X1_2510 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6120_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16274_));
AOI21X1 AOI21X1_2511 ( .A(u2__abc_52138_new_n16275_), .B(u2__abc_52138_new_n16269_), .C(rst), .Y(u2__0root_452_0__416_));
AOI21X1 AOI21X1_2512 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6108_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16282_));
AOI21X1 AOI21X1_2513 ( .A(u2__abc_52138_new_n16283_), .B(u2__abc_52138_new_n16277_), .C(rst), .Y(u2__0root_452_0__417_));
AOI21X1 AOI21X1_2514 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6115_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16289_));
AOI21X1 AOI21X1_2515 ( .A(u2__abc_52138_new_n16290_), .B(u2__abc_52138_new_n16285_), .C(rst), .Y(u2__0root_452_0__418_));
AOI21X1 AOI21X1_2516 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6103_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16297_));
AOI21X1 AOI21X1_2517 ( .A(u2__abc_52138_new_n16298_), .B(u2__abc_52138_new_n16292_), .C(rst), .Y(u2__0root_452_0__419_));
AOI21X1 AOI21X1_2518 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6096_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16305_));
AOI21X1 AOI21X1_2519 ( .A(u2__abc_52138_new_n16306_), .B(u2__abc_52138_new_n16300_), .C(rst), .Y(u2__0root_452_0__420_));
AOI21X1 AOI21X1_252 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3408_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6900_));
AOI21X1 AOI21X1_2520 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6084_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16313_));
AOI21X1 AOI21X1_2521 ( .A(u2__abc_52138_new_n16314_), .B(u2__abc_52138_new_n16308_), .C(rst), .Y(u2__0root_452_0__421_));
AOI21X1 AOI21X1_2522 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6089_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16320_));
AOI21X1 AOI21X1_2523 ( .A(u2__abc_52138_new_n16321_), .B(u2__abc_52138_new_n16316_), .C(rst), .Y(u2__0root_452_0__422_));
AOI21X1 AOI21X1_2524 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6049_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16328_));
AOI21X1 AOI21X1_2525 ( .A(u2__abc_52138_new_n16329_), .B(u2__abc_52138_new_n16323_), .C(rst), .Y(u2__0root_452_0__423_));
AOI21X1 AOI21X1_2526 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6052_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16336_));
AOI21X1 AOI21X1_2527 ( .A(u2__abc_52138_new_n16337_), .B(u2__abc_52138_new_n16331_), .C(rst), .Y(u2__0root_452_0__424_));
AOI21X1 AOI21X1_2528 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6036_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16344_));
AOI21X1 AOI21X1_2529 ( .A(u2__abc_52138_new_n16345_), .B(u2__abc_52138_new_n16339_), .C(rst), .Y(u2__0root_452_0__425_));
AOI21X1 AOI21X1_253 ( .A(u2__abc_52138_new_n6901_), .B(u2__abc_52138_new_n6894_), .C(rst), .Y(u2__0remHi_451_0__37_));
AOI21X1 AOI21X1_2530 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6043_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16351_));
AOI21X1 AOI21X1_2531 ( .A(u2__abc_52138_new_n16352_), .B(u2__abc_52138_new_n16347_), .C(rst), .Y(u2__0root_452_0__426_));
AOI21X1 AOI21X1_2532 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6077_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16359_));
AOI21X1 AOI21X1_2533 ( .A(u2__abc_52138_new_n16360_), .B(u2__abc_52138_new_n16354_), .C(rst), .Y(u2__0root_452_0__427_));
AOI21X1 AOI21X1_2534 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6070_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16367_));
AOI21X1 AOI21X1_2535 ( .A(u2__abc_52138_new_n16368_), .B(u2__abc_52138_new_n16362_), .C(rst), .Y(u2__0root_452_0__428_));
AOI21X1 AOI21X1_2536 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6058_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16375_));
AOI21X1 AOI21X1_2537 ( .A(u2__abc_52138_new_n16376_), .B(u2__abc_52138_new_n16370_), .C(rst), .Y(u2__0root_452_0__429_));
AOI21X1 AOI21X1_2538 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6063_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16382_));
AOI21X1 AOI21X1_2539 ( .A(u2__abc_52138_new_n16383_), .B(u2__abc_52138_new_n16378_), .C(rst), .Y(u2__0root_452_0__430_));
AOI21X1 AOI21X1_254 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3348_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6911_));
AOI21X1 AOI21X1_2540 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6012_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16390_));
AOI21X1 AOI21X1_2541 ( .A(u2__abc_52138_new_n16391_), .B(u2__abc_52138_new_n16385_), .C(rst), .Y(u2__0root_452_0__431_));
AOI21X1 AOI21X1_2542 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6015_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16398_));
AOI21X1 AOI21X1_2543 ( .A(u2__abc_52138_new_n16399_), .B(u2__abc_52138_new_n16393_), .C(rst), .Y(u2__0root_452_0__432_));
AOI21X1 AOI21X1_2544 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6023_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16406_));
AOI21X1 AOI21X1_2545 ( .A(u2__abc_52138_new_n16407_), .B(u2__abc_52138_new_n16401_), .C(rst), .Y(u2__0root_452_0__433_));
AOI21X1 AOI21X1_2546 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6026_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16413_));
AOI21X1 AOI21X1_2547 ( .A(u2__abc_52138_new_n16414_), .B(u2__abc_52138_new_n16409_), .C(rst), .Y(u2__0root_452_0__434_));
AOI21X1 AOI21X1_2548 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6005_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16421_));
AOI21X1 AOI21X1_2549 ( .A(u2__abc_52138_new_n16422_), .B(u2__abc_52138_new_n16416_), .C(rst), .Y(u2__0root_452_0__435_));
AOI21X1 AOI21X1_255 ( .A(u2__abc_52138_new_n6912_), .B(u2__abc_52138_new_n6903_), .C(rst), .Y(u2__0remHi_451_0__38_));
AOI21X1 AOI21X1_2550 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5998_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16429_));
AOI21X1 AOI21X1_2551 ( .A(u2__abc_52138_new_n16430_), .B(u2__abc_52138_new_n16424_), .C(rst), .Y(u2__0root_452_0__436_));
AOI21X1 AOI21X1_2552 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5989_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16437_));
AOI21X1 AOI21X1_2553 ( .A(u2__abc_52138_new_n16438_), .B(u2__abc_52138_new_n16432_), .C(rst), .Y(u2__0root_452_0__437_));
AOI21X1 AOI21X1_2554 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5994_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16444_));
AOI21X1 AOI21X1_2555 ( .A(u2__abc_52138_new_n16445_), .B(u2__abc_52138_new_n16440_), .C(rst), .Y(u2__0root_452_0__438_));
AOI21X1 AOI21X1_2556 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5969_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16452_));
AOI21X1 AOI21X1_2557 ( .A(u2__abc_52138_new_n16453_), .B(u2__abc_52138_new_n16447_), .C(rst), .Y(u2__0root_452_0__439_));
AOI21X1 AOI21X1_2558 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6414_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16460_));
AOI21X1 AOI21X1_2559 ( .A(u2__abc_52138_new_n16461_), .B(u2__abc_52138_new_n16455_), .C(rst), .Y(u2__0root_452_0__440_));
AOI21X1 AOI21X1_256 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3353_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6919_));
AOI21X1 AOI21X1_2560 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5976_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16468_));
AOI21X1 AOI21X1_2561 ( .A(u2__abc_52138_new_n16469_), .B(u2__abc_52138_new_n16463_), .C(rst), .Y(u2__0root_452_0__441_));
AOI21X1 AOI21X1_2562 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5979_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16475_));
AOI21X1 AOI21X1_2563 ( .A(u2__abc_52138_new_n16476_), .B(u2__abc_52138_new_n16471_), .C(rst), .Y(u2__0root_452_0__442_));
AOI21X1 AOI21X1_2564 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5962_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16483_));
AOI21X1 AOI21X1_2565 ( .A(u2__abc_52138_new_n16484_), .B(u2__abc_52138_new_n16478_), .C(rst), .Y(u2__0root_452_0__443_));
AOI21X1 AOI21X1_2566 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5955_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16491_));
AOI21X1 AOI21X1_2567 ( .A(u2__abc_52138_new_n16492_), .B(u2__abc_52138_new_n16486_), .C(rst), .Y(u2__0root_452_0__444_));
AOI21X1 AOI21X1_2568 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5946_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16499_));
AOI21X1 AOI21X1_2569 ( .A(u2__abc_52138_new_n16500_), .B(u2__abc_52138_new_n16494_), .C(rst), .Y(u2__0root_452_0__445_));
AOI21X1 AOI21X1_257 ( .A(u2__abc_52138_new_n6920_), .B(u2__abc_52138_new_n6914_), .C(rst), .Y(u2__0remHi_451_0__39_));
AOI21X1 AOI21X1_2570 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5949_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16506_));
AOI21X1 AOI21X1_2571 ( .A(u2__abc_52138_new_n16507_), .B(u2__abc_52138_new_n16502_), .C(rst), .Y(u2__0root_452_0__446_));
AOI21X1 AOI21X1_2572 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3010_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16514_));
AOI21X1 AOI21X1_2573 ( .A(u2__abc_52138_new_n16515_), .B(u2__abc_52138_new_n16509_), .C(rst), .Y(u2__0root_452_0__447_));
AOI21X1 AOI21X1_2574 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3005_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16522_));
AOI21X1 AOI21X1_2575 ( .A(u2__abc_52138_new_n16523_), .B(u2__abc_52138_new_n16517_), .C(rst), .Y(u2__0root_452_0__448_));
AOI21X1 AOI21X1_2576 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n2997_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16530_));
AOI21X1 AOI21X1_2577 ( .A(u2__abc_52138_new_n16531_), .B(u2__abc_52138_new_n16525_), .C(rst), .Y(u2__0root_452_0__449_));
AOI21X1 AOI21X1_2578 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6446_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n16537_));
AOI21X1 AOI21X1_2579 ( .A(u2__abc_52138_new_n16538_), .B(u2__abc_52138_new_n16533_), .C(rst), .Y(u2__0root_452_0__450_));
AOI21X1 AOI21X1_258 ( .A(u2__abc_52138_new_n6934_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6935_));
AOI21X1 AOI21X1_259 ( .A(u2__abc_52138_new_n6936_), .B(u2__abc_52138_new_n6922_), .C(rst), .Y(u2__0remHi_451_0__40_));
AOI21X1 AOI21X1_26 ( .A(u2__abc_52138_new_n3447_), .B(u2__abc_52138_new_n3407_), .C(u2__abc_52138_new_n3448_), .Y(u2__abc_52138_new_n3449_));
AOI21X1 AOI21X1_260 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3342_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6943_));
AOI21X1 AOI21X1_261 ( .A(u2__abc_52138_new_n6944_), .B(u2__abc_52138_new_n6938_), .C(rst), .Y(u2__0remHi_451_0__41_));
AOI21X1 AOI21X1_262 ( .A(u2__abc_52138_new_n6939_), .B(u2__abc_52138_new_n3354_), .C(u2__abc_52138_new_n6947_), .Y(u2__abc_52138_new_n6948_));
AOI21X1 AOI21X1_263 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3376_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6952_));
AOI21X1 AOI21X1_264 ( .A(u2__abc_52138_new_n6953_), .B(u2__abc_52138_new_n6946_), .C(rst), .Y(u2__0remHi_451_0__42_));
AOI21X1 AOI21X1_265 ( .A(u2__abc_52138_new_n6957_), .B(u2__abc_52138_new_n6958_), .C(u2__abc_52138_new_n6959_), .Y(u2__abc_52138_new_n6960_));
AOI21X1 AOI21X1_266 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3371_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6962_));
AOI21X1 AOI21X1_267 ( .A(u2__abc_52138_new_n6963_), .B(u2__abc_52138_new_n6955_), .C(rst), .Y(u2__0remHi_451_0__43_));
AOI21X1 AOI21X1_268 ( .A(u2__abc_52138_new_n6929_), .B(u2__abc_52138_new_n3425_), .C(u2__abc_52138_new_n6970_), .Y(u2__abc_52138_new_n6971_));
AOI21X1 AOI21X1_269 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3360_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6976_));
AOI21X1 AOI21X1_27 ( .A(u2__abc_52138_new_n3441_), .B(u2__abc_52138_new_n3431_), .C(u2__abc_52138_new_n3450_), .Y(u2__abc_52138_new_n3451_));
AOI21X1 AOI21X1_270 ( .A(u2__abc_52138_new_n6977_), .B(u2__abc_52138_new_n6965_), .C(rst), .Y(u2__0remHi_451_0__44_));
AOI21X1 AOI21X1_271 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3365_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6984_));
AOI21X1 AOI21X1_272 ( .A(u2__abc_52138_new_n6985_), .B(u2__abc_52138_new_n6979_), .C(rst), .Y(u2__0remHi_451_0__45_));
AOI21X1 AOI21X1_273 ( .A(u2__abc_52138_new_n6973_), .B(u2__abc_52138_new_n6989_), .C(u2__abc_52138_new_n6988_), .Y(u2__abc_52138_new_n6990_));
AOI21X1 AOI21X1_274 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3305_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n6994_));
AOI21X1 AOI21X1_275 ( .A(u2__abc_52138_new_n6995_), .B(u2__abc_52138_new_n6987_), .C(rst), .Y(u2__0remHi_451_0__46_));
AOI21X1 AOI21X1_276 ( .A(u2__abc_52138_new_n6990_), .B(u2__abc_52138_new_n3361_), .C(u2__abc_52138_new_n6998_), .Y(u2__abc_52138_new_n6999_));
AOI21X1 AOI21X1_277 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3298_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7003_));
AOI21X1 AOI21X1_278 ( .A(u2__abc_52138_new_n7004_), .B(u2__abc_52138_new_n6997_), .C(rst), .Y(u2__0remHi_451_0__47_));
AOI21X1 AOI21X1_279 ( .A(u2__abc_52138_new_n6970_), .B(u2__abc_52138_new_n3426_), .C(u2__abc_52138_new_n7008_), .Y(u2__abc_52138_new_n7009_));
AOI21X1 AOI21X1_28 ( .A(u2__abc_52138_new_n3453_), .B(u2__abc_52138_new_n3352_), .C(u2__abc_52138_new_n3454_), .Y(u2__abc_52138_new_n3455_));
AOI21X1 AOI21X1_280 ( .A(u2__abc_52138_new_n3368_), .B(u2__abc_52138_new_n7007_), .C(u2__abc_52138_new_n7010_), .Y(u2__abc_52138_new_n7011_));
AOI21X1 AOI21X1_281 ( .A(u2__abc_52138_new_n7017_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7018_));
AOI21X1 AOI21X1_282 ( .A(u2__abc_52138_new_n7019_), .B(u2__abc_52138_new_n7006_), .C(rst), .Y(u2__0remHi_451_0__48_));
AOI21X1 AOI21X1_283 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3292_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7026_));
AOI21X1 AOI21X1_284 ( .A(u2__abc_52138_new_n7027_), .B(u2__abc_52138_new_n7021_), .C(rst), .Y(u2__0remHi_451_0__49_));
AOI21X1 AOI21X1_285 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3329_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7039_));
AOI21X1 AOI21X1_286 ( .A(u2__abc_52138_new_n7040_), .B(u2__abc_52138_new_n7029_), .C(rst), .Y(u2__0remHi_451_0__50_));
AOI21X1 AOI21X1_287 ( .A(u2__abc_52138_new_n3296_), .B(u2__abc_52138_new_n7043_), .C(u2__abc_52138_new_n7044_), .Y(u2__abc_52138_new_n7045_));
AOI21X1 AOI21X1_288 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3324_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7047_));
AOI21X1 AOI21X1_289 ( .A(u2__abc_52138_new_n7048_), .B(u2__abc_52138_new_n7042_), .C(rst), .Y(u2__0remHi_451_0__51_));
AOI21X1 AOI21X1_29 ( .A(u2__abc_52138_new_n3459_), .B(u2__abc_52138_new_n3426_), .C(u2__abc_52138_new_n3466_), .Y(u2__abc_52138_new_n3467_));
AOI21X1 AOI21X1_290 ( .A(u2__abc_52138_new_n7012_), .B(u2__abc_52138_new_n3310_), .C(u2__abc_52138_new_n7055_), .Y(u2__abc_52138_new_n7056_));
AOI21X1 AOI21X1_291 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3313_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7061_));
AOI21X1 AOI21X1_292 ( .A(u2__abc_52138_new_n7062_), .B(u2__abc_52138_new_n7050_), .C(rst), .Y(u2__0remHi_451_0__52_));
AOI21X1 AOI21X1_293 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3318_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7069_));
AOI21X1 AOI21X1_294 ( .A(u2__abc_52138_new_n7070_), .B(u2__abc_52138_new_n7064_), .C(rst), .Y(u2__0remHi_451_0__53_));
AOI21X1 AOI21X1_295 ( .A(u2__abc_52138_new_n7058_), .B(u2__abc_52138_new_n7075_), .C(u2__abc_52138_new_n7073_), .Y(u2__abc_52138_new_n7076_));
AOI21X1 AOI21X1_296 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3253_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7080_));
AOI21X1 AOI21X1_297 ( .A(u2__abc_52138_new_n7081_), .B(u2__abc_52138_new_n7072_), .C(rst), .Y(u2__0remHi_451_0__54_));
AOI21X1 AOI21X1_298 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3258_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7089_));
AOI21X1 AOI21X1_299 ( .A(u2__abc_52138_new_n7090_), .B(u2__abc_52138_new_n7083_), .C(rst), .Y(u2__0remHi_451_0__55_));
AOI21X1 AOI21X1_3 ( .A(_abc_65734_new_n1492_), .B(_abc_65734_new_n1494_), .C(_abc_65734_new_n1483_), .Y(_abc_65734_new_n1495_));
AOI21X1 AOI21X1_30 ( .A(u2__abc_52138_new_n3469_), .B(u2__abc_52138_new_n3470_), .C(u2__abc_52138_new_n3301_), .Y(u2__abc_52138_new_n3471_));
AOI21X1 AOI21X1_300 ( .A(u2__abc_52138_new_n3321_), .B(u2__abc_52138_new_n7095_), .C(u2__abc_52138_new_n7096_), .Y(u2__abc_52138_new_n7097_));
AOI21X1 AOI21X1_301 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3242_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7105_));
AOI21X1 AOI21X1_302 ( .A(u2__abc_52138_new_n7106_), .B(u2__abc_52138_new_n7092_), .C(rst), .Y(u2__0remHi_451_0__56_));
AOI21X1 AOI21X1_303 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3247_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7113_));
AOI21X1 AOI21X1_304 ( .A(u2__abc_52138_new_n7114_), .B(u2__abc_52138_new_n7108_), .C(rst), .Y(u2__0remHi_451_0__57_));
AOI21X1 AOI21X1_305 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3281_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7122_));
AOI21X1 AOI21X1_306 ( .A(u2__abc_52138_new_n7123_), .B(u2__abc_52138_new_n7116_), .C(rst), .Y(u2__0remHi_451_0__58_));
AOI21X1 AOI21X1_307 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3276_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7131_));
AOI21X1 AOI21X1_308 ( .A(u2__abc_52138_new_n7132_), .B(u2__abc_52138_new_n7125_), .C(rst), .Y(u2__0remHi_451_0__59_));
AOI21X1 AOI21X1_309 ( .A(u2__abc_52138_new_n7136_), .B(u2__abc_52138_new_n3250_), .C(u2__abc_52138_new_n7137_), .Y(u2__abc_52138_new_n7138_));
AOI21X1 AOI21X1_31 ( .A(u2__abc_52138_new_n3481_), .B(u2__abc_52138_new_n3317_), .C(u2__abc_52138_new_n3482_), .Y(u2__abc_52138_new_n3483_));
AOI21X1 AOI21X1_310 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3265_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7146_));
AOI21X1 AOI21X1_311 ( .A(u2__abc_52138_new_n7147_), .B(u2__abc_52138_new_n7134_), .C(rst), .Y(u2__0remHi_451_0__60_));
AOI21X1 AOI21X1_312 ( .A(u2__abc_52138_new_n3275_), .B(u2__abc_52138_new_n3277_), .C(u2__abc_52138_new_n7150_), .Y(u2__abc_52138_new_n7151_));
AOI21X1 AOI21X1_313 ( .A(u2__abc_52138_new_n7140_), .B(u2__abc_52138_new_n3280_), .C(u2__abc_52138_new_n3278_), .Y(u2__abc_52138_new_n7152_));
AOI21X1 AOI21X1_314 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3268_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7156_));
AOI21X1 AOI21X1_315 ( .A(u2__abc_52138_new_n7157_), .B(u2__abc_52138_new_n7149_), .C(rst), .Y(u2__0remHi_451_0__61_));
AOI21X1 AOI21X1_316 ( .A(u2__abc_52138_new_n7160_), .B(u2__abc_52138_new_n3267_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n7162_));
AOI21X1 AOI21X1_317 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3834_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7165_));
AOI21X1 AOI21X1_318 ( .A(u2__abc_52138_new_n7166_), .B(u2__abc_52138_new_n7159_), .C(rst), .Y(u2__0remHi_451_0__62_));
AOI21X1 AOI21X1_319 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3839_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7173_));
AOI21X1 AOI21X1_32 ( .A(u2__abc_52138_new_n3476_), .B(u2__abc_52138_new_n3333_), .C(u2__abc_52138_new_n3484_), .Y(u2__abc_52138_new_n3485_));
AOI21X1 AOI21X1_320 ( .A(u2__abc_52138_new_n7174_), .B(u2__abc_52138_new_n7168_), .C(rst), .Y(u2__0remHi_451_0__63_));
AOI21X1 AOI21X1_321 ( .A(u2__abc_52138_new_n7178_), .B(u2__abc_52138_new_n3273_), .C(u2__abc_52138_new_n7179_), .Y(u2__abc_52138_new_n7180_));
AOI21X1 AOI21X1_322 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3845_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7191_));
AOI21X1 AOI21X1_323 ( .A(u2__abc_52138_new_n7192_), .B(u2__abc_52138_new_n7176_), .C(rst), .Y(u2__0remHi_451_0__64_));
AOI21X1 AOI21X1_324 ( .A(u2__abc_52138_new_n3841_), .B(u2__abc_52138_new_n7195_), .C(u2__abc_52138_new_n7196_), .Y(u2__abc_52138_new_n7197_));
AOI21X1 AOI21X1_325 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3850_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7199_));
AOI21X1 AOI21X1_326 ( .A(u2__abc_52138_new_n7200_), .B(u2__abc_52138_new_n7194_), .C(rst), .Y(u2__0remHi_451_0__65_));
AOI21X1 AOI21X1_327 ( .A(u2__abc_52138_new_n7185_), .B(u2__abc_52138_new_n3842_), .C(u2__abc_52138_new_n7203_), .Y(u2__abc_52138_new_n7204_));
AOI21X1 AOI21X1_328 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3864_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7208_));
AOI21X1 AOI21X1_329 ( .A(u2__abc_52138_new_n7209_), .B(u2__abc_52138_new_n7202_), .C(rst), .Y(u2__0remHi_451_0__66_));
AOI21X1 AOI21X1_33 ( .A(u2__abc_52138_new_n3488_), .B(u2__abc_52138_new_n3257_), .C(u2__abc_52138_new_n3489_), .Y(u2__abc_52138_new_n3490_));
AOI21X1 AOI21X1_330 ( .A(u2__abc_52138_new_n7213_), .B(u2__abc_52138_new_n7214_), .C(u2__abc_52138_new_n7215_), .Y(u2__abc_52138_new_n7216_));
AOI21X1 AOI21X1_331 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3883_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7218_));
AOI21X1 AOI21X1_332 ( .A(u2__abc_52138_new_n7219_), .B(u2__abc_52138_new_n7211_), .C(rst), .Y(u2__0remHi_451_0__67_));
AOI21X1 AOI21X1_333 ( .A(u2__abc_52138_new_n7224_), .B(u2__abc_52138_new_n3851_), .C(u2__abc_52138_new_n7212_), .Y(u2__abc_52138_new_n7225_));
AOI21X1 AOI21X1_334 ( .A(u2__abc_52138_new_n7185_), .B(u2__abc_52138_new_n3854_), .C(u2__abc_52138_new_n7226_), .Y(u2__abc_52138_new_n7227_));
AOI21X1 AOI21X1_335 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3888_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7231_));
AOI21X1 AOI21X1_336 ( .A(u2__abc_52138_new_n7232_), .B(u2__abc_52138_new_n7221_), .C(rst), .Y(u2__0remHi_451_0__68_));
AOI21X1 AOI21X1_337 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3858_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7239_));
AOI21X1 AOI21X1_338 ( .A(u2__abc_52138_new_n7240_), .B(u2__abc_52138_new_n7234_), .C(rst), .Y(u2__0remHi_451_0__69_));
AOI21X1 AOI21X1_339 ( .A(u2__abc_52138_new_n3855_), .B(u2__abc_52138_new_n7244_), .C(u2__abc_52138_new_n7245_), .Y(u2__abc_52138_new_n7246_));
AOI21X1 AOI21X1_34 ( .A(u2__abc_52138_new_n3493_), .B(u2__abc_52138_new_n3486_), .C(u2__abc_52138_new_n3498_), .Y(u2__abc_52138_new_n3499_));
AOI21X1 AOI21X1_340 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3786_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7248_));
AOI21X1 AOI21X1_341 ( .A(u2__abc_52138_new_n7249_), .B(u2__abc_52138_new_n7242_), .C(rst), .Y(u2__0remHi_451_0__70_));
AOI21X1 AOI21X1_342 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3791_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7258_));
AOI21X1 AOI21X1_343 ( .A(u2__abc_52138_new_n7259_), .B(u2__abc_52138_new_n7251_), .C(rst), .Y(u2__0remHi_451_0__71_));
AOI21X1 AOI21X1_344 ( .A(u2__abc_52138_new_n7226_), .B(u2__abc_52138_new_n3867_), .C(u2__abc_52138_new_n7266_), .Y(u2__abc_52138_new_n7267_));
AOI21X1 AOI21X1_345 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3799_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7276_));
AOI21X1 AOI21X1_346 ( .A(u2__abc_52138_new_n7277_), .B(u2__abc_52138_new_n7261_), .C(rst), .Y(u2__0remHi_451_0__72_));
AOI21X1 AOI21X1_347 ( .A(u2__abc_52138_new_n3795_), .B(u2__abc_52138_new_n7280_), .C(u2__abc_52138_new_n7281_), .Y(u2__abc_52138_new_n7282_));
AOI21X1 AOI21X1_348 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3804_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7284_));
AOI21X1 AOI21X1_349 ( .A(u2__abc_52138_new_n7285_), .B(u2__abc_52138_new_n7279_), .C(rst), .Y(u2__0remHi_451_0__73_));
AOI21X1 AOI21X1_35 ( .A(u2__abc_52138_new_n3468_), .B(u2__abc_52138_new_n3424_), .C(u2__abc_52138_new_n3500_), .Y(u2__abc_52138_new_n3501_));
AOI21X1 AOI21X1_350 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3824_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7294_));
AOI21X1 AOI21X1_351 ( .A(u2__abc_52138_new_n7295_), .B(u2__abc_52138_new_n7287_), .C(rst), .Y(u2__0remHi_451_0__74_));
AOI21X1 AOI21X1_352 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3819_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7304_));
AOI21X1 AOI21X1_353 ( .A(u2__abc_52138_new_n7305_), .B(u2__abc_52138_new_n7297_), .C(rst), .Y(u2__0remHi_451_0__75_));
AOI21X1 AOI21X1_354 ( .A(u2__abc_52138_new_n7311_), .B(u2__abc_52138_new_n7309_), .C(u2__abc_52138_new_n7312_), .Y(u2__abc_52138_new_n7313_));
AOI21X1 AOI21X1_355 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3808_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7321_));
AOI21X1 AOI21X1_356 ( .A(u2__abc_52138_new_n7322_), .B(u2__abc_52138_new_n7307_), .C(rst), .Y(u2__0remHi_451_0__76_));
AOI21X1 AOI21X1_357 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3813_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7331_));
AOI21X1 AOI21X1_358 ( .A(u2__abc_52138_new_n7332_), .B(u2__abc_52138_new_n7324_), .C(rst), .Y(u2__0remHi_451_0__77_));
AOI21X1 AOI21X1_359 ( .A(u2__abc_52138_new_n7337_), .B(u2__abc_52138_new_n7335_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n7338_));
AOI21X1 AOI21X1_36 ( .A(u2__abc_52138_new_n3874_), .B(u2__abc_52138_new_n3838_), .C(u2__abc_52138_new_n3875_), .Y(u2__abc_52138_new_n3876_));
AOI21X1 AOI21X1_360 ( .A(u2__abc_52138_new_n3808_), .B(u2__abc_52138_new_n6498_), .C(u2__abc_52138_new_n7338_), .Y(u2__abc_52138_new_n7339_));
AOI21X1 AOI21X1_361 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3740_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7340_));
AOI21X1 AOI21X1_362 ( .A(u2__abc_52138_new_n7341_), .B(u2__abc_52138_new_n7334_), .C(rst), .Y(u2__0remHi_451_0__78_));
AOI21X1 AOI21X1_363 ( .A(u2__abc_52138_new_n3817_), .B(u2__abc_52138_new_n7344_), .C(u2__abc_52138_new_n7345_), .Y(u2__abc_52138_new_n7346_));
AOI21X1 AOI21X1_364 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3745_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7348_));
AOI21X1 AOI21X1_365 ( .A(u2__abc_52138_new_n7349_), .B(u2__abc_52138_new_n7343_), .C(rst), .Y(u2__0remHi_451_0__79_));
AOI21X1 AOI21X1_366 ( .A(u2__abc_52138_new_n7357_), .B(u2__abc_52138_new_n3825_), .C(u2__abc_52138_new_n3820_), .Y(u2__abc_52138_new_n7358_));
AOI21X1 AOI21X1_367 ( .A(u2__abc_52138_new_n3809_), .B(u2__abc_52138_new_n7352_), .C(u2__abc_52138_new_n3814_), .Y(u2__abc_52138_new_n7359_));
AOI21X1 AOI21X1_368 ( .A(u2__abc_52138_new_n7185_), .B(u2__abc_52138_new_n3869_), .C(u2__abc_52138_new_n7362_), .Y(u2__abc_52138_new_n7363_));
AOI21X1 AOI21X1_369 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3751_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7367_));
AOI21X1 AOI21X1_37 ( .A(u2__abc_52138_new_n3877_), .B(u2__abc_52138_new_n3849_), .C(u2__abc_52138_new_n3878_), .Y(u2__abc_52138_new_n3879_));
AOI21X1 AOI21X1_370 ( .A(u2__abc_52138_new_n7368_), .B(u2__abc_52138_new_n7351_), .C(rst), .Y(u2__0remHi_451_0__80_));
AOI21X1 AOI21X1_371 ( .A(u2__abc_52138_new_n7371_), .B(u2__abc_52138_new_n7372_), .C(u2__abc_52138_new_n7373_), .Y(u2__abc_52138_new_n7374_));
AOI21X1 AOI21X1_372 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3756_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7376_));
AOI21X1 AOI21X1_373 ( .A(u2__abc_52138_new_n7377_), .B(u2__abc_52138_new_n7370_), .C(rst), .Y(u2__0remHi_451_0__81_));
AOI21X1 AOI21X1_374 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3779_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7386_));
AOI21X1 AOI21X1_375 ( .A(u2__abc_52138_new_n7387_), .B(u2__abc_52138_new_n7379_), .C(rst), .Y(u2__0remHi_451_0__82_));
AOI21X1 AOI21X1_376 ( .A(u2__abc_52138_new_n3758_), .B(u2__abc_52138_new_n7391_), .C(u2__abc_52138_new_n7392_), .Y(u2__abc_52138_new_n7393_));
AOI21X1 AOI21X1_377 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3774_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7395_));
AOI21X1 AOI21X1_378 ( .A(u2__abc_52138_new_n7396_), .B(u2__abc_52138_new_n7389_), .C(rst), .Y(u2__0remHi_451_0__83_));
AOI21X1 AOI21X1_379 ( .A(u2__abc_52138_new_n7403_), .B(u2__abc_52138_new_n7380_), .C(u2__abc_52138_new_n7404_), .Y(u2__abc_52138_new_n7405_));
AOI21X1 AOI21X1_38 ( .A(u2__abc_52138_new_n3886_), .B(u2__abc_52138_new_n3882_), .C(u2__abc_52138_new_n3885_), .Y(u2__abc_52138_new_n3887_));
AOI21X1 AOI21X1_380 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3763_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7413_));
AOI21X1 AOI21X1_381 ( .A(u2__abc_52138_new_n7414_), .B(u2__abc_52138_new_n7398_), .C(rst), .Y(u2__0remHi_451_0__84_));
AOI21X1 AOI21X1_382 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3768_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7421_));
AOI21X1 AOI21X1_383 ( .A(u2__abc_52138_new_n7422_), .B(u2__abc_52138_new_n7416_), .C(rst), .Y(u2__0remHi_451_0__85_));
AOI21X1 AOI21X1_384 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3730_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7432_));
AOI21X1 AOI21X1_385 ( .A(u2__abc_52138_new_n7433_), .B(u2__abc_52138_new_n7424_), .C(rst), .Y(u2__0remHi_451_0__86_));
AOI21X1 AOI21X1_386 ( .A(u2__abc_52138_new_n7437_), .B(u2__abc_52138_new_n7438_), .C(u2__abc_52138_new_n7439_), .Y(u2__abc_52138_new_n7440_));
AOI21X1 AOI21X1_387 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3724_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7442_));
AOI21X1 AOI21X1_388 ( .A(u2__abc_52138_new_n7443_), .B(u2__abc_52138_new_n7435_), .C(rst), .Y(u2__0remHi_451_0__87_));
AOI21X1 AOI21X1_389 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3715_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7458_));
AOI21X1 AOI21X1_39 ( .A(u2__abc_52138_new_n3880_), .B(u2__abc_52138_new_n3867_), .C(u2__abc_52138_new_n3893_), .Y(u2__abc_52138_new_n3894_));
AOI21X1 AOI21X1_390 ( .A(u2__abc_52138_new_n7459_), .B(u2__abc_52138_new_n7445_), .C(rst), .Y(u2__0remHi_451_0__88_));
AOI21X1 AOI21X1_391 ( .A(u2__abc_52138_new_n7462_), .B(u2__abc_52138_new_n7464_), .C(u2__abc_52138_new_n7465_), .Y(u2__abc_52138_new_n7466_));
AOI21X1 AOI21X1_392 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3720_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7468_));
AOI21X1 AOI21X1_393 ( .A(u2__abc_52138_new_n7469_), .B(u2__abc_52138_new_n7461_), .C(rst), .Y(u2__0remHi_451_0__89_));
AOI21X1 AOI21X1_394 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3706_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7479_));
AOI21X1 AOI21X1_395 ( .A(u2__abc_52138_new_n7480_), .B(u2__abc_52138_new_n7471_), .C(rst), .Y(u2__0remHi_451_0__90_));
AOI21X1 AOI21X1_396 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3704_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7487_));
AOI21X1 AOI21X1_397 ( .A(u2__abc_52138_new_n7488_), .B(u2__abc_52138_new_n7482_), .C(rst), .Y(u2__0remHi_451_0__91_));
AOI21X1 AOI21X1_398 ( .A(u2__abc_52138_new_n7495_), .B(u2__abc_52138_new_n7496_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n7497_));
AOI21X1 AOI21X1_399 ( .A(u2__abc_52138_new_n3706_), .B(u2__abc_52138_new_n6498_), .C(u2__abc_52138_new_n7497_), .Y(u2__abc_52138_new_n7498_));
AOI21X1 AOI21X1_4 ( .A(u1__abc_51895_new_n329_), .B(u1__abc_51895_new_n375_), .C(u1__abc_51895_new_n278_), .Y(aNan));
AOI21X1 AOI21X1_40 ( .A(u2__abc_52138_new_n3895_), .B(u2__abc_52138_new_n3789_), .C(u2__abc_52138_new_n3794_), .Y(u2__abc_52138_new_n3896_));
AOI21X1 AOI21X1_400 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3693_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7499_));
AOI21X1 AOI21X1_401 ( .A(u2__abc_52138_new_n7500_), .B(u2__abc_52138_new_n7490_), .C(rst), .Y(u2__0remHi_451_0__92_));
AOI21X1 AOI21X1_402 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3698_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7508_));
AOI21X1 AOI21X1_403 ( .A(u2__abc_52138_new_n7509_), .B(u2__abc_52138_new_n7502_), .C(rst), .Y(u2__0remHi_451_0__93_));
AOI21X1 AOI21X1_404 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3660_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7518_));
AOI21X1 AOI21X1_405 ( .A(u2__abc_52138_new_n7519_), .B(u2__abc_52138_new_n7511_), .C(rst), .Y(u2__0remHi_451_0__94_));
AOI21X1 AOI21X1_406 ( .A(u2__abc_52138_new_n7514_), .B(u2__abc_52138_new_n3694_), .C(u2__abc_52138_new_n7522_), .Y(u2__abc_52138_new_n7523_));
AOI21X1 AOI21X1_407 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3655_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7527_));
AOI21X1 AOI21X1_408 ( .A(u2__abc_52138_new_n7528_), .B(u2__abc_52138_new_n7521_), .C(rst), .Y(u2__0remHi_451_0__95_));
AOI21X1 AOI21X1_409 ( .A(u2__abc_52138_new_n7535_), .B(u2__abc_52138_new_n3712_), .C(u2__abc_52138_new_n7537_), .Y(u2__abc_52138_new_n7538_));
AOI21X1 AOI21X1_41 ( .A(u2__abc_52138_new_n3897_), .B(u2__abc_52138_new_n3803_), .C(u2__abc_52138_new_n3898_), .Y(u2__abc_52138_new_n3899_));
AOI21X1 AOI21X1_410 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n3642_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7547_));
AOI21X1 AOI21X1_411 ( .A(u2__abc_52138_new_n7548_), .B(u2__abc_52138_new_n7530_), .C(rst), .Y(u2__0remHi_451_0__96_));
AOI21X1 AOI21X1_412 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3647_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7555_));
AOI21X1 AOI21X1_413 ( .A(u2__abc_52138_new_n7556_), .B(u2__abc_52138_new_n7550_), .C(rst), .Y(u2__0remHi_451_0__97_));
AOI21X1 AOI21X1_414 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3683_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7565_));
AOI21X1 AOI21X1_415 ( .A(u2__abc_52138_new_n7566_), .B(u2__abc_52138_new_n7558_), .C(rst), .Y(u2__0remHi_451_0__98_));
AOI21X1 AOI21X1_416 ( .A(u2__abc_52138_new_n7561_), .B(u2__abc_52138_new_n3942_), .C(u2__abc_52138_new_n3643_), .Y(u2__abc_52138_new_n7571_));
AOI21X1 AOI21X1_417 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3678_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7575_));
AOI21X1 AOI21X1_418 ( .A(u2__abc_52138_new_n7576_), .B(u2__abc_52138_new_n7568_), .C(rst), .Y(u2__0remHi_451_0__99_));
AOI21X1 AOI21X1_419 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3667_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7593_));
AOI21X1 AOI21X1_42 ( .A(u2__abc_52138_new_n3901_), .B(u2__abc_52138_new_n3827_), .C(u2__abc_52138_new_n3822_), .Y(u2__abc_52138_new_n3902_));
AOI21X1 AOI21X1_420 ( .A(u2__abc_52138_new_n7594_), .B(u2__abc_52138_new_n7578_), .C(rst), .Y(u2__0remHi_451_0__100_));
AOI21X1 AOI21X1_421 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3672_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7601_));
AOI21X1 AOI21X1_422 ( .A(u2__abc_52138_new_n7602_), .B(u2__abc_52138_new_n7596_), .C(rst), .Y(u2__0remHi_451_0__101_));
AOI21X1 AOI21X1_423 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3612_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7612_));
AOI21X1 AOI21X1_424 ( .A(u2__abc_52138_new_n7613_), .B(u2__abc_52138_new_n7604_), .C(rst), .Y(u2__0remHi_451_0__102_));
AOI21X1 AOI21X1_425 ( .A(u2__abc_52138_new_n7616_), .B(u2__abc_52138_new_n7617_), .C(u2__abc_52138_new_n7618_), .Y(u2__abc_52138_new_n7619_));
AOI21X1 AOI21X1_426 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3610_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7621_));
AOI21X1 AOI21X1_427 ( .A(u2__abc_52138_new_n7622_), .B(u2__abc_52138_new_n7615_), .C(rst), .Y(u2__0remHi_451_0__103_));
AOI21X1 AOI21X1_428 ( .A(u2__abc_52138_new_n7626_), .B(u2__abc_52138_new_n7605_), .C(u2__abc_52138_new_n7627_), .Y(u2__abc_52138_new_n7628_));
AOI21X1 AOI21X1_429 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3599_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7638_));
AOI21X1 AOI21X1_43 ( .A(u2__abc_52138_new_n3811_), .B(u2__abc_52138_new_n3903_), .C(u2__abc_52138_new_n3816_), .Y(u2__abc_52138_new_n3904_));
AOI21X1 AOI21X1_430 ( .A(u2__abc_52138_new_n7639_), .B(u2__abc_52138_new_n7624_), .C(rst), .Y(u2__0remHi_451_0__104_));
AOI21X1 AOI21X1_431 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3604_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7647_));
AOI21X1 AOI21X1_432 ( .A(u2__abc_52138_new_n7648_), .B(u2__abc_52138_new_n7641_), .C(rst), .Y(u2__0remHi_451_0__105_));
AOI21X1 AOI21X1_433 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3634_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7658_));
AOI21X1 AOI21X1_434 ( .A(u2__abc_52138_new_n7659_), .B(u2__abc_52138_new_n7650_), .C(rst), .Y(u2__0remHi_451_0__106_));
AOI21X1 AOI21X1_435 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3632_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7666_));
AOI21X1 AOI21X1_436 ( .A(u2__abc_52138_new_n7667_), .B(u2__abc_52138_new_n7661_), .C(rst), .Y(u2__0remHi_451_0__107_));
AOI21X1 AOI21X1_437 ( .A(u2__abc_52138_new_n7677_), .B(u2__abc_52138_new_n7675_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n7678_));
AOI21X1 AOI21X1_438 ( .A(u2__abc_52138_new_n3634_), .B(u2__abc_52138_new_n6498_), .C(u2__abc_52138_new_n7678_), .Y(u2__abc_52138_new_n7679_));
AOI21X1 AOI21X1_439 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3621_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7680_));
AOI21X1 AOI21X1_44 ( .A(u2__abc_52138_new_n3900_), .B(u2__abc_52138_new_n3830_), .C(u2__abc_52138_new_n3905_), .Y(u2__abc_52138_new_n3906_));
AOI21X1 AOI21X1_440 ( .A(u2__abc_52138_new_n7681_), .B(u2__abc_52138_new_n7669_), .C(rst), .Y(u2__0remHi_451_0__108_));
AOI21X1 AOI21X1_441 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3626_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7689_));
AOI21X1 AOI21X1_442 ( .A(u2__abc_52138_new_n7690_), .B(u2__abc_52138_new_n7683_), .C(rst), .Y(u2__0remHi_451_0__109_));
AOI21X1 AOI21X1_443 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3552_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7699_));
AOI21X1 AOI21X1_444 ( .A(u2__abc_52138_new_n7700_), .B(u2__abc_52138_new_n7692_), .C(rst), .Y(u2__0remHi_451_0__110_));
AOI21X1 AOI21X1_445 ( .A(u2__abc_52138_new_n7704_), .B(u2__abc_52138_new_n7706_), .C(u2__abc_52138_new_n7707_), .Y(u2__abc_52138_new_n7708_));
AOI21X1 AOI21X1_446 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3557_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7710_));
AOI21X1 AOI21X1_447 ( .A(u2__abc_52138_new_n7711_), .B(u2__abc_52138_new_n7702_), .C(rst), .Y(u2__0remHi_451_0__111_));
AOI21X1 AOI21X1_448 ( .A(u2__abc_52138_new_n7673_), .B(u2__abc_52138_new_n3640_), .C(u2__abc_52138_new_n7716_), .Y(u2__abc_52138_new_n7717_));
AOI21X1 AOI21X1_449 ( .A(u2__abc_52138_new_n7629_), .B(u2__abc_52138_new_n7715_), .C(u2__abc_52138_new_n7718_), .Y(u2__abc_52138_new_n7719_));
AOI21X1 AOI21X1_45 ( .A(u2__abc_52138_new_n3908_), .B(u2__abc_52138_new_n3744_), .C(u2__abc_52138_new_n3909_), .Y(u2__abc_52138_new_n3910_));
AOI21X1 AOI21X1_450 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3563_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7725_));
AOI21X1 AOI21X1_451 ( .A(u2__abc_52138_new_n7726_), .B(u2__abc_52138_new_n7713_), .C(rst), .Y(u2__0remHi_451_0__112_));
AOI21X1 AOI21X1_452 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3568_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7734_));
AOI21X1 AOI21X1_453 ( .A(u2__abc_52138_new_n7735_), .B(u2__abc_52138_new_n7728_), .C(rst), .Y(u2__0remHi_451_0__113_));
AOI21X1 AOI21X1_454 ( .A(u2__abc_52138_new_n7721_), .B(u2__abc_52138_new_n3560_), .C(u2__abc_52138_new_n7738_), .Y(u2__abc_52138_new_n7739_));
AOI21X1 AOI21X1_455 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3590_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7745_));
AOI21X1 AOI21X1_456 ( .A(u2__abc_52138_new_n7746_), .B(u2__abc_52138_new_n7737_), .C(rst), .Y(u2__0remHi_451_0__114_));
AOI21X1 AOI21X1_457 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3585_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7753_));
AOI21X1 AOI21X1_458 ( .A(u2__abc_52138_new_n7754_), .B(u2__abc_52138_new_n7748_), .C(rst), .Y(u2__0remHi_451_0__115_));
AOI21X1 AOI21X1_459 ( .A(u2__abc_52138_new_n7721_), .B(u2__abc_52138_new_n3572_), .C(u2__abc_52138_new_n7760_), .Y(u2__abc_52138_new_n7761_));
AOI21X1 AOI21X1_46 ( .A(u2__abc_52138_new_n3911_), .B(u2__abc_52138_new_n3755_), .C(u2__abc_52138_new_n3912_), .Y(u2__abc_52138_new_n3913_));
AOI21X1 AOI21X1_460 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3573_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7767_));
AOI21X1 AOI21X1_461 ( .A(u2__abc_52138_new_n7768_), .B(u2__abc_52138_new_n7756_), .C(rst), .Y(u2__0remHi_451_0__116_));
AOI21X1 AOI21X1_462 ( .A(u2__abc_52138_new_n7771_), .B(u2__abc_52138_new_n7772_), .C(u2__abc_52138_new_n7773_), .Y(u2__abc_52138_new_n7774_));
AOI21X1 AOI21X1_463 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3580_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7776_));
AOI21X1 AOI21X1_464 ( .A(u2__abc_52138_new_n7777_), .B(u2__abc_52138_new_n7770_), .C(rst), .Y(u2__0remHi_451_0__117_));
AOI21X1 AOI21X1_465 ( .A(u2__abc_52138_new_n7785_), .B(u2__abc_52138_new_n7783_), .C(u2__abc_52138_new_n7786_), .Y(u2__abc_52138_new_n7787_));
AOI21X1 AOI21X1_466 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3508_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7797_));
AOI21X1 AOI21X1_467 ( .A(u2__abc_52138_new_n7798_), .B(u2__abc_52138_new_n7791_), .C(rst), .Y(u2__0remHi_451_0__119_));
AOI21X1 AOI21X1_468 ( .A(u2__abc_52138_new_n7810_), .B(u2__abc_52138_new_n3507_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n7812_));
AOI21X1 AOI21X1_469 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3518_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7815_));
AOI21X1 AOI21X1_47 ( .A(u2__abc_52138_new_n3914_), .B(u2__abc_52138_new_n3783_), .C(u2__abc_52138_new_n3921_), .Y(u2__abc_52138_new_n3922_));
AOI21X1 AOI21X1_470 ( .A(u2__abc_52138_new_n7816_), .B(u2__abc_52138_new_n7800_), .C(rst), .Y(u2__0remHi_451_0__120_));
AOI21X1 AOI21X1_471 ( .A(u2__abc_52138_new_n7819_), .B(u2__abc_52138_new_n7820_), .C(u2__abc_52138_new_n7821_), .Y(u2__abc_52138_new_n7822_));
AOI21X1 AOI21X1_472 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3523_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7824_));
AOI21X1 AOI21X1_473 ( .A(u2__abc_52138_new_n7825_), .B(u2__abc_52138_new_n7818_), .C(rst), .Y(u2__0remHi_451_0__121_));
AOI21X1 AOI21X1_474 ( .A(u2__abc_52138_new_n7828_), .B(u2__abc_52138_new_n7832_), .C(u2__abc_52138_new_n7833_), .Y(u2__abc_52138_new_n7834_));
AOI21X1 AOI21X1_475 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3542_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7836_));
AOI21X1 AOI21X1_476 ( .A(u2__abc_52138_new_n7837_), .B(u2__abc_52138_new_n7827_), .C(rst), .Y(u2__0remHi_451_0__122_));
AOI21X1 AOI21X1_477 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3540_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7845_));
AOI21X1 AOI21X1_478 ( .A(u2__abc_52138_new_n7846_), .B(u2__abc_52138_new_n7839_), .C(rst), .Y(u2__0remHi_451_0__123_));
AOI21X1 AOI21X1_479 ( .A(u2__abc_52138_new_n7829_), .B(u2__abc_52138_new_n3526_), .C(u2__abc_52138_new_n7849_), .Y(u2__abc_52138_new_n7850_));
AOI21X1 AOI21X1_48 ( .A(u2__abc_52138_new_n3726_), .B(u2__abc_52138_new_n3733_), .C(u2__abc_52138_new_n3728_), .Y(u2__abc_52138_new_n3923_));
AOI21X1 AOI21X1_480 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n3532_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7867_));
AOI21X1 AOI21X1_481 ( .A(u2__abc_52138_new_n7868_), .B(u2__abc_52138_new_n7861_), .C(rst), .Y(u2__0remHi_451_0__125_));
AOI21X1 AOI21X1_482 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4715_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7876_));
AOI21X1 AOI21X1_483 ( .A(u2__abc_52138_new_n7877_), .B(u2__abc_52138_new_n7870_), .C(rst), .Y(u2__0remHi_451_0__126_));
AOI21X1 AOI21X1_484 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4721_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7884_));
AOI21X1 AOI21X1_485 ( .A(u2__abc_52138_new_n7885_), .B(u2__abc_52138_new_n7879_), .C(rst), .Y(u2__0remHi_451_0__127_));
AOI21X1 AOI21X1_486 ( .A(u2__abc_52138_new_n7808_), .B(u2__abc_52138_new_n6489_), .C(u2__abc_52138_new_n7895_), .Y(u2__abc_52138_new_n7896_));
AOI21X1 AOI21X1_487 ( .A(u2__abc_52138_new_n7539_), .B(u2__abc_52138_new_n7892_), .C(u2__abc_52138_new_n7897_), .Y(u2__abc_52138_new_n7898_));
AOI21X1 AOI21X1_488 ( .A(u2__abc_52138_new_n2991_), .B(u2__abc_52138_new_n7905_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7906_));
AOI21X1 AOI21X1_489 ( .A(u2__abc_52138_new_n7907_), .B(u2__abc_52138_new_n7887_), .C(rst), .Y(u2__0remHi_451_0__128_));
AOI21X1 AOI21X1_49 ( .A(u2__abc_52138_new_n3712_), .B(u2__abc_52138_new_n3927_), .C(u2__abc_52138_new_n3935_), .Y(u2__abc_52138_new_n3936_));
AOI21X1 AOI21X1_490 ( .A(u2__abc_52138_new_n4724_), .B(u2__abc_52138_new_n7910_), .C(u2__abc_52138_new_n7911_), .Y(u2__abc_52138_new_n7912_));
AOI21X1 AOI21X1_491 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4729_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7914_));
AOI21X1 AOI21X1_492 ( .A(u2__abc_52138_new_n7915_), .B(u2__abc_52138_new_n7909_), .C(rst), .Y(u2__0remHi_451_0__129_));
AOI21X1 AOI21X1_493 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4776_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7924_));
AOI21X1 AOI21X1_494 ( .A(u2__abc_52138_new_n7925_), .B(u2__abc_52138_new_n7917_), .C(rst), .Y(u2__0remHi_451_0__130_));
AOI21X1 AOI21X1_495 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4746_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7934_));
AOI21X1 AOI21X1_496 ( .A(u2__abc_52138_new_n7935_), .B(u2__abc_52138_new_n7927_), .C(rst), .Y(u2__0remHi_451_0__131_));
AOI21X1 AOI21X1_497 ( .A(u2__abc_52138_new_n7939_), .B(u2__abc_52138_new_n7918_), .C(u2__abc_52138_new_n7941_), .Y(u2__abc_52138_new_n7942_));
AOI21X1 AOI21X1_498 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4735_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7950_));
AOI21X1 AOI21X1_499 ( .A(u2__abc_52138_new_n7951_), .B(u2__abc_52138_new_n7937_), .C(rst), .Y(u2__0remHi_451_0__132_));
AOI21X1 AOI21X1_5 ( .A(u2__abc_52138_new_n2979_), .B(u2__abc_52138_new_n2965_), .C(rst), .Y(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_2_));
AOI21X1 AOI21X1_50 ( .A(u2__abc_52138_new_n3907_), .B(u2__abc_52138_new_n3785_), .C(u2__abc_52138_new_n3937_), .Y(u2__abc_52138_new_n3938_));
AOI21X1 AOI21X1_500 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4740_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7958_));
AOI21X1 AOI21X1_501 ( .A(u2__abc_52138_new_n7959_), .B(u2__abc_52138_new_n7953_), .C(rst), .Y(u2__0remHi_451_0__133_));
AOI21X1 AOI21X1_502 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4679_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7969_));
AOI21X1 AOI21X1_503 ( .A(u2__abc_52138_new_n7970_), .B(u2__abc_52138_new_n7961_), .C(rst), .Y(u2__0remHi_451_0__134_));
AOI21X1 AOI21X1_504 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4684_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7977_));
AOI21X1 AOI21X1_505 ( .A(u2__abc_52138_new_n7978_), .B(u2__abc_52138_new_n7972_), .C(rst), .Y(u2__0remHi_451_0__135_));
AOI21X1 AOI21X1_506 ( .A(u2__abc_52138_new_n7984_), .B(u2__abc_52138_new_n4741_), .C(u2__abc_52138_new_n4780_), .Y(u2__abc_52138_new_n7985_));
AOI21X1 AOI21X1_507 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4668_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n7995_));
AOI21X1 AOI21X1_508 ( .A(u2__abc_52138_new_n7996_), .B(u2__abc_52138_new_n7980_), .C(rst), .Y(u2__0remHi_451_0__136_));
AOI21X1 AOI21X1_509 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4673_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8003_));
AOI21X1 AOI21X1_51 ( .A(u2__abc_52138_new_n3940_), .B(u2__abc_52138_new_n3654_), .C(u2__abc_52138_new_n3939_), .Y(u2__abc_52138_new_n3941_));
AOI21X1 AOI21X1_510 ( .A(u2__abc_52138_new_n8004_), .B(u2__abc_52138_new_n7998_), .C(rst), .Y(u2__0remHi_451_0__137_));
AOI21X1 AOI21X1_511 ( .A(u2__abc_52138_new_n7999_), .B(u2__abc_52138_new_n4685_), .C(u2__abc_52138_new_n8007_), .Y(u2__abc_52138_new_n8008_));
AOI21X1 AOI21X1_512 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4707_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8016_));
AOI21X1 AOI21X1_513 ( .A(u2__abc_52138_new_n8017_), .B(u2__abc_52138_new_n8006_), .C(rst), .Y(u2__0remHi_451_0__138_));
AOI21X1 AOI21X1_514 ( .A(u2__abc_52138_new_n8021_), .B(u2__abc_52138_new_n8022_), .C(u2__abc_52138_new_n8023_), .Y(u2__abc_52138_new_n8024_));
AOI21X1 AOI21X1_515 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4702_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8026_));
AOI21X1 AOI21X1_516 ( .A(u2__abc_52138_new_n8027_), .B(u2__abc_52138_new_n8019_), .C(rst), .Y(u2__0remHi_451_0__139_));
AOI21X1 AOI21X1_517 ( .A(u2__abc_52138_new_n8010_), .B(u2__abc_52138_new_n4674_), .C(u2__abc_52138_new_n4789_), .Y(u2__abc_52138_new_n8032_));
AOI21X1 AOI21X1_518 ( .A(u2__abc_52138_new_n7988_), .B(u2__abc_52138_new_n4688_), .C(u2__abc_52138_new_n8033_), .Y(u2__abc_52138_new_n8034_));
AOI21X1 AOI21X1_519 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4691_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8040_));
AOI21X1 AOI21X1_52 ( .A(u2__abc_52138_new_n3949_), .B(u2__abc_52138_new_n3677_), .C(u2__abc_52138_new_n3948_), .Y(u2__abc_52138_new_n3950_));
AOI21X1 AOI21X1_520 ( .A(u2__abc_52138_new_n8041_), .B(u2__abc_52138_new_n8029_), .C(rst), .Y(u2__0remHi_451_0__140_));
AOI21X1 AOI21X1_521 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4696_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8048_));
AOI21X1 AOI21X1_522 ( .A(u2__abc_52138_new_n8049_), .B(u2__abc_52138_new_n8043_), .C(rst), .Y(u2__0remHi_451_0__141_));
AOI21X1 AOI21X1_523 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4658_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8057_));
AOI21X1 AOI21X1_524 ( .A(u2__abc_52138_new_n8058_), .B(u2__abc_52138_new_n8051_), .C(rst), .Y(u2__0remHi_451_0__142_));
AOI21X1 AOI21X1_525 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4652_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8065_));
AOI21X1 AOI21X1_526 ( .A(u2__abc_52138_new_n8066_), .B(u2__abc_52138_new_n8060_), .C(rst), .Y(u2__0remHi_451_0__143_));
AOI21X1 AOI21X1_527 ( .A(u2__abc_52138_new_n8074_), .B(u2__abc_52138_new_n4699_), .C(u2__abc_52138_new_n8075_), .Y(u2__abc_52138_new_n8076_));
AOI21X1 AOI21X1_528 ( .A(u2__abc_52138_new_n8072_), .B(u2__abc_52138_new_n8071_), .C(u2__abc_52138_new_n8077_), .Y(u2__abc_52138_new_n8078_));
AOI21X1 AOI21X1_529 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4644_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8088_));
AOI21X1 AOI21X1_53 ( .A(u2__abc_52138_new_n3951_), .B(u2__abc_52138_new_n3671_), .C(u2__abc_52138_new_n3952_), .Y(u2__abc_52138_new_n3953_));
AOI21X1 AOI21X1_530 ( .A(u2__abc_52138_new_n8089_), .B(u2__abc_52138_new_n8068_), .C(rst), .Y(u2__0remHi_451_0__144_));
AOI21X1 AOI21X1_531 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4649_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8097_));
AOI21X1 AOI21X1_532 ( .A(u2__abc_52138_new_n8098_), .B(u2__abc_52138_new_n8091_), .C(rst), .Y(u2__0remHi_451_0__145_));
AOI21X1 AOI21X1_533 ( .A(u2__abc_52138_new_n8093_), .B(u2__abc_52138_new_n4657_), .C(u2__abc_52138_new_n4653_), .Y(u2__abc_52138_new_n8102_));
AOI21X1 AOI21X1_534 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4637_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8108_));
AOI21X1 AOI21X1_535 ( .A(u2__abc_52138_new_n8109_), .B(u2__abc_52138_new_n8100_), .C(rst), .Y(u2__0remHi_451_0__146_));
AOI21X1 AOI21X1_536 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4632_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8117_));
AOI21X1 AOI21X1_537 ( .A(u2__abc_52138_new_n8118_), .B(u2__abc_52138_new_n8111_), .C(rst), .Y(u2__0remHi_451_0__147_));
AOI21X1 AOI21X1_538 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4621_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8128_));
AOI21X1 AOI21X1_539 ( .A(u2__abc_52138_new_n8129_), .B(u2__abc_52138_new_n8120_), .C(rst), .Y(u2__0remHi_451_0__148_));
AOI21X1 AOI21X1_54 ( .A(u2__abc_52138_new_n3946_), .B(u2__abc_52138_new_n3687_), .C(u2__abc_52138_new_n3954_), .Y(u2__abc_52138_new_n3955_));
AOI21X1 AOI21X1_540 ( .A(u2__abc_52138_new_n8132_), .B(u2__abc_52138_new_n8133_), .C(u2__abc_52138_new_n8134_), .Y(u2__abc_52138_new_n8135_));
AOI21X1 AOI21X1_541 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4626_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8137_));
AOI21X1 AOI21X1_542 ( .A(u2__abc_52138_new_n8138_), .B(u2__abc_52138_new_n8131_), .C(rst), .Y(u2__0remHi_451_0__149_));
AOI21X1 AOI21X1_543 ( .A(u2__abc_52138_new_n8147_), .B(u2__abc_52138_new_n8145_), .C(u2__abc_52138_new_n8148_), .Y(u2__abc_52138_new_n8149_));
AOI21X1 AOI21X1_544 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4586_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8158_));
AOI21X1 AOI21X1_545 ( .A(u2__abc_52138_new_n8159_), .B(u2__abc_52138_new_n8153_), .C(rst), .Y(u2__0remHi_451_0__151_));
AOI21X1 AOI21X1_546 ( .A(u2__abc_52138_new_n8167_), .B(u2__abc_52138_new_n4641_), .C(u2__abc_52138_new_n8168_), .Y(u2__abc_52138_new_n8169_));
AOI21X1 AOI21X1_547 ( .A(u2__abc_52138_new_n8080_), .B(u2__abc_52138_new_n8078_), .C(u2__abc_52138_new_n4761_), .Y(u2__abc_52138_new_n8171_));
AOI21X1 AOI21X1_548 ( .A(u2__abc_52138_new_n8174_), .B(u2__abc_52138_new_n8172_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8175_));
AOI21X1 AOI21X1_549 ( .A(u2__abc_52138_new_n4591_), .B(u2__abc_52138_new_n6498_), .C(u2__abc_52138_new_n8175_), .Y(u2__abc_52138_new_n8176_));
AOI21X1 AOI21X1_55 ( .A(u2__abc_52138_new_n3640_), .B(u2__abc_52138_new_n3961_), .C(u2__abc_52138_new_n3968_), .Y(u2__abc_52138_new_n3969_));
AOI21X1 AOI21X1_550 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4575_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8177_));
AOI21X1 AOI21X1_551 ( .A(u2__abc_52138_new_n8178_), .B(u2__abc_52138_new_n8161_), .C(rst), .Y(u2__0remHi_451_0__152_));
AOI21X1 AOI21X1_552 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4580_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8185_));
AOI21X1 AOI21X1_553 ( .A(u2__abc_52138_new_n8186_), .B(u2__abc_52138_new_n8180_), .C(rst), .Y(u2__0remHi_451_0__153_));
AOI21X1 AOI21X1_554 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4612_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8195_));
AOI21X1 AOI21X1_555 ( .A(u2__abc_52138_new_n8196_), .B(u2__abc_52138_new_n8188_), .C(rst), .Y(u2__0remHi_451_0__154_));
AOI21X1 AOI21X1_556 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4607_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8203_));
AOI21X1 AOI21X1_557 ( .A(u2__abc_52138_new_n8204_), .B(u2__abc_52138_new_n8198_), .C(rst), .Y(u2__0remHi_451_0__155_));
AOI21X1 AOI21X1_558 ( .A(u2__abc_52138_new_n8207_), .B(u2__abc_52138_new_n4583_), .C(u2__abc_52138_new_n8208_), .Y(u2__abc_52138_new_n8209_));
AOI21X1 AOI21X1_559 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4603_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8225_));
AOI21X1 AOI21X1_56 ( .A(u2__abc_52138_new_n3972_), .B(u2__abc_52138_new_n3556_), .C(u2__abc_52138_new_n3973_), .Y(u2__abc_52138_new_n3974_));
AOI21X1 AOI21X1_560 ( .A(u2__abc_52138_new_n8226_), .B(u2__abc_52138_new_n8220_), .C(rst), .Y(u2__0remHi_451_0__157_));
AOI21X1 AOI21X1_561 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4541_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8235_));
AOI21X1 AOI21X1_562 ( .A(u2__abc_52138_new_n8236_), .B(u2__abc_52138_new_n8228_), .C(rst), .Y(u2__0remHi_451_0__158_));
AOI21X1 AOI21X1_563 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n8243_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8244_));
AOI21X1 AOI21X1_564 ( .A(u2__abc_52138_new_n8245_), .B(u2__abc_52138_new_n8238_), .C(rst), .Y(u2__0remHi_451_0__159_));
AOI21X1 AOI21X1_565 ( .A(u2__abc_52138_new_n8249_), .B(u2__abc_52138_new_n4606_), .C(u2__abc_52138_new_n8250_), .Y(u2__abc_52138_new_n8251_));
AOI21X1 AOI21X1_566 ( .A(u2__abc_52138_new_n4618_), .B(u2__abc_52138_new_n8170_), .C(u2__abc_52138_new_n8253_), .Y(u2__abc_52138_new_n8254_));
AOI21X1 AOI21X1_567 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4527_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8264_));
AOI21X1 AOI21X1_568 ( .A(u2__abc_52138_new_n8265_), .B(u2__abc_52138_new_n8247_), .C(rst), .Y(u2__0remHi_451_0__160_));
AOI21X1 AOI21X1_569 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4532_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8272_));
AOI21X1 AOI21X1_57 ( .A(u2__abc_52138_new_n3978_), .B(u2__abc_52138_new_n3594_), .C(u2__abc_52138_new_n3985_), .Y(u2__abc_52138_new_n3986_));
AOI21X1 AOI21X1_570 ( .A(u2__abc_52138_new_n8273_), .B(u2__abc_52138_new_n8267_), .C(rst), .Y(u2__0remHi_451_0__161_));
AOI21X1 AOI21X1_571 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4566_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8285_));
AOI21X1 AOI21X1_572 ( .A(u2__abc_52138_new_n8286_), .B(u2__abc_52138_new_n8275_), .C(rst), .Y(u2__0remHi_451_0__162_));
AOI21X1 AOI21X1_573 ( .A(u2__abc_52138_new_n8290_), .B(u2__abc_52138_new_n8291_), .C(u2__abc_52138_new_n8292_), .Y(u2__abc_52138_new_n8293_));
AOI21X1 AOI21X1_574 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4561_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8295_));
AOI21X1 AOI21X1_575 ( .A(u2__abc_52138_new_n8296_), .B(u2__abc_52138_new_n8288_), .C(rst), .Y(u2__0remHi_451_0__163_));
AOI21X1 AOI21X1_576 ( .A(u2__abc_52138_new_n8279_), .B(u2__abc_52138_new_n4533_), .C(u2__abc_52138_new_n4833_), .Y(u2__abc_52138_new_n8300_));
AOI21X1 AOI21X1_577 ( .A(u2__abc_52138_new_n8256_), .B(u2__abc_52138_new_n4547_), .C(u2__abc_52138_new_n8301_), .Y(u2__abc_52138_new_n8302_));
AOI21X1 AOI21X1_578 ( .A(u2__abc_52138_new_n8304_), .B(u2__abc_52138_new_n8305_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8306_));
AOI21X1 AOI21X1_579 ( .A(u2__abc_52138_new_n4566_), .B(u2__abc_52138_new_n6498_), .C(u2__abc_52138_new_n8306_), .Y(u2__abc_52138_new_n8307_));
AOI21X1 AOI21X1_58 ( .A(u2__abc_52138_new_n3995_), .B(u2__abc_52138_new_n3991_), .C(u2__abc_52138_new_n3993_), .Y(u2__abc_52138_new_n3996_));
AOI21X1 AOI21X1_580 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4550_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8308_));
AOI21X1 AOI21X1_581 ( .A(u2__abc_52138_new_n8309_), .B(u2__abc_52138_new_n8298_), .C(rst), .Y(u2__0remHi_451_0__164_));
AOI21X1 AOI21X1_582 ( .A(u2__abc_52138_new_n8312_), .B(u2__abc_52138_new_n8313_), .C(u2__abc_52138_new_n8314_), .Y(u2__abc_52138_new_n8315_));
AOI21X1 AOI21X1_583 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4555_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8317_));
AOI21X1 AOI21X1_584 ( .A(u2__abc_52138_new_n8318_), .B(u2__abc_52138_new_n8311_), .C(rst), .Y(u2__0remHi_451_0__165_));
AOI21X1 AOI21X1_585 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4517_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8327_));
AOI21X1 AOI21X1_586 ( .A(u2__abc_52138_new_n8328_), .B(u2__abc_52138_new_n8320_), .C(rst), .Y(u2__0remHi_451_0__166_));
AOI21X1 AOI21X1_587 ( .A(u2__abc_52138_new_n8323_), .B(u2__abc_52138_new_n4551_), .C(u2__abc_52138_new_n8331_), .Y(u2__abc_52138_new_n8332_));
AOI21X1 AOI21X1_588 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4514_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8336_));
AOI21X1 AOI21X1_589 ( .A(u2__abc_52138_new_n8337_), .B(u2__abc_52138_new_n8330_), .C(rst), .Y(u2__0remHi_451_0__167_));
AOI21X1 AOI21X1_59 ( .A(u2__abc_52138_new_n3990_), .B(u2__abc_52138_new_n3548_), .C(u2__abc_52138_new_n3997_), .Y(u2__abc_52138_new_n3998_));
AOI21X1 AOI21X1_590 ( .A(u2__abc_52138_new_n8301_), .B(u2__abc_52138_new_n4570_), .C(u2__abc_52138_new_n8340_), .Y(u2__abc_52138_new_n8341_));
AOI21X1 AOI21X1_591 ( .A(u2__abc_52138_new_n8345_), .B(u2__abc_52138_new_n4521_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8348_));
AOI21X1 AOI21X1_592 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4503_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8351_));
AOI21X1 AOI21X1_593 ( .A(u2__abc_52138_new_n8352_), .B(u2__abc_52138_new_n8339_), .C(rst), .Y(u2__0remHi_451_0__168_));
AOI21X1 AOI21X1_594 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4508_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8359_));
AOI21X1 AOI21X1_595 ( .A(u2__abc_52138_new_n8360_), .B(u2__abc_52138_new_n8354_), .C(rst), .Y(u2__0remHi_451_0__169_));
AOI21X1 AOI21X1_596 ( .A(u2__abc_52138_new_n8355_), .B(u2__abc_52138_new_n4515_), .C(u2__abc_52138_new_n8363_), .Y(u2__abc_52138_new_n8364_));
AOI21X1 AOI21X1_597 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4496_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8370_));
AOI21X1 AOI21X1_598 ( .A(u2__abc_52138_new_n8371_), .B(u2__abc_52138_new_n8362_), .C(rst), .Y(u2__0remHi_451_0__170_));
AOI21X1 AOI21X1_599 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4491_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8378_));
AOI21X1 AOI21X1_6 ( .A(u2__abc_52138_new_n3073_), .B(u2__abc_52138_new_n3076_), .C(u2__abc_52138_new_n3075_), .Y(u2__abc_52138_new_n3077_));
AOI21X1 AOI21X1_60 ( .A(u2__abc_52138_new_n3970_), .B(u2__abc_52138_new_n3596_), .C(u2__abc_52138_new_n3999_), .Y(u2__abc_52138_new_n4000_));
AOI21X1 AOI21X1_600 ( .A(u2__abc_52138_new_n8379_), .B(u2__abc_52138_new_n8373_), .C(rst), .Y(u2__0remHi_451_0__171_));
AOI21X1 AOI21X1_601 ( .A(u2__abc_52138_new_n8383_), .B(u2__abc_52138_new_n4498_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8386_));
AOI21X1 AOI21X1_602 ( .A(u2__abc_52138_new_n8385_), .B(u2__abc_52138_new_n8386_), .C(u2__abc_52138_new_n8387_), .Y(u2__abc_52138_new_n8388_));
AOI21X1 AOI21X1_603 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4485_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8397_));
AOI21X1 AOI21X1_604 ( .A(u2__abc_52138_new_n8398_), .B(u2__abc_52138_new_n8392_), .C(rst), .Y(u2__0remHi_451_0__173_));
AOI21X1 AOI21X1_605 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4465_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8406_));
AOI21X1 AOI21X1_606 ( .A(u2__abc_52138_new_n8407_), .B(u2__abc_52138_new_n8400_), .C(rst), .Y(u2__0remHi_451_0__174_));
AOI21X1 AOI21X1_607 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4471_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8414_));
AOI21X1 AOI21X1_608 ( .A(u2__abc_52138_new_n8415_), .B(u2__abc_52138_new_n8409_), .C(rst), .Y(u2__0remHi_451_0__175_));
AOI21X1 AOI21X1_609 ( .A(u2__abc_52138_new_n8421_), .B(u2__abc_52138_new_n4755_), .C(u2__abc_52138_new_n8427_), .Y(u2__abc_52138_new_n8428_));
AOI21X1 AOI21X1_61 ( .A(u2__abc_52138_new_n3502_), .B(u2__abc_52138_new_n3871_), .C(u2__abc_52138_new_n4001_), .Y(u2__abc_52138_new_n4002_));
AOI21X1 AOI21X1_610 ( .A(u2__abc_52138_new_n8432_), .B(u2__abc_52138_new_n4467_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8433_));
AOI21X1 AOI21X1_611 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4454_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8436_));
AOI21X1 AOI21X1_612 ( .A(u2__abc_52138_new_n8437_), .B(u2__abc_52138_new_n8417_), .C(rst), .Y(u2__0remHi_451_0__176_));
AOI21X1 AOI21X1_613 ( .A(u2__abc_52138_new_n4474_), .B(u2__abc_52138_new_n8440_), .C(u2__abc_52138_new_n8441_), .Y(u2__abc_52138_new_n8442_));
AOI21X1 AOI21X1_614 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4459_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8444_));
AOI21X1 AOI21X1_615 ( .A(u2__abc_52138_new_n8445_), .B(u2__abc_52138_new_n8439_), .C(rst), .Y(u2__0remHi_451_0__177_));
AOI21X1 AOI21X1_616 ( .A(u2__abc_52138_new_n8456_), .B(u2__abc_52138_new_n8454_), .C(u2__abc_52138_new_n8457_), .Y(u2__abc_52138_new_n8458_));
AOI21X1 AOI21X1_617 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4442_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8467_));
AOI21X1 AOI21X1_618 ( .A(u2__abc_52138_new_n8468_), .B(u2__abc_52138_new_n8462_), .C(rst), .Y(u2__0remHi_451_0__179_));
AOI21X1 AOI21X1_619 ( .A(u2__abc_52138_new_n4462_), .B(u2__abc_52138_new_n8451_), .C(u2__abc_52138_new_n8471_), .Y(u2__abc_52138_new_n8472_));
AOI21X1 AOI21X1_62 ( .A(u2__abc_52138_new_n4767_), .B(u2__abc_52138_new_n4720_), .C(u2__abc_52138_new_n4768_), .Y(u2__abc_52138_new_n4769_));
AOI21X1 AOI21X1_620 ( .A(u2__abc_52138_new_n8474_), .B(u2__abc_52138_new_n4449_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8477_));
AOI21X1 AOI21X1_621 ( .A(u2__abc_52138_new_n8476_), .B(u2__abc_52138_new_n8477_), .C(u2__abc_52138_new_n8478_), .Y(u2__abc_52138_new_n8479_));
AOI21X1 AOI21X1_622 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4436_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8488_));
AOI21X1 AOI21X1_623 ( .A(u2__abc_52138_new_n8489_), .B(u2__abc_52138_new_n8483_), .C(rst), .Y(u2__0remHi_451_0__181_));
AOI21X1 AOI21X1_624 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4384_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8497_));
AOI21X1 AOI21X1_625 ( .A(u2__abc_52138_new_n8498_), .B(u2__abc_52138_new_n8491_), .C(rst), .Y(u2__0remHi_451_0__182_));
AOI21X1 AOI21X1_626 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4389_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8505_));
AOI21X1 AOI21X1_627 ( .A(u2__abc_52138_new_n8506_), .B(u2__abc_52138_new_n8500_), .C(rst), .Y(u2__0remHi_451_0__183_));
AOI21X1 AOI21X1_628 ( .A(u2__abc_52138_new_n4439_), .B(u2__abc_52138_new_n8509_), .C(u2__abc_52138_new_n8512_), .Y(u2__abc_52138_new_n8513_));
AOI21X1 AOI21X1_629 ( .A(u2__abc_52138_new_n8516_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n8517_), .Y(u2__abc_52138_new_n8518_));
AOI21X1 AOI21X1_63 ( .A(u2__abc_52138_new_n4771_), .B(u2__abc_52138_new_n4728_), .C(u2__abc_52138_new_n4772_), .Y(u2__abc_52138_new_n4773_));
AOI21X1 AOI21X1_630 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4400_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8528_));
AOI21X1 AOI21X1_631 ( .A(u2__abc_52138_new_n8529_), .B(u2__abc_52138_new_n8522_), .C(rst), .Y(u2__0remHi_451_0__185_));
AOI21X1 AOI21X1_632 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4423_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8539_));
AOI21X1 AOI21X1_633 ( .A(u2__abc_52138_new_n8540_), .B(u2__abc_52138_new_n8531_), .C(rst), .Y(u2__0remHi_451_0__186_));
AOI21X1 AOI21X1_634 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4418_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8548_));
AOI21X1 AOI21X1_635 ( .A(u2__abc_52138_new_n8549_), .B(u2__abc_52138_new_n8542_), .C(rst), .Y(u2__0remHi_451_0__187_));
AOI21X1 AOI21X1_636 ( .A(u2__abc_52138_new_n8532_), .B(u2__abc_52138_new_n4403_), .C(u2__abc_52138_new_n8552_), .Y(u2__abc_52138_new_n8553_));
AOI21X1 AOI21X1_637 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4407_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8561_));
AOI21X1 AOI21X1_638 ( .A(u2__abc_52138_new_n8562_), .B(u2__abc_52138_new_n8551_), .C(rst), .Y(u2__0remHi_451_0__188_));
AOI21X1 AOI21X1_639 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4412_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8569_));
AOI21X1 AOI21X1_64 ( .A(u2__abc_52138_new_n4774_), .B(u2__abc_52138_new_n4766_), .C(u2__abc_52138_new_n4783_), .Y(u2__abc_52138_new_n4784_));
AOI21X1 AOI21X1_640 ( .A(u2__abc_52138_new_n8570_), .B(u2__abc_52138_new_n8564_), .C(rst), .Y(u2__0remHi_451_0__189_));
AOI21X1 AOI21X1_641 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4364_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8578_));
AOI21X1 AOI21X1_642 ( .A(u2__abc_52138_new_n8579_), .B(u2__abc_52138_new_n8572_), .C(rst), .Y(u2__0remHi_451_0__190_));
AOI21X1 AOI21X1_643 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4369_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8586_));
AOI21X1 AOI21X1_644 ( .A(u2__abc_52138_new_n8587_), .B(u2__abc_52138_new_n8581_), .C(rst), .Y(u2__0remHi_451_0__191_));
AOI21X1 AOI21X1_645 ( .A(u2__abc_52138_new_n8596_), .B(u2__abc_52138_new_n4413_), .C(u2__abc_52138_new_n4872_), .Y(u2__abc_52138_new_n8597_));
AOI21X1 AOI21X1_646 ( .A(u2__abc_52138_new_n8429_), .B(u2__abc_52138_new_n4754_), .C(u2__abc_52138_new_n8599_), .Y(u2__abc_52138_new_n8600_));
AOI21X1 AOI21X1_647 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4354_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8611_));
AOI21X1 AOI21X1_648 ( .A(u2__abc_52138_new_n8612_), .B(u2__abc_52138_new_n8589_), .C(rst), .Y(u2__0remHi_451_0__192_));
AOI21X1 AOI21X1_649 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4360_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8619_));
AOI21X1 AOI21X1_65 ( .A(u2__abc_52138_new_n4786_), .B(u2__abc_52138_new_n4683_), .C(u2__abc_52138_new_n4787_), .Y(u2__abc_52138_new_n4788_));
AOI21X1 AOI21X1_650 ( .A(u2__abc_52138_new_n8620_), .B(u2__abc_52138_new_n8614_), .C(rst), .Y(u2__0remHi_451_0__193_));
AOI21X1 AOI21X1_651 ( .A(u2__abc_52138_new_n8615_), .B(u2__abc_52138_new_n4374_), .C(u2__abc_52138_new_n4370_), .Y(u2__abc_52138_new_n8623_));
AOI21X1 AOI21X1_652 ( .A(u2__abc_52138_new_n8625_), .B(u2__abc_52138_new_n8626_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8627_));
AOI21X1 AOI21X1_653 ( .A(u2__abc_52138_new_n4354_), .B(u2__abc_52138_new_n6498_), .C(u2__abc_52138_new_n8627_), .Y(u2__abc_52138_new_n8628_));
AOI21X1 AOI21X1_654 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4349_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8629_));
AOI21X1 AOI21X1_655 ( .A(u2__abc_52138_new_n8630_), .B(u2__abc_52138_new_n8622_), .C(rst), .Y(u2__0remHi_451_0__194_));
AOI21X1 AOI21X1_656 ( .A(u2__abc_52138_new_n4883_), .B(u2__abc_52138_new_n8633_), .C(u2__abc_52138_new_n8634_), .Y(u2__abc_52138_new_n8635_));
AOI21X1 AOI21X1_657 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4344_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8637_));
AOI21X1 AOI21X1_658 ( .A(u2__abc_52138_new_n8638_), .B(u2__abc_52138_new_n8632_), .C(rst), .Y(u2__0remHi_451_0__195_));
AOI21X1 AOI21X1_659 ( .A(u2__abc_52138_new_n4355_), .B(u2__abc_52138_new_n4361_), .C(u2__abc_52138_new_n4881_), .Y(u2__abc_52138_new_n8642_));
AOI21X1 AOI21X1_66 ( .A(u2__abc_52138_new_n4792_), .B(u2__abc_52138_new_n4711_), .C(u2__abc_52138_new_n4798_), .Y(u2__abc_52138_new_n4799_));
AOI21X1 AOI21X1_660 ( .A(u2__abc_52138_new_n8603_), .B(u2__abc_52138_new_n4377_), .C(u2__abc_52138_new_n8643_), .Y(u2__abc_52138_new_n8644_));
AOI21X1 AOI21X1_661 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4333_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8650_));
AOI21X1 AOI21X1_662 ( .A(u2__abc_52138_new_n8651_), .B(u2__abc_52138_new_n8640_), .C(rst), .Y(u2__0remHi_451_0__196_));
AOI21X1 AOI21X1_663 ( .A(u2__abc_52138_new_n8654_), .B(u2__abc_52138_new_n8655_), .C(u2__abc_52138_new_n8656_), .Y(u2__abc_52138_new_n8657_));
AOI21X1 AOI21X1_664 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4338_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8659_));
AOI21X1 AOI21X1_665 ( .A(u2__abc_52138_new_n8660_), .B(u2__abc_52138_new_n8653_), .C(rst), .Y(u2__0remHi_451_0__197_));
AOI21X1 AOI21X1_666 ( .A(u2__abc_52138_new_n8670_), .B(u2__abc_52138_new_n8668_), .C(u2__abc_52138_new_n8671_), .Y(u2__abc_52138_new_n8672_));
AOI21X1 AOI21X1_667 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4302_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8681_));
AOI21X1 AOI21X1_668 ( .A(u2__abc_52138_new_n8682_), .B(u2__abc_52138_new_n8676_), .C(rst), .Y(u2__0remHi_451_0__199_));
AOI21X1 AOI21X1_669 ( .A(u2__abc_52138_new_n8663_), .B(u2__abc_52138_new_n4339_), .C(u2__abc_52138_new_n4892_), .Y(u2__abc_52138_new_n8689_));
AOI21X1 AOI21X1_67 ( .A(u2__abc_52138_new_n4654_), .B(u2__abc_52138_new_n4661_), .C(u2__abc_52138_new_n4656_), .Y(u2__abc_52138_new_n4801_));
AOI21X1 AOI21X1_670 ( .A(u2__abc_52138_new_n8694_), .B(u2__abc_52138_new_n8692_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8695_));
AOI21X1 AOI21X1_671 ( .A(u2__abc_52138_new_n4307_), .B(u2__abc_52138_new_n6498_), .C(u2__abc_52138_new_n8695_), .Y(u2__abc_52138_new_n8696_));
AOI21X1 AOI21X1_672 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4291_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8697_));
AOI21X1 AOI21X1_673 ( .A(u2__abc_52138_new_n8698_), .B(u2__abc_52138_new_n8684_), .C(rst), .Y(u2__0remHi_451_0__200_));
AOI21X1 AOI21X1_674 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4296_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8705_));
AOI21X1 AOI21X1_675 ( .A(u2__abc_52138_new_n8706_), .B(u2__abc_52138_new_n8700_), .C(rst), .Y(u2__0remHi_451_0__201_));
AOI21X1 AOI21X1_676 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4905_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8715_));
AOI21X1 AOI21X1_677 ( .A(u2__abc_52138_new_n8716_), .B(u2__abc_52138_new_n8708_), .C(rst), .Y(u2__0remHi_451_0__202_));
AOI21X1 AOI21X1_678 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4323_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8723_));
AOI21X1 AOI21X1_679 ( .A(u2__abc_52138_new_n8724_), .B(u2__abc_52138_new_n8718_), .C(rst), .Y(u2__0remHi_451_0__203_));
AOI21X1 AOI21X1_68 ( .A(u2__abc_52138_new_n4810_), .B(u2__abc_52138_new_n4625_), .C(u2__abc_52138_new_n4811_), .Y(u2__abc_52138_new_n4812_));
AOI21X1 AOI21X1_680 ( .A(u2__abc_52138_new_n8727_), .B(u2__abc_52138_new_n4299_), .C(u2__abc_52138_new_n8728_), .Y(u2__abc_52138_new_n8729_));
AOI21X1 AOI21X1_681 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4319_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8745_));
AOI21X1 AOI21X1_682 ( .A(u2__abc_52138_new_n8746_), .B(u2__abc_52138_new_n8740_), .C(rst), .Y(u2__0remHi_451_0__205_));
AOI21X1 AOI21X1_683 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4254_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8755_));
AOI21X1 AOI21X1_684 ( .A(u2__abc_52138_new_n8756_), .B(u2__abc_52138_new_n8748_), .C(rst), .Y(u2__0remHi_451_0__206_));
AOI21X1 AOI21X1_685 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4259_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8763_));
AOI21X1 AOI21X1_686 ( .A(u2__abc_52138_new_n8764_), .B(u2__abc_52138_new_n8758_), .C(rst), .Y(u2__0remHi_451_0__207_));
AOI21X1 AOI21X1_687 ( .A(u2__abc_52138_new_n8770_), .B(u2__abc_52138_new_n4322_), .C(u2__abc_52138_new_n8771_), .Y(u2__abc_52138_new_n8772_));
AOI21X1 AOI21X1_688 ( .A(u2__abc_52138_new_n8777_), .B(u2__abc_52138_new_n4256_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n8778_));
AOI21X1 AOI21X1_689 ( .A(u2__abc_52138_new_n8778_), .B(u2__abc_52138_new_n8776_), .C(u2__abc_52138_new_n8779_), .Y(u2__abc_52138_new_n8780_));
AOI21X1 AOI21X1_69 ( .A(u2__abc_52138_new_n4805_), .B(u2__abc_52138_new_n4641_), .C(u2__abc_52138_new_n4813_), .Y(u2__abc_52138_new_n4814_));
AOI21X1 AOI21X1_690 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4248_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8789_));
AOI21X1 AOI21X1_691 ( .A(u2__abc_52138_new_n8790_), .B(u2__abc_52138_new_n8784_), .C(rst), .Y(u2__0remHi_451_0__209_));
AOI21X1 AOI21X1_692 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4280_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8798_));
AOI21X1 AOI21X1_693 ( .A(u2__abc_52138_new_n8799_), .B(u2__abc_52138_new_n8792_), .C(rst), .Y(u2__0remHi_451_0__210_));
AOI21X1 AOI21X1_694 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4275_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8807_));
AOI21X1 AOI21X1_695 ( .A(u2__abc_52138_new_n8808_), .B(u2__abc_52138_new_n8801_), .C(rst), .Y(u2__0remHi_451_0__211_));
AOI21X1 AOI21X1_696 ( .A(u2__abc_52138_new_n8812_), .B(u2__abc_52138_new_n8811_), .C(u2__abc_52138_new_n8813_), .Y(u2__abc_52138_new_n8814_));
AOI21X1 AOI21X1_697 ( .A(u2__abc_52138_new_n8819_), .B(u2__abc_52138_new_n8817_), .C(u2__abc_52138_new_n8820_), .Y(u2__abc_52138_new_n8821_));
AOI21X1 AOI21X1_698 ( .A(u2__abc_52138_new_n4279_), .B(u2__abc_52138_new_n8826_), .C(u2__abc_52138_new_n8827_), .Y(u2__abc_52138_new_n8828_));
AOI21X1 AOI21X1_699 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4269_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8830_));
AOI21X1 AOI21X1_7 ( .A(u2__abc_52138_new_n3084_), .B(u2__abc_52138_new_n3080_), .C(u2__abc_52138_new_n3083_), .Y(u2__abc_52138_new_n3085_));
AOI21X1 AOI21X1_70 ( .A(u2__abc_52138_new_n4815_), .B(u2__abc_52138_new_n4821_), .C(u2__abc_52138_new_n4827_), .Y(u2__abc_52138_new_n4828_));
AOI21X1 AOI21X1_700 ( .A(u2__abc_52138_new_n8831_), .B(u2__abc_52138_new_n8825_), .C(rst), .Y(u2__0remHi_451_0__213_));
AOI21X1 AOI21X1_701 ( .A(u2__abc_52138_new_n4268_), .B(u2__abc_52138_new_n8835_), .C(u2__abc_52138_new_n8836_), .Y(u2__abc_52138_new_n8837_));
AOI21X1 AOI21X1_702 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4207_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8839_));
AOI21X1 AOI21X1_703 ( .A(u2__abc_52138_new_n8840_), .B(u2__abc_52138_new_n8833_), .C(rst), .Y(u2__0remHi_451_0__214_));
AOI21X1 AOI21X1_704 ( .A(u2__abc_52138_new_n8835_), .B(u2__abc_52138_new_n4268_), .C(u2__abc_52138_new_n4265_), .Y(u2__abc_52138_new_n8843_));
AOI21X1 AOI21X1_705 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4212_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8847_));
AOI21X1 AOI21X1_706 ( .A(u2__abc_52138_new_n8848_), .B(u2__abc_52138_new_n8842_), .C(rst), .Y(u2__0remHi_451_0__215_));
AOI21X1 AOI21X1_707 ( .A(u2__abc_52138_new_n4923_), .B(u2__abc_52138_new_n4265_), .C(u2__abc_52138_new_n4270_), .Y(u2__abc_52138_new_n8855_));
AOI21X1 AOI21X1_708 ( .A(u2__abc_52138_new_n8851_), .B(u2__abc_52138_new_n8853_), .C(u2__abc_52138_new_n8856_), .Y(u2__abc_52138_new_n8857_));
AOI21X1 AOI21X1_709 ( .A(u2__abc_52138_new_n8859_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n8860_), .Y(u2__abc_52138_new_n8861_));
AOI21X1 AOI21X1_71 ( .A(u2__abc_52138_new_n4800_), .B(u2__abc_52138_new_n4762_), .C(u2__abc_52138_new_n4829_), .Y(u2__abc_52138_new_n4830_));
AOI21X1 AOI21X1_710 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4201_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8871_));
AOI21X1 AOI21X1_711 ( .A(u2__abc_52138_new_n8872_), .B(u2__abc_52138_new_n8865_), .C(rst), .Y(u2__0remHi_451_0__217_));
AOI21X1 AOI21X1_712 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4235_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8881_));
AOI21X1 AOI21X1_713 ( .A(u2__abc_52138_new_n8882_), .B(u2__abc_52138_new_n8874_), .C(rst), .Y(u2__0remHi_451_0__218_));
AOI21X1 AOI21X1_714 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4228_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8890_));
AOI21X1 AOI21X1_715 ( .A(u2__abc_52138_new_n8891_), .B(u2__abc_52138_new_n8884_), .C(rst), .Y(u2__0remHi_451_0__219_));
AOI21X1 AOI21X1_716 ( .A(u2__abc_52138_new_n8875_), .B(u2__abc_52138_new_n4928_), .C(u2__abc_52138_new_n8896_), .Y(u2__abc_52138_new_n8897_));
AOI21X1 AOI21X1_717 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4219_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8904_));
AOI21X1 AOI21X1_718 ( .A(u2__abc_52138_new_n8905_), .B(u2__abc_52138_new_n8893_), .C(rst), .Y(u2__0remHi_451_0__220_));
AOI21X1 AOI21X1_719 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4224_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8912_));
AOI21X1 AOI21X1_72 ( .A(u2__abc_52138_new_n4544_), .B(u2__abc_52138_new_n4537_), .C(u2__abc_52138_new_n4538_), .Y(u2__abc_52138_new_n4832_));
AOI21X1 AOI21X1_720 ( .A(u2__abc_52138_new_n8913_), .B(u2__abc_52138_new_n8907_), .C(rst), .Y(u2__0remHi_451_0__221_));
AOI21X1 AOI21X1_721 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4164_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8922_));
AOI21X1 AOI21X1_722 ( .A(u2__abc_52138_new_n8923_), .B(u2__abc_52138_new_n8915_), .C(rst), .Y(u2__0remHi_451_0__222_));
AOI21X1 AOI21X1_723 ( .A(u2__abc_52138_new_n8918_), .B(u2__abc_52138_new_n4220_), .C(u2__abc_52138_new_n8926_), .Y(u2__abc_52138_new_n8927_));
AOI21X1 AOI21X1_724 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4159_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8931_));
AOI21X1 AOI21X1_725 ( .A(u2__abc_52138_new_n8932_), .B(u2__abc_52138_new_n8925_), .C(rst), .Y(u2__0remHi_451_0__223_));
AOI21X1 AOI21X1_726 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4148_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8951_));
AOI21X1 AOI21X1_727 ( .A(u2__abc_52138_new_n8952_), .B(u2__abc_52138_new_n8934_), .C(rst), .Y(u2__0remHi_451_0__224_));
AOI21X1 AOI21X1_728 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4153_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8959_));
AOI21X1 AOI21X1_729 ( .A(u2__abc_52138_new_n8960_), .B(u2__abc_52138_new_n8954_), .C(rst), .Y(u2__0remHi_451_0__225_));
AOI21X1 AOI21X1_73 ( .A(u2__abc_52138_new_n4836_), .B(u2__abc_52138_new_n4570_), .C(u2__abc_52138_new_n4843_), .Y(u2__abc_52138_new_n4844_));
AOI21X1 AOI21X1_730 ( .A(u2__abc_52138_new_n8947_), .B(u2__abc_52138_new_n4167_), .C(u2__abc_52138_new_n8963_), .Y(u2__abc_52138_new_n8964_));
AOI21X1 AOI21X1_731 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4185_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8968_));
AOI21X1 AOI21X1_732 ( .A(u2__abc_52138_new_n8969_), .B(u2__abc_52138_new_n8962_), .C(rst), .Y(u2__0remHi_451_0__226_));
AOI21X1 AOI21X1_733 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4180_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8976_));
AOI21X1 AOI21X1_734 ( .A(u2__abc_52138_new_n8977_), .B(u2__abc_52138_new_n8971_), .C(rst), .Y(u2__0remHi_451_0__227_));
AOI21X1 AOI21X1_735 ( .A(u2__abc_52138_new_n8963_), .B(u2__abc_52138_new_n4156_), .C(u2__abc_52138_new_n8980_), .Y(u2__abc_52138_new_n8981_));
AOI21X1 AOI21X1_736 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4176_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n8997_));
AOI21X1 AOI21X1_737 ( .A(u2__abc_52138_new_n8998_), .B(u2__abc_52138_new_n8992_), .C(rst), .Y(u2__0remHi_451_0__229_));
AOI21X1 AOI21X1_738 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4138_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9007_));
AOI21X1 AOI21X1_739 ( .A(u2__abc_52138_new_n9008_), .B(u2__abc_52138_new_n9000_), .C(rst), .Y(u2__0remHi_451_0__230_));
AOI21X1 AOI21X1_74 ( .A(u2__abc_52138_new_n4850_), .B(u2__abc_52138_new_n4755_), .C(u2__abc_52138_new_n4855_), .Y(u2__abc_52138_new_n4856_));
AOI21X1 AOI21X1_740 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4134_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9015_));
AOI21X1 AOI21X1_741 ( .A(u2__abc_52138_new_n9016_), .B(u2__abc_52138_new_n9010_), .C(rst), .Y(u2__0remHi_451_0__231_));
AOI21X1 AOI21X1_742 ( .A(u2__abc_52138_new_n9020_), .B(u2__abc_52138_new_n4177_), .C(u2__abc_52138_new_n4954_), .Y(u2__abc_52138_new_n9021_));
AOI21X1 AOI21X1_743 ( .A(u2__abc_52138_new_n9002_), .B(u2__abc_52138_new_n9019_), .C(u2__abc_52138_new_n9022_), .Y(u2__abc_52138_new_n9023_));
AOI21X1 AOI21X1_744 ( .A(u2__abc_52138_new_n9027_), .B(u2__abc_52138_new_n9025_), .C(u2__abc_52138_new_n9028_), .Y(u2__abc_52138_new_n9029_));
AOI21X1 AOI21X1_745 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4130_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9039_));
AOI21X1 AOI21X1_746 ( .A(u2__abc_52138_new_n9040_), .B(u2__abc_52138_new_n9033_), .C(rst), .Y(u2__0remHi_451_0__233_));
AOI21X1 AOI21X1_747 ( .A(u2__abc_52138_new_n9035_), .B(u2__abc_52138_new_n4137_), .C(u2__abc_52138_new_n4135_), .Y(u2__abc_52138_new_n9043_));
AOI21X1 AOI21X1_748 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4117_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9049_));
AOI21X1 AOI21X1_749 ( .A(u2__abc_52138_new_n9050_), .B(u2__abc_52138_new_n9042_), .C(rst), .Y(u2__0remHi_451_0__234_));
AOI21X1 AOI21X1_75 ( .A(u2__abc_52138_new_n4462_), .B(u2__abc_52138_new_n4859_), .C(u2__abc_52138_new_n4860_), .Y(u2__abc_52138_new_n4861_));
AOI21X1 AOI21X1_750 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4112_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9057_));
AOI21X1 AOI21X1_751 ( .A(u2__abc_52138_new_n9058_), .B(u2__abc_52138_new_n9052_), .C(rst), .Y(u2__0remHi_451_0__235_));
AOI21X1 AOI21X1_752 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4101_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9068_));
AOI21X1 AOI21X1_753 ( .A(u2__abc_52138_new_n9069_), .B(u2__abc_52138_new_n9060_), .C(rst), .Y(u2__0remHi_451_0__236_));
AOI21X1 AOI21X1_754 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4106_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9076_));
AOI21X1 AOI21X1_755 ( .A(u2__abc_52138_new_n9077_), .B(u2__abc_52138_new_n9071_), .C(rst), .Y(u2__0remHi_451_0__237_));
AOI21X1 AOI21X1_756 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4052_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9085_));
AOI21X1 AOI21X1_757 ( .A(u2__abc_52138_new_n9086_), .B(u2__abc_52138_new_n9079_), .C(rst), .Y(u2__0remHi_451_0__238_));
AOI21X1 AOI21X1_758 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4057_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9093_));
AOI21X1 AOI21X1_759 ( .A(u2__abc_52138_new_n9094_), .B(u2__abc_52138_new_n9088_), .C(rst), .Y(u2__0remHi_451_0__239_));
AOI21X1 AOI21X1_76 ( .A(u2__abc_52138_new_n4864_), .B(u2__abc_52138_new_n4439_), .C(u2__abc_52138_new_n4863_), .Y(u2__abc_52138_new_n4865_));
AOI21X1 AOI21X1_760 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4063_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9111_));
AOI21X1 AOI21X1_761 ( .A(u2__abc_52138_new_n9112_), .B(u2__abc_52138_new_n9096_), .C(rst), .Y(u2__0remHi_451_0__240_));
AOI21X1 AOI21X1_762 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4068_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9120_));
AOI21X1 AOI21X1_763 ( .A(u2__abc_52138_new_n9121_), .B(u2__abc_52138_new_n9114_), .C(rst), .Y(u2__0remHi_451_0__241_));
AOI21X1 AOI21X1_764 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4092_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9130_));
AOI21X1 AOI21X1_765 ( .A(u2__abc_52138_new_n9131_), .B(u2__abc_52138_new_n9123_), .C(rst), .Y(u2__0remHi_451_0__242_));
AOI21X1 AOI21X1_766 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4085_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9139_));
AOI21X1 AOI21X1_767 ( .A(u2__abc_52138_new_n9140_), .B(u2__abc_52138_new_n9133_), .C(rst), .Y(u2__0remHi_451_0__243_));
AOI21X1 AOI21X1_768 ( .A(u2__abc_52138_new_n9124_), .B(u2__abc_52138_new_n4071_), .C(u2__abc_52138_new_n9144_), .Y(u2__abc_52138_new_n9145_));
AOI21X1 AOI21X1_769 ( .A(u2__abc_52138_new_n9107_), .B(u2__abc_52138_new_n4073_), .C(u2__abc_52138_new_n9146_), .Y(u2__abc_52138_new_n9147_));
AOI21X1 AOI21X1_77 ( .A(u2__abc_52138_new_n4868_), .B(u2__abc_52138_new_n4403_), .C(u2__abc_52138_new_n4869_), .Y(u2__abc_52138_new_n4870_));
AOI21X1 AOI21X1_770 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4076_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9151_));
AOI21X1 AOI21X1_771 ( .A(u2__abc_52138_new_n9152_), .B(u2__abc_52138_new_n9142_), .C(rst), .Y(u2__0remHi_451_0__244_));
AOI21X1 AOI21X1_772 ( .A(u2__abc_52138_new_n4089_), .B(u2__abc_52138_new_n9155_), .C(u2__abc_52138_new_n9156_), .Y(u2__abc_52138_new_n9157_));
AOI21X1 AOI21X1_773 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4081_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9159_));
AOI21X1 AOI21X1_774 ( .A(u2__abc_52138_new_n9160_), .B(u2__abc_52138_new_n9154_), .C(rst), .Y(u2__0remHi_451_0__245_));
AOI21X1 AOI21X1_775 ( .A(u2__abc_52138_new_n9163_), .B(u2__abc_52138_new_n9165_), .C(u2__abc_52138_new_n9166_), .Y(u2__abc_52138_new_n9167_));
AOI21X1 AOI21X1_776 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4005_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9169_));
AOI21X1 AOI21X1_777 ( .A(u2__abc_52138_new_n9170_), .B(u2__abc_52138_new_n9162_), .C(rst), .Y(u2__0remHi_451_0__246_));
AOI21X1 AOI21X1_778 ( .A(u2__abc_52138_new_n9165_), .B(u2__abc_52138_new_n4077_), .C(u2__abc_52138_new_n9173_), .Y(u2__abc_52138_new_n9174_));
AOI21X1 AOI21X1_779 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4010_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9178_));
AOI21X1 AOI21X1_78 ( .A(u2__abc_52138_new_n4871_), .B(u2__abc_52138_new_n4415_), .C(u2__abc_52138_new_n4873_), .Y(u2__abc_52138_new_n4874_));
AOI21X1 AOI21X1_780 ( .A(u2__abc_52138_new_n9179_), .B(u2__abc_52138_new_n9172_), .C(rst), .Y(u2__0remHi_451_0__247_));
AOI21X1 AOI21X1_781 ( .A(u2__abc_52138_new_n4084_), .B(u2__abc_52138_new_n9183_), .C(u2__abc_52138_new_n9184_), .Y(u2__abc_52138_new_n9185_));
AOI21X1 AOI21X1_782 ( .A(u2__abc_52138_new_n9188_), .B(u2__abc_52138_new_n4007_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n9190_));
AOI21X1 AOI21X1_783 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4016_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9193_));
AOI21X1 AOI21X1_784 ( .A(u2__abc_52138_new_n9194_), .B(u2__abc_52138_new_n9181_), .C(rst), .Y(u2__0remHi_451_0__248_));
AOI21X1 AOI21X1_785 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4021_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9201_));
AOI21X1 AOI21X1_786 ( .A(u2__abc_52138_new_n9202_), .B(u2__abc_52138_new_n9196_), .C(rst), .Y(u2__0remHi_451_0__249_));
AOI21X1 AOI21X1_787 ( .A(u2__abc_52138_new_n9205_), .B(u2__abc_52138_new_n9209_), .C(u2__abc_52138_new_n9210_), .Y(u2__abc_52138_new_n9211_));
AOI21X1 AOI21X1_788 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4044_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9213_));
AOI21X1 AOI21X1_789 ( .A(u2__abc_52138_new_n9214_), .B(u2__abc_52138_new_n9204_), .C(rst), .Y(u2__0remHi_451_0__250_));
AOI21X1 AOI21X1_79 ( .A(u2__abc_52138_new_n4857_), .B(u2__abc_52138_new_n4754_), .C(u2__abc_52138_new_n4877_), .Y(u2__abc_52138_new_n4878_));
AOI21X1 AOI21X1_790 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4039_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9222_));
AOI21X1 AOI21X1_791 ( .A(u2__abc_52138_new_n9223_), .B(u2__abc_52138_new_n9216_), .C(rst), .Y(u2__0remHi_451_0__251_));
AOI21X1 AOI21X1_792 ( .A(u2__abc_52138_new_n9206_), .B(u2__abc_52138_new_n4024_), .C(u2__abc_52138_new_n9227_), .Y(u2__abc_52138_new_n9228_));
AOI21X1 AOI21X1_793 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4028_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9235_));
AOI21X1 AOI21X1_794 ( .A(u2__abc_52138_new_n9236_), .B(u2__abc_52138_new_n9225_), .C(rst), .Y(u2__0remHi_451_0__252_));
AOI21X1 AOI21X1_795 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n4031_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9243_));
AOI21X1 AOI21X1_796 ( .A(u2__abc_52138_new_n9244_), .B(u2__abc_52138_new_n9238_), .C(rst), .Y(u2__0remHi_451_0__253_));
AOI21X1 AOI21X1_797 ( .A(u2__abc_52138_new_n9229_), .B(u2__abc_52138_new_n4047_), .C(u2__abc_52138_new_n9247_), .Y(u2__abc_52138_new_n9248_));
AOI21X1 AOI21X1_798 ( .A(u2__abc_52138_new_n9249_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n9250_), .Y(u2__abc_52138_new_n9251_));
AOI21X1 AOI21X1_799 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5688_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9260_));
AOI21X1 AOI21X1_8 ( .A(u2__abc_52138_new_n3088_), .B(u2__abc_52138_new_n3057_), .C(u2__abc_52138_new_n3089_), .Y(u2__abc_52138_new_n3090_));
AOI21X1 AOI21X1_80 ( .A(u2__abc_52138_new_n4371_), .B(u2__abc_52138_new_n4367_), .C(u2__abc_52138_new_n4373_), .Y(u2__abc_52138_new_n4885_));
AOI21X1 AOI21X1_800 ( .A(u2__abc_52138_new_n9261_), .B(u2__abc_52138_new_n9255_), .C(rst), .Y(u2__0remHi_451_0__255_));
AOI21X1 AOI21X1_801 ( .A(u2__abc_52138_new_n9247_), .B(u2__abc_52138_new_n4036_), .C(u2__abc_52138_new_n9271_), .Y(u2__abc_52138_new_n9272_));
AOI21X1 AOI21X1_802 ( .A(u2__abc_52138_new_n8942_), .B(u2__abc_52138_new_n9267_), .C(u2__abc_52138_new_n9274_), .Y(u2__abc_52138_new_n9275_));
AOI21X1 AOI21X1_803 ( .A(u2__abc_52138_new_n4982_), .B(u2__abc_52138_new_n9186_), .C(u2__abc_52138_new_n9276_), .Y(u2__abc_52138_new_n9277_));
AOI21X1 AOI21X1_804 ( .A(u2__abc_52138_new_n9266_), .B(u2__abc_52138_new_n9278_), .C(u2__abc_52138_new_n9279_), .Y(u2__abc_52138_new_n9280_));
AOI21X1 AOI21X1_805 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5697_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9282_));
AOI21X1 AOI21X1_806 ( .A(u2__abc_52138_new_n9283_), .B(u2__abc_52138_new_n9263_), .C(rst), .Y(u2__0remHi_451_0__256_));
AOI21X1 AOI21X1_807 ( .A(u2__abc_52138_new_n9286_), .B(u2__abc_52138_new_n9289_), .C(u2__abc_52138_new_n9290_), .Y(u2__abc_52138_new_n9291_));
AOI21X1 AOI21X1_808 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5702_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9293_));
AOI21X1 AOI21X1_809 ( .A(u2__abc_52138_new_n9294_), .B(u2__abc_52138_new_n9285_), .C(rst), .Y(u2__0remHi_451_0__257_));
AOI21X1 AOI21X1_81 ( .A(u2__abc_52138_new_n4357_), .B(u2__abc_52138_new_n4359_), .C(u2__abc_52138_new_n4882_), .Y(u2__abc_52138_new_n4886_));
AOI21X1 AOI21X1_810 ( .A(u2__abc_52138_new_n5701_), .B(u2__abc_52138_new_n9298_), .C(u2__abc_52138_new_n9299_), .Y(u2__abc_52138_new_n9300_));
AOI21X1 AOI21X1_811 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5720_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9302_));
AOI21X1 AOI21X1_812 ( .A(u2__abc_52138_new_n9303_), .B(u2__abc_52138_new_n9296_), .C(rst), .Y(u2__0remHi_451_0__258_));
AOI21X1 AOI21X1_813 ( .A(u2__abc_52138_new_n5706_), .B(u2__abc_52138_new_n9308_), .C(u2__abc_52138_new_n9309_), .Y(u2__abc_52138_new_n9310_));
AOI21X1 AOI21X1_814 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5725_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9312_));
AOI21X1 AOI21X1_815 ( .A(u2__abc_52138_new_n9313_), .B(u2__abc_52138_new_n9305_), .C(rst), .Y(u2__0remHi_451_0__259_));
AOI21X1 AOI21X1_816 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5709_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9327_));
AOI21X1 AOI21X1_817 ( .A(u2__abc_52138_new_n9328_), .B(u2__abc_52138_new_n9315_), .C(rst), .Y(u2__0remHi_451_0__260_));
AOI21X1 AOI21X1_818 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5714_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9335_));
AOI21X1 AOI21X1_819 ( .A(u2__abc_52138_new_n9336_), .B(u2__abc_52138_new_n9330_), .C(rst), .Y(u2__0remHi_451_0__261_));
AOI21X1 AOI21X1_82 ( .A(u2__abc_52138_new_n4887_), .B(u2__abc_52138_new_n4353_), .C(u2__abc_52138_new_n4895_), .Y(u2__abc_52138_new_n4896_));
AOI21X1 AOI21X1_820 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5676_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9347_));
AOI21X1 AOI21X1_821 ( .A(u2__abc_52138_new_n9348_), .B(u2__abc_52138_new_n9338_), .C(rst), .Y(u2__0remHi_451_0__262_));
AOI21X1 AOI21X1_822 ( .A(u2__abc_52138_new_n5718_), .B(u2__abc_52138_new_n9352_), .C(u2__abc_52138_new_n9353_), .Y(u2__abc_52138_new_n9354_));
AOI21X1 AOI21X1_823 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5681_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9356_));
AOI21X1 AOI21X1_824 ( .A(u2__abc_52138_new_n9357_), .B(u2__abc_52138_new_n9350_), .C(rst), .Y(u2__0remHi_451_0__263_));
AOI21X1 AOI21X1_825 ( .A(u2__abc_52138_new_n5718_), .B(u2__abc_52138_new_n5710_), .C(u2__abc_52138_new_n5715_), .Y(u2__abc_52138_new_n9361_));
AOI21X1 AOI21X1_826 ( .A(u2__abc_52138_new_n5731_), .B(u2__abc_52138_new_n9319_), .C(u2__abc_52138_new_n9362_), .Y(u2__abc_52138_new_n9363_));
AOI21X1 AOI21X1_827 ( .A(u2__abc_52138_new_n5678_), .B(u2__abc_52138_new_n9364_), .C(u2__abc_52138_new_n9365_), .Y(u2__abc_52138_new_n9366_));
AOI21X1 AOI21X1_828 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5663_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9368_));
AOI21X1 AOI21X1_829 ( .A(u2__abc_52138_new_n9369_), .B(u2__abc_52138_new_n9359_), .C(rst), .Y(u2__0remHi_451_0__264_));
AOI21X1 AOI21X1_83 ( .A(u2__abc_52138_new_n4897_), .B(u2__abc_52138_new_n4903_), .C(u2__abc_52138_new_n4911_), .Y(u2__abc_52138_new_n4912_));
AOI21X1 AOI21X1_830 ( .A(u2__abc_52138_new_n5683_), .B(u2__abc_52138_new_n9374_), .C(u2__abc_52138_new_n9375_), .Y(u2__abc_52138_new_n9376_));
AOI21X1 AOI21X1_831 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5668_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9378_));
AOI21X1 AOI21X1_832 ( .A(u2__abc_52138_new_n9379_), .B(u2__abc_52138_new_n9371_), .C(rst), .Y(u2__0remHi_451_0__265_));
AOI21X1 AOI21X1_833 ( .A(u2__abc_52138_new_n5683_), .B(u2__abc_52138_new_n5677_), .C(u2__abc_52138_new_n5682_), .Y(u2__abc_52138_new_n9382_));
AOI21X1 AOI21X1_834 ( .A(u2__abc_52138_new_n5667_), .B(u2__abc_52138_new_n9383_), .C(u2__abc_52138_new_n9384_), .Y(u2__abc_52138_new_n9385_));
AOI21X1 AOI21X1_835 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5651_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9387_));
AOI21X1 AOI21X1_836 ( .A(u2__abc_52138_new_n9388_), .B(u2__abc_52138_new_n9381_), .C(rst), .Y(u2__0remHi_451_0__266_));
AOI21X1 AOI21X1_837 ( .A(u2__abc_52138_new_n5672_), .B(u2__abc_52138_new_n9392_), .C(u2__abc_52138_new_n9393_), .Y(u2__abc_52138_new_n9394_));
AOI21X1 AOI21X1_838 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5656_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9396_));
AOI21X1 AOI21X1_839 ( .A(u2__abc_52138_new_n9397_), .B(u2__abc_52138_new_n9390_), .C(rst), .Y(u2__0remHi_451_0__267_));
AOI21X1 AOI21X1_84 ( .A(u2__abc_52138_new_n4914_), .B(u2__abc_52138_new_n4258_), .C(u2__abc_52138_new_n4915_), .Y(u2__abc_52138_new_n4916_));
AOI21X1 AOI21X1_840 ( .A(u2__abc_52138_new_n9391_), .B(u2__abc_52138_new_n9400_), .C(u2__abc_52138_new_n5671_), .Y(u2__abc_52138_new_n9401_));
AOI21X1 AOI21X1_841 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5642_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9406_));
AOI21X1 AOI21X1_842 ( .A(u2__abc_52138_new_n9407_), .B(u2__abc_52138_new_n9399_), .C(rst), .Y(u2__0remHi_451_0__268_));
AOI21X1 AOI21X1_843 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5647_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9414_));
AOI21X1 AOI21X1_844 ( .A(u2__abc_52138_new_n9415_), .B(u2__abc_52138_new_n9409_), .C(rst), .Y(u2__0remHi_451_0__269_));
AOI21X1 AOI21X1_845 ( .A(u2__abc_52138_new_n5644_), .B(u2__abc_52138_new_n9422_), .C(u2__abc_52138_new_n9423_), .Y(u2__abc_52138_new_n9424_));
AOI21X1 AOI21X1_846 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5606_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9426_));
AOI21X1 AOI21X1_847 ( .A(u2__abc_52138_new_n9427_), .B(u2__abc_52138_new_n9417_), .C(rst), .Y(u2__0remHi_451_0__270_));
AOI21X1 AOI21X1_848 ( .A(u2__abc_52138_new_n5649_), .B(u2__abc_52138_new_n9431_), .C(u2__abc_52138_new_n9432_), .Y(u2__abc_52138_new_n9433_));
AOI21X1 AOI21X1_849 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5611_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9435_));
AOI21X1 AOI21X1_85 ( .A(u2__abc_52138_new_n4917_), .B(u2__abc_52138_new_n4247_), .C(u2__abc_52138_new_n4918_), .Y(u2__abc_52138_new_n4919_));
AOI21X1 AOI21X1_850 ( .A(u2__abc_52138_new_n9436_), .B(u2__abc_52138_new_n9429_), .C(rst), .Y(u2__0remHi_451_0__271_));
AOI21X1 AOI21X1_851 ( .A(u2__abc_52138_new_n5649_), .B(u2__abc_52138_new_n5643_), .C(u2__abc_52138_new_n5648_), .Y(u2__abc_52138_new_n9440_));
AOI21X1 AOI21X1_852 ( .A(u2__abc_52138_new_n9439_), .B(u2__abc_52138_new_n5662_), .C(u2__abc_52138_new_n9442_), .Y(u2__abc_52138_new_n9443_));
AOI21X1 AOI21X1_853 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5595_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9453_));
AOI21X1 AOI21X1_854 ( .A(u2__abc_52138_new_n9454_), .B(u2__abc_52138_new_n9438_), .C(rst), .Y(u2__0remHi_451_0__272_));
AOI21X1 AOI21X1_855 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5600_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9461_));
AOI21X1 AOI21X1_856 ( .A(u2__abc_52138_new_n9462_), .B(u2__abc_52138_new_n9456_), .C(rst), .Y(u2__0remHi_451_0__273_));
AOI21X1 AOI21X1_857 ( .A(u2__abc_52138_new_n5599_), .B(u2__abc_52138_new_n9467_), .C(u2__abc_52138_new_n9468_), .Y(u2__abc_52138_new_n9469_));
AOI21X1 AOI21X1_858 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n9471_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9472_));
AOI21X1 AOI21X1_859 ( .A(u2__abc_52138_new_n9473_), .B(u2__abc_52138_new_n9464_), .C(rst), .Y(u2__0remHi_451_0__274_));
AOI21X1 AOI21X1_86 ( .A(u2__abc_52138_new_n4921_), .B(u2__abc_52138_new_n4283_), .C(u2__abc_52138_new_n4278_), .Y(u2__abc_52138_new_n4922_));
AOI21X1 AOI21X1_860 ( .A(u2__abc_52138_new_n5604_), .B(u2__abc_52138_new_n9477_), .C(u2__abc_52138_new_n9478_), .Y(u2__abc_52138_new_n9479_));
AOI21X1 AOI21X1_861 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5630_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9481_));
AOI21X1 AOI21X1_862 ( .A(u2__abc_52138_new_n9482_), .B(u2__abc_52138_new_n9475_), .C(rst), .Y(u2__0remHi_451_0__275_));
AOI21X1 AOI21X1_863 ( .A(u2__abc_52138_new_n5604_), .B(u2__abc_52138_new_n5596_), .C(u2__abc_52138_new_n5601_), .Y(u2__abc_52138_new_n9486_));
AOI21X1 AOI21X1_864 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5618_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9496_));
AOI21X1 AOI21X1_865 ( .A(u2__abc_52138_new_n9497_), .B(u2__abc_52138_new_n9484_), .C(rst), .Y(u2__0remHi_451_0__276_));
AOI21X1 AOI21X1_866 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5623_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9504_));
AOI21X1 AOI21X1_867 ( .A(u2__abc_52138_new_n9505_), .B(u2__abc_52138_new_n9499_), .C(rst), .Y(u2__0remHi_451_0__277_));
AOI21X1 AOI21X1_868 ( .A(u2__abc_52138_new_n5622_), .B(u2__abc_52138_new_n9511_), .C(u2__abc_52138_new_n9512_), .Y(u2__abc_52138_new_n9513_));
AOI21X1 AOI21X1_869 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5559_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9515_));
AOI21X1 AOI21X1_87 ( .A(u2__abc_52138_new_n4920_), .B(u2__abc_52138_new_n4286_), .C(u2__abc_52138_new_n4926_), .Y(u2__abc_52138_new_n4927_));
AOI21X1 AOI21X1_870 ( .A(u2__abc_52138_new_n9516_), .B(u2__abc_52138_new_n9507_), .C(rst), .Y(u2__0remHi_451_0__278_));
AOI21X1 AOI21X1_871 ( .A(u2__abc_52138_new_n5627_), .B(u2__abc_52138_new_n9520_), .C(u2__abc_52138_new_n9521_), .Y(u2__abc_52138_new_n9522_));
AOI21X1 AOI21X1_872 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5564_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9524_));
AOI21X1 AOI21X1_873 ( .A(u2__abc_52138_new_n9525_), .B(u2__abc_52138_new_n9518_), .C(rst), .Y(u2__0remHi_451_0__279_));
AOI21X1 AOI21X1_874 ( .A(u2__abc_52138_new_n5627_), .B(u2__abc_52138_new_n5619_), .C(u2__abc_52138_new_n5624_), .Y(u2__abc_52138_new_n9529_));
AOI21X1 AOI21X1_875 ( .A(u2__abc_52138_new_n9488_), .B(u2__abc_52138_new_n5636_), .C(u2__abc_52138_new_n9530_), .Y(u2__abc_52138_new_n9531_));
AOI21X1 AOI21X1_876 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5548_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9538_));
AOI21X1 AOI21X1_877 ( .A(u2__abc_52138_new_n9539_), .B(u2__abc_52138_new_n9527_), .C(rst), .Y(u2__0remHi_451_0__280_));
AOI21X1 AOI21X1_878 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5553_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9546_));
AOI21X1 AOI21X1_879 ( .A(u2__abc_52138_new_n9547_), .B(u2__abc_52138_new_n9541_), .C(rst), .Y(u2__0remHi_451_0__281_));
AOI21X1 AOI21X1_88 ( .A(u2__abc_52138_new_n4934_), .B(u2__abc_52138_new_n4938_), .C(u2__abc_52138_new_n4936_), .Y(u2__abc_52138_new_n4939_));
AOI21X1 AOI21X1_880 ( .A(u2__abc_52138_new_n5552_), .B(u2__abc_52138_new_n9552_), .C(u2__abc_52138_new_n9553_), .Y(u2__abc_52138_new_n9554_));
AOI21X1 AOI21X1_881 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5582_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9556_));
AOI21X1 AOI21X1_882 ( .A(u2__abc_52138_new_n9557_), .B(u2__abc_52138_new_n9549_), .C(rst), .Y(u2__0remHi_451_0__282_));
AOI21X1 AOI21X1_883 ( .A(u2__abc_52138_new_n5557_), .B(u2__abc_52138_new_n9561_), .C(u2__abc_52138_new_n9562_), .Y(u2__abc_52138_new_n9563_));
AOI21X1 AOI21X1_884 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5587_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9565_));
AOI21X1 AOI21X1_885 ( .A(u2__abc_52138_new_n9566_), .B(u2__abc_52138_new_n9559_), .C(rst), .Y(u2__0remHi_451_0__283_));
AOI21X1 AOI21X1_886 ( .A(u2__abc_52138_new_n9532_), .B(u2__abc_52138_new_n5570_), .C(u2__abc_52138_new_n9572_), .Y(u2__abc_52138_new_n9573_));
AOI21X1 AOI21X1_887 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5571_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9580_));
AOI21X1 AOI21X1_888 ( .A(u2__abc_52138_new_n9581_), .B(u2__abc_52138_new_n9568_), .C(rst), .Y(u2__0remHi_451_0__284_));
AOI21X1 AOI21X1_889 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5576_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9589_));
AOI21X1 AOI21X1_89 ( .A(u2__abc_52138_new_n4933_), .B(u2__abc_52138_new_n4239_), .C(u2__abc_52138_new_n4940_), .Y(u2__abc_52138_new_n4941_));
AOI21X1 AOI21X1_890 ( .A(u2__abc_52138_new_n9590_), .B(u2__abc_52138_new_n9583_), .C(rst), .Y(u2__0remHi_451_0__285_));
AOI21X1 AOI21X1_891 ( .A(u2__abc_52138_new_n5575_), .B(u2__abc_52138_new_n9596_), .C(u2__abc_52138_new_n9597_), .Y(u2__abc_52138_new_n9598_));
AOI21X1 AOI21X1_892 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5513_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9600_));
AOI21X1 AOI21X1_893 ( .A(u2__abc_52138_new_n9601_), .B(u2__abc_52138_new_n9592_), .C(rst), .Y(u2__0remHi_451_0__286_));
AOI21X1 AOI21X1_894 ( .A(u2__abc_52138_new_n5580_), .B(u2__abc_52138_new_n9605_), .C(u2__abc_52138_new_n9606_), .Y(u2__abc_52138_new_n9607_));
AOI21X1 AOI21X1_895 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5518_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9609_));
AOI21X1 AOI21X1_896 ( .A(u2__abc_52138_new_n9610_), .B(u2__abc_52138_new_n9603_), .C(rst), .Y(u2__0remHi_451_0__287_));
AOI21X1 AOI21X1_897 ( .A(u2__abc_52138_new_n5593_), .B(u2__abc_52138_new_n9572_), .C(u2__abc_52138_new_n9616_), .Y(u2__abc_52138_new_n9617_));
AOI21X1 AOI21X1_898 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5502_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9628_));
AOI21X1 AOI21X1_899 ( .A(u2__abc_52138_new_n9629_), .B(u2__abc_52138_new_n9612_), .C(rst), .Y(u2__0remHi_451_0__288_));
AOI21X1 AOI21X1_9 ( .A(u2__abc_52138_new_n3065_), .B(u2__abc_52138_new_n3078_), .C(u2__abc_52138_new_n3091_), .Y(u2__abc_52138_new_n3092_));
AOI21X1 AOI21X1_90 ( .A(u2__abc_52138_new_n4913_), .B(u2__abc_52138_new_n4288_), .C(u2__abc_52138_new_n4942_), .Y(u2__abc_52138_new_n4943_));
AOI21X1 AOI21X1_900 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5507_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9636_));
AOI21X1 AOI21X1_901 ( .A(u2__abc_52138_new_n9637_), .B(u2__abc_52138_new_n9631_), .C(rst), .Y(u2__0remHi_451_0__289_));
AOI21X1 AOI21X1_902 ( .A(u2__abc_52138_new_n5506_), .B(u2__abc_52138_new_n9642_), .C(u2__abc_52138_new_n9643_), .Y(u2__abc_52138_new_n9644_));
AOI21X1 AOI21X1_903 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n9646_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9647_));
AOI21X1 AOI21X1_904 ( .A(u2__abc_52138_new_n9648_), .B(u2__abc_52138_new_n9639_), .C(rst), .Y(u2__0remHi_451_0__290_));
AOI21X1 AOI21X1_905 ( .A(u2__abc_52138_new_n5511_), .B(u2__abc_52138_new_n9652_), .C(u2__abc_52138_new_n9653_), .Y(u2__abc_52138_new_n9654_));
AOI21X1 AOI21X1_906 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5537_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9656_));
AOI21X1 AOI21X1_907 ( .A(u2__abc_52138_new_n9657_), .B(u2__abc_52138_new_n9650_), .C(rst), .Y(u2__0remHi_451_0__291_));
AOI21X1 AOI21X1_908 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5525_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9672_));
AOI21X1 AOI21X1_909 ( .A(u2__abc_52138_new_n9673_), .B(u2__abc_52138_new_n9659_), .C(rst), .Y(u2__0remHi_451_0__292_));
AOI21X1 AOI21X1_91 ( .A(u2__abc_52138_new_n4944_), .B(u2__abc_52138_new_n4950_), .C(u2__abc_52138_new_n4957_), .Y(u2__abc_52138_new_n4958_));
AOI21X1 AOI21X1_910 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5530_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9680_));
AOI21X1 AOI21X1_911 ( .A(u2__abc_52138_new_n9681_), .B(u2__abc_52138_new_n9675_), .C(rst), .Y(u2__0remHi_451_0__293_));
AOI21X1 AOI21X1_912 ( .A(u2__abc_52138_new_n5529_), .B(u2__abc_52138_new_n9687_), .C(u2__abc_52138_new_n9688_), .Y(u2__abc_52138_new_n9689_));
AOI21X1 AOI21X1_913 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5457_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9691_));
AOI21X1 AOI21X1_914 ( .A(u2__abc_52138_new_n9692_), .B(u2__abc_52138_new_n9683_), .C(rst), .Y(u2__0remHi_451_0__294_));
AOI21X1 AOI21X1_915 ( .A(u2__abc_52138_new_n5534_), .B(u2__abc_52138_new_n9696_), .C(u2__abc_52138_new_n9697_), .Y(u2__abc_52138_new_n9698_));
AOI21X1 AOI21X1_916 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5460_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9700_));
AOI21X1 AOI21X1_917 ( .A(u2__abc_52138_new_n9701_), .B(u2__abc_52138_new_n9694_), .C(rst), .Y(u2__0remHi_451_0__295_));
AOI21X1 AOI21X1_918 ( .A(u2__abc_52138_new_n5534_), .B(u2__abc_52138_new_n5526_), .C(u2__abc_52138_new_n5531_), .Y(u2__abc_52138_new_n9705_));
AOI21X1 AOI21X1_919 ( .A(u2__abc_52138_new_n9664_), .B(u2__abc_52138_new_n5543_), .C(u2__abc_52138_new_n9706_), .Y(u2__abc_52138_new_n9707_));
AOI21X1 AOI21X1_92 ( .A(u2__abc_52138_new_n4962_), .B(u2__abc_52138_new_n4959_), .C(u2__abc_52138_new_n4963_), .Y(u2__abc_52138_new_n4964_));
AOI21X1 AOI21X1_920 ( .A(u2__abc_52138_new_n5459_), .B(u2__abc_52138_new_n9708_), .C(u2__abc_52138_new_n9709_), .Y(u2__abc_52138_new_n9710_));
AOI21X1 AOI21X1_921 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5466_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9712_));
AOI21X1 AOI21X1_922 ( .A(u2__abc_52138_new_n9713_), .B(u2__abc_52138_new_n9703_), .C(rst), .Y(u2__0remHi_451_0__296_));
AOI21X1 AOI21X1_923 ( .A(u2__abc_52138_new_n5464_), .B(u2__abc_52138_new_n9718_), .C(u2__abc_52138_new_n9719_), .Y(u2__abc_52138_new_n9720_));
AOI21X1 AOI21X1_924 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5471_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9722_));
AOI21X1 AOI21X1_925 ( .A(u2__abc_52138_new_n9723_), .B(u2__abc_52138_new_n9715_), .C(rst), .Y(u2__0remHi_451_0__297_));
AOI21X1 AOI21X1_926 ( .A(u2__abc_52138_new_n5470_), .B(u2__abc_52138_new_n9728_), .C(u2__abc_52138_new_n9729_), .Y(u2__abc_52138_new_n9730_));
AOI21X1 AOI21X1_927 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5489_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9732_));
AOI21X1 AOI21X1_928 ( .A(u2__abc_52138_new_n9733_), .B(u2__abc_52138_new_n9725_), .C(rst), .Y(u2__0remHi_451_0__298_));
AOI21X1 AOI21X1_929 ( .A(u2__abc_52138_new_n5475_), .B(u2__abc_52138_new_n9737_), .C(u2__abc_52138_new_n9738_), .Y(u2__abc_52138_new_n9739_));
AOI21X1 AOI21X1_93 ( .A(u2__abc_52138_new_n4965_), .B(u2__abc_52138_new_n4109_), .C(u2__abc_52138_new_n4966_), .Y(u2__abc_52138_new_n4967_));
AOI21X1 AOI21X1_930 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5494_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9741_));
AOI21X1 AOI21X1_931 ( .A(u2__abc_52138_new_n9742_), .B(u2__abc_52138_new_n9735_), .C(rst), .Y(u2__0remHi_451_0__299_));
AOI21X1 AOI21X1_932 ( .A(u2__abc_52138_new_n5475_), .B(u2__abc_52138_new_n5467_), .C(u2__abc_52138_new_n5472_), .Y(u2__abc_52138_new_n9745_));
AOI21X1 AOI21X1_933 ( .A(u2__abc_52138_new_n9708_), .B(u2__abc_52138_new_n5477_), .C(u2__abc_52138_new_n9746_), .Y(u2__abc_52138_new_n9747_));
AOI21X1 AOI21X1_934 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5478_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9754_));
AOI21X1 AOI21X1_935 ( .A(u2__abc_52138_new_n9755_), .B(u2__abc_52138_new_n9744_), .C(rst), .Y(u2__0remHi_451_0__300_));
AOI21X1 AOI21X1_936 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5483_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9762_));
AOI21X1 AOI21X1_937 ( .A(u2__abc_52138_new_n9763_), .B(u2__abc_52138_new_n9757_), .C(rst), .Y(u2__0remHi_451_0__301_));
AOI21X1 AOI21X1_938 ( .A(u2__abc_52138_new_n5482_), .B(u2__abc_52138_new_n9770_), .C(u2__abc_52138_new_n9771_), .Y(u2__abc_52138_new_n9772_));
AOI21X1 AOI21X1_939 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5409_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9774_));
AOI21X1 AOI21X1_94 ( .A(u2__abc_52138_new_n4978_), .B(u2__abc_52138_new_n4036_), .C(u2__abc_52138_new_n4977_), .Y(u2__abc_52138_new_n4979_));
AOI21X1 AOI21X1_940 ( .A(u2__abc_52138_new_n9775_), .B(u2__abc_52138_new_n9765_), .C(rst), .Y(u2__0remHi_451_0__302_));
AOI21X1 AOI21X1_941 ( .A(u2__abc_52138_new_n5487_), .B(u2__abc_52138_new_n9779_), .C(u2__abc_52138_new_n9780_), .Y(u2__abc_52138_new_n9781_));
AOI21X1 AOI21X1_942 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5414_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9783_));
AOI21X1 AOI21X1_943 ( .A(u2__abc_52138_new_n9784_), .B(u2__abc_52138_new_n9777_), .C(rst), .Y(u2__0remHi_451_0__303_));
AOI21X1 AOI21X1_944 ( .A(u2__abc_52138_new_n5487_), .B(u2__abc_52138_new_n5479_), .C(u2__abc_52138_new_n5484_), .Y(u2__abc_52138_new_n9790_));
AOI21X1 AOI21X1_945 ( .A(u2__abc_52138_new_n5411_), .B(u2__abc_52138_new_n9794_), .C(u2__abc_52138_new_n9795_), .Y(u2__abc_52138_new_n9796_));
AOI21X1 AOI21X1_946 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5418_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9798_));
AOI21X1 AOI21X1_947 ( .A(u2__abc_52138_new_n9799_), .B(u2__abc_52138_new_n9786_), .C(rst), .Y(u2__0remHi_451_0__304_));
AOI21X1 AOI21X1_948 ( .A(u2__abc_52138_new_n5416_), .B(u2__abc_52138_new_n9804_), .C(u2__abc_52138_new_n9805_), .Y(u2__abc_52138_new_n9806_));
AOI21X1 AOI21X1_949 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5423_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9808_));
AOI21X1 AOI21X1_95 ( .A(u2__abc_52138_new_n4976_), .B(u2__abc_52138_new_n4971_), .C(u2__abc_52138_new_n4980_), .Y(u2__abc_52138_new_n4981_));
AOI21X1 AOI21X1_950 ( .A(u2__abc_52138_new_n9809_), .B(u2__abc_52138_new_n9801_), .C(rst), .Y(u2__0remHi_451_0__305_));
AOI21X1 AOI21X1_951 ( .A(u2__abc_52138_new_n5416_), .B(u2__abc_52138_new_n5410_), .C(u2__abc_52138_new_n5415_), .Y(u2__abc_52138_new_n9812_));
AOI21X1 AOI21X1_952 ( .A(u2__abc_52138_new_n5422_), .B(u2__abc_52138_new_n9813_), .C(u2__abc_52138_new_n9814_), .Y(u2__abc_52138_new_n9815_));
AOI21X1 AOI21X1_953 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5446_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9817_));
AOI21X1 AOI21X1_954 ( .A(u2__abc_52138_new_n9818_), .B(u2__abc_52138_new_n9811_), .C(rst), .Y(u2__0remHi_451_0__306_));
AOI21X1 AOI21X1_955 ( .A(u2__abc_52138_new_n5427_), .B(u2__abc_52138_new_n9822_), .C(u2__abc_52138_new_n9823_), .Y(u2__abc_52138_new_n9824_));
AOI21X1 AOI21X1_956 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5441_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9826_));
AOI21X1 AOI21X1_957 ( .A(u2__abc_52138_new_n9827_), .B(u2__abc_52138_new_n9820_), .C(rst), .Y(u2__0remHi_451_0__307_));
AOI21X1 AOI21X1_958 ( .A(u2__abc_52138_new_n5427_), .B(u2__abc_52138_new_n5419_), .C(u2__abc_52138_new_n5424_), .Y(u2__abc_52138_new_n9831_));
AOI21X1 AOI21X1_959 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5430_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9840_));
AOI21X1 AOI21X1_96 ( .A(u2__abc_52138_new_n4984_), .B(u2__abc_52138_new_n4071_), .C(u2__abc_52138_new_n4985_), .Y(u2__abc_52138_new_n4986_));
AOI21X1 AOI21X1_960 ( .A(u2__abc_52138_new_n9841_), .B(u2__abc_52138_new_n9829_), .C(rst), .Y(u2__0remHi_451_0__308_));
AOI21X1 AOI21X1_961 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5435_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9850_));
AOI21X1 AOI21X1_962 ( .A(u2__abc_52138_new_n9851_), .B(u2__abc_52138_new_n9843_), .C(rst), .Y(u2__0remHi_451_0__309_));
AOI21X1 AOI21X1_963 ( .A(u2__abc_52138_new_n5434_), .B(u2__abc_52138_new_n9854_), .C(u2__abc_52138_new_n9855_), .Y(u2__abc_52138_new_n9856_));
AOI21X1 AOI21X1_964 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n9858_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9859_));
AOI21X1 AOI21X1_965 ( .A(u2__abc_52138_new_n9860_), .B(u2__abc_52138_new_n9853_), .C(rst), .Y(u2__0remHi_451_0__310_));
AOI21X1 AOI21X1_966 ( .A(u2__abc_52138_new_n5439_), .B(u2__abc_52138_new_n9864_), .C(u2__abc_52138_new_n9865_), .Y(u2__abc_52138_new_n9866_));
AOI21X1 AOI21X1_967 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5380_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9868_));
AOI21X1 AOI21X1_968 ( .A(u2__abc_52138_new_n9869_), .B(u2__abc_52138_new_n9862_), .C(rst), .Y(u2__0remHi_451_0__311_));
AOI21X1 AOI21X1_969 ( .A(u2__abc_52138_new_n5445_), .B(u2__abc_52138_new_n5447_), .C(u2__abc_52138_new_n5442_), .Y(u2__abc_52138_new_n9872_));
AOI21X1 AOI21X1_97 ( .A(u2__abc_52138_new_n4084_), .B(u2__abc_52138_new_n4990_), .C(u2__abc_52138_new_n4988_), .Y(u2__abc_52138_new_n4991_));
AOI21X1 AOI21X1_970 ( .A(u2__abc_52138_new_n5439_), .B(u2__abc_52138_new_n5431_), .C(u2__abc_52138_new_n5436_), .Y(u2__abc_52138_new_n9873_));
AOI21X1 AOI21X1_971 ( .A(u2__abc_52138_new_n5452_), .B(u2__abc_52138_new_n9832_), .C(u2__abc_52138_new_n9874_), .Y(u2__abc_52138_new_n9875_));
AOI21X1 AOI21X1_972 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5368_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9882_));
AOI21X1 AOI21X1_973 ( .A(u2__abc_52138_new_n9883_), .B(u2__abc_52138_new_n9871_), .C(rst), .Y(u2__0remHi_451_0__312_));
AOI21X1 AOI21X1_974 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5373_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9890_));
AOI21X1 AOI21X1_975 ( .A(u2__abc_52138_new_n9891_), .B(u2__abc_52138_new_n9885_), .C(rst), .Y(u2__0remHi_451_0__313_));
AOI21X1 AOI21X1_976 ( .A(u2__abc_52138_new_n5372_), .B(u2__abc_52138_new_n9897_), .C(u2__abc_52138_new_n9898_), .Y(u2__abc_52138_new_n9899_));
AOI21X1 AOI21X1_977 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5818_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9901_));
AOI21X1 AOI21X1_978 ( .A(u2__abc_52138_new_n9902_), .B(u2__abc_52138_new_n9893_), .C(rst), .Y(u2__0remHi_451_0__314_));
AOI21X1 AOI21X1_979 ( .A(u2__abc_52138_new_n5377_), .B(u2__abc_52138_new_n9906_), .C(u2__abc_52138_new_n9907_), .Y(u2__abc_52138_new_n9908_));
AOI21X1 AOI21X1_98 ( .A(u2__abc_52138_new_n4970_), .B(u2__abc_52138_new_n4098_), .C(u2__abc_52138_new_n4994_), .Y(u2__abc_52138_new_n4995_));
AOI21X1 AOI21X1_980 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5399_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9910_));
AOI21X1 AOI21X1_981 ( .A(u2__abc_52138_new_n9911_), .B(u2__abc_52138_new_n9904_), .C(rst), .Y(u2__0remHi_451_0__315_));
AOI21X1 AOI21X1_982 ( .A(u2__abc_52138_new_n5810_), .B(u2__abc_52138_new_n5369_), .C(u2__abc_52138_new_n5374_), .Y(u2__abc_52138_new_n9915_));
AOI21X1 AOI21X1_983 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5387_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9925_));
AOI21X1 AOI21X1_984 ( .A(u2__abc_52138_new_n9926_), .B(u2__abc_52138_new_n9913_), .C(rst), .Y(u2__0remHi_451_0__316_));
AOI21X1 AOI21X1_985 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5392_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9933_));
AOI21X1 AOI21X1_986 ( .A(u2__abc_52138_new_n9934_), .B(u2__abc_52138_new_n9928_), .C(rst), .Y(u2__0remHi_451_0__317_));
AOI21X1 AOI21X1_987 ( .A(u2__abc_52138_new_n5391_), .B(u2__abc_52138_new_n9940_), .C(u2__abc_52138_new_n9941_), .Y(u2__abc_52138_new_n9942_));
AOI21X1 AOI21X1_988 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5343_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9944_));
AOI21X1 AOI21X1_989 ( .A(u2__abc_52138_new_n9945_), .B(u2__abc_52138_new_n9936_), .C(rst), .Y(u2__0remHi_451_0__318_));
AOI21X1 AOI21X1_99 ( .A(u2__abc_52138_new_n4879_), .B(u2__abc_52138_new_n4381_), .C(u2__abc_52138_new_n4996_), .Y(u2__abc_52138_new_n4997_));
AOI21X1 AOI21X1_990 ( .A(u2__abc_52138_new_n5396_), .B(u2__abc_52138_new_n9949_), .C(u2__abc_52138_new_n9950_), .Y(u2__abc_52138_new_n9951_));
AOI21X1 AOI21X1_991 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5346_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9953_));
AOI21X1 AOI21X1_992 ( .A(u2__abc_52138_new_n9954_), .B(u2__abc_52138_new_n9947_), .C(rst), .Y(u2__0remHi_451_0__319_));
AOI21X1 AOI21X1_993 ( .A(u2__abc_52138_new_n9960_), .B(u2__abc_52138_new_n9938_), .C(u2__abc_52138_new_n9961_), .Y(u2__abc_52138_new_n9962_));
AOI21X1 AOI21X1_994 ( .A(u2__abc_52138_new_n9959_), .B(u2__abc_52138_new_n5454_), .C(u2__abc_52138_new_n9963_), .Y(u2__abc_52138_new_n9964_));
AOI21X1 AOI21X1_995 ( .A(u2__abc_52138_new_n5345_), .B(u2__abc_52138_new_n9968_), .C(u2__abc_52138_new_n9969_), .Y(u2__abc_52138_new_n9970_));
AOI21X1 AOI21X1_996 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5352_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9972_));
AOI21X1 AOI21X1_997 ( .A(u2__abc_52138_new_n9973_), .B(u2__abc_52138_new_n9956_), .C(rst), .Y(u2__0remHi_451_0__320_));
AOI21X1 AOI21X1_998 ( .A(u2__abc_52138_new_n5350_), .B(u2__abc_52138_new_n9977_), .C(u2__abc_52138_new_n9978_), .Y(u2__abc_52138_new_n9979_));
AOI21X1 AOI21X1_999 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n5357_), .C(u2__abc_52138_new_n6505_), .Y(u2__abc_52138_new_n9981_));
AOI22X1 AOI22X1_1 ( .A(_abc_65734_new_n1456_), .B(_abc_65734_new_n1459_), .C(_abc_65734_new_n753_), .D(_abc_65734_new_n1457_), .Y(\o[227] ));
AOI22X1 AOI22X1_10 ( .A(u2__abc_52138_new_n11386_), .B(u2__abc_52138_new_n11387_), .C(u2__abc_52138_new_n2981_), .D(u2__abc_52138_new_n11389_), .Y(u2__0cnt_7_0__2_));
AOI22X1 AOI22X1_100 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_116_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11792_));
AOI22X1 AOI22X1_101 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_117_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11795_));
AOI22X1 AOI22X1_102 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_118_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11798_));
AOI22X1 AOI22X1_103 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_119_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11801_));
AOI22X1 AOI22X1_104 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_120_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11804_));
AOI22X1 AOI22X1_105 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_121_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11807_));
AOI22X1 AOI22X1_106 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_122_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11810_));
AOI22X1 AOI22X1_107 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_123_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11813_));
AOI22X1 AOI22X1_108 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_124_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11816_));
AOI22X1 AOI22X1_109 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_125_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11819_));
AOI22X1 AOI22X1_11 ( .A(u2__abc_52138_new_n7779_), .B(u2__abc_52138_new_n2994_), .C(u2__abc_52138_new_n2981_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11508_));
AOI22X1 AOI22X1_110 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_126_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11822_));
AOI22X1 AOI22X1_111 ( .A(u2_remLo_127_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_129_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11824_));
AOI22X1 AOI22X1_112 ( .A(u2_remLo_129_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11825_));
AOI22X1 AOI22X1_113 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_128_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11828_));
AOI22X1 AOI22X1_114 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_130_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11837_));
AOI22X1 AOI22X1_115 ( .A(1'h0), .B(u2__abc_52138_new_n11717_), .C(u2__abc_52138_new_n11840_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11841_));
AOI22X1 AOI22X1_116 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_132_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11844_));
AOI22X1 AOI22X1_117 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_133_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11847_));
AOI22X1 AOI22X1_118 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_134_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11850_));
AOI22X1 AOI22X1_119 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_135_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11853_));
AOI22X1 AOI22X1_12 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_30_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11510_));
AOI22X1 AOI22X1_120 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_136_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11856_));
AOI22X1 AOI22X1_121 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_137_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11859_));
AOI22X1 AOI22X1_122 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_138_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11862_));
AOI22X1 AOI22X1_123 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_139_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11865_));
AOI22X1 AOI22X1_124 ( .A(u2_remLo_140_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_142_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11867_));
AOI22X1 AOI22X1_125 ( .A(u2_remLo_142_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11868_));
AOI22X1 AOI22X1_126 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_141_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11871_));
AOI22X1 AOI22X1_127 ( .A(fracta1_0_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_142_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11874_));
AOI22X1 AOI22X1_128 ( .A(fracta1_1_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_143_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11877_));
AOI22X1 AOI22X1_129 ( .A(fracta1_2_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_144_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11880_));
AOI22X1 AOI22X1_13 ( .A(u2_remLo_32_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_34_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11518_));
AOI22X1 AOI22X1_130 ( .A(fracta1_3_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_145_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11883_));
AOI22X1 AOI22X1_131 ( .A(fracta1_4_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_146_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11886_));
AOI22X1 AOI22X1_132 ( .A(fracta1_5_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_147_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11889_));
AOI22X1 AOI22X1_133 ( .A(fracta1_6_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_148_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11892_));
AOI22X1 AOI22X1_134 ( .A(fracta1_7_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_149_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11895_));
AOI22X1 AOI22X1_135 ( .A(fracta1_8_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_150_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11898_));
AOI22X1 AOI22X1_136 ( .A(fracta1_9_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_151_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11901_));
AOI22X1 AOI22X1_137 ( .A(fracta1_10_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_152_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11904_));
AOI22X1 AOI22X1_138 ( .A(fracta1_11_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_153_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11907_));
AOI22X1 AOI22X1_139 ( .A(fracta1_12_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_154_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11910_));
AOI22X1 AOI22X1_14 ( .A(u2_remLo_34_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11519_));
AOI22X1 AOI22X1_140 ( .A(fracta1_13_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_155_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11913_));
AOI22X1 AOI22X1_141 ( .A(fracta1_14_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_156_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11916_));
AOI22X1 AOI22X1_142 ( .A(fracta1_15_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_157_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11919_));
AOI22X1 AOI22X1_143 ( .A(u2_remLo_158_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_160_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11921_));
AOI22X1 AOI22X1_144 ( .A(u2_remLo_160_), .B(u2__abc_52138_new_n2994_), .C(fracta1_16_), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11922_));
AOI22X1 AOI22X1_145 ( .A(u2_remLo_159_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_161_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11924_));
AOI22X1 AOI22X1_146 ( .A(u2_remLo_161_), .B(u2__abc_52138_new_n2994_), .C(fracta1_17_), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11925_));
AOI22X1 AOI22X1_147 ( .A(fracta1_18_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_160_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11928_));
AOI22X1 AOI22X1_148 ( .A(fracta1_20_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_162_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11937_));
AOI22X1 AOI22X1_149 ( .A(fracta1_21_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_163_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11940_));
AOI22X1 AOI22X1_15 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_33_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11522_));
AOI22X1 AOI22X1_150 ( .A(fracta1_22_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_164_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11943_));
AOI22X1 AOI22X1_151 ( .A(fracta1_23_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_165_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11946_));
AOI22X1 AOI22X1_152 ( .A(fracta1_24_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_166_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11949_));
AOI22X1 AOI22X1_153 ( .A(fracta1_25_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_167_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11952_));
AOI22X1 AOI22X1_154 ( .A(fracta1_26_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_168_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11955_));
AOI22X1 AOI22X1_155 ( .A(fracta1_27_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_169_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11958_));
AOI22X1 AOI22X1_156 ( .A(fracta1_28_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_170_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11961_));
AOI22X1 AOI22X1_157 ( .A(fracta1_29_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_171_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11964_));
AOI22X1 AOI22X1_158 ( .A(fracta1_30_), .B(u2__abc_52138_new_n11717_), .C(u2__abc_52138_new_n11967_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11968_));
AOI22X1 AOI22X1_159 ( .A(fracta1_31_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_173_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11971_));
AOI22X1 AOI22X1_16 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_35_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11531_));
AOI22X1 AOI22X1_160 ( .A(fracta1_32_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_174_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11974_));
AOI22X1 AOI22X1_161 ( .A(fracta1_33_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_175_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11977_));
AOI22X1 AOI22X1_162 ( .A(fracta1_34_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_176_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11980_));
AOI22X1 AOI22X1_163 ( .A(fracta1_35_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_177_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11983_));
AOI22X1 AOI22X1_164 ( .A(fracta1_36_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_178_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11986_));
AOI22X1 AOI22X1_165 ( .A(fracta1_37_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_179_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11989_));
AOI22X1 AOI22X1_166 ( .A(fracta1_38_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_180_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11992_));
AOI22X1 AOI22X1_167 ( .A(fracta1_39_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_181_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11995_));
AOI22X1 AOI22X1_168 ( .A(fracta1_40_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_182_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11998_));
AOI22X1 AOI22X1_169 ( .A(fracta1_41_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_183_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12001_));
AOI22X1 AOI22X1_17 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_36_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11534_));
AOI22X1 AOI22X1_170 ( .A(fracta1_42_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_184_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12004_));
AOI22X1 AOI22X1_171 ( .A(fracta1_43_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_185_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12007_));
AOI22X1 AOI22X1_172 ( .A(fracta1_44_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_186_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12010_));
AOI22X1 AOI22X1_173 ( .A(fracta1_45_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_187_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12013_));
AOI22X1 AOI22X1_174 ( .A(fracta1_46_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_188_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12016_));
AOI22X1 AOI22X1_175 ( .A(fracta1_47_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_189_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12019_));
AOI22X1 AOI22X1_176 ( .A(fracta1_48_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_190_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12022_));
AOI22X1 AOI22X1_177 ( .A(u2_remLo_191_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_193_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n12024_));
AOI22X1 AOI22X1_178 ( .A(u2_remLo_193_), .B(u2__abc_52138_new_n2994_), .C(fracta1_49_), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n12025_));
AOI22X1 AOI22X1_179 ( .A(fracta1_50_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_192_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12028_));
AOI22X1 AOI22X1_18 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_37_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11537_));
AOI22X1 AOI22X1_180 ( .A(fracta1_52_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_194_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12037_));
AOI22X1 AOI22X1_181 ( .A(fracta1_53_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_195_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12040_));
AOI22X1 AOI22X1_182 ( .A(fracta1_54_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_196_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12043_));
AOI22X1 AOI22X1_183 ( .A(fracta1_55_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_197_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12046_));
AOI22X1 AOI22X1_184 ( .A(fracta1_56_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_198_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12049_));
AOI22X1 AOI22X1_185 ( .A(fracta1_57_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_199_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12052_));
AOI22X1 AOI22X1_186 ( .A(u2_remLo_200_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_202_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n12054_));
AOI22X1 AOI22X1_187 ( .A(u2_remLo_202_), .B(u2__abc_52138_new_n2994_), .C(fracta1_58_), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n12055_));
AOI22X1 AOI22X1_188 ( .A(fracta1_59_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_201_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12058_));
AOI22X1 AOI22X1_189 ( .A(fracta1_61_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_203_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12067_));
AOI22X1 AOI22X1_19 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_38_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11540_));
AOI22X1 AOI22X1_190 ( .A(fracta1_62_), .B(u2__abc_52138_new_n11717_), .C(u2__abc_52138_new_n12070_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12071_));
AOI22X1 AOI22X1_191 ( .A(fracta1_63_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_205_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12074_));
AOI22X1 AOI22X1_192 ( .A(fracta1_64_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_206_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12077_));
AOI22X1 AOI22X1_193 ( .A(fracta1_65_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_207_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12080_));
AOI22X1 AOI22X1_194 ( .A(fracta1_66_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_208_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12083_));
AOI22X1 AOI22X1_195 ( .A(fracta1_67_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_209_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12086_));
AOI22X1 AOI22X1_196 ( .A(fracta1_68_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_210_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12089_));
AOI22X1 AOI22X1_197 ( .A(fracta1_69_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_211_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12092_));
AOI22X1 AOI22X1_198 ( .A(fracta1_70_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_212_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12095_));
AOI22X1 AOI22X1_199 ( .A(fracta1_71_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_213_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12098_));
AOI22X1 AOI22X1_2 ( .A(_abc_65734_new_n1464_), .B(_abc_65734_new_n1471_), .C(_abc_65734_new_n1474_), .D(_abc_65734_new_n1472_), .Y(_abc_65734_new_n1475_));
AOI22X1 AOI22X1_20 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_39_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11543_));
AOI22X1 AOI22X1_200 ( .A(fracta1_72_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_214_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12101_));
AOI22X1 AOI22X1_201 ( .A(fracta1_73_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_215_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12104_));
AOI22X1 AOI22X1_202 ( .A(fracta1_74_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_216_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12107_));
AOI22X1 AOI22X1_203 ( .A(fracta1_75_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_217_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12110_));
AOI22X1 AOI22X1_204 ( .A(fracta1_76_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_218_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12113_));
AOI22X1 AOI22X1_205 ( .A(fracta1_77_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_219_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12116_));
AOI22X1 AOI22X1_206 ( .A(fracta1_78_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_220_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12119_));
AOI22X1 AOI22X1_207 ( .A(fracta1_79_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_221_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12122_));
AOI22X1 AOI22X1_208 ( .A(fracta1_80_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_222_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12125_));
AOI22X1 AOI22X1_209 ( .A(u2_remLo_223_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_225_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n12127_));
AOI22X1 AOI22X1_21 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_40_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11546_));
AOI22X1 AOI22X1_210 ( .A(u2_remLo_225_), .B(u2__abc_52138_new_n2994_), .C(fracta1_81_), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n12128_));
AOI22X1 AOI22X1_211 ( .A(u2_remLo_224_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_226_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n12130_));
AOI22X1 AOI22X1_212 ( .A(u2_remLo_226_), .B(u2__abc_52138_new_n2994_), .C(fracta1_82_), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n12131_));
AOI22X1 AOI22X1_213 ( .A(fracta1_85_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_227_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12146_));
AOI22X1 AOI22X1_214 ( .A(fracta1_86_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_228_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12149_));
AOI22X1 AOI22X1_215 ( .A(fracta1_87_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_229_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12152_));
AOI22X1 AOI22X1_216 ( .A(fracta1_88_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_230_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12155_));
AOI22X1 AOI22X1_217 ( .A(fracta1_89_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_231_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12158_));
AOI22X1 AOI22X1_218 ( .A(fracta1_90_), .B(u2__abc_52138_new_n11717_), .C(u2__abc_52138_new_n12161_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12162_));
AOI22X1 AOI22X1_219 ( .A(fracta1_91_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_233_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12165_));
AOI22X1 AOI22X1_22 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_41_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11549_));
AOI22X1 AOI22X1_220 ( .A(fracta1_92_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_234_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12168_));
AOI22X1 AOI22X1_221 ( .A(fracta1_93_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_235_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12171_));
AOI22X1 AOI22X1_222 ( .A(fracta1_94_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_236_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12174_));
AOI22X1 AOI22X1_223 ( .A(fracta1_95_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_237_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12177_));
AOI22X1 AOI22X1_224 ( .A(u2_remLo_238_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_240_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n12179_));
AOI22X1 AOI22X1_225 ( .A(u2_remLo_240_), .B(u2__abc_52138_new_n2994_), .C(fracta1_96_), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n12180_));
AOI22X1 AOI22X1_226 ( .A(fracta1_97_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_239_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12183_));
AOI22X1 AOI22X1_227 ( .A(fracta1_98_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_240_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12186_));
AOI22X1 AOI22X1_228 ( .A(fracta1_99_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_241_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12189_));
AOI22X1 AOI22X1_229 ( .A(fracta1_100_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_242_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12192_));
AOI22X1 AOI22X1_23 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_42_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11552_));
AOI22X1 AOI22X1_230 ( .A(fracta1_101_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_243_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12195_));
AOI22X1 AOI22X1_231 ( .A(fracta1_102_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_244_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12198_));
AOI22X1 AOI22X1_232 ( .A(fracta1_103_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_245_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12201_));
AOI22X1 AOI22X1_233 ( .A(fracta1_104_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_246_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12204_));
AOI22X1 AOI22X1_234 ( .A(fracta1_105_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_247_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12207_));
AOI22X1 AOI22X1_235 ( .A(fracta1_106_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_248_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12210_));
AOI22X1 AOI22X1_236 ( .A(fracta1_107_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_249_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12213_));
AOI22X1 AOI22X1_237 ( .A(fracta1_108_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_250_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12216_));
AOI22X1 AOI22X1_238 ( .A(fracta1_109_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_251_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12219_));
AOI22X1 AOI22X1_239 ( .A(fracta1_110_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_252_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12222_));
AOI22X1 AOI22X1_24 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_43_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11555_));
AOI22X1 AOI22X1_240 ( .A(fracta1_111_), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_253_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12225_));
AOI22X1 AOI22X1_241 ( .A(fracta1_112_), .B(u2__abc_52138_new_n11717_), .C(u2__abc_52138_new_n12228_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n12229_));
AOI22X1 AOI22X1_242 ( .A(u2_remLo_255_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_257_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n12231_));
AOI22X1 AOI22X1_243 ( .A(u2_remLo_257_), .B(u2__abc_52138_new_n2994_), .C(fracta1_113_), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n12232_));
AOI22X1 AOI22X1_25 ( .A(u2_remLo_44_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_46_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11557_));
AOI22X1 AOI22X1_26 ( .A(u2_remLo_46_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11558_));
AOI22X1 AOI22X1_27 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_45_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11561_));
AOI22X1 AOI22X1_28 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_47_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11570_));
AOI22X1 AOI22X1_29 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_48_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11573_));
AOI22X1 AOI22X1_3 ( .A(u2__abc_52138_new_n2963_), .B(u2__abc_52138_new_n2982_), .C(u2__abc_52138_new_n2981_), .D(u2__abc_52138_new_n2984_), .Y(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_0_));
AOI22X1 AOI22X1_30 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_49_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11576_));
AOI22X1 AOI22X1_31 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_50_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11579_));
AOI22X1 AOI22X1_32 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_51_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11582_));
AOI22X1 AOI22X1_33 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_52_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11585_));
AOI22X1 AOI22X1_34 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_53_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11588_));
AOI22X1 AOI22X1_35 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_54_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11591_));
AOI22X1 AOI22X1_36 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_55_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11594_));
AOI22X1 AOI22X1_37 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_56_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11597_));
AOI22X1 AOI22X1_38 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_57_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11600_));
AOI22X1 AOI22X1_39 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_58_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11603_));
AOI22X1 AOI22X1_4 ( .A(u2__abc_52138_new_n5368_), .B(u2_o_312_), .C(u2__abc_52138_new_n5814_), .D(u2__abc_52138_new_n5813_), .Y(u2__abc_52138_new_n5815_));
AOI22X1 AOI22X1_40 ( .A(u2_remLo_59_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_61_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11605_));
AOI22X1 AOI22X1_41 ( .A(u2_remLo_61_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11606_));
AOI22X1 AOI22X1_42 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_60_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11609_));
AOI22X1 AOI22X1_43 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_61_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11612_));
AOI22X1 AOI22X1_44 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_62_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11615_));
AOI22X1 AOI22X1_45 ( .A(u2_remLo_63_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_65_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11617_));
AOI22X1 AOI22X1_46 ( .A(u2_remLo_65_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11618_));
AOI22X1 AOI22X1_47 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_64_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11621_));
AOI22X1 AOI22X1_48 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_66_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11630_));
AOI22X1 AOI22X1_49 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_67_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11633_));
AOI22X1 AOI22X1_5 ( .A(u2__abc_52138_new_n5872_), .B(u2__abc_52138_new_n5873_), .C(u2__abc_52138_new_n5876_), .D(u2__abc_52138_new_n5240_), .Y(u2__abc_52138_new_n5877_));
AOI22X1 AOI22X1_50 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_68_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11636_));
AOI22X1 AOI22X1_51 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_69_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11639_));
AOI22X1 AOI22X1_52 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_70_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11642_));
AOI22X1 AOI22X1_53 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_71_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11645_));
AOI22X1 AOI22X1_54 ( .A(u2_remLo_72_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_74_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11647_));
AOI22X1 AOI22X1_55 ( .A(u2_remLo_74_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11648_));
AOI22X1 AOI22X1_56 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_73_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11651_));
AOI22X1 AOI22X1_57 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_75_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11660_));
AOI22X1 AOI22X1_58 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_76_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11663_));
AOI22X1 AOI22X1_59 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_77_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11666_));
AOI22X1 AOI22X1_6 ( .A(u2__abc_52138_new_n6479_), .B(u2__abc_52138_new_n6497_), .C(u2__abc_52138_new_n6450_), .D(u2__abc_52138_new_n6442_), .Y(u2__abc_52138_new_n6498_));
AOI22X1 AOI22X1_60 ( .A(u2_remLo_78_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_80_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11668_));
AOI22X1 AOI22X1_61 ( .A(u2_remLo_80_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11669_));
AOI22X1 AOI22X1_62 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_79_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11672_));
AOI22X1 AOI22X1_63 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_80_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11675_));
AOI22X1 AOI22X1_64 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_81_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11678_));
AOI22X1 AOI22X1_65 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_82_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11681_));
AOI22X1 AOI22X1_66 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_83_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11684_));
AOI22X1 AOI22X1_67 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_84_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11687_));
AOI22X1 AOI22X1_68 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_85_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11690_));
AOI22X1 AOI22X1_69 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_86_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11693_));
AOI22X1 AOI22X1_7 ( .A(u2__abc_52138_new_n3082_), .B(u2__abc_52138_new_n6559_), .C(u2__abc_52138_new_n6465_), .D(u2__abc_52138_new_n6542_), .Y(u2__abc_52138_new_n6560_));
AOI22X1 AOI22X1_70 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_87_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11696_));
AOI22X1 AOI22X1_71 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_88_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11699_));
AOI22X1 AOI22X1_72 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_89_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11702_));
AOI22X1 AOI22X1_73 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_90_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11705_));
AOI22X1 AOI22X1_74 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_91_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11708_));
AOI22X1 AOI22X1_75 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_92_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11711_));
AOI22X1 AOI22X1_76 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_93_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11714_));
AOI22X1 AOI22X1_77 ( .A(1'h0), .B(u2__abc_52138_new_n11717_), .C(u2__abc_52138_new_n11718_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11719_));
AOI22X1 AOI22X1_78 ( .A(u2_remLo_95_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_97_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11721_));
AOI22X1 AOI22X1_79 ( .A(u2_remLo_97_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11722_));
AOI22X1 AOI22X1_8 ( .A(u2__abc_52138_new_n4109_), .B(u2__abc_52138_new_n9102_), .C(u2__abc_52138_new_n4122_), .D(u2__abc_52138_new_n9100_), .Y(u2__abc_52138_new_n9103_));
AOI22X1 AOI22X1_80 ( .A(1'h0), .B(u2__abc_52138_new_n11717_), .C(u2__abc_52138_new_n11725_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11726_));
AOI22X1 AOI22X1_81 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_98_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11735_));
AOI22X1 AOI22X1_82 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_99_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11738_));
AOI22X1 AOI22X1_83 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_100_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11741_));
AOI22X1 AOI22X1_84 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_101_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11744_));
AOI22X1 AOI22X1_85 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_102_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11747_));
AOI22X1 AOI22X1_86 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_103_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11750_));
AOI22X1 AOI22X1_87 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_104_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11753_));
AOI22X1 AOI22X1_88 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_105_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11756_));
AOI22X1 AOI22X1_89 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_106_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11759_));
AOI22X1 AOI22X1_9 ( .A(u2__abc_52138_new_n5887_), .B(u2__abc_52138_new_n10524_), .C(u2__abc_52138_new_n10505_), .D(u2__abc_52138_new_n10525_), .Y(u2__abc_52138_new_n10526_));
AOI22X1 AOI22X1_90 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_107_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11762_));
AOI22X1 AOI22X1_91 ( .A(u2_remLo_108_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_110_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11764_));
AOI22X1 AOI22X1_92 ( .A(u2_remLo_110_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11765_));
AOI22X1 AOI22X1_93 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_109_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11768_));
AOI22X1 AOI22X1_94 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_110_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11771_));
AOI22X1 AOI22X1_95 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_111_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11774_));
AOI22X1 AOI22X1_96 ( .A(u2_remLo_112_), .B(u2__abc_52138_new_n11509_), .C(u2_remLo_114_), .D(u2__abc_52138_new_n11412_), .Y(u2__abc_52138_new_n11776_));
AOI22X1 AOI22X1_97 ( .A(u2_remLo_114_), .B(u2__abc_52138_new_n2994_), .C(1'h0), .D(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11777_));
AOI22X1 AOI22X1_98 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_113_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11780_));
AOI22X1 AOI22X1_99 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .C(u2_remLo_115_), .D(u2__abc_52138_new_n11509_), .Y(u2__abc_52138_new_n11789_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_0_), .Q(u2_state_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(u2__0root_452_0__6_), .Q(sqrto_5_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk), .D(u2__0root_452_0__96_), .Q(sqrto_95_));
DFFPOSX1 DFFPOSX1_1000 ( .CLK(clk), .D(u2__0remHi_451_0__93_), .Q(u2_remHi_93_));
DFFPOSX1 DFFPOSX1_1001 ( .CLK(clk), .D(u2__0remHi_451_0__94_), .Q(u2_remHi_94_));
DFFPOSX1 DFFPOSX1_1002 ( .CLK(clk), .D(u2__0remHi_451_0__95_), .Q(u2_remHi_95_));
DFFPOSX1 DFFPOSX1_1003 ( .CLK(clk), .D(u2__0remHi_451_0__96_), .Q(u2_remHi_96_));
DFFPOSX1 DFFPOSX1_1004 ( .CLK(clk), .D(u2__0remHi_451_0__97_), .Q(u2_remHi_97_));
DFFPOSX1 DFFPOSX1_1005 ( .CLK(clk), .D(u2__0remHi_451_0__98_), .Q(u2_remHi_98_));
DFFPOSX1 DFFPOSX1_1006 ( .CLK(clk), .D(u2__0remHi_451_0__99_), .Q(u2_remHi_99_));
DFFPOSX1 DFFPOSX1_1007 ( .CLK(clk), .D(u2__0remHi_451_0__100_), .Q(u2_remHi_100_));
DFFPOSX1 DFFPOSX1_1008 ( .CLK(clk), .D(u2__0remHi_451_0__101_), .Q(u2_remHi_101_));
DFFPOSX1 DFFPOSX1_1009 ( .CLK(clk), .D(u2__0remHi_451_0__102_), .Q(u2_remHi_102_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk), .D(u2__0root_452_0__97_), .Q(sqrto_96_));
DFFPOSX1 DFFPOSX1_1010 ( .CLK(clk), .D(u2__0remHi_451_0__103_), .Q(u2_remHi_103_));
DFFPOSX1 DFFPOSX1_1011 ( .CLK(clk), .D(u2__0remHi_451_0__104_), .Q(u2_remHi_104_));
DFFPOSX1 DFFPOSX1_1012 ( .CLK(clk), .D(u2__0remHi_451_0__105_), .Q(u2_remHi_105_));
DFFPOSX1 DFFPOSX1_1013 ( .CLK(clk), .D(u2__0remHi_451_0__106_), .Q(u2_remHi_106_));
DFFPOSX1 DFFPOSX1_1014 ( .CLK(clk), .D(u2__0remHi_451_0__107_), .Q(u2_remHi_107_));
DFFPOSX1 DFFPOSX1_1015 ( .CLK(clk), .D(u2__0remHi_451_0__108_), .Q(u2_remHi_108_));
DFFPOSX1 DFFPOSX1_1016 ( .CLK(clk), .D(u2__0remHi_451_0__109_), .Q(u2_remHi_109_));
DFFPOSX1 DFFPOSX1_1017 ( .CLK(clk), .D(u2__0remHi_451_0__110_), .Q(u2_remHi_110_));
DFFPOSX1 DFFPOSX1_1018 ( .CLK(clk), .D(u2__0remHi_451_0__111_), .Q(u2_remHi_111_));
DFFPOSX1 DFFPOSX1_1019 ( .CLK(clk), .D(u2__0remHi_451_0__112_), .Q(u2_remHi_112_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk), .D(u2__0root_452_0__98_), .Q(sqrto_97_));
DFFPOSX1 DFFPOSX1_1020 ( .CLK(clk), .D(u2__0remHi_451_0__113_), .Q(u2_remHi_113_));
DFFPOSX1 DFFPOSX1_1021 ( .CLK(clk), .D(u2__0remHi_451_0__114_), .Q(u2_remHi_114_));
DFFPOSX1 DFFPOSX1_1022 ( .CLK(clk), .D(u2__0remHi_451_0__115_), .Q(u2_remHi_115_));
DFFPOSX1 DFFPOSX1_1023 ( .CLK(clk), .D(u2__0remHi_451_0__116_), .Q(u2_remHi_116_));
DFFPOSX1 DFFPOSX1_1024 ( .CLK(clk), .D(u2__0remHi_451_0__117_), .Q(u2_remHi_117_));
DFFPOSX1 DFFPOSX1_1025 ( .CLK(clk), .D(u2__0remHi_451_0__118_), .Q(u2_remHi_118_));
DFFPOSX1 DFFPOSX1_1026 ( .CLK(clk), .D(u2__0remHi_451_0__119_), .Q(u2_remHi_119_));
DFFPOSX1 DFFPOSX1_1027 ( .CLK(clk), .D(u2__0remHi_451_0__120_), .Q(u2_remHi_120_));
DFFPOSX1 DFFPOSX1_1028 ( .CLK(clk), .D(u2__0remHi_451_0__121_), .Q(u2_remHi_121_));
DFFPOSX1 DFFPOSX1_1029 ( .CLK(clk), .D(u2__0remHi_451_0__122_), .Q(u2_remHi_122_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk), .D(u2__0root_452_0__99_), .Q(sqrto_98_));
DFFPOSX1 DFFPOSX1_1030 ( .CLK(clk), .D(u2__0remHi_451_0__123_), .Q(u2_remHi_123_));
DFFPOSX1 DFFPOSX1_1031 ( .CLK(clk), .D(u2__0remHi_451_0__124_), .Q(u2_remHi_124_));
DFFPOSX1 DFFPOSX1_1032 ( .CLK(clk), .D(u2__0remHi_451_0__125_), .Q(u2_remHi_125_));
DFFPOSX1 DFFPOSX1_1033 ( .CLK(clk), .D(u2__0remHi_451_0__126_), .Q(u2_remHi_126_));
DFFPOSX1 DFFPOSX1_1034 ( .CLK(clk), .D(u2__0remHi_451_0__127_), .Q(u2_remHi_127_));
DFFPOSX1 DFFPOSX1_1035 ( .CLK(clk), .D(u2__0remHi_451_0__128_), .Q(u2_remHi_128_));
DFFPOSX1 DFFPOSX1_1036 ( .CLK(clk), .D(u2__0remHi_451_0__129_), .Q(u2_remHi_129_));
DFFPOSX1 DFFPOSX1_1037 ( .CLK(clk), .D(u2__0remHi_451_0__130_), .Q(u2_remHi_130_));
DFFPOSX1 DFFPOSX1_1038 ( .CLK(clk), .D(u2__0remHi_451_0__131_), .Q(u2_remHi_131_));
DFFPOSX1 DFFPOSX1_1039 ( .CLK(clk), .D(u2__0remHi_451_0__132_), .Q(u2_remHi_132_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk), .D(u2__0root_452_0__100_), .Q(sqrto_99_));
DFFPOSX1 DFFPOSX1_1040 ( .CLK(clk), .D(u2__0remHi_451_0__133_), .Q(u2_remHi_133_));
DFFPOSX1 DFFPOSX1_1041 ( .CLK(clk), .D(u2__0remHi_451_0__134_), .Q(u2_remHi_134_));
DFFPOSX1 DFFPOSX1_1042 ( .CLK(clk), .D(u2__0remHi_451_0__135_), .Q(u2_remHi_135_));
DFFPOSX1 DFFPOSX1_1043 ( .CLK(clk), .D(u2__0remHi_451_0__136_), .Q(u2_remHi_136_));
DFFPOSX1 DFFPOSX1_1044 ( .CLK(clk), .D(u2__0remHi_451_0__137_), .Q(u2_remHi_137_));
DFFPOSX1 DFFPOSX1_1045 ( .CLK(clk), .D(u2__0remHi_451_0__138_), .Q(u2_remHi_138_));
DFFPOSX1 DFFPOSX1_1046 ( .CLK(clk), .D(u2__0remHi_451_0__139_), .Q(u2_remHi_139_));
DFFPOSX1 DFFPOSX1_1047 ( .CLK(clk), .D(u2__0remHi_451_0__140_), .Q(u2_remHi_140_));
DFFPOSX1 DFFPOSX1_1048 ( .CLK(clk), .D(u2__0remHi_451_0__141_), .Q(u2_remHi_141_));
DFFPOSX1 DFFPOSX1_1049 ( .CLK(clk), .D(u2__0remHi_451_0__142_), .Q(u2_remHi_142_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk), .D(u2__0root_452_0__101_), .Q(sqrto_100_));
DFFPOSX1 DFFPOSX1_1050 ( .CLK(clk), .D(u2__0remHi_451_0__143_), .Q(u2_remHi_143_));
DFFPOSX1 DFFPOSX1_1051 ( .CLK(clk), .D(u2__0remHi_451_0__144_), .Q(u2_remHi_144_));
DFFPOSX1 DFFPOSX1_1052 ( .CLK(clk), .D(u2__0remHi_451_0__145_), .Q(u2_remHi_145_));
DFFPOSX1 DFFPOSX1_1053 ( .CLK(clk), .D(u2__0remHi_451_0__146_), .Q(u2_remHi_146_));
DFFPOSX1 DFFPOSX1_1054 ( .CLK(clk), .D(u2__0remHi_451_0__147_), .Q(u2_remHi_147_));
DFFPOSX1 DFFPOSX1_1055 ( .CLK(clk), .D(u2__0remHi_451_0__148_), .Q(u2_remHi_148_));
DFFPOSX1 DFFPOSX1_1056 ( .CLK(clk), .D(u2__0remHi_451_0__149_), .Q(u2_remHi_149_));
DFFPOSX1 DFFPOSX1_1057 ( .CLK(clk), .D(u2__0remHi_451_0__150_), .Q(u2_remHi_150_));
DFFPOSX1 DFFPOSX1_1058 ( .CLK(clk), .D(u2__0remHi_451_0__151_), .Q(u2_remHi_151_));
DFFPOSX1 DFFPOSX1_1059 ( .CLK(clk), .D(u2__0remHi_451_0__152_), .Q(u2_remHi_152_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk), .D(u2__0root_452_0__102_), .Q(sqrto_101_));
DFFPOSX1 DFFPOSX1_1060 ( .CLK(clk), .D(u2__0remHi_451_0__153_), .Q(u2_remHi_153_));
DFFPOSX1 DFFPOSX1_1061 ( .CLK(clk), .D(u2__0remHi_451_0__154_), .Q(u2_remHi_154_));
DFFPOSX1 DFFPOSX1_1062 ( .CLK(clk), .D(u2__0remHi_451_0__155_), .Q(u2_remHi_155_));
DFFPOSX1 DFFPOSX1_1063 ( .CLK(clk), .D(u2__0remHi_451_0__156_), .Q(u2_remHi_156_));
DFFPOSX1 DFFPOSX1_1064 ( .CLK(clk), .D(u2__0remHi_451_0__157_), .Q(u2_remHi_157_));
DFFPOSX1 DFFPOSX1_1065 ( .CLK(clk), .D(u2__0remHi_451_0__158_), .Q(u2_remHi_158_));
DFFPOSX1 DFFPOSX1_1066 ( .CLK(clk), .D(u2__0remHi_451_0__159_), .Q(u2_remHi_159_));
DFFPOSX1 DFFPOSX1_1067 ( .CLK(clk), .D(u2__0remHi_451_0__160_), .Q(u2_remHi_160_));
DFFPOSX1 DFFPOSX1_1068 ( .CLK(clk), .D(u2__0remHi_451_0__161_), .Q(u2_remHi_161_));
DFFPOSX1 DFFPOSX1_1069 ( .CLK(clk), .D(u2__0remHi_451_0__162_), .Q(u2_remHi_162_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk), .D(u2__0root_452_0__103_), .Q(sqrto_102_));
DFFPOSX1 DFFPOSX1_1070 ( .CLK(clk), .D(u2__0remHi_451_0__163_), .Q(u2_remHi_163_));
DFFPOSX1 DFFPOSX1_1071 ( .CLK(clk), .D(u2__0remHi_451_0__164_), .Q(u2_remHi_164_));
DFFPOSX1 DFFPOSX1_1072 ( .CLK(clk), .D(u2__0remHi_451_0__165_), .Q(u2_remHi_165_));
DFFPOSX1 DFFPOSX1_1073 ( .CLK(clk), .D(u2__0remHi_451_0__166_), .Q(u2_remHi_166_));
DFFPOSX1 DFFPOSX1_1074 ( .CLK(clk), .D(u2__0remHi_451_0__167_), .Q(u2_remHi_167_));
DFFPOSX1 DFFPOSX1_1075 ( .CLK(clk), .D(u2__0remHi_451_0__168_), .Q(u2_remHi_168_));
DFFPOSX1 DFFPOSX1_1076 ( .CLK(clk), .D(u2__0remHi_451_0__169_), .Q(u2_remHi_169_));
DFFPOSX1 DFFPOSX1_1077 ( .CLK(clk), .D(u2__0remHi_451_0__170_), .Q(u2_remHi_170_));
DFFPOSX1 DFFPOSX1_1078 ( .CLK(clk), .D(u2__0remHi_451_0__171_), .Q(u2_remHi_171_));
DFFPOSX1 DFFPOSX1_1079 ( .CLK(clk), .D(u2__0remHi_451_0__172_), .Q(u2_remHi_172_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk), .D(u2__0root_452_0__104_), .Q(sqrto_103_));
DFFPOSX1 DFFPOSX1_1080 ( .CLK(clk), .D(u2__0remHi_451_0__173_), .Q(u2_remHi_173_));
DFFPOSX1 DFFPOSX1_1081 ( .CLK(clk), .D(u2__0remHi_451_0__174_), .Q(u2_remHi_174_));
DFFPOSX1 DFFPOSX1_1082 ( .CLK(clk), .D(u2__0remHi_451_0__175_), .Q(u2_remHi_175_));
DFFPOSX1 DFFPOSX1_1083 ( .CLK(clk), .D(u2__0remHi_451_0__176_), .Q(u2_remHi_176_));
DFFPOSX1 DFFPOSX1_1084 ( .CLK(clk), .D(u2__0remHi_451_0__177_), .Q(u2_remHi_177_));
DFFPOSX1 DFFPOSX1_1085 ( .CLK(clk), .D(u2__0remHi_451_0__178_), .Q(u2_remHi_178_));
DFFPOSX1 DFFPOSX1_1086 ( .CLK(clk), .D(u2__0remHi_451_0__179_), .Q(u2_remHi_179_));
DFFPOSX1 DFFPOSX1_1087 ( .CLK(clk), .D(u2__0remHi_451_0__180_), .Q(u2_remHi_180_));
DFFPOSX1 DFFPOSX1_1088 ( .CLK(clk), .D(u2__0remHi_451_0__181_), .Q(u2_remHi_181_));
DFFPOSX1 DFFPOSX1_1089 ( .CLK(clk), .D(u2__0remHi_451_0__182_), .Q(u2_remHi_182_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk), .D(u2__0root_452_0__105_), .Q(sqrto_104_));
DFFPOSX1 DFFPOSX1_1090 ( .CLK(clk), .D(u2__0remHi_451_0__183_), .Q(u2_remHi_183_));
DFFPOSX1 DFFPOSX1_1091 ( .CLK(clk), .D(u2__0remHi_451_0__184_), .Q(u2_remHi_184_));
DFFPOSX1 DFFPOSX1_1092 ( .CLK(clk), .D(u2__0remHi_451_0__185_), .Q(u2_remHi_185_));
DFFPOSX1 DFFPOSX1_1093 ( .CLK(clk), .D(u2__0remHi_451_0__186_), .Q(u2_remHi_186_));
DFFPOSX1 DFFPOSX1_1094 ( .CLK(clk), .D(u2__0remHi_451_0__187_), .Q(u2_remHi_187_));
DFFPOSX1 DFFPOSX1_1095 ( .CLK(clk), .D(u2__0remHi_451_0__188_), .Q(u2_remHi_188_));
DFFPOSX1 DFFPOSX1_1096 ( .CLK(clk), .D(u2__0remHi_451_0__189_), .Q(u2_remHi_189_));
DFFPOSX1 DFFPOSX1_1097 ( .CLK(clk), .D(u2__0remHi_451_0__190_), .Q(u2_remHi_190_));
DFFPOSX1 DFFPOSX1_1098 ( .CLK(clk), .D(u2__0remHi_451_0__191_), .Q(u2_remHi_191_));
DFFPOSX1 DFFPOSX1_1099 ( .CLK(clk), .D(u2__0remHi_451_0__192_), .Q(u2_remHi_192_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(u2__0root_452_0__7_), .Q(sqrto_6_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk), .D(u2__0root_452_0__106_), .Q(sqrto_105_));
DFFPOSX1 DFFPOSX1_1100 ( .CLK(clk), .D(u2__0remHi_451_0__193_), .Q(u2_remHi_193_));
DFFPOSX1 DFFPOSX1_1101 ( .CLK(clk), .D(u2__0remHi_451_0__194_), .Q(u2_remHi_194_));
DFFPOSX1 DFFPOSX1_1102 ( .CLK(clk), .D(u2__0remHi_451_0__195_), .Q(u2_remHi_195_));
DFFPOSX1 DFFPOSX1_1103 ( .CLK(clk), .D(u2__0remHi_451_0__196_), .Q(u2_remHi_196_));
DFFPOSX1 DFFPOSX1_1104 ( .CLK(clk), .D(u2__0remHi_451_0__197_), .Q(u2_remHi_197_));
DFFPOSX1 DFFPOSX1_1105 ( .CLK(clk), .D(u2__0remHi_451_0__198_), .Q(u2_remHi_198_));
DFFPOSX1 DFFPOSX1_1106 ( .CLK(clk), .D(u2__0remHi_451_0__199_), .Q(u2_remHi_199_));
DFFPOSX1 DFFPOSX1_1107 ( .CLK(clk), .D(u2__0remHi_451_0__200_), .Q(u2_remHi_200_));
DFFPOSX1 DFFPOSX1_1108 ( .CLK(clk), .D(u2__0remHi_451_0__201_), .Q(u2_remHi_201_));
DFFPOSX1 DFFPOSX1_1109 ( .CLK(clk), .D(u2__0remHi_451_0__202_), .Q(u2_remHi_202_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk), .D(u2__0root_452_0__107_), .Q(sqrto_106_));
DFFPOSX1 DFFPOSX1_1110 ( .CLK(clk), .D(u2__0remHi_451_0__203_), .Q(u2_remHi_203_));
DFFPOSX1 DFFPOSX1_1111 ( .CLK(clk), .D(u2__0remHi_451_0__204_), .Q(u2_remHi_204_));
DFFPOSX1 DFFPOSX1_1112 ( .CLK(clk), .D(u2__0remHi_451_0__205_), .Q(u2_remHi_205_));
DFFPOSX1 DFFPOSX1_1113 ( .CLK(clk), .D(u2__0remHi_451_0__206_), .Q(u2_remHi_206_));
DFFPOSX1 DFFPOSX1_1114 ( .CLK(clk), .D(u2__0remHi_451_0__207_), .Q(u2_remHi_207_));
DFFPOSX1 DFFPOSX1_1115 ( .CLK(clk), .D(u2__0remHi_451_0__208_), .Q(u2_remHi_208_));
DFFPOSX1 DFFPOSX1_1116 ( .CLK(clk), .D(u2__0remHi_451_0__209_), .Q(u2_remHi_209_));
DFFPOSX1 DFFPOSX1_1117 ( .CLK(clk), .D(u2__0remHi_451_0__210_), .Q(u2_remHi_210_));
DFFPOSX1 DFFPOSX1_1118 ( .CLK(clk), .D(u2__0remHi_451_0__211_), .Q(u2_remHi_211_));
DFFPOSX1 DFFPOSX1_1119 ( .CLK(clk), .D(u2__0remHi_451_0__212_), .Q(u2_remHi_212_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk), .D(u2__0root_452_0__108_), .Q(sqrto_107_));
DFFPOSX1 DFFPOSX1_1120 ( .CLK(clk), .D(u2__0remHi_451_0__213_), .Q(u2_remHi_213_));
DFFPOSX1 DFFPOSX1_1121 ( .CLK(clk), .D(u2__0remHi_451_0__214_), .Q(u2_remHi_214_));
DFFPOSX1 DFFPOSX1_1122 ( .CLK(clk), .D(u2__0remHi_451_0__215_), .Q(u2_remHi_215_));
DFFPOSX1 DFFPOSX1_1123 ( .CLK(clk), .D(u2__0remHi_451_0__216_), .Q(u2_remHi_216_));
DFFPOSX1 DFFPOSX1_1124 ( .CLK(clk), .D(u2__0remHi_451_0__217_), .Q(u2_remHi_217_));
DFFPOSX1 DFFPOSX1_1125 ( .CLK(clk), .D(u2__0remHi_451_0__218_), .Q(u2_remHi_218_));
DFFPOSX1 DFFPOSX1_1126 ( .CLK(clk), .D(u2__0remHi_451_0__219_), .Q(u2_remHi_219_));
DFFPOSX1 DFFPOSX1_1127 ( .CLK(clk), .D(u2__0remHi_451_0__220_), .Q(u2_remHi_220_));
DFFPOSX1 DFFPOSX1_1128 ( .CLK(clk), .D(u2__0remHi_451_0__221_), .Q(u2_remHi_221_));
DFFPOSX1 DFFPOSX1_1129 ( .CLK(clk), .D(u2__0remHi_451_0__222_), .Q(u2_remHi_222_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk), .D(u2__0root_452_0__109_), .Q(sqrto_108_));
DFFPOSX1 DFFPOSX1_1130 ( .CLK(clk), .D(u2__0remHi_451_0__223_), .Q(u2_remHi_223_));
DFFPOSX1 DFFPOSX1_1131 ( .CLK(clk), .D(u2__0remHi_451_0__224_), .Q(u2_remHi_224_));
DFFPOSX1 DFFPOSX1_1132 ( .CLK(clk), .D(u2__0remHi_451_0__225_), .Q(u2_remHi_225_));
DFFPOSX1 DFFPOSX1_1133 ( .CLK(clk), .D(u2__0remHi_451_0__226_), .Q(u2_remHi_226_));
DFFPOSX1 DFFPOSX1_1134 ( .CLK(clk), .D(u2__0remHi_451_0__227_), .Q(u2_remHi_227_));
DFFPOSX1 DFFPOSX1_1135 ( .CLK(clk), .D(u2__0remHi_451_0__228_), .Q(u2_remHi_228_));
DFFPOSX1 DFFPOSX1_1136 ( .CLK(clk), .D(u2__0remHi_451_0__229_), .Q(u2_remHi_229_));
DFFPOSX1 DFFPOSX1_1137 ( .CLK(clk), .D(u2__0remHi_451_0__230_), .Q(u2_remHi_230_));
DFFPOSX1 DFFPOSX1_1138 ( .CLK(clk), .D(u2__0remHi_451_0__231_), .Q(u2_remHi_231_));
DFFPOSX1 DFFPOSX1_1139 ( .CLK(clk), .D(u2__0remHi_451_0__232_), .Q(u2_remHi_232_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk), .D(u2__0root_452_0__110_), .Q(sqrto_109_));
DFFPOSX1 DFFPOSX1_1140 ( .CLK(clk), .D(u2__0remHi_451_0__233_), .Q(u2_remHi_233_));
DFFPOSX1 DFFPOSX1_1141 ( .CLK(clk), .D(u2__0remHi_451_0__234_), .Q(u2_remHi_234_));
DFFPOSX1 DFFPOSX1_1142 ( .CLK(clk), .D(u2__0remHi_451_0__235_), .Q(u2_remHi_235_));
DFFPOSX1 DFFPOSX1_1143 ( .CLK(clk), .D(u2__0remHi_451_0__236_), .Q(u2_remHi_236_));
DFFPOSX1 DFFPOSX1_1144 ( .CLK(clk), .D(u2__0remHi_451_0__237_), .Q(u2_remHi_237_));
DFFPOSX1 DFFPOSX1_1145 ( .CLK(clk), .D(u2__0remHi_451_0__238_), .Q(u2_remHi_238_));
DFFPOSX1 DFFPOSX1_1146 ( .CLK(clk), .D(u2__0remHi_451_0__239_), .Q(u2_remHi_239_));
DFFPOSX1 DFFPOSX1_1147 ( .CLK(clk), .D(u2__0remHi_451_0__240_), .Q(u2_remHi_240_));
DFFPOSX1 DFFPOSX1_1148 ( .CLK(clk), .D(u2__0remHi_451_0__241_), .Q(u2_remHi_241_));
DFFPOSX1 DFFPOSX1_1149 ( .CLK(clk), .D(u2__0remHi_451_0__242_), .Q(u2_remHi_242_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk), .D(u2__0root_452_0__111_), .Q(sqrto_110_));
DFFPOSX1 DFFPOSX1_1150 ( .CLK(clk), .D(u2__0remHi_451_0__243_), .Q(u2_remHi_243_));
DFFPOSX1 DFFPOSX1_1151 ( .CLK(clk), .D(u2__0remHi_451_0__244_), .Q(u2_remHi_244_));
DFFPOSX1 DFFPOSX1_1152 ( .CLK(clk), .D(u2__0remHi_451_0__245_), .Q(u2_remHi_245_));
DFFPOSX1 DFFPOSX1_1153 ( .CLK(clk), .D(u2__0remHi_451_0__246_), .Q(u2_remHi_246_));
DFFPOSX1 DFFPOSX1_1154 ( .CLK(clk), .D(u2__0remHi_451_0__247_), .Q(u2_remHi_247_));
DFFPOSX1 DFFPOSX1_1155 ( .CLK(clk), .D(u2__0remHi_451_0__248_), .Q(u2_remHi_248_));
DFFPOSX1 DFFPOSX1_1156 ( .CLK(clk), .D(u2__0remHi_451_0__249_), .Q(u2_remHi_249_));
DFFPOSX1 DFFPOSX1_1157 ( .CLK(clk), .D(u2__0remHi_451_0__250_), .Q(u2_remHi_250_));
DFFPOSX1 DFFPOSX1_1158 ( .CLK(clk), .D(u2__0remHi_451_0__251_), .Q(u2_remHi_251_));
DFFPOSX1 DFFPOSX1_1159 ( .CLK(clk), .D(u2__0remHi_451_0__252_), .Q(u2_remHi_252_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk), .D(u2__0root_452_0__112_), .Q(sqrto_111_));
DFFPOSX1 DFFPOSX1_1160 ( .CLK(clk), .D(u2__0remHi_451_0__253_), .Q(u2_remHi_253_));
DFFPOSX1 DFFPOSX1_1161 ( .CLK(clk), .D(u2__0remHi_451_0__254_), .Q(u2_remHi_254_));
DFFPOSX1 DFFPOSX1_1162 ( .CLK(clk), .D(u2__0remHi_451_0__255_), .Q(u2_remHi_255_));
DFFPOSX1 DFFPOSX1_1163 ( .CLK(clk), .D(u2__0remHi_451_0__256_), .Q(u2_remHi_256_));
DFFPOSX1 DFFPOSX1_1164 ( .CLK(clk), .D(u2__0remHi_451_0__257_), .Q(u2_remHi_257_));
DFFPOSX1 DFFPOSX1_1165 ( .CLK(clk), .D(u2__0remHi_451_0__258_), .Q(u2_remHi_258_));
DFFPOSX1 DFFPOSX1_1166 ( .CLK(clk), .D(u2__0remHi_451_0__259_), .Q(u2_remHi_259_));
DFFPOSX1 DFFPOSX1_1167 ( .CLK(clk), .D(u2__0remHi_451_0__260_), .Q(u2_remHi_260_));
DFFPOSX1 DFFPOSX1_1168 ( .CLK(clk), .D(u2__0remHi_451_0__261_), .Q(u2_remHi_261_));
DFFPOSX1 DFFPOSX1_1169 ( .CLK(clk), .D(u2__0remHi_451_0__262_), .Q(u2_remHi_262_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk), .D(u2__0root_452_0__113_), .Q(sqrto_112_));
DFFPOSX1 DFFPOSX1_1170 ( .CLK(clk), .D(u2__0remHi_451_0__263_), .Q(u2_remHi_263_));
DFFPOSX1 DFFPOSX1_1171 ( .CLK(clk), .D(u2__0remHi_451_0__264_), .Q(u2_remHi_264_));
DFFPOSX1 DFFPOSX1_1172 ( .CLK(clk), .D(u2__0remHi_451_0__265_), .Q(u2_remHi_265_));
DFFPOSX1 DFFPOSX1_1173 ( .CLK(clk), .D(u2__0remHi_451_0__266_), .Q(u2_remHi_266_));
DFFPOSX1 DFFPOSX1_1174 ( .CLK(clk), .D(u2__0remHi_451_0__267_), .Q(u2_remHi_267_));
DFFPOSX1 DFFPOSX1_1175 ( .CLK(clk), .D(u2__0remHi_451_0__268_), .Q(u2_remHi_268_));
DFFPOSX1 DFFPOSX1_1176 ( .CLK(clk), .D(u2__0remHi_451_0__269_), .Q(u2_remHi_269_));
DFFPOSX1 DFFPOSX1_1177 ( .CLK(clk), .D(u2__0remHi_451_0__270_), .Q(u2_remHi_270_));
DFFPOSX1 DFFPOSX1_1178 ( .CLK(clk), .D(u2__0remHi_451_0__271_), .Q(u2_remHi_271_));
DFFPOSX1 DFFPOSX1_1179 ( .CLK(clk), .D(u2__0remHi_451_0__272_), .Q(u2_remHi_272_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk), .D(u2__0root_452_0__114_), .Q(sqrto_113_));
DFFPOSX1 DFFPOSX1_1180 ( .CLK(clk), .D(u2__0remHi_451_0__273_), .Q(u2_remHi_273_));
DFFPOSX1 DFFPOSX1_1181 ( .CLK(clk), .D(u2__0remHi_451_0__274_), .Q(u2_remHi_274_));
DFFPOSX1 DFFPOSX1_1182 ( .CLK(clk), .D(u2__0remHi_451_0__275_), .Q(u2_remHi_275_));
DFFPOSX1 DFFPOSX1_1183 ( .CLK(clk), .D(u2__0remHi_451_0__276_), .Q(u2_remHi_276_));
DFFPOSX1 DFFPOSX1_1184 ( .CLK(clk), .D(u2__0remHi_451_0__277_), .Q(u2_remHi_277_));
DFFPOSX1 DFFPOSX1_1185 ( .CLK(clk), .D(u2__0remHi_451_0__278_), .Q(u2_remHi_278_));
DFFPOSX1 DFFPOSX1_1186 ( .CLK(clk), .D(u2__0remHi_451_0__279_), .Q(u2_remHi_279_));
DFFPOSX1 DFFPOSX1_1187 ( .CLK(clk), .D(u2__0remHi_451_0__280_), .Q(u2_remHi_280_));
DFFPOSX1 DFFPOSX1_1188 ( .CLK(clk), .D(u2__0remHi_451_0__281_), .Q(u2_remHi_281_));
DFFPOSX1 DFFPOSX1_1189 ( .CLK(clk), .D(u2__0remHi_451_0__282_), .Q(u2_remHi_282_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk), .D(u2__0root_452_0__115_), .Q(sqrto_114_));
DFFPOSX1 DFFPOSX1_1190 ( .CLK(clk), .D(u2__0remHi_451_0__283_), .Q(u2_remHi_283_));
DFFPOSX1 DFFPOSX1_1191 ( .CLK(clk), .D(u2__0remHi_451_0__284_), .Q(u2_remHi_284_));
DFFPOSX1 DFFPOSX1_1192 ( .CLK(clk), .D(u2__0remHi_451_0__285_), .Q(u2_remHi_285_));
DFFPOSX1 DFFPOSX1_1193 ( .CLK(clk), .D(u2__0remHi_451_0__286_), .Q(u2_remHi_286_));
DFFPOSX1 DFFPOSX1_1194 ( .CLK(clk), .D(u2__0remHi_451_0__287_), .Q(u2_remHi_287_));
DFFPOSX1 DFFPOSX1_1195 ( .CLK(clk), .D(u2__0remHi_451_0__288_), .Q(u2_remHi_288_));
DFFPOSX1 DFFPOSX1_1196 ( .CLK(clk), .D(u2__0remHi_451_0__289_), .Q(u2_remHi_289_));
DFFPOSX1 DFFPOSX1_1197 ( .CLK(clk), .D(u2__0remHi_451_0__290_), .Q(u2_remHi_290_));
DFFPOSX1 DFFPOSX1_1198 ( .CLK(clk), .D(u2__0remHi_451_0__291_), .Q(u2_remHi_291_));
DFFPOSX1 DFFPOSX1_1199 ( .CLK(clk), .D(u2__0remHi_451_0__292_), .Q(u2_remHi_292_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(u2__0root_452_0__8_), .Q(sqrto_7_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk), .D(u2__0root_452_0__116_), .Q(sqrto_115_));
DFFPOSX1 DFFPOSX1_1200 ( .CLK(clk), .D(u2__0remHi_451_0__293_), .Q(u2_remHi_293_));
DFFPOSX1 DFFPOSX1_1201 ( .CLK(clk), .D(u2__0remHi_451_0__294_), .Q(u2_remHi_294_));
DFFPOSX1 DFFPOSX1_1202 ( .CLK(clk), .D(u2__0remHi_451_0__295_), .Q(u2_remHi_295_));
DFFPOSX1 DFFPOSX1_1203 ( .CLK(clk), .D(u2__0remHi_451_0__296_), .Q(u2_remHi_296_));
DFFPOSX1 DFFPOSX1_1204 ( .CLK(clk), .D(u2__0remHi_451_0__297_), .Q(u2_remHi_297_));
DFFPOSX1 DFFPOSX1_1205 ( .CLK(clk), .D(u2__0remHi_451_0__298_), .Q(u2_remHi_298_));
DFFPOSX1 DFFPOSX1_1206 ( .CLK(clk), .D(u2__0remHi_451_0__299_), .Q(u2_remHi_299_));
DFFPOSX1 DFFPOSX1_1207 ( .CLK(clk), .D(u2__0remHi_451_0__300_), .Q(u2_remHi_300_));
DFFPOSX1 DFFPOSX1_1208 ( .CLK(clk), .D(u2__0remHi_451_0__301_), .Q(u2_remHi_301_));
DFFPOSX1 DFFPOSX1_1209 ( .CLK(clk), .D(u2__0remHi_451_0__302_), .Q(u2_remHi_302_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk), .D(u2__0root_452_0__117_), .Q(sqrto_116_));
DFFPOSX1 DFFPOSX1_1210 ( .CLK(clk), .D(u2__0remHi_451_0__303_), .Q(u2_remHi_303_));
DFFPOSX1 DFFPOSX1_1211 ( .CLK(clk), .D(u2__0remHi_451_0__304_), .Q(u2_remHi_304_));
DFFPOSX1 DFFPOSX1_1212 ( .CLK(clk), .D(u2__0remHi_451_0__305_), .Q(u2_remHi_305_));
DFFPOSX1 DFFPOSX1_1213 ( .CLK(clk), .D(u2__0remHi_451_0__306_), .Q(u2_remHi_306_));
DFFPOSX1 DFFPOSX1_1214 ( .CLK(clk), .D(u2__0remHi_451_0__307_), .Q(u2_remHi_307_));
DFFPOSX1 DFFPOSX1_1215 ( .CLK(clk), .D(u2__0remHi_451_0__308_), .Q(u2_remHi_308_));
DFFPOSX1 DFFPOSX1_1216 ( .CLK(clk), .D(u2__0remHi_451_0__309_), .Q(u2_remHi_309_));
DFFPOSX1 DFFPOSX1_1217 ( .CLK(clk), .D(u2__0remHi_451_0__310_), .Q(u2_remHi_310_));
DFFPOSX1 DFFPOSX1_1218 ( .CLK(clk), .D(u2__0remHi_451_0__311_), .Q(u2_remHi_311_));
DFFPOSX1 DFFPOSX1_1219 ( .CLK(clk), .D(u2__0remHi_451_0__312_), .Q(u2_remHi_312_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk), .D(u2__0root_452_0__118_), .Q(sqrto_117_));
DFFPOSX1 DFFPOSX1_1220 ( .CLK(clk), .D(u2__0remHi_451_0__313_), .Q(u2_remHi_313_));
DFFPOSX1 DFFPOSX1_1221 ( .CLK(clk), .D(u2__0remHi_451_0__314_), .Q(u2_remHi_314_));
DFFPOSX1 DFFPOSX1_1222 ( .CLK(clk), .D(u2__0remHi_451_0__315_), .Q(u2_remHi_315_));
DFFPOSX1 DFFPOSX1_1223 ( .CLK(clk), .D(u2__0remHi_451_0__316_), .Q(u2_remHi_316_));
DFFPOSX1 DFFPOSX1_1224 ( .CLK(clk), .D(u2__0remHi_451_0__317_), .Q(u2_remHi_317_));
DFFPOSX1 DFFPOSX1_1225 ( .CLK(clk), .D(u2__0remHi_451_0__318_), .Q(u2_remHi_318_));
DFFPOSX1 DFFPOSX1_1226 ( .CLK(clk), .D(u2__0remHi_451_0__319_), .Q(u2_remHi_319_));
DFFPOSX1 DFFPOSX1_1227 ( .CLK(clk), .D(u2__0remHi_451_0__320_), .Q(u2_remHi_320_));
DFFPOSX1 DFFPOSX1_1228 ( .CLK(clk), .D(u2__0remHi_451_0__321_), .Q(u2_remHi_321_));
DFFPOSX1 DFFPOSX1_1229 ( .CLK(clk), .D(u2__0remHi_451_0__322_), .Q(u2_remHi_322_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk), .D(u2__0root_452_0__119_), .Q(sqrto_118_));
DFFPOSX1 DFFPOSX1_1230 ( .CLK(clk), .D(u2__0remHi_451_0__323_), .Q(u2_remHi_323_));
DFFPOSX1 DFFPOSX1_1231 ( .CLK(clk), .D(u2__0remHi_451_0__324_), .Q(u2_remHi_324_));
DFFPOSX1 DFFPOSX1_1232 ( .CLK(clk), .D(u2__0remHi_451_0__325_), .Q(u2_remHi_325_));
DFFPOSX1 DFFPOSX1_1233 ( .CLK(clk), .D(u2__0remHi_451_0__326_), .Q(u2_remHi_326_));
DFFPOSX1 DFFPOSX1_1234 ( .CLK(clk), .D(u2__0remHi_451_0__327_), .Q(u2_remHi_327_));
DFFPOSX1 DFFPOSX1_1235 ( .CLK(clk), .D(u2__0remHi_451_0__328_), .Q(u2_remHi_328_));
DFFPOSX1 DFFPOSX1_1236 ( .CLK(clk), .D(u2__0remHi_451_0__329_), .Q(u2_remHi_329_));
DFFPOSX1 DFFPOSX1_1237 ( .CLK(clk), .D(u2__0remHi_451_0__330_), .Q(u2_remHi_330_));
DFFPOSX1 DFFPOSX1_1238 ( .CLK(clk), .D(u2__0remHi_451_0__331_), .Q(u2_remHi_331_));
DFFPOSX1 DFFPOSX1_1239 ( .CLK(clk), .D(u2__0remHi_451_0__332_), .Q(u2_remHi_332_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk), .D(u2__0root_452_0__120_), .Q(sqrto_119_));
DFFPOSX1 DFFPOSX1_1240 ( .CLK(clk), .D(u2__0remHi_451_0__333_), .Q(u2_remHi_333_));
DFFPOSX1 DFFPOSX1_1241 ( .CLK(clk), .D(u2__0remHi_451_0__334_), .Q(u2_remHi_334_));
DFFPOSX1 DFFPOSX1_1242 ( .CLK(clk), .D(u2__0remHi_451_0__335_), .Q(u2_remHi_335_));
DFFPOSX1 DFFPOSX1_1243 ( .CLK(clk), .D(u2__0remHi_451_0__336_), .Q(u2_remHi_336_));
DFFPOSX1 DFFPOSX1_1244 ( .CLK(clk), .D(u2__0remHi_451_0__337_), .Q(u2_remHi_337_));
DFFPOSX1 DFFPOSX1_1245 ( .CLK(clk), .D(u2__0remHi_451_0__338_), .Q(u2_remHi_338_));
DFFPOSX1 DFFPOSX1_1246 ( .CLK(clk), .D(u2__0remHi_451_0__339_), .Q(u2_remHi_339_));
DFFPOSX1 DFFPOSX1_1247 ( .CLK(clk), .D(u2__0remHi_451_0__340_), .Q(u2_remHi_340_));
DFFPOSX1 DFFPOSX1_1248 ( .CLK(clk), .D(u2__0remHi_451_0__341_), .Q(u2_remHi_341_));
DFFPOSX1 DFFPOSX1_1249 ( .CLK(clk), .D(u2__0remHi_451_0__342_), .Q(u2_remHi_342_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk), .D(u2__0root_452_0__121_), .Q(sqrto_120_));
DFFPOSX1 DFFPOSX1_1250 ( .CLK(clk), .D(u2__0remHi_451_0__343_), .Q(u2_remHi_343_));
DFFPOSX1 DFFPOSX1_1251 ( .CLK(clk), .D(u2__0remHi_451_0__344_), .Q(u2_remHi_344_));
DFFPOSX1 DFFPOSX1_1252 ( .CLK(clk), .D(u2__0remHi_451_0__345_), .Q(u2_remHi_345_));
DFFPOSX1 DFFPOSX1_1253 ( .CLK(clk), .D(u2__0remHi_451_0__346_), .Q(u2_remHi_346_));
DFFPOSX1 DFFPOSX1_1254 ( .CLK(clk), .D(u2__0remHi_451_0__347_), .Q(u2_remHi_347_));
DFFPOSX1 DFFPOSX1_1255 ( .CLK(clk), .D(u2__0remHi_451_0__348_), .Q(u2_remHi_348_));
DFFPOSX1 DFFPOSX1_1256 ( .CLK(clk), .D(u2__0remHi_451_0__349_), .Q(u2_remHi_349_));
DFFPOSX1 DFFPOSX1_1257 ( .CLK(clk), .D(u2__0remHi_451_0__350_), .Q(u2_remHi_350_));
DFFPOSX1 DFFPOSX1_1258 ( .CLK(clk), .D(u2__0remHi_451_0__351_), .Q(u2_remHi_351_));
DFFPOSX1 DFFPOSX1_1259 ( .CLK(clk), .D(u2__0remHi_451_0__352_), .Q(u2_remHi_352_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk), .D(u2__0root_452_0__122_), .Q(sqrto_121_));
DFFPOSX1 DFFPOSX1_1260 ( .CLK(clk), .D(u2__0remHi_451_0__353_), .Q(u2_remHi_353_));
DFFPOSX1 DFFPOSX1_1261 ( .CLK(clk), .D(u2__0remHi_451_0__354_), .Q(u2_remHi_354_));
DFFPOSX1 DFFPOSX1_1262 ( .CLK(clk), .D(u2__0remHi_451_0__355_), .Q(u2_remHi_355_));
DFFPOSX1 DFFPOSX1_1263 ( .CLK(clk), .D(u2__0remHi_451_0__356_), .Q(u2_remHi_356_));
DFFPOSX1 DFFPOSX1_1264 ( .CLK(clk), .D(u2__0remHi_451_0__357_), .Q(u2_remHi_357_));
DFFPOSX1 DFFPOSX1_1265 ( .CLK(clk), .D(u2__0remHi_451_0__358_), .Q(u2_remHi_358_));
DFFPOSX1 DFFPOSX1_1266 ( .CLK(clk), .D(u2__0remHi_451_0__359_), .Q(u2_remHi_359_));
DFFPOSX1 DFFPOSX1_1267 ( .CLK(clk), .D(u2__0remHi_451_0__360_), .Q(u2_remHi_360_));
DFFPOSX1 DFFPOSX1_1268 ( .CLK(clk), .D(u2__0remHi_451_0__361_), .Q(u2_remHi_361_));
DFFPOSX1 DFFPOSX1_1269 ( .CLK(clk), .D(u2__0remHi_451_0__362_), .Q(u2_remHi_362_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk), .D(u2__0root_452_0__123_), .Q(sqrto_122_));
DFFPOSX1 DFFPOSX1_1270 ( .CLK(clk), .D(u2__0remHi_451_0__363_), .Q(u2_remHi_363_));
DFFPOSX1 DFFPOSX1_1271 ( .CLK(clk), .D(u2__0remHi_451_0__364_), .Q(u2_remHi_364_));
DFFPOSX1 DFFPOSX1_1272 ( .CLK(clk), .D(u2__0remHi_451_0__365_), .Q(u2_remHi_365_));
DFFPOSX1 DFFPOSX1_1273 ( .CLK(clk), .D(u2__0remHi_451_0__366_), .Q(u2_remHi_366_));
DFFPOSX1 DFFPOSX1_1274 ( .CLK(clk), .D(u2__0remHi_451_0__367_), .Q(u2_remHi_367_));
DFFPOSX1 DFFPOSX1_1275 ( .CLK(clk), .D(u2__0remHi_451_0__368_), .Q(u2_remHi_368_));
DFFPOSX1 DFFPOSX1_1276 ( .CLK(clk), .D(u2__0remHi_451_0__369_), .Q(u2_remHi_369_));
DFFPOSX1 DFFPOSX1_1277 ( .CLK(clk), .D(u2__0remHi_451_0__370_), .Q(u2_remHi_370_));
DFFPOSX1 DFFPOSX1_1278 ( .CLK(clk), .D(u2__0remHi_451_0__371_), .Q(u2_remHi_371_));
DFFPOSX1 DFFPOSX1_1279 ( .CLK(clk), .D(u2__0remHi_451_0__372_), .Q(u2_remHi_372_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk), .D(u2__0root_452_0__124_), .Q(sqrto_123_));
DFFPOSX1 DFFPOSX1_1280 ( .CLK(clk), .D(u2__0remHi_451_0__373_), .Q(u2_remHi_373_));
DFFPOSX1 DFFPOSX1_1281 ( .CLK(clk), .D(u2__0remHi_451_0__374_), .Q(u2_remHi_374_));
DFFPOSX1 DFFPOSX1_1282 ( .CLK(clk), .D(u2__0remHi_451_0__375_), .Q(u2_remHi_375_));
DFFPOSX1 DFFPOSX1_1283 ( .CLK(clk), .D(u2__0remHi_451_0__376_), .Q(u2_remHi_376_));
DFFPOSX1 DFFPOSX1_1284 ( .CLK(clk), .D(u2__0remHi_451_0__377_), .Q(u2_remHi_377_));
DFFPOSX1 DFFPOSX1_1285 ( .CLK(clk), .D(u2__0remHi_451_0__378_), .Q(u2_remHi_378_));
DFFPOSX1 DFFPOSX1_1286 ( .CLK(clk), .D(u2__0remHi_451_0__379_), .Q(u2_remHi_379_));
DFFPOSX1 DFFPOSX1_1287 ( .CLK(clk), .D(u2__0remHi_451_0__380_), .Q(u2_remHi_380_));
DFFPOSX1 DFFPOSX1_1288 ( .CLK(clk), .D(u2__0remHi_451_0__381_), .Q(u2_remHi_381_));
DFFPOSX1 DFFPOSX1_1289 ( .CLK(clk), .D(u2__0remHi_451_0__382_), .Q(u2_remHi_382_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk), .D(u2__0root_452_0__125_), .Q(sqrto_124_));
DFFPOSX1 DFFPOSX1_1290 ( .CLK(clk), .D(u2__0remHi_451_0__383_), .Q(u2_remHi_383_));
DFFPOSX1 DFFPOSX1_1291 ( .CLK(clk), .D(u2__0remHi_451_0__384_), .Q(u2_remHi_384_));
DFFPOSX1 DFFPOSX1_1292 ( .CLK(clk), .D(u2__0remHi_451_0__385_), .Q(u2_remHi_385_));
DFFPOSX1 DFFPOSX1_1293 ( .CLK(clk), .D(u2__0remHi_451_0__386_), .Q(u2_remHi_386_));
DFFPOSX1 DFFPOSX1_1294 ( .CLK(clk), .D(u2__0remHi_451_0__387_), .Q(u2_remHi_387_));
DFFPOSX1 DFFPOSX1_1295 ( .CLK(clk), .D(u2__0remHi_451_0__388_), .Q(u2_remHi_388_));
DFFPOSX1 DFFPOSX1_1296 ( .CLK(clk), .D(u2__0remHi_451_0__389_), .Q(u2_remHi_389_));
DFFPOSX1 DFFPOSX1_1297 ( .CLK(clk), .D(u2__0remHi_451_0__390_), .Q(u2_remHi_390_));
DFFPOSX1 DFFPOSX1_1298 ( .CLK(clk), .D(u2__0remHi_451_0__391_), .Q(u2_remHi_391_));
DFFPOSX1 DFFPOSX1_1299 ( .CLK(clk), .D(u2__0remHi_451_0__392_), .Q(u2_remHi_392_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(u2__0root_452_0__9_), .Q(sqrto_8_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk), .D(u2__0root_452_0__126_), .Q(sqrto_125_));
DFFPOSX1 DFFPOSX1_1300 ( .CLK(clk), .D(u2__0remHi_451_0__393_), .Q(u2_remHi_393_));
DFFPOSX1 DFFPOSX1_1301 ( .CLK(clk), .D(u2__0remHi_451_0__394_), .Q(u2_remHi_394_));
DFFPOSX1 DFFPOSX1_1302 ( .CLK(clk), .D(u2__0remHi_451_0__395_), .Q(u2_remHi_395_));
DFFPOSX1 DFFPOSX1_1303 ( .CLK(clk), .D(u2__0remHi_451_0__396_), .Q(u2_remHi_396_));
DFFPOSX1 DFFPOSX1_1304 ( .CLK(clk), .D(u2__0remHi_451_0__397_), .Q(u2_remHi_397_));
DFFPOSX1 DFFPOSX1_1305 ( .CLK(clk), .D(u2__0remHi_451_0__398_), .Q(u2_remHi_398_));
DFFPOSX1 DFFPOSX1_1306 ( .CLK(clk), .D(u2__0remHi_451_0__399_), .Q(u2_remHi_399_));
DFFPOSX1 DFFPOSX1_1307 ( .CLK(clk), .D(u2__0remHi_451_0__400_), .Q(u2_remHi_400_));
DFFPOSX1 DFFPOSX1_1308 ( .CLK(clk), .D(u2__0remHi_451_0__401_), .Q(u2_remHi_401_));
DFFPOSX1 DFFPOSX1_1309 ( .CLK(clk), .D(u2__0remHi_451_0__402_), .Q(u2_remHi_402_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk), .D(u2__0root_452_0__127_), .Q(sqrto_126_));
DFFPOSX1 DFFPOSX1_1310 ( .CLK(clk), .D(u2__0remHi_451_0__403_), .Q(u2_remHi_403_));
DFFPOSX1 DFFPOSX1_1311 ( .CLK(clk), .D(u2__0remHi_451_0__404_), .Q(u2_remHi_404_));
DFFPOSX1 DFFPOSX1_1312 ( .CLK(clk), .D(u2__0remHi_451_0__405_), .Q(u2_remHi_405_));
DFFPOSX1 DFFPOSX1_1313 ( .CLK(clk), .D(u2__0remHi_451_0__406_), .Q(u2_remHi_406_));
DFFPOSX1 DFFPOSX1_1314 ( .CLK(clk), .D(u2__0remHi_451_0__407_), .Q(u2_remHi_407_));
DFFPOSX1 DFFPOSX1_1315 ( .CLK(clk), .D(u2__0remHi_451_0__408_), .Q(u2_remHi_408_));
DFFPOSX1 DFFPOSX1_1316 ( .CLK(clk), .D(u2__0remHi_451_0__409_), .Q(u2_remHi_409_));
DFFPOSX1 DFFPOSX1_1317 ( .CLK(clk), .D(u2__0remHi_451_0__410_), .Q(u2_remHi_410_));
DFFPOSX1 DFFPOSX1_1318 ( .CLK(clk), .D(u2__0remHi_451_0__411_), .Q(u2_remHi_411_));
DFFPOSX1 DFFPOSX1_1319 ( .CLK(clk), .D(u2__0remHi_451_0__412_), .Q(u2_remHi_412_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk), .D(u2__0root_452_0__128_), .Q(sqrto_127_));
DFFPOSX1 DFFPOSX1_1320 ( .CLK(clk), .D(u2__0remHi_451_0__413_), .Q(u2_remHi_413_));
DFFPOSX1 DFFPOSX1_1321 ( .CLK(clk), .D(u2__0remHi_451_0__414_), .Q(u2_remHi_414_));
DFFPOSX1 DFFPOSX1_1322 ( .CLK(clk), .D(u2__0remHi_451_0__415_), .Q(u2_remHi_415_));
DFFPOSX1 DFFPOSX1_1323 ( .CLK(clk), .D(u2__0remHi_451_0__416_), .Q(u2_remHi_416_));
DFFPOSX1 DFFPOSX1_1324 ( .CLK(clk), .D(u2__0remHi_451_0__417_), .Q(u2_remHi_417_));
DFFPOSX1 DFFPOSX1_1325 ( .CLK(clk), .D(u2__0remHi_451_0__418_), .Q(u2_remHi_418_));
DFFPOSX1 DFFPOSX1_1326 ( .CLK(clk), .D(u2__0remHi_451_0__419_), .Q(u2_remHi_419_));
DFFPOSX1 DFFPOSX1_1327 ( .CLK(clk), .D(u2__0remHi_451_0__420_), .Q(u2_remHi_420_));
DFFPOSX1 DFFPOSX1_1328 ( .CLK(clk), .D(u2__0remHi_451_0__421_), .Q(u2_remHi_421_));
DFFPOSX1 DFFPOSX1_1329 ( .CLK(clk), .D(u2__0remHi_451_0__422_), .Q(u2_remHi_422_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk), .D(u2__0root_452_0__129_), .Q(sqrto_128_));
DFFPOSX1 DFFPOSX1_1330 ( .CLK(clk), .D(u2__0remHi_451_0__423_), .Q(u2_remHi_423_));
DFFPOSX1 DFFPOSX1_1331 ( .CLK(clk), .D(u2__0remHi_451_0__424_), .Q(u2_remHi_424_));
DFFPOSX1 DFFPOSX1_1332 ( .CLK(clk), .D(u2__0remHi_451_0__425_), .Q(u2_remHi_425_));
DFFPOSX1 DFFPOSX1_1333 ( .CLK(clk), .D(u2__0remHi_451_0__426_), .Q(u2_remHi_426_));
DFFPOSX1 DFFPOSX1_1334 ( .CLK(clk), .D(u2__0remHi_451_0__427_), .Q(u2_remHi_427_));
DFFPOSX1 DFFPOSX1_1335 ( .CLK(clk), .D(u2__0remHi_451_0__428_), .Q(u2_remHi_428_));
DFFPOSX1 DFFPOSX1_1336 ( .CLK(clk), .D(u2__0remHi_451_0__429_), .Q(u2_remHi_429_));
DFFPOSX1 DFFPOSX1_1337 ( .CLK(clk), .D(u2__0remHi_451_0__430_), .Q(u2_remHi_430_));
DFFPOSX1 DFFPOSX1_1338 ( .CLK(clk), .D(u2__0remHi_451_0__431_), .Q(u2_remHi_431_));
DFFPOSX1 DFFPOSX1_1339 ( .CLK(clk), .D(u2__0remHi_451_0__432_), .Q(u2_remHi_432_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk), .D(u2__0root_452_0__130_), .Q(sqrto_129_));
DFFPOSX1 DFFPOSX1_1340 ( .CLK(clk), .D(u2__0remHi_451_0__433_), .Q(u2_remHi_433_));
DFFPOSX1 DFFPOSX1_1341 ( .CLK(clk), .D(u2__0remHi_451_0__434_), .Q(u2_remHi_434_));
DFFPOSX1 DFFPOSX1_1342 ( .CLK(clk), .D(u2__0remHi_451_0__435_), .Q(u2_remHi_435_));
DFFPOSX1 DFFPOSX1_1343 ( .CLK(clk), .D(u2__0remHi_451_0__436_), .Q(u2_remHi_436_));
DFFPOSX1 DFFPOSX1_1344 ( .CLK(clk), .D(u2__0remHi_451_0__437_), .Q(u2_remHi_437_));
DFFPOSX1 DFFPOSX1_1345 ( .CLK(clk), .D(u2__0remHi_451_0__438_), .Q(u2_remHi_438_));
DFFPOSX1 DFFPOSX1_1346 ( .CLK(clk), .D(u2__0remHi_451_0__439_), .Q(u2_remHi_439_));
DFFPOSX1 DFFPOSX1_1347 ( .CLK(clk), .D(u2__0remHi_451_0__440_), .Q(u2_remHi_440_));
DFFPOSX1 DFFPOSX1_1348 ( .CLK(clk), .D(u2__0remHi_451_0__441_), .Q(u2_remHi_441_));
DFFPOSX1 DFFPOSX1_1349 ( .CLK(clk), .D(u2__0remHi_451_0__442_), .Q(u2_remHi_442_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk), .D(u2__0root_452_0__131_), .Q(sqrto_130_));
DFFPOSX1 DFFPOSX1_1350 ( .CLK(clk), .D(u2__0remHi_451_0__443_), .Q(u2_remHi_443_));
DFFPOSX1 DFFPOSX1_1351 ( .CLK(clk), .D(u2__0remHi_451_0__444_), .Q(u2_remHi_444_));
DFFPOSX1 DFFPOSX1_1352 ( .CLK(clk), .D(u2__0remHi_451_0__445_), .Q(u2_remHi_445_));
DFFPOSX1 DFFPOSX1_1353 ( .CLK(clk), .D(u2__0remHi_451_0__446_), .Q(u2_remHi_446_));
DFFPOSX1 DFFPOSX1_1354 ( .CLK(clk), .D(u2__0remHi_451_0__447_), .Q(u2_remHi_447_));
DFFPOSX1 DFFPOSX1_1355 ( .CLK(clk), .D(u2__0remHi_451_0__448_), .Q(u2_remHi_448_));
DFFPOSX1 DFFPOSX1_1356 ( .CLK(clk), .D(u2__0remHi_451_0__449_), .Q(u2_remHi_449_));
DFFPOSX1 DFFPOSX1_1357 ( .CLK(clk), .D(u2__0cnt_7_0__0_), .Q(u2_cnt_0_));
DFFPOSX1 DFFPOSX1_1358 ( .CLK(clk), .D(u2__0cnt_7_0__1_), .Q(u2_cnt_1_));
DFFPOSX1 DFFPOSX1_1359 ( .CLK(clk), .D(u2__0cnt_7_0__2_), .Q(u2_cnt_2_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk), .D(u2__0root_452_0__132_), .Q(sqrto_131_));
DFFPOSX1 DFFPOSX1_1360 ( .CLK(clk), .D(u2__0cnt_7_0__3_), .Q(u2_cnt_3_));
DFFPOSX1 DFFPOSX1_1361 ( .CLK(clk), .D(u2__0cnt_7_0__4_), .Q(u2_cnt_4_));
DFFPOSX1 DFFPOSX1_1362 ( .CLK(clk), .D(u2__0cnt_7_0__5_), .Q(u2_cnt_5_));
DFFPOSX1 DFFPOSX1_1363 ( .CLK(clk), .D(u2__0cnt_7_0__6_), .Q(u2_cnt_6_));
DFFPOSX1 DFFPOSX1_1364 ( .CLK(clk), .D(u2__0cnt_7_0__7_), .Q(u2_cnt_7_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk), .D(u2__0root_452_0__133_), .Q(sqrto_132_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk), .D(u2__0root_452_0__134_), .Q(sqrto_133_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk), .D(u2__0root_452_0__135_), .Q(sqrto_134_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(u2__0root_452_0__10_), .Q(sqrto_9_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk), .D(u2__0root_452_0__136_), .Q(sqrto_135_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk), .D(u2__0root_452_0__137_), .Q(sqrto_136_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk), .D(u2__0root_452_0__138_), .Q(sqrto_137_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk), .D(u2__0root_452_0__139_), .Q(sqrto_138_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk), .D(u2__0root_452_0__140_), .Q(sqrto_139_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk), .D(u2__0root_452_0__141_), .Q(sqrto_140_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk), .D(u2__0root_452_0__142_), .Q(sqrto_141_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk), .D(u2__0root_452_0__143_), .Q(sqrto_142_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk), .D(u2__0root_452_0__144_), .Q(sqrto_143_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk), .D(u2__0root_452_0__145_), .Q(sqrto_144_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(u2__0root_452_0__11_), .Q(sqrto_10_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk), .D(u2__0root_452_0__146_), .Q(sqrto_145_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk), .D(u2__0root_452_0__147_), .Q(sqrto_146_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk), .D(u2__0root_452_0__148_), .Q(sqrto_147_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk), .D(u2__0root_452_0__149_), .Q(sqrto_148_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk), .D(u2__0root_452_0__150_), .Q(sqrto_149_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk), .D(u2__0root_452_0__151_), .Q(sqrto_150_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk), .D(u2__0root_452_0__152_), .Q(sqrto_151_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk), .D(u2__0root_452_0__153_), .Q(sqrto_152_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk), .D(u2__0root_452_0__154_), .Q(sqrto_153_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk), .D(u2__0root_452_0__155_), .Q(sqrto_154_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(u2__0root_452_0__12_), .Q(sqrto_11_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk), .D(u2__0root_452_0__156_), .Q(sqrto_155_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk), .D(u2__0root_452_0__157_), .Q(sqrto_156_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk), .D(u2__0root_452_0__158_), .Q(sqrto_157_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk), .D(u2__0root_452_0__159_), .Q(sqrto_158_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk), .D(u2__0root_452_0__160_), .Q(sqrto_159_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk), .D(u2__0root_452_0__161_), .Q(sqrto_160_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk), .D(u2__0root_452_0__162_), .Q(sqrto_161_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk), .D(u2__0root_452_0__163_), .Q(sqrto_162_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk), .D(u2__0root_452_0__164_), .Q(sqrto_163_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk), .D(u2__0root_452_0__165_), .Q(sqrto_164_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(u2__0root_452_0__13_), .Q(sqrto_12_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk), .D(u2__0root_452_0__166_), .Q(sqrto_165_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk), .D(u2__0root_452_0__167_), .Q(sqrto_166_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk), .D(u2__0root_452_0__168_), .Q(sqrto_167_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk), .D(u2__0root_452_0__169_), .Q(sqrto_168_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk), .D(u2__0root_452_0__170_), .Q(sqrto_169_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk), .D(u2__0root_452_0__171_), .Q(sqrto_170_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk), .D(u2__0root_452_0__172_), .Q(sqrto_171_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk), .D(u2__0root_452_0__173_), .Q(sqrto_172_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk), .D(u2__0root_452_0__174_), .Q(sqrto_173_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk), .D(u2__0root_452_0__175_), .Q(sqrto_174_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(u2__0root_452_0__14_), .Q(sqrto_13_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk), .D(u2__0root_452_0__176_), .Q(sqrto_175_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk), .D(u2__0root_452_0__177_), .Q(sqrto_176_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk), .D(u2__0root_452_0__178_), .Q(sqrto_177_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk), .D(u2__0root_452_0__179_), .Q(sqrto_178_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk), .D(u2__0root_452_0__180_), .Q(sqrto_179_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk), .D(u2__0root_452_0__181_), .Q(sqrto_180_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk), .D(u2__0root_452_0__182_), .Q(sqrto_181_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk), .D(u2__0root_452_0__183_), .Q(sqrto_182_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk), .D(u2__0root_452_0__184_), .Q(sqrto_183_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk), .D(u2__0root_452_0__185_), .Q(sqrto_184_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(u2__0root_452_0__15_), .Q(sqrto_14_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk), .D(u2__0root_452_0__186_), .Q(sqrto_185_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk), .D(u2__0root_452_0__187_), .Q(sqrto_186_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk), .D(u2__0root_452_0__188_), .Q(sqrto_187_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk), .D(u2__0root_452_0__189_), .Q(sqrto_188_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk), .D(u2__0root_452_0__190_), .Q(sqrto_189_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk), .D(u2__0root_452_0__191_), .Q(sqrto_190_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk), .D(u2__0root_452_0__192_), .Q(sqrto_191_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk), .D(u2__0root_452_0__193_), .Q(sqrto_192_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk), .D(u2__0root_452_0__194_), .Q(sqrto_193_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk), .D(u2__0root_452_0__195_), .Q(sqrto_194_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_1_), .Q(done));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(u2__0root_452_0__16_), .Q(sqrto_15_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk), .D(u2__0root_452_0__196_), .Q(sqrto_195_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk), .D(u2__0root_452_0__197_), .Q(sqrto_196_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk), .D(u2__0root_452_0__198_), .Q(sqrto_197_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk), .D(u2__0root_452_0__199_), .Q(sqrto_198_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk), .D(u2__0root_452_0__200_), .Q(sqrto_199_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk), .D(u2__0root_452_0__201_), .Q(sqrto_200_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk), .D(u2__0root_452_0__202_), .Q(sqrto_201_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk), .D(u2__0root_452_0__203_), .Q(sqrto_202_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk), .D(u2__0root_452_0__204_), .Q(sqrto_203_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk), .D(u2__0root_452_0__205_), .Q(sqrto_204_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(u2__0root_452_0__17_), .Q(sqrto_16_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk), .D(u2__0root_452_0__206_), .Q(sqrto_205_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk), .D(u2__0root_452_0__207_), .Q(sqrto_206_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk), .D(u2__0root_452_0__208_), .Q(sqrto_207_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk), .D(u2__0root_452_0__209_), .Q(sqrto_208_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk), .D(u2__0root_452_0__210_), .Q(sqrto_209_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk), .D(u2__0root_452_0__211_), .Q(sqrto_210_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk), .D(u2__0root_452_0__212_), .Q(sqrto_211_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk), .D(u2__0root_452_0__213_), .Q(sqrto_212_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk), .D(u2__0root_452_0__214_), .Q(sqrto_213_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk), .D(u2__0root_452_0__215_), .Q(sqrto_214_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(u2__0root_452_0__18_), .Q(sqrto_17_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk), .D(u2__0root_452_0__216_), .Q(sqrto_215_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk), .D(u2__0root_452_0__217_), .Q(sqrto_216_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk), .D(u2__0root_452_0__218_), .Q(sqrto_217_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk), .D(u2__0root_452_0__219_), .Q(sqrto_218_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk), .D(u2__0root_452_0__220_), .Q(sqrto_219_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk), .D(u2__0root_452_0__221_), .Q(sqrto_220_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk), .D(u2__0root_452_0__222_), .Q(sqrto_221_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk), .D(u2__0root_452_0__223_), .Q(sqrto_222_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk), .D(u2__0root_452_0__224_), .Q(sqrto_223_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk), .D(u2__0root_452_0__225_), .Q(sqrto_224_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(u2__0root_452_0__19_), .Q(sqrto_18_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk), .D(u2__0root_452_0__226_), .Q(sqrto_225_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk), .D(u2__0root_452_0__227_), .Q(u2_o_226_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk), .D(u2__0root_452_0__228_), .Q(u2_o_227_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk), .D(u2__0root_452_0__229_), .Q(u2_o_228_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk), .D(u2__0root_452_0__230_), .Q(u2_o_229_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk), .D(u2__0root_452_0__231_), .Q(u2_o_230_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk), .D(u2__0root_452_0__232_), .Q(u2_o_231_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk), .D(u2__0root_452_0__233_), .Q(u2_o_232_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk), .D(u2__0root_452_0__234_), .Q(u2_o_233_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk), .D(u2__0root_452_0__235_), .Q(u2_o_234_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(u2__0root_452_0__20_), .Q(sqrto_19_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk), .D(u2__0root_452_0__236_), .Q(u2_o_235_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk), .D(u2__0root_452_0__237_), .Q(u2_o_236_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk), .D(u2__0root_452_0__238_), .Q(u2_o_237_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk), .D(u2__0root_452_0__239_), .Q(u2_o_238_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk), .D(u2__0root_452_0__240_), .Q(u2_o_239_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk), .D(u2__0root_452_0__241_), .Q(u2_o_240_));
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk), .D(u2__0root_452_0__242_), .Q(u2_o_241_));
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk), .D(u2__0root_452_0__243_), .Q(u2_o_242_));
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk), .D(u2__0root_452_0__244_), .Q(u2_o_243_));
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk), .D(u2__0root_452_0__245_), .Q(u2_o_244_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(u2__0root_452_0__21_), .Q(sqrto_20_));
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk), .D(u2__0root_452_0__246_), .Q(u2_o_245_));
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk), .D(u2__0root_452_0__247_), .Q(u2_o_246_));
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk), .D(u2__0root_452_0__248_), .Q(u2_o_247_));
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk), .D(u2__0root_452_0__249_), .Q(u2_o_248_));
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk), .D(u2__0root_452_0__250_), .Q(u2_o_249_));
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk), .D(u2__0root_452_0__251_), .Q(u2_o_250_));
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk), .D(u2__0root_452_0__252_), .Q(u2_o_251_));
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk), .D(u2__0root_452_0__253_), .Q(u2_o_252_));
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk), .D(u2__0root_452_0__254_), .Q(u2_o_253_));
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk), .D(u2__0root_452_0__255_), .Q(u2_o_254_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(u2__0root_452_0__22_), .Q(sqrto_21_));
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk), .D(u2__0root_452_0__256_), .Q(u2_o_255_));
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk), .D(u2__0root_452_0__257_), .Q(u2_o_256_));
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk), .D(u2__0root_452_0__258_), .Q(u2_o_257_));
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk), .D(u2__0root_452_0__259_), .Q(u2_o_258_));
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk), .D(u2__0root_452_0__260_), .Q(u2_o_259_));
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk), .D(u2__0root_452_0__261_), .Q(u2_o_260_));
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk), .D(u2__0root_452_0__262_), .Q(u2_o_261_));
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk), .D(u2__0root_452_0__263_), .Q(u2_o_262_));
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk), .D(u2__0root_452_0__264_), .Q(u2_o_263_));
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk), .D(u2__0root_452_0__265_), .Q(u2_o_264_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(u2__0root_452_0__23_), .Q(sqrto_22_));
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk), .D(u2__0root_452_0__266_), .Q(u2_o_265_));
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk), .D(u2__0root_452_0__267_), .Q(u2_o_266_));
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk), .D(u2__0root_452_0__268_), .Q(u2_o_267_));
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk), .D(u2__0root_452_0__269_), .Q(u2_o_268_));
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk), .D(u2__0root_452_0__270_), .Q(u2_o_269_));
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk), .D(u2__0root_452_0__271_), .Q(u2_o_270_));
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk), .D(u2__0root_452_0__272_), .Q(u2_o_271_));
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk), .D(u2__0root_452_0__273_), .Q(u2_o_272_));
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk), .D(u2__0root_452_0__274_), .Q(u2_o_273_));
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk), .D(u2__0root_452_0__275_), .Q(u2_o_274_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(u2__0root_452_0__24_), .Q(sqrto_23_));
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk), .D(u2__0root_452_0__276_), .Q(u2_o_275_));
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk), .D(u2__0root_452_0__277_), .Q(u2_o_276_));
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk), .D(u2__0root_452_0__278_), .Q(u2_o_277_));
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk), .D(u2__0root_452_0__279_), .Q(u2_o_278_));
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk), .D(u2__0root_452_0__280_), .Q(u2_o_279_));
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk), .D(u2__0root_452_0__281_), .Q(u2_o_280_));
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk), .D(u2__0root_452_0__282_), .Q(u2_o_281_));
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk), .D(u2__0root_452_0__283_), .Q(u2_o_282_));
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk), .D(u2__0root_452_0__284_), .Q(u2_o_283_));
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk), .D(u2__0root_452_0__285_), .Q(u2_o_284_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(u2__0root_452_0__25_), .Q(sqrto_24_));
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk), .D(u2__0root_452_0__286_), .Q(u2_o_285_));
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk), .D(u2__0root_452_0__287_), .Q(u2_o_286_));
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk), .D(u2__0root_452_0__288_), .Q(u2_o_287_));
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk), .D(u2__0root_452_0__289_), .Q(u2_o_288_));
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk), .D(u2__0root_452_0__290_), .Q(u2_o_289_));
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk), .D(u2__0root_452_0__291_), .Q(u2_o_290_));
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk), .D(u2__0root_452_0__292_), .Q(u2_o_291_));
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk), .D(u2__0root_452_0__293_), .Q(u2_o_292_));
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk), .D(u2__0root_452_0__294_), .Q(u2_o_293_));
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk), .D(u2__0root_452_0__295_), .Q(u2_o_294_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_2_), .Q(u2_state_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(u2__0root_452_0__26_), .Q(sqrto_25_));
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk), .D(u2__0root_452_0__296_), .Q(u2_o_295_));
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk), .D(u2__0root_452_0__297_), .Q(u2_o_296_));
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk), .D(u2__0root_452_0__298_), .Q(u2_o_297_));
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk), .D(u2__0root_452_0__299_), .Q(u2_o_298_));
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk), .D(u2__0root_452_0__300_), .Q(u2_o_299_));
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk), .D(u2__0root_452_0__301_), .Q(u2_o_300_));
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk), .D(u2__0root_452_0__302_), .Q(u2_o_301_));
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk), .D(u2__0root_452_0__303_), .Q(u2_o_302_));
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk), .D(u2__0root_452_0__304_), .Q(u2_o_303_));
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk), .D(u2__0root_452_0__305_), .Q(u2_o_304_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(u2__0root_452_0__27_), .Q(sqrto_26_));
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk), .D(u2__0root_452_0__306_), .Q(u2_o_305_));
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk), .D(u2__0root_452_0__307_), .Q(u2_o_306_));
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk), .D(u2__0root_452_0__308_), .Q(u2_o_307_));
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk), .D(u2__0root_452_0__309_), .Q(u2_o_308_));
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk), .D(u2__0root_452_0__310_), .Q(u2_o_309_));
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk), .D(u2__0root_452_0__311_), .Q(u2_o_310_));
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk), .D(u2__0root_452_0__312_), .Q(u2_o_311_));
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk), .D(u2__0root_452_0__313_), .Q(u2_o_312_));
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk), .D(u2__0root_452_0__314_), .Q(u2_o_313_));
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk), .D(u2__0root_452_0__315_), .Q(u2_o_314_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(u2__0root_452_0__28_), .Q(sqrto_27_));
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk), .D(u2__0root_452_0__316_), .Q(u2_o_315_));
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk), .D(u2__0root_452_0__317_), .Q(u2_o_316_));
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk), .D(u2__0root_452_0__318_), .Q(u2_o_317_));
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk), .D(u2__0root_452_0__319_), .Q(u2_o_318_));
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk), .D(u2__0root_452_0__320_), .Q(u2_o_319_));
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk), .D(u2__0root_452_0__321_), .Q(u2_o_320_));
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk), .D(u2__0root_452_0__322_), .Q(u2_o_321_));
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk), .D(u2__0root_452_0__323_), .Q(u2_o_322_));
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk), .D(u2__0root_452_0__324_), .Q(u2_o_323_));
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk), .D(u2__0root_452_0__325_), .Q(u2_o_324_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(u2__0root_452_0__29_), .Q(sqrto_28_));
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk), .D(u2__0root_452_0__326_), .Q(u2_o_325_));
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk), .D(u2__0root_452_0__327_), .Q(u2_o_326_));
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk), .D(u2__0root_452_0__328_), .Q(u2_o_327_));
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk), .D(u2__0root_452_0__329_), .Q(u2_o_328_));
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk), .D(u2__0root_452_0__330_), .Q(u2_o_329_));
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk), .D(u2__0root_452_0__331_), .Q(u2_o_330_));
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk), .D(u2__0root_452_0__332_), .Q(u2_o_331_));
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk), .D(u2__0root_452_0__333_), .Q(u2_o_332_));
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk), .D(u2__0root_452_0__334_), .Q(u2_o_333_));
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk), .D(u2__0root_452_0__335_), .Q(u2_o_334_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(u2__0root_452_0__30_), .Q(sqrto_29_));
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk), .D(u2__0root_452_0__336_), .Q(u2_o_335_));
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk), .D(u2__0root_452_0__337_), .Q(u2_o_336_));
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk), .D(u2__0root_452_0__338_), .Q(u2_o_337_));
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk), .D(u2__0root_452_0__339_), .Q(u2_o_338_));
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk), .D(u2__0root_452_0__340_), .Q(u2_o_339_));
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk), .D(u2__0root_452_0__341_), .Q(u2_o_340_));
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk), .D(u2__0root_452_0__342_), .Q(u2_o_341_));
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk), .D(u2__0root_452_0__343_), .Q(u2_o_342_));
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk), .D(u2__0root_452_0__344_), .Q(u2_o_343_));
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk), .D(u2__0root_452_0__345_), .Q(u2_o_344_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(u2__0root_452_0__31_), .Q(sqrto_30_));
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk), .D(u2__0root_452_0__346_), .Q(u2_o_345_));
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk), .D(u2__0root_452_0__347_), .Q(u2_o_346_));
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk), .D(u2__0root_452_0__348_), .Q(u2_o_347_));
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk), .D(u2__0root_452_0__349_), .Q(u2_o_348_));
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk), .D(u2__0root_452_0__350_), .Q(u2_o_349_));
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk), .D(u2__0root_452_0__351_), .Q(u2_o_350_));
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk), .D(u2__0root_452_0__352_), .Q(u2_o_351_));
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk), .D(u2__0root_452_0__353_), .Q(u2_o_352_));
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk), .D(u2__0root_452_0__354_), .Q(u2_o_353_));
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk), .D(u2__0root_452_0__355_), .Q(u2_o_354_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(u2__0root_452_0__32_), .Q(sqrto_31_));
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk), .D(u2__0root_452_0__356_), .Q(u2_o_355_));
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk), .D(u2__0root_452_0__357_), .Q(u2_o_356_));
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk), .D(u2__0root_452_0__358_), .Q(u2_o_357_));
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk), .D(u2__0root_452_0__359_), .Q(u2_o_358_));
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk), .D(u2__0root_452_0__360_), .Q(u2_o_359_));
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk), .D(u2__0root_452_0__361_), .Q(u2_o_360_));
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk), .D(u2__0root_452_0__362_), .Q(u2_o_361_));
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk), .D(u2__0root_452_0__363_), .Q(u2_o_362_));
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk), .D(u2__0root_452_0__364_), .Q(u2_o_363_));
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk), .D(u2__0root_452_0__365_), .Q(u2_o_364_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(u2__0root_452_0__33_), .Q(sqrto_32_));
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk), .D(u2__0root_452_0__366_), .Q(u2_o_365_));
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk), .D(u2__0root_452_0__367_), .Q(u2_o_366_));
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk), .D(u2__0root_452_0__368_), .Q(u2_o_367_));
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk), .D(u2__0root_452_0__369_), .Q(u2_o_368_));
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk), .D(u2__0root_452_0__370_), .Q(u2_o_369_));
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk), .D(u2__0root_452_0__371_), .Q(u2_o_370_));
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk), .D(u2__0root_452_0__372_), .Q(u2_o_371_));
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk), .D(u2__0root_452_0__373_), .Q(u2_o_372_));
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk), .D(u2__0root_452_0__374_), .Q(u2_o_373_));
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk), .D(u2__0root_452_0__375_), .Q(u2_o_374_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(u2__0root_452_0__34_), .Q(sqrto_33_));
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk), .D(u2__0root_452_0__376_), .Q(u2_o_375_));
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk), .D(u2__0root_452_0__377_), .Q(u2_o_376_));
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk), .D(u2__0root_452_0__378_), .Q(u2_o_377_));
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk), .D(u2__0root_452_0__379_), .Q(u2_o_378_));
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk), .D(u2__0root_452_0__380_), .Q(u2_o_379_));
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk), .D(u2__0root_452_0__381_), .Q(u2_o_380_));
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk), .D(u2__0root_452_0__382_), .Q(u2_o_381_));
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk), .D(u2__0root_452_0__383_), .Q(u2_o_382_));
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk), .D(u2__0root_452_0__384_), .Q(u2_o_383_));
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk), .D(u2__0root_452_0__385_), .Q(u2_o_384_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(u2__0root_452_0__35_), .Q(sqrto_34_));
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk), .D(u2__0root_452_0__386_), .Q(u2_o_385_));
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk), .D(u2__0root_452_0__387_), .Q(u2_o_386_));
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk), .D(u2__0root_452_0__388_), .Q(u2_o_387_));
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk), .D(u2__0root_452_0__389_), .Q(u2_o_388_));
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk), .D(u2__0root_452_0__390_), .Q(u2_o_389_));
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk), .D(u2__0root_452_0__391_), .Q(u2_o_390_));
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk), .D(u2__0root_452_0__392_), .Q(u2_o_391_));
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk), .D(u2__0root_452_0__393_), .Q(u2_o_392_));
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk), .D(u2__0root_452_0__394_), .Q(u2_o_393_));
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk), .D(u2__0root_452_0__395_), .Q(u2_o_394_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(u2__0root_452_0__0_), .Q(u2_root_0_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(u2__0root_452_0__36_), .Q(sqrto_35_));
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk), .D(u2__0root_452_0__396_), .Q(u2_o_395_));
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk), .D(u2__0root_452_0__397_), .Q(u2_o_396_));
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk), .D(u2__0root_452_0__398_), .Q(u2_o_397_));
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk), .D(u2__0root_452_0__399_), .Q(u2_o_398_));
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk), .D(u2__0root_452_0__400_), .Q(u2_o_399_));
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk), .D(u2__0root_452_0__401_), .Q(u2_o_400_));
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk), .D(u2__0root_452_0__402_), .Q(u2_o_401_));
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk), .D(u2__0root_452_0__403_), .Q(u2_o_402_));
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk), .D(u2__0root_452_0__404_), .Q(u2_o_403_));
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk), .D(u2__0root_452_0__405_), .Q(u2_o_404_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(u2__0root_452_0__37_), .Q(sqrto_36_));
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk), .D(u2__0root_452_0__406_), .Q(u2_o_405_));
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk), .D(u2__0root_452_0__407_), .Q(u2_o_406_));
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk), .D(u2__0root_452_0__408_), .Q(u2_o_407_));
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk), .D(u2__0root_452_0__409_), .Q(u2_o_408_));
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk), .D(u2__0root_452_0__410_), .Q(u2_o_409_));
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk), .D(u2__0root_452_0__411_), .Q(u2_o_410_));
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk), .D(u2__0root_452_0__412_), .Q(u2_o_411_));
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk), .D(u2__0root_452_0__413_), .Q(u2_o_412_));
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk), .D(u2__0root_452_0__414_), .Q(u2_o_413_));
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk), .D(u2__0root_452_0__415_), .Q(u2_o_414_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(u2__0root_452_0__38_), .Q(sqrto_37_));
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk), .D(u2__0root_452_0__416_), .Q(u2_o_415_));
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk), .D(u2__0root_452_0__417_), .Q(u2_o_416_));
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk), .D(u2__0root_452_0__418_), .Q(u2_o_417_));
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk), .D(u2__0root_452_0__419_), .Q(u2_o_418_));
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk), .D(u2__0root_452_0__420_), .Q(u2_o_419_));
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk), .D(u2__0root_452_0__421_), .Q(u2_o_420_));
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk), .D(u2__0root_452_0__422_), .Q(u2_o_421_));
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk), .D(u2__0root_452_0__423_), .Q(u2_o_422_));
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk), .D(u2__0root_452_0__424_), .Q(u2_o_423_));
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk), .D(u2__0root_452_0__425_), .Q(u2_o_424_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(u2__0root_452_0__39_), .Q(sqrto_38_));
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk), .D(u2__0root_452_0__426_), .Q(u2_o_425_));
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk), .D(u2__0root_452_0__427_), .Q(u2_o_426_));
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk), .D(u2__0root_452_0__428_), .Q(u2_o_427_));
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk), .D(u2__0root_452_0__429_), .Q(u2_o_428_));
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk), .D(u2__0root_452_0__430_), .Q(u2_o_429_));
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk), .D(u2__0root_452_0__431_), .Q(u2_o_430_));
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk), .D(u2__0root_452_0__432_), .Q(u2_o_431_));
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk), .D(u2__0root_452_0__433_), .Q(u2_o_432_));
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk), .D(u2__0root_452_0__434_), .Q(u2_o_433_));
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk), .D(u2__0root_452_0__435_), .Q(u2_o_434_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(u2__0root_452_0__40_), .Q(sqrto_39_));
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk), .D(u2__0root_452_0__436_), .Q(u2_o_435_));
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk), .D(u2__0root_452_0__437_), .Q(u2_o_436_));
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk), .D(u2__0root_452_0__438_), .Q(u2_o_437_));
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk), .D(u2__0root_452_0__439_), .Q(u2_o_438_));
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk), .D(u2__0root_452_0__440_), .Q(u2_o_439_));
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk), .D(u2__0root_452_0__441_), .Q(u2_o_440_));
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk), .D(u2__0root_452_0__442_), .Q(u2_o_441_));
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk), .D(u2__0root_452_0__443_), .Q(u2_o_442_));
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk), .D(u2__0root_452_0__444_), .Q(u2_o_443_));
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk), .D(u2__0root_452_0__445_), .Q(u2_o_444_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(u2__0root_452_0__41_), .Q(sqrto_40_));
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk), .D(u2__0root_452_0__446_), .Q(u2_o_445_));
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk), .D(u2__0root_452_0__447_), .Q(u2_o_446_));
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk), .D(u2__0root_452_0__448_), .Q(u2_o_447_));
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk), .D(u2__0root_452_0__449_), .Q(u2_o_448_));
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk), .D(u2__0root_452_0__450_), .Q(u2_o_449_));
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk), .D(u2__0remLo_451_0__0_), .Q(u2_remLo_0_));
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk), .D(u2__0remLo_451_0__1_), .Q(u2_remLo_1_));
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk), .D(u2__0remLo_451_0__2_), .Q(u2_remLo_2_));
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk), .D(u2__0remLo_451_0__3_), .Q(u2_remLo_3_));
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk), .D(u2__0remLo_451_0__4_), .Q(u2_remLo_4_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(u2__0root_452_0__42_), .Q(sqrto_41_));
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk), .D(u2__0remLo_451_0__5_), .Q(u2_remLo_5_));
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk), .D(u2__0remLo_451_0__6_), .Q(u2_remLo_6_));
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk), .D(u2__0remLo_451_0__7_), .Q(u2_remLo_7_));
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk), .D(u2__0remLo_451_0__8_), .Q(u2_remLo_8_));
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk), .D(u2__0remLo_451_0__9_), .Q(u2_remLo_9_));
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk), .D(u2__0remLo_451_0__10_), .Q(u2_remLo_10_));
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk), .D(u2__0remLo_451_0__11_), .Q(u2_remLo_11_));
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk), .D(u2__0remLo_451_0__12_), .Q(u2_remLo_12_));
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk), .D(u2__0remLo_451_0__13_), .Q(u2_remLo_13_));
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk), .D(u2__0remLo_451_0__14_), .Q(u2_remLo_14_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(u2__0root_452_0__43_), .Q(sqrto_42_));
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk), .D(u2__0remLo_451_0__15_), .Q(u2_remLo_15_));
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk), .D(u2__0remLo_451_0__16_), .Q(u2_remLo_16_));
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk), .D(u2__0remLo_451_0__17_), .Q(u2_remLo_17_));
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk), .D(u2__0remLo_451_0__18_), .Q(u2_remLo_18_));
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk), .D(u2__0remLo_451_0__19_), .Q(u2_remLo_19_));
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk), .D(u2__0remLo_451_0__20_), .Q(u2_remLo_20_));
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk), .D(u2__0remLo_451_0__21_), .Q(u2_remLo_21_));
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk), .D(u2__0remLo_451_0__22_), .Q(u2_remLo_22_));
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk), .D(u2__0remLo_451_0__23_), .Q(u2_remLo_23_));
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk), .D(u2__0remLo_451_0__24_), .Q(u2_remLo_24_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(u2__0root_452_0__44_), .Q(sqrto_43_));
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk), .D(u2__0remLo_451_0__25_), .Q(u2_remLo_25_));
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk), .D(u2__0remLo_451_0__26_), .Q(u2_remLo_26_));
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk), .D(u2__0remLo_451_0__27_), .Q(u2_remLo_27_));
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk), .D(u2__0remLo_451_0__28_), .Q(u2_remLo_28_));
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk), .D(u2__0remLo_451_0__29_), .Q(u2_remLo_29_));
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk), .D(u2__0remLo_451_0__30_), .Q(u2_remLo_30_));
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk), .D(u2__0remLo_451_0__31_), .Q(u2_remLo_31_));
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk), .D(u2__0remLo_451_0__32_), .Q(u2_remLo_32_));
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk), .D(u2__0remLo_451_0__33_), .Q(u2_remLo_33_));
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk), .D(u2__0remLo_451_0__34_), .Q(u2_remLo_34_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(u2__0root_452_0__45_), .Q(sqrto_44_));
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk), .D(u2__0remLo_451_0__35_), .Q(u2_remLo_35_));
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk), .D(u2__0remLo_451_0__36_), .Q(u2_remLo_36_));
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk), .D(u2__0remLo_451_0__37_), .Q(u2_remLo_37_));
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk), .D(u2__0remLo_451_0__38_), .Q(u2_remLo_38_));
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk), .D(u2__0remLo_451_0__39_), .Q(u2_remLo_39_));
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk), .D(u2__0remLo_451_0__40_), .Q(u2_remLo_40_));
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk), .D(u2__0remLo_451_0__41_), .Q(u2_remLo_41_));
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk), .D(u2__0remLo_451_0__42_), .Q(u2_remLo_42_));
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk), .D(u2__0remLo_451_0__43_), .Q(u2_remLo_43_));
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk), .D(u2__0remLo_451_0__44_), .Q(u2_remLo_44_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(u2__0root_452_0__1_), .Q(sqrto_0_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(u2__0root_452_0__46_), .Q(sqrto_45_));
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk), .D(u2__0remLo_451_0__45_), .Q(u2_remLo_45_));
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk), .D(u2__0remLo_451_0__46_), .Q(u2_remLo_46_));
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk), .D(u2__0remLo_451_0__47_), .Q(u2_remLo_47_));
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk), .D(u2__0remLo_451_0__48_), .Q(u2_remLo_48_));
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk), .D(u2__0remLo_451_0__49_), .Q(u2_remLo_49_));
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk), .D(u2__0remLo_451_0__50_), .Q(u2_remLo_50_));
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk), .D(u2__0remLo_451_0__51_), .Q(u2_remLo_51_));
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk), .D(u2__0remLo_451_0__52_), .Q(u2_remLo_52_));
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk), .D(u2__0remLo_451_0__53_), .Q(u2_remLo_53_));
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk), .D(u2__0remLo_451_0__54_), .Q(u2_remLo_54_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(u2__0root_452_0__47_), .Q(sqrto_46_));
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk), .D(u2__0remLo_451_0__55_), .Q(u2_remLo_55_));
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk), .D(u2__0remLo_451_0__56_), .Q(u2_remLo_56_));
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk), .D(u2__0remLo_451_0__57_), .Q(u2_remLo_57_));
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk), .D(u2__0remLo_451_0__58_), .Q(u2_remLo_58_));
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk), .D(u2__0remLo_451_0__59_), .Q(u2_remLo_59_));
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk), .D(u2__0remLo_451_0__60_), .Q(u2_remLo_60_));
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk), .D(u2__0remLo_451_0__61_), .Q(u2_remLo_61_));
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk), .D(u2__0remLo_451_0__62_), .Q(u2_remLo_62_));
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk), .D(u2__0remLo_451_0__63_), .Q(u2_remLo_63_));
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk), .D(u2__0remLo_451_0__64_), .Q(u2_remLo_64_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(u2__0root_452_0__48_), .Q(sqrto_47_));
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk), .D(u2__0remLo_451_0__65_), .Q(u2_remLo_65_));
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk), .D(u2__0remLo_451_0__66_), .Q(u2_remLo_66_));
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk), .D(u2__0remLo_451_0__67_), .Q(u2_remLo_67_));
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk), .D(u2__0remLo_451_0__68_), .Q(u2_remLo_68_));
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk), .D(u2__0remLo_451_0__69_), .Q(u2_remLo_69_));
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk), .D(u2__0remLo_451_0__70_), .Q(u2_remLo_70_));
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk), .D(u2__0remLo_451_0__71_), .Q(u2_remLo_71_));
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk), .D(u2__0remLo_451_0__72_), .Q(u2_remLo_72_));
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk), .D(u2__0remLo_451_0__73_), .Q(u2_remLo_73_));
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk), .D(u2__0remLo_451_0__74_), .Q(u2_remLo_74_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(u2__0root_452_0__49_), .Q(sqrto_48_));
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk), .D(u2__0remLo_451_0__75_), .Q(u2_remLo_75_));
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk), .D(u2__0remLo_451_0__76_), .Q(u2_remLo_76_));
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk), .D(u2__0remLo_451_0__77_), .Q(u2_remLo_77_));
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk), .D(u2__0remLo_451_0__78_), .Q(u2_remLo_78_));
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk), .D(u2__0remLo_451_0__79_), .Q(u2_remLo_79_));
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk), .D(u2__0remLo_451_0__80_), .Q(u2_remLo_80_));
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk), .D(u2__0remLo_451_0__81_), .Q(u2_remLo_81_));
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk), .D(u2__0remLo_451_0__82_), .Q(u2_remLo_82_));
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk), .D(u2__0remLo_451_0__83_), .Q(u2_remLo_83_));
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk), .D(u2__0remLo_451_0__84_), .Q(u2_remLo_84_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(u2__0root_452_0__50_), .Q(sqrto_49_));
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk), .D(u2__0remLo_451_0__85_), .Q(u2_remLo_85_));
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk), .D(u2__0remLo_451_0__86_), .Q(u2_remLo_86_));
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk), .D(u2__0remLo_451_0__87_), .Q(u2_remLo_87_));
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk), .D(u2__0remLo_451_0__88_), .Q(u2_remLo_88_));
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk), .D(u2__0remLo_451_0__89_), .Q(u2_remLo_89_));
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk), .D(u2__0remLo_451_0__90_), .Q(u2_remLo_90_));
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk), .D(u2__0remLo_451_0__91_), .Q(u2_remLo_91_));
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk), .D(u2__0remLo_451_0__92_), .Q(u2_remLo_92_));
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk), .D(u2__0remLo_451_0__93_), .Q(u2_remLo_93_));
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk), .D(u2__0remLo_451_0__94_), .Q(u2_remLo_94_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(u2__0root_452_0__51_), .Q(sqrto_50_));
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk), .D(u2__0remLo_451_0__95_), .Q(u2_remLo_95_));
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk), .D(u2__0remLo_451_0__96_), .Q(u2_remLo_96_));
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk), .D(u2__0remLo_451_0__97_), .Q(u2_remLo_97_));
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk), .D(u2__0remLo_451_0__98_), .Q(u2_remLo_98_));
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk), .D(u2__0remLo_451_0__99_), .Q(u2_remLo_99_));
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk), .D(u2__0remLo_451_0__100_), .Q(u2_remLo_100_));
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk), .D(u2__0remLo_451_0__101_), .Q(u2_remLo_101_));
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk), .D(u2__0remLo_451_0__102_), .Q(u2_remLo_102_));
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk), .D(u2__0remLo_451_0__103_), .Q(u2_remLo_103_));
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk), .D(u2__0remLo_451_0__104_), .Q(u2_remLo_104_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(u2__0root_452_0__52_), .Q(sqrto_51_));
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk), .D(u2__0remLo_451_0__105_), .Q(u2_remLo_105_));
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk), .D(u2__0remLo_451_0__106_), .Q(u2_remLo_106_));
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk), .D(u2__0remLo_451_0__107_), .Q(u2_remLo_107_));
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk), .D(u2__0remLo_451_0__108_), .Q(u2_remLo_108_));
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk), .D(u2__0remLo_451_0__109_), .Q(u2_remLo_109_));
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk), .D(u2__0remLo_451_0__110_), .Q(u2_remLo_110_));
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk), .D(u2__0remLo_451_0__111_), .Q(u2_remLo_111_));
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk), .D(u2__0remLo_451_0__112_), .Q(u2_remLo_112_));
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk), .D(u2__0remLo_451_0__113_), .Q(u2_remLo_113_));
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk), .D(u2__0remLo_451_0__114_), .Q(u2_remLo_114_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(u2__0root_452_0__53_), .Q(sqrto_52_));
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk), .D(u2__0remLo_451_0__115_), .Q(u2_remLo_115_));
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk), .D(u2__0remLo_451_0__116_), .Q(u2_remLo_116_));
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk), .D(u2__0remLo_451_0__117_), .Q(u2_remLo_117_));
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk), .D(u2__0remLo_451_0__118_), .Q(u2_remLo_118_));
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk), .D(u2__0remLo_451_0__119_), .Q(u2_remLo_119_));
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk), .D(u2__0remLo_451_0__120_), .Q(u2_remLo_120_));
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk), .D(u2__0remLo_451_0__121_), .Q(u2_remLo_121_));
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk), .D(u2__0remLo_451_0__122_), .Q(u2_remLo_122_));
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk), .D(u2__0remLo_451_0__123_), .Q(u2_remLo_123_));
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk), .D(u2__0remLo_451_0__124_), .Q(u2_remLo_124_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(u2__0root_452_0__54_), .Q(sqrto_53_));
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk), .D(u2__0remLo_451_0__125_), .Q(u2_remLo_125_));
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk), .D(u2__0remLo_451_0__126_), .Q(u2_remLo_126_));
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk), .D(u2__0remLo_451_0__127_), .Q(u2_remLo_127_));
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk), .D(u2__0remLo_451_0__128_), .Q(u2_remLo_128_));
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk), .D(u2__0remLo_451_0__129_), .Q(u2_remLo_129_));
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk), .D(u2__0remLo_451_0__130_), .Q(u2_remLo_130_));
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk), .D(u2__0remLo_451_0__131_), .Q(u2_remLo_131_));
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk), .D(u2__0remLo_451_0__132_), .Q(u2_remLo_132_));
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk), .D(u2__0remLo_451_0__133_), .Q(u2_remLo_133_));
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk), .D(u2__0remLo_451_0__134_), .Q(u2_remLo_134_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(u2__0root_452_0__55_), .Q(sqrto_54_));
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk), .D(u2__0remLo_451_0__135_), .Q(u2_remLo_135_));
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk), .D(u2__0remLo_451_0__136_), .Q(u2_remLo_136_));
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk), .D(u2__0remLo_451_0__137_), .Q(u2_remLo_137_));
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk), .D(u2__0remLo_451_0__138_), .Q(u2_remLo_138_));
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk), .D(u2__0remLo_451_0__139_), .Q(u2_remLo_139_));
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk), .D(u2__0remLo_451_0__140_), .Q(u2_remLo_140_));
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk), .D(u2__0remLo_451_0__141_), .Q(u2_remLo_141_));
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk), .D(u2__0remLo_451_0__142_), .Q(u2_remLo_142_));
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk), .D(u2__0remLo_451_0__143_), .Q(u2_remLo_143_));
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk), .D(u2__0remLo_451_0__144_), .Q(u2_remLo_144_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(u2__0root_452_0__2_), .Q(sqrto_1_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(u2__0root_452_0__56_), .Q(sqrto_55_));
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk), .D(u2__0remLo_451_0__145_), .Q(u2_remLo_145_));
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk), .D(u2__0remLo_451_0__146_), .Q(u2_remLo_146_));
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk), .D(u2__0remLo_451_0__147_), .Q(u2_remLo_147_));
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk), .D(u2__0remLo_451_0__148_), .Q(u2_remLo_148_));
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk), .D(u2__0remLo_451_0__149_), .Q(u2_remLo_149_));
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk), .D(u2__0remLo_451_0__150_), .Q(u2_remLo_150_));
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk), .D(u2__0remLo_451_0__151_), .Q(u2_remLo_151_));
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk), .D(u2__0remLo_451_0__152_), .Q(u2_remLo_152_));
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk), .D(u2__0remLo_451_0__153_), .Q(u2_remLo_153_));
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk), .D(u2__0remLo_451_0__154_), .Q(u2_remLo_154_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(u2__0root_452_0__57_), .Q(sqrto_56_));
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk), .D(u2__0remLo_451_0__155_), .Q(u2_remLo_155_));
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk), .D(u2__0remLo_451_0__156_), .Q(u2_remLo_156_));
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk), .D(u2__0remLo_451_0__157_), .Q(u2_remLo_157_));
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk), .D(u2__0remLo_451_0__158_), .Q(u2_remLo_158_));
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk), .D(u2__0remLo_451_0__159_), .Q(u2_remLo_159_));
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk), .D(u2__0remLo_451_0__160_), .Q(u2_remLo_160_));
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk), .D(u2__0remLo_451_0__161_), .Q(u2_remLo_161_));
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk), .D(u2__0remLo_451_0__162_), .Q(u2_remLo_162_));
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk), .D(u2__0remLo_451_0__163_), .Q(u2_remLo_163_));
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk), .D(u2__0remLo_451_0__164_), .Q(u2_remLo_164_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(u2__0root_452_0__58_), .Q(sqrto_57_));
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk), .D(u2__0remLo_451_0__165_), .Q(u2_remLo_165_));
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk), .D(u2__0remLo_451_0__166_), .Q(u2_remLo_166_));
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk), .D(u2__0remLo_451_0__167_), .Q(u2_remLo_167_));
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk), .D(u2__0remLo_451_0__168_), .Q(u2_remLo_168_));
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk), .D(u2__0remLo_451_0__169_), .Q(u2_remLo_169_));
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk), .D(u2__0remLo_451_0__170_), .Q(u2_remLo_170_));
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk), .D(u2__0remLo_451_0__171_), .Q(u2_remLo_171_));
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk), .D(u2__0remLo_451_0__172_), .Q(u2_remLo_172_));
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk), .D(u2__0remLo_451_0__173_), .Q(u2_remLo_173_));
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk), .D(u2__0remLo_451_0__174_), .Q(u2_remLo_174_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(u2__0root_452_0__59_), .Q(sqrto_58_));
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk), .D(u2__0remLo_451_0__175_), .Q(u2_remLo_175_));
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk), .D(u2__0remLo_451_0__176_), .Q(u2_remLo_176_));
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk), .D(u2__0remLo_451_0__177_), .Q(u2_remLo_177_));
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk), .D(u2__0remLo_451_0__178_), .Q(u2_remLo_178_));
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk), .D(u2__0remLo_451_0__179_), .Q(u2_remLo_179_));
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk), .D(u2__0remLo_451_0__180_), .Q(u2_remLo_180_));
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk), .D(u2__0remLo_451_0__181_), .Q(u2_remLo_181_));
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk), .D(u2__0remLo_451_0__182_), .Q(u2_remLo_182_));
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk), .D(u2__0remLo_451_0__183_), .Q(u2_remLo_183_));
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk), .D(u2__0remLo_451_0__184_), .Q(u2_remLo_184_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(u2__0root_452_0__60_), .Q(sqrto_59_));
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk), .D(u2__0remLo_451_0__185_), .Q(u2_remLo_185_));
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk), .D(u2__0remLo_451_0__186_), .Q(u2_remLo_186_));
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk), .D(u2__0remLo_451_0__187_), .Q(u2_remLo_187_));
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk), .D(u2__0remLo_451_0__188_), .Q(u2_remLo_188_));
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk), .D(u2__0remLo_451_0__189_), .Q(u2_remLo_189_));
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk), .D(u2__0remLo_451_0__190_), .Q(u2_remLo_190_));
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk), .D(u2__0remLo_451_0__191_), .Q(u2_remLo_191_));
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk), .D(u2__0remLo_451_0__192_), .Q(u2_remLo_192_));
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk), .D(u2__0remLo_451_0__193_), .Q(u2_remLo_193_));
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk), .D(u2__0remLo_451_0__194_), .Q(u2_remLo_194_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk), .D(u2__0root_452_0__61_), .Q(sqrto_60_));
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk), .D(u2__0remLo_451_0__195_), .Q(u2_remLo_195_));
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk), .D(u2__0remLo_451_0__196_), .Q(u2_remLo_196_));
DFFPOSX1 DFFPOSX1_652 ( .CLK(clk), .D(u2__0remLo_451_0__197_), .Q(u2_remLo_197_));
DFFPOSX1 DFFPOSX1_653 ( .CLK(clk), .D(u2__0remLo_451_0__198_), .Q(u2_remLo_198_));
DFFPOSX1 DFFPOSX1_654 ( .CLK(clk), .D(u2__0remLo_451_0__199_), .Q(u2_remLo_199_));
DFFPOSX1 DFFPOSX1_655 ( .CLK(clk), .D(u2__0remLo_451_0__200_), .Q(u2_remLo_200_));
DFFPOSX1 DFFPOSX1_656 ( .CLK(clk), .D(u2__0remLo_451_0__201_), .Q(u2_remLo_201_));
DFFPOSX1 DFFPOSX1_657 ( .CLK(clk), .D(u2__0remLo_451_0__202_), .Q(u2_remLo_202_));
DFFPOSX1 DFFPOSX1_658 ( .CLK(clk), .D(u2__0remLo_451_0__203_), .Q(u2_remLo_203_));
DFFPOSX1 DFFPOSX1_659 ( .CLK(clk), .D(u2__0remLo_451_0__204_), .Q(u2_remLo_204_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk), .D(u2__0root_452_0__62_), .Q(sqrto_61_));
DFFPOSX1 DFFPOSX1_660 ( .CLK(clk), .D(u2__0remLo_451_0__205_), .Q(u2_remLo_205_));
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk), .D(u2__0remLo_451_0__206_), .Q(u2_remLo_206_));
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk), .D(u2__0remLo_451_0__207_), .Q(u2_remLo_207_));
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk), .D(u2__0remLo_451_0__208_), .Q(u2_remLo_208_));
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk), .D(u2__0remLo_451_0__209_), .Q(u2_remLo_209_));
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk), .D(u2__0remLo_451_0__210_), .Q(u2_remLo_210_));
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk), .D(u2__0remLo_451_0__211_), .Q(u2_remLo_211_));
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk), .D(u2__0remLo_451_0__212_), .Q(u2_remLo_212_));
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk), .D(u2__0remLo_451_0__213_), .Q(u2_remLo_213_));
DFFPOSX1 DFFPOSX1_669 ( .CLK(clk), .D(u2__0remLo_451_0__214_), .Q(u2_remLo_214_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk), .D(u2__0root_452_0__63_), .Q(sqrto_62_));
DFFPOSX1 DFFPOSX1_670 ( .CLK(clk), .D(u2__0remLo_451_0__215_), .Q(u2_remLo_215_));
DFFPOSX1 DFFPOSX1_671 ( .CLK(clk), .D(u2__0remLo_451_0__216_), .Q(u2_remLo_216_));
DFFPOSX1 DFFPOSX1_672 ( .CLK(clk), .D(u2__0remLo_451_0__217_), .Q(u2_remLo_217_));
DFFPOSX1 DFFPOSX1_673 ( .CLK(clk), .D(u2__0remLo_451_0__218_), .Q(u2_remLo_218_));
DFFPOSX1 DFFPOSX1_674 ( .CLK(clk), .D(u2__0remLo_451_0__219_), .Q(u2_remLo_219_));
DFFPOSX1 DFFPOSX1_675 ( .CLK(clk), .D(u2__0remLo_451_0__220_), .Q(u2_remLo_220_));
DFFPOSX1 DFFPOSX1_676 ( .CLK(clk), .D(u2__0remLo_451_0__221_), .Q(u2_remLo_221_));
DFFPOSX1 DFFPOSX1_677 ( .CLK(clk), .D(u2__0remLo_451_0__222_), .Q(u2_remLo_222_));
DFFPOSX1 DFFPOSX1_678 ( .CLK(clk), .D(u2__0remLo_451_0__223_), .Q(u2_remLo_223_));
DFFPOSX1 DFFPOSX1_679 ( .CLK(clk), .D(u2__0remLo_451_0__224_), .Q(u2_remLo_224_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk), .D(u2__0root_452_0__64_), .Q(sqrto_63_));
DFFPOSX1 DFFPOSX1_680 ( .CLK(clk), .D(u2__0remLo_451_0__225_), .Q(u2_remLo_225_));
DFFPOSX1 DFFPOSX1_681 ( .CLK(clk), .D(u2__0remLo_451_0__226_), .Q(u2_remLo_226_));
DFFPOSX1 DFFPOSX1_682 ( .CLK(clk), .D(u2__0remLo_451_0__227_), .Q(u2_remLo_227_));
DFFPOSX1 DFFPOSX1_683 ( .CLK(clk), .D(u2__0remLo_451_0__228_), .Q(u2_remLo_228_));
DFFPOSX1 DFFPOSX1_684 ( .CLK(clk), .D(u2__0remLo_451_0__229_), .Q(u2_remLo_229_));
DFFPOSX1 DFFPOSX1_685 ( .CLK(clk), .D(u2__0remLo_451_0__230_), .Q(u2_remLo_230_));
DFFPOSX1 DFFPOSX1_686 ( .CLK(clk), .D(u2__0remLo_451_0__231_), .Q(u2_remLo_231_));
DFFPOSX1 DFFPOSX1_687 ( .CLK(clk), .D(u2__0remLo_451_0__232_), .Q(u2_remLo_232_));
DFFPOSX1 DFFPOSX1_688 ( .CLK(clk), .D(u2__0remLo_451_0__233_), .Q(u2_remLo_233_));
DFFPOSX1 DFFPOSX1_689 ( .CLK(clk), .D(u2__0remLo_451_0__234_), .Q(u2_remLo_234_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk), .D(u2__0root_452_0__65_), .Q(sqrto_64_));
DFFPOSX1 DFFPOSX1_690 ( .CLK(clk), .D(u2__0remLo_451_0__235_), .Q(u2_remLo_235_));
DFFPOSX1 DFFPOSX1_691 ( .CLK(clk), .D(u2__0remLo_451_0__236_), .Q(u2_remLo_236_));
DFFPOSX1 DFFPOSX1_692 ( .CLK(clk), .D(u2__0remLo_451_0__237_), .Q(u2_remLo_237_));
DFFPOSX1 DFFPOSX1_693 ( .CLK(clk), .D(u2__0remLo_451_0__238_), .Q(u2_remLo_238_));
DFFPOSX1 DFFPOSX1_694 ( .CLK(clk), .D(u2__0remLo_451_0__239_), .Q(u2_remLo_239_));
DFFPOSX1 DFFPOSX1_695 ( .CLK(clk), .D(u2__0remLo_451_0__240_), .Q(u2_remLo_240_));
DFFPOSX1 DFFPOSX1_696 ( .CLK(clk), .D(u2__0remLo_451_0__241_), .Q(u2_remLo_241_));
DFFPOSX1 DFFPOSX1_697 ( .CLK(clk), .D(u2__0remLo_451_0__242_), .Q(u2_remLo_242_));
DFFPOSX1 DFFPOSX1_698 ( .CLK(clk), .D(u2__0remLo_451_0__243_), .Q(u2_remLo_243_));
DFFPOSX1 DFFPOSX1_699 ( .CLK(clk), .D(u2__0remLo_451_0__244_), .Q(u2_remLo_244_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(u2__0root_452_0__3_), .Q(sqrto_2_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk), .D(u2__0root_452_0__66_), .Q(sqrto_65_));
DFFPOSX1 DFFPOSX1_700 ( .CLK(clk), .D(u2__0remLo_451_0__245_), .Q(u2_remLo_245_));
DFFPOSX1 DFFPOSX1_701 ( .CLK(clk), .D(u2__0remLo_451_0__246_), .Q(u2_remLo_246_));
DFFPOSX1 DFFPOSX1_702 ( .CLK(clk), .D(u2__0remLo_451_0__247_), .Q(u2_remLo_247_));
DFFPOSX1 DFFPOSX1_703 ( .CLK(clk), .D(u2__0remLo_451_0__248_), .Q(u2_remLo_248_));
DFFPOSX1 DFFPOSX1_704 ( .CLK(clk), .D(u2__0remLo_451_0__249_), .Q(u2_remLo_249_));
DFFPOSX1 DFFPOSX1_705 ( .CLK(clk), .D(u2__0remLo_451_0__250_), .Q(u2_remLo_250_));
DFFPOSX1 DFFPOSX1_706 ( .CLK(clk), .D(u2__0remLo_451_0__251_), .Q(u2_remLo_251_));
DFFPOSX1 DFFPOSX1_707 ( .CLK(clk), .D(u2__0remLo_451_0__252_), .Q(u2_remLo_252_));
DFFPOSX1 DFFPOSX1_708 ( .CLK(clk), .D(u2__0remLo_451_0__253_), .Q(u2_remLo_253_));
DFFPOSX1 DFFPOSX1_709 ( .CLK(clk), .D(u2__0remLo_451_0__254_), .Q(u2_remLo_254_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk), .D(u2__0root_452_0__67_), .Q(sqrto_66_));
DFFPOSX1 DFFPOSX1_710 ( .CLK(clk), .D(u2__0remLo_451_0__255_), .Q(u2_remLo_255_));
DFFPOSX1 DFFPOSX1_711 ( .CLK(clk), .D(u2__0remLo_451_0__256_), .Q(u2_remLo_256_));
DFFPOSX1 DFFPOSX1_712 ( .CLK(clk), .D(u2__0remLo_451_0__257_), .Q(u2_remLo_257_));
DFFPOSX1 DFFPOSX1_713 ( .CLK(clk), .D(u2__0remLo_451_0__258_), .Q(u2_remLo_258_));
DFFPOSX1 DFFPOSX1_714 ( .CLK(clk), .D(u2__0remLo_451_0__259_), .Q(u2_remLo_259_));
DFFPOSX1 DFFPOSX1_715 ( .CLK(clk), .D(u2__0remLo_451_0__260_), .Q(u2_remLo_260_));
DFFPOSX1 DFFPOSX1_716 ( .CLK(clk), .D(u2__0remLo_451_0__261_), .Q(u2_remLo_261_));
DFFPOSX1 DFFPOSX1_717 ( .CLK(clk), .D(u2__0remLo_451_0__262_), .Q(u2_remLo_262_));
DFFPOSX1 DFFPOSX1_718 ( .CLK(clk), .D(u2__0remLo_451_0__263_), .Q(u2_remLo_263_));
DFFPOSX1 DFFPOSX1_719 ( .CLK(clk), .D(u2__0remLo_451_0__264_), .Q(u2_remLo_264_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk), .D(u2__0root_452_0__68_), .Q(sqrto_67_));
DFFPOSX1 DFFPOSX1_720 ( .CLK(clk), .D(u2__0remLo_451_0__265_), .Q(u2_remLo_265_));
DFFPOSX1 DFFPOSX1_721 ( .CLK(clk), .D(u2__0remLo_451_0__266_), .Q(u2_remLo_266_));
DFFPOSX1 DFFPOSX1_722 ( .CLK(clk), .D(u2__0remLo_451_0__267_), .Q(u2_remLo_267_));
DFFPOSX1 DFFPOSX1_723 ( .CLK(clk), .D(u2__0remLo_451_0__268_), .Q(u2_remLo_268_));
DFFPOSX1 DFFPOSX1_724 ( .CLK(clk), .D(u2__0remLo_451_0__269_), .Q(u2_remLo_269_));
DFFPOSX1 DFFPOSX1_725 ( .CLK(clk), .D(u2__0remLo_451_0__270_), .Q(u2_remLo_270_));
DFFPOSX1 DFFPOSX1_726 ( .CLK(clk), .D(u2__0remLo_451_0__271_), .Q(u2_remLo_271_));
DFFPOSX1 DFFPOSX1_727 ( .CLK(clk), .D(u2__0remLo_451_0__272_), .Q(u2_remLo_272_));
DFFPOSX1 DFFPOSX1_728 ( .CLK(clk), .D(u2__0remLo_451_0__273_), .Q(u2_remLo_273_));
DFFPOSX1 DFFPOSX1_729 ( .CLK(clk), .D(u2__0remLo_451_0__274_), .Q(u2_remLo_274_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk), .D(u2__0root_452_0__69_), .Q(sqrto_68_));
DFFPOSX1 DFFPOSX1_730 ( .CLK(clk), .D(u2__0remLo_451_0__275_), .Q(u2_remLo_275_));
DFFPOSX1 DFFPOSX1_731 ( .CLK(clk), .D(u2__0remLo_451_0__276_), .Q(u2_remLo_276_));
DFFPOSX1 DFFPOSX1_732 ( .CLK(clk), .D(u2__0remLo_451_0__277_), .Q(u2_remLo_277_));
DFFPOSX1 DFFPOSX1_733 ( .CLK(clk), .D(u2__0remLo_451_0__278_), .Q(u2_remLo_278_));
DFFPOSX1 DFFPOSX1_734 ( .CLK(clk), .D(u2__0remLo_451_0__279_), .Q(u2_remLo_279_));
DFFPOSX1 DFFPOSX1_735 ( .CLK(clk), .D(u2__0remLo_451_0__280_), .Q(u2_remLo_280_));
DFFPOSX1 DFFPOSX1_736 ( .CLK(clk), .D(u2__0remLo_451_0__281_), .Q(u2_remLo_281_));
DFFPOSX1 DFFPOSX1_737 ( .CLK(clk), .D(u2__0remLo_451_0__282_), .Q(u2_remLo_282_));
DFFPOSX1 DFFPOSX1_738 ( .CLK(clk), .D(u2__0remLo_451_0__283_), .Q(u2_remLo_283_));
DFFPOSX1 DFFPOSX1_739 ( .CLK(clk), .D(u2__0remLo_451_0__284_), .Q(u2_remLo_284_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk), .D(u2__0root_452_0__70_), .Q(sqrto_69_));
DFFPOSX1 DFFPOSX1_740 ( .CLK(clk), .D(u2__0remLo_451_0__285_), .Q(u2_remLo_285_));
DFFPOSX1 DFFPOSX1_741 ( .CLK(clk), .D(u2__0remLo_451_0__286_), .Q(u2_remLo_286_));
DFFPOSX1 DFFPOSX1_742 ( .CLK(clk), .D(u2__0remLo_451_0__287_), .Q(u2_remLo_287_));
DFFPOSX1 DFFPOSX1_743 ( .CLK(clk), .D(u2__0remLo_451_0__288_), .Q(u2_remLo_288_));
DFFPOSX1 DFFPOSX1_744 ( .CLK(clk), .D(u2__0remLo_451_0__289_), .Q(u2_remLo_289_));
DFFPOSX1 DFFPOSX1_745 ( .CLK(clk), .D(u2__0remLo_451_0__290_), .Q(u2_remLo_290_));
DFFPOSX1 DFFPOSX1_746 ( .CLK(clk), .D(u2__0remLo_451_0__291_), .Q(u2_remLo_291_));
DFFPOSX1 DFFPOSX1_747 ( .CLK(clk), .D(u2__0remLo_451_0__292_), .Q(u2_remLo_292_));
DFFPOSX1 DFFPOSX1_748 ( .CLK(clk), .D(u2__0remLo_451_0__293_), .Q(u2_remLo_293_));
DFFPOSX1 DFFPOSX1_749 ( .CLK(clk), .D(u2__0remLo_451_0__294_), .Q(u2_remLo_294_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk), .D(u2__0root_452_0__71_), .Q(sqrto_70_));
DFFPOSX1 DFFPOSX1_750 ( .CLK(clk), .D(u2__0remLo_451_0__295_), .Q(u2_remLo_295_));
DFFPOSX1 DFFPOSX1_751 ( .CLK(clk), .D(u2__0remLo_451_0__296_), .Q(u2_remLo_296_));
DFFPOSX1 DFFPOSX1_752 ( .CLK(clk), .D(u2__0remLo_451_0__297_), .Q(u2_remLo_297_));
DFFPOSX1 DFFPOSX1_753 ( .CLK(clk), .D(u2__0remLo_451_0__298_), .Q(u2_remLo_298_));
DFFPOSX1 DFFPOSX1_754 ( .CLK(clk), .D(u2__0remLo_451_0__299_), .Q(u2_remLo_299_));
DFFPOSX1 DFFPOSX1_755 ( .CLK(clk), .D(u2__0remLo_451_0__300_), .Q(u2_remLo_300_));
DFFPOSX1 DFFPOSX1_756 ( .CLK(clk), .D(u2__0remLo_451_0__301_), .Q(u2_remLo_301_));
DFFPOSX1 DFFPOSX1_757 ( .CLK(clk), .D(u2__0remLo_451_0__302_), .Q(u2_remLo_302_));
DFFPOSX1 DFFPOSX1_758 ( .CLK(clk), .D(u2__0remLo_451_0__303_), .Q(u2_remLo_303_));
DFFPOSX1 DFFPOSX1_759 ( .CLK(clk), .D(u2__0remLo_451_0__304_), .Q(u2_remLo_304_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk), .D(u2__0root_452_0__72_), .Q(sqrto_71_));
DFFPOSX1 DFFPOSX1_760 ( .CLK(clk), .D(u2__0remLo_451_0__305_), .Q(u2_remLo_305_));
DFFPOSX1 DFFPOSX1_761 ( .CLK(clk), .D(u2__0remLo_451_0__306_), .Q(u2_remLo_306_));
DFFPOSX1 DFFPOSX1_762 ( .CLK(clk), .D(u2__0remLo_451_0__307_), .Q(u2_remLo_307_));
DFFPOSX1 DFFPOSX1_763 ( .CLK(clk), .D(u2__0remLo_451_0__308_), .Q(u2_remLo_308_));
DFFPOSX1 DFFPOSX1_764 ( .CLK(clk), .D(u2__0remLo_451_0__309_), .Q(u2_remLo_309_));
DFFPOSX1 DFFPOSX1_765 ( .CLK(clk), .D(u2__0remLo_451_0__310_), .Q(u2_remLo_310_));
DFFPOSX1 DFFPOSX1_766 ( .CLK(clk), .D(u2__0remLo_451_0__311_), .Q(u2_remLo_311_));
DFFPOSX1 DFFPOSX1_767 ( .CLK(clk), .D(u2__0remLo_451_0__312_), .Q(u2_remLo_312_));
DFFPOSX1 DFFPOSX1_768 ( .CLK(clk), .D(u2__0remLo_451_0__313_), .Q(u2_remLo_313_));
DFFPOSX1 DFFPOSX1_769 ( .CLK(clk), .D(u2__0remLo_451_0__314_), .Q(u2_remLo_314_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk), .D(u2__0root_452_0__73_), .Q(sqrto_72_));
DFFPOSX1 DFFPOSX1_770 ( .CLK(clk), .D(u2__0remLo_451_0__315_), .Q(u2_remLo_315_));
DFFPOSX1 DFFPOSX1_771 ( .CLK(clk), .D(u2__0remLo_451_0__316_), .Q(u2_remLo_316_));
DFFPOSX1 DFFPOSX1_772 ( .CLK(clk), .D(u2__0remLo_451_0__317_), .Q(u2_remLo_317_));
DFFPOSX1 DFFPOSX1_773 ( .CLK(clk), .D(u2__0remLo_451_0__318_), .Q(u2_remLo_318_));
DFFPOSX1 DFFPOSX1_774 ( .CLK(clk), .D(u2__0remLo_451_0__319_), .Q(u2_remLo_319_));
DFFPOSX1 DFFPOSX1_775 ( .CLK(clk), .D(u2__0remLo_451_0__320_), .Q(u2_remLo_320_));
DFFPOSX1 DFFPOSX1_776 ( .CLK(clk), .D(u2__0remLo_451_0__321_), .Q(u2_remLo_321_));
DFFPOSX1 DFFPOSX1_777 ( .CLK(clk), .D(u2__0remLo_451_0__322_), .Q(u2_remLo_322_));
DFFPOSX1 DFFPOSX1_778 ( .CLK(clk), .D(u2__0remLo_451_0__323_), .Q(u2_remLo_323_));
DFFPOSX1 DFFPOSX1_779 ( .CLK(clk), .D(u2__0remLo_451_0__324_), .Q(u2_remLo_324_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk), .D(u2__0root_452_0__74_), .Q(sqrto_73_));
DFFPOSX1 DFFPOSX1_780 ( .CLK(clk), .D(u2__0remLo_451_0__325_), .Q(u2_remLo_325_));
DFFPOSX1 DFFPOSX1_781 ( .CLK(clk), .D(u2__0remLo_451_0__326_), .Q(u2_remLo_326_));
DFFPOSX1 DFFPOSX1_782 ( .CLK(clk), .D(u2__0remLo_451_0__327_), .Q(u2_remLo_327_));
DFFPOSX1 DFFPOSX1_783 ( .CLK(clk), .D(u2__0remLo_451_0__328_), .Q(u2_remLo_328_));
DFFPOSX1 DFFPOSX1_784 ( .CLK(clk), .D(u2__0remLo_451_0__329_), .Q(u2_remLo_329_));
DFFPOSX1 DFFPOSX1_785 ( .CLK(clk), .D(u2__0remLo_451_0__330_), .Q(u2_remLo_330_));
DFFPOSX1 DFFPOSX1_786 ( .CLK(clk), .D(u2__0remLo_451_0__331_), .Q(u2_remLo_331_));
DFFPOSX1 DFFPOSX1_787 ( .CLK(clk), .D(u2__0remLo_451_0__332_), .Q(u2_remLo_332_));
DFFPOSX1 DFFPOSX1_788 ( .CLK(clk), .D(u2__0remLo_451_0__333_), .Q(u2_remLo_333_));
DFFPOSX1 DFFPOSX1_789 ( .CLK(clk), .D(u2__0remLo_451_0__334_), .Q(u2_remLo_334_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk), .D(u2__0root_452_0__75_), .Q(sqrto_74_));
DFFPOSX1 DFFPOSX1_790 ( .CLK(clk), .D(u2__0remLo_451_0__335_), .Q(u2_remLo_335_));
DFFPOSX1 DFFPOSX1_791 ( .CLK(clk), .D(u2__0remLo_451_0__336_), .Q(u2_remLo_336_));
DFFPOSX1 DFFPOSX1_792 ( .CLK(clk), .D(u2__0remLo_451_0__337_), .Q(u2_remLo_337_));
DFFPOSX1 DFFPOSX1_793 ( .CLK(clk), .D(u2__0remLo_451_0__338_), .Q(u2_remLo_338_));
DFFPOSX1 DFFPOSX1_794 ( .CLK(clk), .D(u2__0remLo_451_0__339_), .Q(u2_remLo_339_));
DFFPOSX1 DFFPOSX1_795 ( .CLK(clk), .D(u2__0remLo_451_0__340_), .Q(u2_remLo_340_));
DFFPOSX1 DFFPOSX1_796 ( .CLK(clk), .D(u2__0remLo_451_0__341_), .Q(u2_remLo_341_));
DFFPOSX1 DFFPOSX1_797 ( .CLK(clk), .D(u2__0remLo_451_0__342_), .Q(u2_remLo_342_));
DFFPOSX1 DFFPOSX1_798 ( .CLK(clk), .D(u2__0remLo_451_0__343_), .Q(u2_remLo_343_));
DFFPOSX1 DFFPOSX1_799 ( .CLK(clk), .D(u2__0remLo_451_0__344_), .Q(u2_remLo_344_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(u2__0root_452_0__4_), .Q(sqrto_3_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk), .D(u2__0root_452_0__76_), .Q(sqrto_75_));
DFFPOSX1 DFFPOSX1_800 ( .CLK(clk), .D(u2__0remLo_451_0__345_), .Q(u2_remLo_345_));
DFFPOSX1 DFFPOSX1_801 ( .CLK(clk), .D(u2__0remLo_451_0__346_), .Q(u2_remLo_346_));
DFFPOSX1 DFFPOSX1_802 ( .CLK(clk), .D(u2__0remLo_451_0__347_), .Q(u2_remLo_347_));
DFFPOSX1 DFFPOSX1_803 ( .CLK(clk), .D(u2__0remLo_451_0__348_), .Q(u2_remLo_348_));
DFFPOSX1 DFFPOSX1_804 ( .CLK(clk), .D(u2__0remLo_451_0__349_), .Q(u2_remLo_349_));
DFFPOSX1 DFFPOSX1_805 ( .CLK(clk), .D(u2__0remLo_451_0__350_), .Q(u2_remLo_350_));
DFFPOSX1 DFFPOSX1_806 ( .CLK(clk), .D(u2__0remLo_451_0__351_), .Q(u2_remLo_351_));
DFFPOSX1 DFFPOSX1_807 ( .CLK(clk), .D(u2__0remLo_451_0__352_), .Q(u2_remLo_352_));
DFFPOSX1 DFFPOSX1_808 ( .CLK(clk), .D(u2__0remLo_451_0__353_), .Q(u2_remLo_353_));
DFFPOSX1 DFFPOSX1_809 ( .CLK(clk), .D(u2__0remLo_451_0__354_), .Q(u2_remLo_354_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk), .D(u2__0root_452_0__77_), .Q(sqrto_76_));
DFFPOSX1 DFFPOSX1_810 ( .CLK(clk), .D(u2__0remLo_451_0__355_), .Q(u2_remLo_355_));
DFFPOSX1 DFFPOSX1_811 ( .CLK(clk), .D(u2__0remLo_451_0__356_), .Q(u2_remLo_356_));
DFFPOSX1 DFFPOSX1_812 ( .CLK(clk), .D(u2__0remLo_451_0__357_), .Q(u2_remLo_357_));
DFFPOSX1 DFFPOSX1_813 ( .CLK(clk), .D(u2__0remLo_451_0__358_), .Q(u2_remLo_358_));
DFFPOSX1 DFFPOSX1_814 ( .CLK(clk), .D(u2__0remLo_451_0__359_), .Q(u2_remLo_359_));
DFFPOSX1 DFFPOSX1_815 ( .CLK(clk), .D(u2__0remLo_451_0__360_), .Q(u2_remLo_360_));
DFFPOSX1 DFFPOSX1_816 ( .CLK(clk), .D(u2__0remLo_451_0__361_), .Q(u2_remLo_361_));
DFFPOSX1 DFFPOSX1_817 ( .CLK(clk), .D(u2__0remLo_451_0__362_), .Q(u2_remLo_362_));
DFFPOSX1 DFFPOSX1_818 ( .CLK(clk), .D(u2__0remLo_451_0__363_), .Q(u2_remLo_363_));
DFFPOSX1 DFFPOSX1_819 ( .CLK(clk), .D(u2__0remLo_451_0__364_), .Q(u2_remLo_364_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk), .D(u2__0root_452_0__78_), .Q(sqrto_77_));
DFFPOSX1 DFFPOSX1_820 ( .CLK(clk), .D(u2__0remLo_451_0__365_), .Q(u2_remLo_365_));
DFFPOSX1 DFFPOSX1_821 ( .CLK(clk), .D(u2__0remLo_451_0__366_), .Q(u2_remLo_366_));
DFFPOSX1 DFFPOSX1_822 ( .CLK(clk), .D(u2__0remLo_451_0__367_), .Q(u2_remLo_367_));
DFFPOSX1 DFFPOSX1_823 ( .CLK(clk), .D(u2__0remLo_451_0__368_), .Q(u2_remLo_368_));
DFFPOSX1 DFFPOSX1_824 ( .CLK(clk), .D(u2__0remLo_451_0__369_), .Q(u2_remLo_369_));
DFFPOSX1 DFFPOSX1_825 ( .CLK(clk), .D(u2__0remLo_451_0__370_), .Q(u2_remLo_370_));
DFFPOSX1 DFFPOSX1_826 ( .CLK(clk), .D(u2__0remLo_451_0__371_), .Q(u2_remLo_371_));
DFFPOSX1 DFFPOSX1_827 ( .CLK(clk), .D(u2__0remLo_451_0__372_), .Q(u2_remLo_372_));
DFFPOSX1 DFFPOSX1_828 ( .CLK(clk), .D(u2__0remLo_451_0__373_), .Q(u2_remLo_373_));
DFFPOSX1 DFFPOSX1_829 ( .CLK(clk), .D(u2__0remLo_451_0__374_), .Q(u2_remLo_374_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk), .D(u2__0root_452_0__79_), .Q(sqrto_78_));
DFFPOSX1 DFFPOSX1_830 ( .CLK(clk), .D(u2__0remLo_451_0__375_), .Q(u2_remLo_375_));
DFFPOSX1 DFFPOSX1_831 ( .CLK(clk), .D(u2__0remLo_451_0__376_), .Q(u2_remLo_376_));
DFFPOSX1 DFFPOSX1_832 ( .CLK(clk), .D(u2__0remLo_451_0__377_), .Q(u2_remLo_377_));
DFFPOSX1 DFFPOSX1_833 ( .CLK(clk), .D(u2__0remLo_451_0__378_), .Q(u2_remLo_378_));
DFFPOSX1 DFFPOSX1_834 ( .CLK(clk), .D(u2__0remLo_451_0__379_), .Q(u2_remLo_379_));
DFFPOSX1 DFFPOSX1_835 ( .CLK(clk), .D(u2__0remLo_451_0__380_), .Q(u2_remLo_380_));
DFFPOSX1 DFFPOSX1_836 ( .CLK(clk), .D(u2__0remLo_451_0__381_), .Q(u2_remLo_381_));
DFFPOSX1 DFFPOSX1_837 ( .CLK(clk), .D(u2__0remLo_451_0__382_), .Q(u2_remLo_382_));
DFFPOSX1 DFFPOSX1_838 ( .CLK(clk), .D(u2__0remLo_451_0__383_), .Q(u2_remLo_383_));
DFFPOSX1 DFFPOSX1_839 ( .CLK(clk), .D(u2__0remLo_451_0__384_), .Q(u2_remLo_384_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk), .D(u2__0root_452_0__80_), .Q(sqrto_79_));
DFFPOSX1 DFFPOSX1_840 ( .CLK(clk), .D(u2__0remLo_451_0__385_), .Q(u2_remLo_385_));
DFFPOSX1 DFFPOSX1_841 ( .CLK(clk), .D(u2__0remLo_451_0__386_), .Q(u2_remLo_386_));
DFFPOSX1 DFFPOSX1_842 ( .CLK(clk), .D(u2__0remLo_451_0__387_), .Q(u2_remLo_387_));
DFFPOSX1 DFFPOSX1_843 ( .CLK(clk), .D(u2__0remLo_451_0__388_), .Q(u2_remLo_388_));
DFFPOSX1 DFFPOSX1_844 ( .CLK(clk), .D(u2__0remLo_451_0__389_), .Q(u2_remLo_389_));
DFFPOSX1 DFFPOSX1_845 ( .CLK(clk), .D(u2__0remLo_451_0__390_), .Q(u2_remLo_390_));
DFFPOSX1 DFFPOSX1_846 ( .CLK(clk), .D(u2__0remLo_451_0__391_), .Q(u2_remLo_391_));
DFFPOSX1 DFFPOSX1_847 ( .CLK(clk), .D(u2__0remLo_451_0__392_), .Q(u2_remLo_392_));
DFFPOSX1 DFFPOSX1_848 ( .CLK(clk), .D(u2__0remLo_451_0__393_), .Q(u2_remLo_393_));
DFFPOSX1 DFFPOSX1_849 ( .CLK(clk), .D(u2__0remLo_451_0__394_), .Q(u2_remLo_394_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk), .D(u2__0root_452_0__81_), .Q(sqrto_80_));
DFFPOSX1 DFFPOSX1_850 ( .CLK(clk), .D(u2__0remLo_451_0__395_), .Q(u2_remLo_395_));
DFFPOSX1 DFFPOSX1_851 ( .CLK(clk), .D(u2__0remLo_451_0__396_), .Q(u2_remLo_396_));
DFFPOSX1 DFFPOSX1_852 ( .CLK(clk), .D(u2__0remLo_451_0__397_), .Q(u2_remLo_397_));
DFFPOSX1 DFFPOSX1_853 ( .CLK(clk), .D(u2__0remLo_451_0__398_), .Q(u2_remLo_398_));
DFFPOSX1 DFFPOSX1_854 ( .CLK(clk), .D(u2__0remLo_451_0__399_), .Q(u2_remLo_399_));
DFFPOSX1 DFFPOSX1_855 ( .CLK(clk), .D(u2__0remLo_451_0__400_), .Q(u2_remLo_400_));
DFFPOSX1 DFFPOSX1_856 ( .CLK(clk), .D(u2__0remLo_451_0__401_), .Q(u2_remLo_401_));
DFFPOSX1 DFFPOSX1_857 ( .CLK(clk), .D(u2__0remLo_451_0__402_), .Q(u2_remLo_402_));
DFFPOSX1 DFFPOSX1_858 ( .CLK(clk), .D(u2__0remLo_451_0__403_), .Q(u2_remLo_403_));
DFFPOSX1 DFFPOSX1_859 ( .CLK(clk), .D(u2__0remLo_451_0__404_), .Q(u2_remLo_404_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk), .D(u2__0root_452_0__82_), .Q(sqrto_81_));
DFFPOSX1 DFFPOSX1_860 ( .CLK(clk), .D(u2__0remLo_451_0__405_), .Q(u2_remLo_405_));
DFFPOSX1 DFFPOSX1_861 ( .CLK(clk), .D(u2__0remLo_451_0__406_), .Q(u2_remLo_406_));
DFFPOSX1 DFFPOSX1_862 ( .CLK(clk), .D(u2__0remLo_451_0__407_), .Q(u2_remLo_407_));
DFFPOSX1 DFFPOSX1_863 ( .CLK(clk), .D(u2__0remLo_451_0__408_), .Q(u2_remLo_408_));
DFFPOSX1 DFFPOSX1_864 ( .CLK(clk), .D(u2__0remLo_451_0__409_), .Q(u2_remLo_409_));
DFFPOSX1 DFFPOSX1_865 ( .CLK(clk), .D(u2__0remLo_451_0__410_), .Q(u2_remLo_410_));
DFFPOSX1 DFFPOSX1_866 ( .CLK(clk), .D(u2__0remLo_451_0__411_), .Q(u2_remLo_411_));
DFFPOSX1 DFFPOSX1_867 ( .CLK(clk), .D(u2__0remLo_451_0__412_), .Q(u2_remLo_412_));
DFFPOSX1 DFFPOSX1_868 ( .CLK(clk), .D(u2__0remLo_451_0__413_), .Q(u2_remLo_413_));
DFFPOSX1 DFFPOSX1_869 ( .CLK(clk), .D(u2__0remLo_451_0__414_), .Q(u2_remLo_414_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk), .D(u2__0root_452_0__83_), .Q(sqrto_82_));
DFFPOSX1 DFFPOSX1_870 ( .CLK(clk), .D(u2__0remLo_451_0__415_), .Q(u2_remLo_415_));
DFFPOSX1 DFFPOSX1_871 ( .CLK(clk), .D(u2__0remLo_451_0__416_), .Q(u2_remLo_416_));
DFFPOSX1 DFFPOSX1_872 ( .CLK(clk), .D(u2__0remLo_451_0__417_), .Q(u2_remLo_417_));
DFFPOSX1 DFFPOSX1_873 ( .CLK(clk), .D(u2__0remLo_451_0__418_), .Q(u2_remLo_418_));
DFFPOSX1 DFFPOSX1_874 ( .CLK(clk), .D(u2__0remLo_451_0__419_), .Q(u2_remLo_419_));
DFFPOSX1 DFFPOSX1_875 ( .CLK(clk), .D(u2__0remLo_451_0__420_), .Q(u2_remLo_420_));
DFFPOSX1 DFFPOSX1_876 ( .CLK(clk), .D(u2__0remLo_451_0__421_), .Q(u2_remLo_421_));
DFFPOSX1 DFFPOSX1_877 ( .CLK(clk), .D(u2__0remLo_451_0__422_), .Q(u2_remLo_422_));
DFFPOSX1 DFFPOSX1_878 ( .CLK(clk), .D(u2__0remLo_451_0__423_), .Q(u2_remLo_423_));
DFFPOSX1 DFFPOSX1_879 ( .CLK(clk), .D(u2__0remLo_451_0__424_), .Q(u2_remLo_424_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk), .D(u2__0root_452_0__84_), .Q(sqrto_83_));
DFFPOSX1 DFFPOSX1_880 ( .CLK(clk), .D(u2__0remLo_451_0__425_), .Q(u2_remLo_425_));
DFFPOSX1 DFFPOSX1_881 ( .CLK(clk), .D(u2__0remLo_451_0__426_), .Q(u2_remLo_426_));
DFFPOSX1 DFFPOSX1_882 ( .CLK(clk), .D(u2__0remLo_451_0__427_), .Q(u2_remLo_427_));
DFFPOSX1 DFFPOSX1_883 ( .CLK(clk), .D(u2__0remLo_451_0__428_), .Q(u2_remLo_428_));
DFFPOSX1 DFFPOSX1_884 ( .CLK(clk), .D(u2__0remLo_451_0__429_), .Q(u2_remLo_429_));
DFFPOSX1 DFFPOSX1_885 ( .CLK(clk), .D(u2__0remLo_451_0__430_), .Q(u2_remLo_430_));
DFFPOSX1 DFFPOSX1_886 ( .CLK(clk), .D(u2__0remLo_451_0__431_), .Q(u2_remLo_431_));
DFFPOSX1 DFFPOSX1_887 ( .CLK(clk), .D(u2__0remLo_451_0__432_), .Q(u2_remLo_432_));
DFFPOSX1 DFFPOSX1_888 ( .CLK(clk), .D(u2__0remLo_451_0__433_), .Q(u2_remLo_433_));
DFFPOSX1 DFFPOSX1_889 ( .CLK(clk), .D(u2__0remLo_451_0__434_), .Q(u2_remLo_434_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk), .D(u2__0root_452_0__85_), .Q(sqrto_84_));
DFFPOSX1 DFFPOSX1_890 ( .CLK(clk), .D(u2__0remLo_451_0__435_), .Q(u2_remLo_435_));
DFFPOSX1 DFFPOSX1_891 ( .CLK(clk), .D(u2__0remLo_451_0__436_), .Q(u2_remLo_436_));
DFFPOSX1 DFFPOSX1_892 ( .CLK(clk), .D(u2__0remLo_451_0__437_), .Q(u2_remLo_437_));
DFFPOSX1 DFFPOSX1_893 ( .CLK(clk), .D(u2__0remLo_451_0__438_), .Q(u2_remLo_438_));
DFFPOSX1 DFFPOSX1_894 ( .CLK(clk), .D(u2__0remLo_451_0__439_), .Q(u2_remLo_439_));
DFFPOSX1 DFFPOSX1_895 ( .CLK(clk), .D(u2__0remLo_451_0__440_), .Q(u2_remLo_440_));
DFFPOSX1 DFFPOSX1_896 ( .CLK(clk), .D(u2__0remLo_451_0__441_), .Q(u2_remLo_441_));
DFFPOSX1 DFFPOSX1_897 ( .CLK(clk), .D(u2__0remLo_451_0__442_), .Q(u2_remLo_442_));
DFFPOSX1 DFFPOSX1_898 ( .CLK(clk), .D(u2__0remLo_451_0__443_), .Q(u2_remLo_443_));
DFFPOSX1 DFFPOSX1_899 ( .CLK(clk), .D(u2__0remLo_451_0__444_), .Q(u2_remLo_444_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(u2__0root_452_0__5_), .Q(sqrto_4_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk), .D(u2__0root_452_0__86_), .Q(sqrto_85_));
DFFPOSX1 DFFPOSX1_900 ( .CLK(clk), .D(u2__0remLo_451_0__445_), .Q(u2_remLo_445_));
DFFPOSX1 DFFPOSX1_901 ( .CLK(clk), .D(u2__0remLo_451_0__446_), .Q(u2_remLo_446_));
DFFPOSX1 DFFPOSX1_902 ( .CLK(clk), .D(u2__0remLo_451_0__447_), .Q(u2_remLo_447_));
DFFPOSX1 DFFPOSX1_903 ( .CLK(clk), .D(u2__0remLo_451_0__448_), .Q(u2_remLo_448_));
DFFPOSX1 DFFPOSX1_904 ( .CLK(clk), .D(u2__0remLo_451_0__449_), .Q(u2_remLo_449_));
DFFPOSX1 DFFPOSX1_905 ( .CLK(clk), .D(u2__0remLo_451_0__450_), .Q(u2_remHiShift_0_));
DFFPOSX1 DFFPOSX1_906 ( .CLK(clk), .D(u2__0remLo_451_0__451_), .Q(u2_remHiShift_1_));
DFFPOSX1 DFFPOSX1_907 ( .CLK(clk), .D(u2__0remHi_451_0__0_), .Q(u2_remHi_0_));
DFFPOSX1 DFFPOSX1_908 ( .CLK(clk), .D(u2__0remHi_451_0__1_), .Q(u2_remHi_1_));
DFFPOSX1 DFFPOSX1_909 ( .CLK(clk), .D(u2__0remHi_451_0__2_), .Q(u2_remHi_2_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk), .D(u2__0root_452_0__87_), .Q(sqrto_86_));
DFFPOSX1 DFFPOSX1_910 ( .CLK(clk), .D(u2__0remHi_451_0__3_), .Q(u2_remHi_3_));
DFFPOSX1 DFFPOSX1_911 ( .CLK(clk), .D(u2__0remHi_451_0__4_), .Q(u2_remHi_4_));
DFFPOSX1 DFFPOSX1_912 ( .CLK(clk), .D(u2__0remHi_451_0__5_), .Q(u2_remHi_5_));
DFFPOSX1 DFFPOSX1_913 ( .CLK(clk), .D(u2__0remHi_451_0__6_), .Q(u2_remHi_6_));
DFFPOSX1 DFFPOSX1_914 ( .CLK(clk), .D(u2__0remHi_451_0__7_), .Q(u2_remHi_7_));
DFFPOSX1 DFFPOSX1_915 ( .CLK(clk), .D(u2__0remHi_451_0__8_), .Q(u2_remHi_8_));
DFFPOSX1 DFFPOSX1_916 ( .CLK(clk), .D(u2__0remHi_451_0__9_), .Q(u2_remHi_9_));
DFFPOSX1 DFFPOSX1_917 ( .CLK(clk), .D(u2__0remHi_451_0__10_), .Q(u2_remHi_10_));
DFFPOSX1 DFFPOSX1_918 ( .CLK(clk), .D(u2__0remHi_451_0__11_), .Q(u2_remHi_11_));
DFFPOSX1 DFFPOSX1_919 ( .CLK(clk), .D(u2__0remHi_451_0__12_), .Q(u2_remHi_12_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk), .D(u2__0root_452_0__88_), .Q(sqrto_87_));
DFFPOSX1 DFFPOSX1_920 ( .CLK(clk), .D(u2__0remHi_451_0__13_), .Q(u2_remHi_13_));
DFFPOSX1 DFFPOSX1_921 ( .CLK(clk), .D(u2__0remHi_451_0__14_), .Q(u2_remHi_14_));
DFFPOSX1 DFFPOSX1_922 ( .CLK(clk), .D(u2__0remHi_451_0__15_), .Q(u2_remHi_15_));
DFFPOSX1 DFFPOSX1_923 ( .CLK(clk), .D(u2__0remHi_451_0__16_), .Q(u2_remHi_16_));
DFFPOSX1 DFFPOSX1_924 ( .CLK(clk), .D(u2__0remHi_451_0__17_), .Q(u2_remHi_17_));
DFFPOSX1 DFFPOSX1_925 ( .CLK(clk), .D(u2__0remHi_451_0__18_), .Q(u2_remHi_18_));
DFFPOSX1 DFFPOSX1_926 ( .CLK(clk), .D(u2__0remHi_451_0__19_), .Q(u2_remHi_19_));
DFFPOSX1 DFFPOSX1_927 ( .CLK(clk), .D(u2__0remHi_451_0__20_), .Q(u2_remHi_20_));
DFFPOSX1 DFFPOSX1_928 ( .CLK(clk), .D(u2__0remHi_451_0__21_), .Q(u2_remHi_21_));
DFFPOSX1 DFFPOSX1_929 ( .CLK(clk), .D(u2__0remHi_451_0__22_), .Q(u2_remHi_22_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk), .D(u2__0root_452_0__89_), .Q(sqrto_88_));
DFFPOSX1 DFFPOSX1_930 ( .CLK(clk), .D(u2__0remHi_451_0__23_), .Q(u2_remHi_23_));
DFFPOSX1 DFFPOSX1_931 ( .CLK(clk), .D(u2__0remHi_451_0__24_), .Q(u2_remHi_24_));
DFFPOSX1 DFFPOSX1_932 ( .CLK(clk), .D(u2__0remHi_451_0__25_), .Q(u2_remHi_25_));
DFFPOSX1 DFFPOSX1_933 ( .CLK(clk), .D(u2__0remHi_451_0__26_), .Q(u2_remHi_26_));
DFFPOSX1 DFFPOSX1_934 ( .CLK(clk), .D(u2__0remHi_451_0__27_), .Q(u2_remHi_27_));
DFFPOSX1 DFFPOSX1_935 ( .CLK(clk), .D(u2__0remHi_451_0__28_), .Q(u2_remHi_28_));
DFFPOSX1 DFFPOSX1_936 ( .CLK(clk), .D(u2__0remHi_451_0__29_), .Q(u2_remHi_29_));
DFFPOSX1 DFFPOSX1_937 ( .CLK(clk), .D(u2__0remHi_451_0__30_), .Q(u2_remHi_30_));
DFFPOSX1 DFFPOSX1_938 ( .CLK(clk), .D(u2__0remHi_451_0__31_), .Q(u2_remHi_31_));
DFFPOSX1 DFFPOSX1_939 ( .CLK(clk), .D(u2__0remHi_451_0__32_), .Q(u2_remHi_32_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk), .D(u2__0root_452_0__90_), .Q(sqrto_89_));
DFFPOSX1 DFFPOSX1_940 ( .CLK(clk), .D(u2__0remHi_451_0__33_), .Q(u2_remHi_33_));
DFFPOSX1 DFFPOSX1_941 ( .CLK(clk), .D(u2__0remHi_451_0__34_), .Q(u2_remHi_34_));
DFFPOSX1 DFFPOSX1_942 ( .CLK(clk), .D(u2__0remHi_451_0__35_), .Q(u2_remHi_35_));
DFFPOSX1 DFFPOSX1_943 ( .CLK(clk), .D(u2__0remHi_451_0__36_), .Q(u2_remHi_36_));
DFFPOSX1 DFFPOSX1_944 ( .CLK(clk), .D(u2__0remHi_451_0__37_), .Q(u2_remHi_37_));
DFFPOSX1 DFFPOSX1_945 ( .CLK(clk), .D(u2__0remHi_451_0__38_), .Q(u2_remHi_38_));
DFFPOSX1 DFFPOSX1_946 ( .CLK(clk), .D(u2__0remHi_451_0__39_), .Q(u2_remHi_39_));
DFFPOSX1 DFFPOSX1_947 ( .CLK(clk), .D(u2__0remHi_451_0__40_), .Q(u2_remHi_40_));
DFFPOSX1 DFFPOSX1_948 ( .CLK(clk), .D(u2__0remHi_451_0__41_), .Q(u2_remHi_41_));
DFFPOSX1 DFFPOSX1_949 ( .CLK(clk), .D(u2__0remHi_451_0__42_), .Q(u2_remHi_42_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk), .D(u2__0root_452_0__91_), .Q(sqrto_90_));
DFFPOSX1 DFFPOSX1_950 ( .CLK(clk), .D(u2__0remHi_451_0__43_), .Q(u2_remHi_43_));
DFFPOSX1 DFFPOSX1_951 ( .CLK(clk), .D(u2__0remHi_451_0__44_), .Q(u2_remHi_44_));
DFFPOSX1 DFFPOSX1_952 ( .CLK(clk), .D(u2__0remHi_451_0__45_), .Q(u2_remHi_45_));
DFFPOSX1 DFFPOSX1_953 ( .CLK(clk), .D(u2__0remHi_451_0__46_), .Q(u2_remHi_46_));
DFFPOSX1 DFFPOSX1_954 ( .CLK(clk), .D(u2__0remHi_451_0__47_), .Q(u2_remHi_47_));
DFFPOSX1 DFFPOSX1_955 ( .CLK(clk), .D(u2__0remHi_451_0__48_), .Q(u2_remHi_48_));
DFFPOSX1 DFFPOSX1_956 ( .CLK(clk), .D(u2__0remHi_451_0__49_), .Q(u2_remHi_49_));
DFFPOSX1 DFFPOSX1_957 ( .CLK(clk), .D(u2__0remHi_451_0__50_), .Q(u2_remHi_50_));
DFFPOSX1 DFFPOSX1_958 ( .CLK(clk), .D(u2__0remHi_451_0__51_), .Q(u2_remHi_51_));
DFFPOSX1 DFFPOSX1_959 ( .CLK(clk), .D(u2__0remHi_451_0__52_), .Q(u2_remHi_52_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk), .D(u2__0root_452_0__92_), .Q(sqrto_91_));
DFFPOSX1 DFFPOSX1_960 ( .CLK(clk), .D(u2__0remHi_451_0__53_), .Q(u2_remHi_53_));
DFFPOSX1 DFFPOSX1_961 ( .CLK(clk), .D(u2__0remHi_451_0__54_), .Q(u2_remHi_54_));
DFFPOSX1 DFFPOSX1_962 ( .CLK(clk), .D(u2__0remHi_451_0__55_), .Q(u2_remHi_55_));
DFFPOSX1 DFFPOSX1_963 ( .CLK(clk), .D(u2__0remHi_451_0__56_), .Q(u2_remHi_56_));
DFFPOSX1 DFFPOSX1_964 ( .CLK(clk), .D(u2__0remHi_451_0__57_), .Q(u2_remHi_57_));
DFFPOSX1 DFFPOSX1_965 ( .CLK(clk), .D(u2__0remHi_451_0__58_), .Q(u2_remHi_58_));
DFFPOSX1 DFFPOSX1_966 ( .CLK(clk), .D(u2__0remHi_451_0__59_), .Q(u2_remHi_59_));
DFFPOSX1 DFFPOSX1_967 ( .CLK(clk), .D(u2__0remHi_451_0__60_), .Q(u2_remHi_60_));
DFFPOSX1 DFFPOSX1_968 ( .CLK(clk), .D(u2__0remHi_451_0__61_), .Q(u2_remHi_61_));
DFFPOSX1 DFFPOSX1_969 ( .CLK(clk), .D(u2__0remHi_451_0__62_), .Q(u2_remHi_62_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk), .D(u2__0root_452_0__93_), .Q(sqrto_92_));
DFFPOSX1 DFFPOSX1_970 ( .CLK(clk), .D(u2__0remHi_451_0__63_), .Q(u2_remHi_63_));
DFFPOSX1 DFFPOSX1_971 ( .CLK(clk), .D(u2__0remHi_451_0__64_), .Q(u2_remHi_64_));
DFFPOSX1 DFFPOSX1_972 ( .CLK(clk), .D(u2__0remHi_451_0__65_), .Q(u2_remHi_65_));
DFFPOSX1 DFFPOSX1_973 ( .CLK(clk), .D(u2__0remHi_451_0__66_), .Q(u2_remHi_66_));
DFFPOSX1 DFFPOSX1_974 ( .CLK(clk), .D(u2__0remHi_451_0__67_), .Q(u2_remHi_67_));
DFFPOSX1 DFFPOSX1_975 ( .CLK(clk), .D(u2__0remHi_451_0__68_), .Q(u2_remHi_68_));
DFFPOSX1 DFFPOSX1_976 ( .CLK(clk), .D(u2__0remHi_451_0__69_), .Q(u2_remHi_69_));
DFFPOSX1 DFFPOSX1_977 ( .CLK(clk), .D(u2__0remHi_451_0__70_), .Q(u2_remHi_70_));
DFFPOSX1 DFFPOSX1_978 ( .CLK(clk), .D(u2__0remHi_451_0__71_), .Q(u2_remHi_71_));
DFFPOSX1 DFFPOSX1_979 ( .CLK(clk), .D(u2__0remHi_451_0__72_), .Q(u2_remHi_72_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk), .D(u2__0root_452_0__94_), .Q(sqrto_93_));
DFFPOSX1 DFFPOSX1_980 ( .CLK(clk), .D(u2__0remHi_451_0__73_), .Q(u2_remHi_73_));
DFFPOSX1 DFFPOSX1_981 ( .CLK(clk), .D(u2__0remHi_451_0__74_), .Q(u2_remHi_74_));
DFFPOSX1 DFFPOSX1_982 ( .CLK(clk), .D(u2__0remHi_451_0__75_), .Q(u2_remHi_75_));
DFFPOSX1 DFFPOSX1_983 ( .CLK(clk), .D(u2__0remHi_451_0__76_), .Q(u2_remHi_76_));
DFFPOSX1 DFFPOSX1_984 ( .CLK(clk), .D(u2__0remHi_451_0__77_), .Q(u2_remHi_77_));
DFFPOSX1 DFFPOSX1_985 ( .CLK(clk), .D(u2__0remHi_451_0__78_), .Q(u2_remHi_78_));
DFFPOSX1 DFFPOSX1_986 ( .CLK(clk), .D(u2__0remHi_451_0__79_), .Q(u2_remHi_79_));
DFFPOSX1 DFFPOSX1_987 ( .CLK(clk), .D(u2__0remHi_451_0__80_), .Q(u2_remHi_80_));
DFFPOSX1 DFFPOSX1_988 ( .CLK(clk), .D(u2__0remHi_451_0__81_), .Q(u2_remHi_81_));
DFFPOSX1 DFFPOSX1_989 ( .CLK(clk), .D(u2__0remHi_451_0__82_), .Q(u2_remHi_82_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk), .D(u2__0root_452_0__95_), .Q(sqrto_94_));
DFFPOSX1 DFFPOSX1_990 ( .CLK(clk), .D(u2__0remHi_451_0__83_), .Q(u2_remHi_83_));
DFFPOSX1 DFFPOSX1_991 ( .CLK(clk), .D(u2__0remHi_451_0__84_), .Q(u2_remHi_84_));
DFFPOSX1 DFFPOSX1_992 ( .CLK(clk), .D(u2__0remHi_451_0__85_), .Q(u2_remHi_85_));
DFFPOSX1 DFFPOSX1_993 ( .CLK(clk), .D(u2__0remHi_451_0__86_), .Q(u2_remHi_86_));
DFFPOSX1 DFFPOSX1_994 ( .CLK(clk), .D(u2__0remHi_451_0__87_), .Q(u2_remHi_87_));
DFFPOSX1 DFFPOSX1_995 ( .CLK(clk), .D(u2__0remHi_451_0__88_), .Q(u2_remHi_88_));
DFFPOSX1 DFFPOSX1_996 ( .CLK(clk), .D(u2__0remHi_451_0__89_), .Q(u2_remHi_89_));
DFFPOSX1 DFFPOSX1_997 ( .CLK(clk), .D(u2__0remHi_451_0__90_), .Q(u2_remHi_90_));
DFFPOSX1 DFFPOSX1_998 ( .CLK(clk), .D(u2__0remHi_451_0__91_), .Q(u2_remHi_91_));
DFFPOSX1 DFFPOSX1_999 ( .CLK(clk), .D(u2__0remHi_451_0__92_), .Q(u2_remHi_92_));
INVX1 INVX1_1 ( .A(aNan), .Y(_abc_65734_new_n753_));
INVX1 INVX1_10 ( .A(sqrto_84_), .Y(_abc_65734_new_n854_));
INVX1 INVX1_100 ( .A(sqrto_174_), .Y(_abc_65734_new_n1124_));
INVX1 INVX1_1000 ( .A(u2_remHi_304_), .Y(u2__abc_52138_new_n5418_));
INVX1 INVX1_1001 ( .A(u2_o_304_), .Y(u2__abc_52138_new_n5420_));
INVX1 INVX1_1002 ( .A(u2_remHi_305_), .Y(u2__abc_52138_new_n5423_));
INVX1 INVX1_1003 ( .A(u2_o_305_), .Y(u2__abc_52138_new_n5425_));
INVX1 INVX1_1004 ( .A(u2_remHi_308_), .Y(u2__abc_52138_new_n5430_));
INVX1 INVX1_1005 ( .A(u2_o_308_), .Y(u2__abc_52138_new_n5432_));
INVX1 INVX1_1006 ( .A(u2_remHi_309_), .Y(u2__abc_52138_new_n5435_));
INVX1 INVX1_1007 ( .A(u2_o_309_), .Y(u2__abc_52138_new_n5437_));
INVX1 INVX1_1008 ( .A(u2_remHi_307_), .Y(u2__abc_52138_new_n5441_));
INVX1 INVX1_1009 ( .A(u2_o_307_), .Y(u2__abc_52138_new_n5443_));
INVX1 INVX1_101 ( .A(sqrto_175_), .Y(_abc_65734_new_n1127_));
INVX1 INVX1_1010 ( .A(u2_remHi_306_), .Y(u2__abc_52138_new_n5446_));
INVX1 INVX1_1011 ( .A(u2_o_306_), .Y(u2__abc_52138_new_n5448_));
INVX1 INVX1_1012 ( .A(u2_o_294_), .Y(u2__abc_52138_new_n5455_));
INVX1 INVX1_1013 ( .A(u2_remHi_294_), .Y(u2__abc_52138_new_n5457_));
INVX1 INVX1_1014 ( .A(u2_remHi_295_), .Y(u2__abc_52138_new_n5460_));
INVX1 INVX1_1015 ( .A(u2_o_295_), .Y(u2__abc_52138_new_n5462_));
INVX1 INVX1_1016 ( .A(u2_remHi_296_), .Y(u2__abc_52138_new_n5466_));
INVX1 INVX1_1017 ( .A(u2_o_296_), .Y(u2__abc_52138_new_n5468_));
INVX1 INVX1_1018 ( .A(u2_remHi_297_), .Y(u2__abc_52138_new_n5471_));
INVX1 INVX1_1019 ( .A(u2_o_297_), .Y(u2__abc_52138_new_n5473_));
INVX1 INVX1_102 ( .A(sqrto_176_), .Y(_abc_65734_new_n1130_));
INVX1 INVX1_1020 ( .A(u2_remHi_300_), .Y(u2__abc_52138_new_n5478_));
INVX1 INVX1_1021 ( .A(u2_o_300_), .Y(u2__abc_52138_new_n5480_));
INVX1 INVX1_1022 ( .A(u2_remHi_301_), .Y(u2__abc_52138_new_n5483_));
INVX1 INVX1_1023 ( .A(u2_o_301_), .Y(u2__abc_52138_new_n5485_));
INVX1 INVX1_1024 ( .A(u2_remHi_298_), .Y(u2__abc_52138_new_n5489_));
INVX1 INVX1_1025 ( .A(u2_o_298_), .Y(u2__abc_52138_new_n5491_));
INVX1 INVX1_1026 ( .A(u2_remHi_299_), .Y(u2__abc_52138_new_n5494_));
INVX1 INVX1_1027 ( .A(u2_o_299_), .Y(u2__abc_52138_new_n5496_));
INVX1 INVX1_1028 ( .A(u2_remHi_288_), .Y(u2__abc_52138_new_n5502_));
INVX1 INVX1_1029 ( .A(u2_o_288_), .Y(u2__abc_52138_new_n5504_));
INVX1 INVX1_103 ( .A(sqrto_177_), .Y(_abc_65734_new_n1133_));
INVX1 INVX1_1030 ( .A(u2_remHi_289_), .Y(u2__abc_52138_new_n5507_));
INVX1 INVX1_1031 ( .A(u2_o_289_), .Y(u2__abc_52138_new_n5509_));
INVX1 INVX1_1032 ( .A(u2_remHi_286_), .Y(u2__abc_52138_new_n5513_));
INVX1 INVX1_1033 ( .A(u2_o_286_), .Y(u2__abc_52138_new_n5515_));
INVX1 INVX1_1034 ( .A(u2_remHi_287_), .Y(u2__abc_52138_new_n5518_));
INVX1 INVX1_1035 ( .A(u2_o_287_), .Y(u2__abc_52138_new_n5520_));
INVX1 INVX1_1036 ( .A(u2_remHi_292_), .Y(u2__abc_52138_new_n5525_));
INVX1 INVX1_1037 ( .A(u2_o_292_), .Y(u2__abc_52138_new_n5527_));
INVX1 INVX1_1038 ( .A(u2_remHi_293_), .Y(u2__abc_52138_new_n5530_));
INVX1 INVX1_1039 ( .A(u2_o_293_), .Y(u2__abc_52138_new_n5532_));
INVX1 INVX1_104 ( .A(sqrto_178_), .Y(_abc_65734_new_n1136_));
INVX1 INVX1_1040 ( .A(u2_remHi_291_), .Y(u2__abc_52138_new_n5537_));
INVX1 INVX1_1041 ( .A(u2_o_291_), .Y(u2__abc_52138_new_n5539_));
INVX1 INVX1_1042 ( .A(u2__abc_52138_new_n5546_), .Y(u2__abc_52138_new_n5547_));
INVX1 INVX1_1043 ( .A(u2_remHi_280_), .Y(u2__abc_52138_new_n5548_));
INVX1 INVX1_1044 ( .A(u2_o_280_), .Y(u2__abc_52138_new_n5550_));
INVX1 INVX1_1045 ( .A(u2_remHi_281_), .Y(u2__abc_52138_new_n5553_));
INVX1 INVX1_1046 ( .A(u2_o_281_), .Y(u2__abc_52138_new_n5555_));
INVX1 INVX1_1047 ( .A(u2_remHi_278_), .Y(u2__abc_52138_new_n5559_));
INVX1 INVX1_1048 ( .A(u2_o_278_), .Y(u2__abc_52138_new_n5561_));
INVX1 INVX1_1049 ( .A(u2_remHi_279_), .Y(u2__abc_52138_new_n5564_));
INVX1 INVX1_105 ( .A(sqrto_179_), .Y(_abc_65734_new_n1139_));
INVX1 INVX1_1050 ( .A(u2_o_279_), .Y(u2__abc_52138_new_n5566_));
INVX1 INVX1_1051 ( .A(u2_remHi_284_), .Y(u2__abc_52138_new_n5571_));
INVX1 INVX1_1052 ( .A(u2_o_284_), .Y(u2__abc_52138_new_n5573_));
INVX1 INVX1_1053 ( .A(u2_remHi_285_), .Y(u2__abc_52138_new_n5576_));
INVX1 INVX1_1054 ( .A(u2_o_285_), .Y(u2__abc_52138_new_n5578_));
INVX1 INVX1_1055 ( .A(u2_remHi_282_), .Y(u2__abc_52138_new_n5582_));
INVX1 INVX1_1056 ( .A(u2_o_282_), .Y(u2__abc_52138_new_n5584_));
INVX1 INVX1_1057 ( .A(u2_remHi_283_), .Y(u2__abc_52138_new_n5587_));
INVX1 INVX1_1058 ( .A(u2_o_283_), .Y(u2__abc_52138_new_n5589_));
INVX1 INVX1_1059 ( .A(u2_remHi_272_), .Y(u2__abc_52138_new_n5595_));
INVX1 INVX1_106 ( .A(sqrto_180_), .Y(_abc_65734_new_n1142_));
INVX1 INVX1_1060 ( .A(u2_o_272_), .Y(u2__abc_52138_new_n5597_));
INVX1 INVX1_1061 ( .A(u2_remHi_273_), .Y(u2__abc_52138_new_n5600_));
INVX1 INVX1_1062 ( .A(u2_o_273_), .Y(u2__abc_52138_new_n5602_));
INVX1 INVX1_1063 ( .A(u2_remHi_270_), .Y(u2__abc_52138_new_n5606_));
INVX1 INVX1_1064 ( .A(u2_o_270_), .Y(u2__abc_52138_new_n5608_));
INVX1 INVX1_1065 ( .A(u2_remHi_271_), .Y(u2__abc_52138_new_n5611_));
INVX1 INVX1_1066 ( .A(u2_o_271_), .Y(u2__abc_52138_new_n5613_));
INVX1 INVX1_1067 ( .A(u2_remHi_276_), .Y(u2__abc_52138_new_n5618_));
INVX1 INVX1_1068 ( .A(u2_o_276_), .Y(u2__abc_52138_new_n5620_));
INVX1 INVX1_1069 ( .A(u2_remHi_277_), .Y(u2__abc_52138_new_n5623_));
INVX1 INVX1_107 ( .A(sqrto_181_), .Y(_abc_65734_new_n1145_));
INVX1 INVX1_1070 ( .A(u2_o_277_), .Y(u2__abc_52138_new_n5625_));
INVX1 INVX1_1071 ( .A(u2_remHi_275_), .Y(u2__abc_52138_new_n5630_));
INVX1 INVX1_1072 ( .A(u2_o_275_), .Y(u2__abc_52138_new_n5632_));
INVX1 INVX1_1073 ( .A(u2__abc_52138_new_n5638_), .Y(u2__abc_52138_new_n5639_));
INVX1 INVX1_1074 ( .A(u2_o_268_), .Y(u2__abc_52138_new_n5640_));
INVX1 INVX1_1075 ( .A(u2_remHi_268_), .Y(u2__abc_52138_new_n5642_));
INVX1 INVX1_1076 ( .A(u2_o_269_), .Y(u2__abc_52138_new_n5645_));
INVX1 INVX1_1077 ( .A(u2_remHi_269_), .Y(u2__abc_52138_new_n5647_));
INVX1 INVX1_1078 ( .A(u2_remHi_266_), .Y(u2__abc_52138_new_n5651_));
INVX1 INVX1_1079 ( .A(u2_o_266_), .Y(u2__abc_52138_new_n5653_));
INVX1 INVX1_108 ( .A(sqrto_182_), .Y(_abc_65734_new_n1148_));
INVX1 INVX1_1080 ( .A(u2_remHi_267_), .Y(u2__abc_52138_new_n5656_));
INVX1 INVX1_1081 ( .A(u2_o_267_), .Y(u2__abc_52138_new_n5658_));
INVX1 INVX1_1082 ( .A(u2_remHi_264_), .Y(u2__abc_52138_new_n5663_));
INVX1 INVX1_1083 ( .A(u2_o_264_), .Y(u2__abc_52138_new_n5665_));
INVX1 INVX1_1084 ( .A(u2_remHi_265_), .Y(u2__abc_52138_new_n5668_));
INVX1 INVX1_1085 ( .A(u2_o_265_), .Y(u2__abc_52138_new_n5670_));
INVX1 INVX1_1086 ( .A(u2_o_262_), .Y(u2__abc_52138_new_n5674_));
INVX1 INVX1_1087 ( .A(u2_remHi_262_), .Y(u2__abc_52138_new_n5676_));
INVX1 INVX1_1088 ( .A(u2_o_263_), .Y(u2__abc_52138_new_n5679_));
INVX1 INVX1_1089 ( .A(u2_remHi_263_), .Y(u2__abc_52138_new_n5681_));
INVX1 INVX1_109 ( .A(sqrto_183_), .Y(_abc_65734_new_n1151_));
INVX1 INVX1_1090 ( .A(u2_o_254_), .Y(u2__abc_52138_new_n5687_));
INVX1 INVX1_1091 ( .A(u2_remHi_255_), .Y(u2__abc_52138_new_n5688_));
INVX1 INVX1_1092 ( .A(u2_remHi_254_), .Y(u2__abc_52138_new_n5691_));
INVX1 INVX1_1093 ( .A(u2_o_255_), .Y(u2__abc_52138_new_n5692_));
INVX1 INVX1_1094 ( .A(u2__abc_52138_new_n5695_), .Y(u2__abc_52138_new_n5696_));
INVX1 INVX1_1095 ( .A(u2_remHi_256_), .Y(u2__abc_52138_new_n5697_));
INVX1 INVX1_1096 ( .A(u2_o_256_), .Y(u2__abc_52138_new_n5699_));
INVX1 INVX1_1097 ( .A(u2_remHi_257_), .Y(u2__abc_52138_new_n5702_));
INVX1 INVX1_1098 ( .A(u2_o_257_), .Y(u2__abc_52138_new_n5704_));
INVX1 INVX1_1099 ( .A(u2_remHi_260_), .Y(u2__abc_52138_new_n5709_));
INVX1 INVX1_11 ( .A(sqrto_85_), .Y(_abc_65734_new_n857_));
INVX1 INVX1_110 ( .A(sqrto_184_), .Y(_abc_65734_new_n1154_));
INVX1 INVX1_1100 ( .A(u2_o_260_), .Y(u2__abc_52138_new_n5711_));
INVX1 INVX1_1101 ( .A(u2_remHi_261_), .Y(u2__abc_52138_new_n5714_));
INVX1 INVX1_1102 ( .A(u2_o_261_), .Y(u2__abc_52138_new_n5716_));
INVX1 INVX1_1103 ( .A(u2_remHi_258_), .Y(u2__abc_52138_new_n5720_));
INVX1 INVX1_1104 ( .A(u2_o_258_), .Y(u2__abc_52138_new_n5722_));
INVX1 INVX1_1105 ( .A(u2_remHi_259_), .Y(u2__abc_52138_new_n5725_));
INVX1 INVX1_1106 ( .A(u2_o_259_), .Y(u2__abc_52138_new_n5727_));
INVX1 INVX1_1107 ( .A(u2__abc_52138_new_n5703_), .Y(u2__abc_52138_new_n5738_));
INVX1 INVX1_1108 ( .A(u2__abc_52138_new_n5726_), .Y(u2__abc_52138_new_n5741_));
INVX1 INVX1_1109 ( .A(u2__abc_52138_new_n5612_), .Y(u2__abc_52138_new_n5756_));
INVX1 INVX1_111 ( .A(sqrto_185_), .Y(_abc_65734_new_n1157_));
INVX1 INVX1_1110 ( .A(u2_o_274_), .Y(u2__abc_52138_new_n5761_));
INVX1 INVX1_1111 ( .A(u2__abc_52138_new_n5565_), .Y(u2__abc_52138_new_n5768_));
INVX1 INVX1_1112 ( .A(u2__abc_52138_new_n5554_), .Y(u2__abc_52138_new_n5770_));
INVX1 INVX1_1113 ( .A(u2__abc_52138_new_n5581_), .Y(u2__abc_52138_new_n5774_));
INVX1 INVX1_1114 ( .A(u2__abc_52138_new_n5577_), .Y(u2__abc_52138_new_n5777_));
INVX1 INVX1_1115 ( .A(u2__abc_52138_new_n5508_), .Y(u2__abc_52138_new_n5782_));
INVX1 INVX1_1116 ( .A(u2__abc_52138_new_n5519_), .Y(u2__abc_52138_new_n5784_));
INVX1 INVX1_1117 ( .A(u2_o_290_), .Y(u2__abc_52138_new_n5787_));
INVX1 INVX1_1118 ( .A(u2__abc_52138_new_n5540_), .Y(u2__abc_52138_new_n5788_));
INVX1 INVX1_1119 ( .A(u2__abc_52138_new_n5472_), .Y(u2__abc_52138_new_n5797_));
INVX1 INVX1_112 ( .A(sqrto_186_), .Y(_abc_65734_new_n1160_));
INVX1 INVX1_1120 ( .A(u2__abc_52138_new_n5488_), .Y(u2__abc_52138_new_n5801_));
INVX1 INVX1_1121 ( .A(u2__abc_52138_new_n5393_), .Y(u2__abc_52138_new_n5808_));
INVX1 INVX1_1122 ( .A(u2__abc_52138_new_n5376_), .Y(u2__abc_52138_new_n5810_));
INVX1 INVX1_1123 ( .A(u2_o_310_), .Y(u2__abc_52138_new_n5811_));
INVX1 INVX1_1124 ( .A(u2__abc_52138_new_n5383_), .Y(u2__abc_52138_new_n5812_));
INVX1 INVX1_1125 ( .A(u2_remHi_314_), .Y(u2__abc_52138_new_n5818_));
INVX1 INVX1_1126 ( .A(u2__abc_52138_new_n5402_), .Y(u2__abc_52138_new_n5820_));
INVX1 INVX1_1127 ( .A(u2__abc_52138_new_n5424_), .Y(u2__abc_52138_new_n5825_));
INVX1 INVX1_1128 ( .A(u2__abc_52138_new_n5358_), .Y(u2__abc_52138_new_n5838_));
INVX1 INVX1_1129 ( .A(u2__abc_52138_new_n5331_), .Y(u2__abc_52138_new_n5843_));
INVX1 INVX1_113 ( .A(sqrto_187_), .Y(_abc_65734_new_n1163_));
INVX1 INVX1_1130 ( .A(u2_o_322_), .Y(u2__abc_52138_new_n5844_));
INVX1 INVX1_1131 ( .A(u2__abc_52138_new_n5291_), .Y(u2__abc_52138_new_n5850_));
INVX1 INVX1_1132 ( .A(u2__abc_52138_new_n5307_), .Y(u2__abc_52138_new_n5854_));
INVX1 INVX1_1133 ( .A(u2__abc_52138_new_n5191_), .Y(u2__abc_52138_new_n5862_));
INVX1 INVX1_1134 ( .A(u2__abc_52138_new_n5224_), .Y(u2__abc_52138_new_n5865_));
INVX1 INVX1_1135 ( .A(u2__abc_52138_new_n5213_), .Y(u2__abc_52138_new_n5868_));
INVX1 INVX1_1136 ( .A(u2__abc_52138_new_n5235_), .Y(u2__abc_52138_new_n5872_));
INVX1 INVX1_1137 ( .A(u2_remHi_334_), .Y(u2__abc_52138_new_n5874_));
INVX1 INVX1_1138 ( .A(u2__abc_52138_new_n5257_), .Y(u2__abc_52138_new_n5878_));
INVX1 INVX1_1139 ( .A(u2__abc_52138_new_n5269_), .Y(u2__abc_52138_new_n5880_));
INVX1 INVX1_114 ( .A(\a[112] ), .Y(_abc_65734_new_n1168_));
INVX1 INVX1_1140 ( .A(u2_remHi_369_), .Y(u2__abc_52138_new_n5886_));
INVX1 INVX1_1141 ( .A(u2_o_366_), .Y(u2__abc_52138_new_n5890_));
INVX1 INVX1_1142 ( .A(u2__abc_52138_new_n5073_), .Y(u2__abc_52138_new_n5894_));
INVX1 INVX1_1143 ( .A(u2__abc_52138_new_n5075_), .Y(u2__abc_52138_new_n5895_));
INVX1 INVX1_1144 ( .A(u2__abc_52138_new_n5132_), .Y(u2__abc_52138_new_n5902_));
INVX1 INVX1_1145 ( .A(u2__abc_52138_new_n5110_), .Y(u2__abc_52138_new_n5903_));
INVX1 INVX1_1146 ( .A(u2__abc_52138_new_n5124_), .Y(u2__abc_52138_new_n5909_));
INVX1 INVX1_1147 ( .A(u2__abc_52138_new_n5127_), .Y(u2__abc_52138_new_n5910_));
INVX1 INVX1_1148 ( .A(u2_o_362_), .Y(u2__abc_52138_new_n5911_));
INVX1 INVX1_1149 ( .A(u2__abc_52138_new_n5129_), .Y(u2__abc_52138_new_n5912_));
INVX1 INVX1_115 ( .A(\a[0] ), .Y(_abc_65734_new_n1169_));
INVX1 INVX1_1150 ( .A(u2__abc_52138_new_n5120_), .Y(u2__abc_52138_new_n5915_));
INVX1 INVX1_1151 ( .A(u2__abc_52138_new_n5140_), .Y(u2__abc_52138_new_n5918_));
INVX1 INVX1_1152 ( .A(u2__abc_52138_new_n5151_), .Y(u2__abc_52138_new_n5920_));
INVX1 INVX1_1153 ( .A(u2_o_378_), .Y(u2__abc_52138_new_n5933_));
INVX1 INVX1_1154 ( .A(u2__abc_52138_new_n5014_), .Y(u2__abc_52138_new_n5934_));
INVX1 INVX1_1155 ( .A(u2_remHi_444_), .Y(u2__abc_52138_new_n5944_));
INVX1 INVX1_1156 ( .A(u2_o_444_), .Y(u2__abc_52138_new_n5946_));
INVX1 INVX1_1157 ( .A(u2_o_445_), .Y(u2__abc_52138_new_n5949_));
INVX1 INVX1_1158 ( .A(u2_remHi_445_), .Y(u2__abc_52138_new_n5951_));
INVX1 INVX1_1159 ( .A(u2_o_443_), .Y(u2__abc_52138_new_n5955_));
INVX1 INVX1_116 ( .A(\a[2] ), .Y(_abc_65734_new_n1173_));
INVX1 INVX1_1160 ( .A(u2_remHi_443_), .Y(u2__abc_52138_new_n5957_));
INVX1 INVX1_1161 ( .A(u2_remHi_442_), .Y(u2__abc_52138_new_n5960_));
INVX1 INVX1_1162 ( .A(u2_o_442_), .Y(u2__abc_52138_new_n5962_));
INVX1 INVX1_1163 ( .A(u2_remHi_438_), .Y(u2__abc_52138_new_n5967_));
INVX1 INVX1_1164 ( .A(u2_o_438_), .Y(u2__abc_52138_new_n5969_));
INVX1 INVX1_1165 ( .A(u2_remHi_440_), .Y(u2__abc_52138_new_n5974_));
INVX1 INVX1_1166 ( .A(u2_o_440_), .Y(u2__abc_52138_new_n5976_));
INVX1 INVX1_1167 ( .A(u2_o_441_), .Y(u2__abc_52138_new_n5979_));
INVX1 INVX1_1168 ( .A(u2_remHi_441_), .Y(u2__abc_52138_new_n5981_));
INVX1 INVX1_1169 ( .A(u2_remHi_436_), .Y(u2__abc_52138_new_n5987_));
INVX1 INVX1_117 ( .A(\a[4] ), .Y(_abc_65734_new_n1178_));
INVX1 INVX1_1170 ( .A(u2_o_436_), .Y(u2__abc_52138_new_n5989_));
INVX1 INVX1_1171 ( .A(u2_remHi_437_), .Y(u2__abc_52138_new_n5992_));
INVX1 INVX1_1172 ( .A(u2_o_437_), .Y(u2__abc_52138_new_n5994_));
INVX1 INVX1_1173 ( .A(u2_o_435_), .Y(u2__abc_52138_new_n5998_));
INVX1 INVX1_1174 ( .A(u2_remHi_435_), .Y(u2__abc_52138_new_n6000_));
INVX1 INVX1_1175 ( .A(u2_remHi_434_), .Y(u2__abc_52138_new_n6003_));
INVX1 INVX1_1176 ( .A(u2_o_434_), .Y(u2__abc_52138_new_n6005_));
INVX1 INVX1_1177 ( .A(u2_remHi_430_), .Y(u2__abc_52138_new_n6010_));
INVX1 INVX1_1178 ( .A(u2_o_430_), .Y(u2__abc_52138_new_n6012_));
INVX1 INVX1_1179 ( .A(u2_o_431_), .Y(u2__abc_52138_new_n6015_));
INVX1 INVX1_118 ( .A(\a[6] ), .Y(_abc_65734_new_n1183_));
INVX1 INVX1_1180 ( .A(u2_remHi_431_), .Y(u2__abc_52138_new_n6017_));
INVX1 INVX1_1181 ( .A(u2_remHi_432_), .Y(u2__abc_52138_new_n6021_));
INVX1 INVX1_1182 ( .A(u2_o_432_), .Y(u2__abc_52138_new_n6023_));
INVX1 INVX1_1183 ( .A(u2_o_433_), .Y(u2__abc_52138_new_n6026_));
INVX1 INVX1_1184 ( .A(u2_remHi_433_), .Y(u2__abc_52138_new_n6028_));
INVX1 INVX1_1185 ( .A(u2__abc_52138_new_n6034_), .Y(u2__abc_52138_new_n6035_));
INVX1 INVX1_1186 ( .A(u2_o_424_), .Y(u2__abc_52138_new_n6036_));
INVX1 INVX1_1187 ( .A(u2_remHi_424_), .Y(u2__abc_52138_new_n6038_));
INVX1 INVX1_1188 ( .A(u2_remHi_425_), .Y(u2__abc_52138_new_n6041_));
INVX1 INVX1_1189 ( .A(u2_o_425_), .Y(u2__abc_52138_new_n6043_));
INVX1 INVX1_119 ( .A(\a[8] ), .Y(_abc_65734_new_n1188_));
INVX1 INVX1_1190 ( .A(u2_remHi_422_), .Y(u2__abc_52138_new_n6047_));
INVX1 INVX1_1191 ( .A(u2_o_422_), .Y(u2__abc_52138_new_n6049_));
INVX1 INVX1_1192 ( .A(u2_o_423_), .Y(u2__abc_52138_new_n6052_));
INVX1 INVX1_1193 ( .A(u2_remHi_423_), .Y(u2__abc_52138_new_n6054_));
INVX1 INVX1_1194 ( .A(u2_o_428_), .Y(u2__abc_52138_new_n6058_));
INVX1 INVX1_1195 ( .A(u2_remHi_428_), .Y(u2__abc_52138_new_n6060_));
INVX1 INVX1_1196 ( .A(u2_o_429_), .Y(u2__abc_52138_new_n6063_));
INVX1 INVX1_1197 ( .A(u2_remHi_429_), .Y(u2__abc_52138_new_n6065_));
INVX1 INVX1_1198 ( .A(u2__abc_52138_new_n6068_), .Y(u2__abc_52138_new_n6069_));
INVX1 INVX1_1199 ( .A(u2_o_427_), .Y(u2__abc_52138_new_n6070_));
INVX1 INVX1_12 ( .A(sqrto_86_), .Y(_abc_65734_new_n860_));
INVX1 INVX1_120 ( .A(\a[10] ), .Y(_abc_65734_new_n1193_));
INVX1 INVX1_1200 ( .A(u2_remHi_427_), .Y(u2__abc_52138_new_n6072_));
INVX1 INVX1_1201 ( .A(u2_remHi_426_), .Y(u2__abc_52138_new_n6075_));
INVX1 INVX1_1202 ( .A(u2_o_426_), .Y(u2__abc_52138_new_n6077_));
INVX1 INVX1_1203 ( .A(u2__abc_52138_new_n6081_), .Y(u2__abc_52138_new_n6082_));
INVX1 INVX1_1204 ( .A(u2_o_420_), .Y(u2__abc_52138_new_n6084_));
INVX1 INVX1_1205 ( .A(u2_remHi_420_), .Y(u2__abc_52138_new_n6086_));
INVX1 INVX1_1206 ( .A(u2_o_421_), .Y(u2__abc_52138_new_n6089_));
INVX1 INVX1_1207 ( .A(u2_remHi_421_), .Y(u2__abc_52138_new_n6091_));
INVX1 INVX1_1208 ( .A(u2__abc_52138_new_n6094_), .Y(u2__abc_52138_new_n6095_));
INVX1 INVX1_1209 ( .A(u2_o_419_), .Y(u2__abc_52138_new_n6096_));
INVX1 INVX1_121 ( .A(\a[12] ), .Y(_abc_65734_new_n1198_));
INVX1 INVX1_1210 ( .A(u2_remHi_419_), .Y(u2__abc_52138_new_n6098_));
INVX1 INVX1_1211 ( .A(u2_remHi_418_), .Y(u2__abc_52138_new_n6101_));
INVX1 INVX1_1212 ( .A(u2_o_418_), .Y(u2__abc_52138_new_n6103_));
INVX1 INVX1_1213 ( .A(u2_o_416_), .Y(u2__abc_52138_new_n6108_));
INVX1 INVX1_1214 ( .A(u2_remHi_416_), .Y(u2__abc_52138_new_n6110_));
INVX1 INVX1_1215 ( .A(u2_remHi_417_), .Y(u2__abc_52138_new_n6113_));
INVX1 INVX1_1216 ( .A(u2_o_417_), .Y(u2__abc_52138_new_n6115_));
INVX1 INVX1_1217 ( .A(u2__abc_52138_new_n6118_), .Y(u2__abc_52138_new_n6119_));
INVX1 INVX1_1218 ( .A(u2_o_415_), .Y(u2__abc_52138_new_n6120_));
INVX1 INVX1_1219 ( .A(u2_remHi_415_), .Y(u2__abc_52138_new_n6122_));
INVX1 INVX1_122 ( .A(\a[14] ), .Y(_abc_65734_new_n1203_));
INVX1 INVX1_1220 ( .A(u2_remHi_414_), .Y(u2__abc_52138_new_n6125_));
INVX1 INVX1_1221 ( .A(u2_o_414_), .Y(u2__abc_52138_new_n6127_));
INVX1 INVX1_1222 ( .A(u2__abc_52138_new_n6132_), .Y(u2__abc_52138_new_n6133_));
INVX1 INVX1_1223 ( .A(u2_remHi_388_), .Y(u2__abc_52138_new_n6136_));
INVX1 INVX1_1224 ( .A(u2_o_388_), .Y(u2__abc_52138_new_n6138_));
INVX1 INVX1_1225 ( .A(u2_remHi_389_), .Y(u2__abc_52138_new_n6141_));
INVX1 INVX1_1226 ( .A(u2_o_389_), .Y(u2__abc_52138_new_n6143_));
INVX1 INVX1_1227 ( .A(u2_o_387_), .Y(u2__abc_52138_new_n6147_));
INVX1 INVX1_1228 ( .A(u2_remHi_387_), .Y(u2__abc_52138_new_n6149_));
INVX1 INVX1_1229 ( .A(u2_remHi_386_), .Y(u2__abc_52138_new_n6152_));
INVX1 INVX1_123 ( .A(\a[16] ), .Y(_abc_65734_new_n1208_));
INVX1 INVX1_1230 ( .A(u2_o_386_), .Y(u2__abc_52138_new_n6154_));
INVX1 INVX1_1231 ( .A(u2__abc_52138_new_n6158_), .Y(u2__abc_52138_new_n6159_));
INVX1 INVX1_1232 ( .A(u2_remHi_384_), .Y(u2__abc_52138_new_n6160_));
INVX1 INVX1_1233 ( .A(u2_o_384_), .Y(u2__abc_52138_new_n6162_));
INVX1 INVX1_1234 ( .A(u2_o_385_), .Y(u2__abc_52138_new_n6165_));
INVX1 INVX1_1235 ( .A(u2_remHi_385_), .Y(u2__abc_52138_new_n6167_));
INVX1 INVX1_1236 ( .A(u2_o_383_), .Y(u2__abc_52138_new_n6171_));
INVX1 INVX1_1237 ( .A(u2_remHi_383_), .Y(u2__abc_52138_new_n6173_));
INVX1 INVX1_1238 ( .A(u2_remHi_382_), .Y(u2__abc_52138_new_n6176_));
INVX1 INVX1_1239 ( .A(u2_o_382_), .Y(u2__abc_52138_new_n6178_));
INVX1 INVX1_124 ( .A(\a[18] ), .Y(_abc_65734_new_n1213_));
INVX1 INVX1_1240 ( .A(u2__abc_52138_new_n6182_), .Y(u2__abc_52138_new_n6183_));
INVX1 INVX1_1241 ( .A(u2_remHi_408_), .Y(u2__abc_52138_new_n6185_));
INVX1 INVX1_1242 ( .A(u2_o_408_), .Y(u2__abc_52138_new_n6187_));
INVX1 INVX1_1243 ( .A(u2_o_409_), .Y(u2__abc_52138_new_n6190_));
INVX1 INVX1_1244 ( .A(u2_remHi_409_), .Y(u2__abc_52138_new_n6192_));
INVX1 INVX1_1245 ( .A(u2_o_407_), .Y(u2__abc_52138_new_n6196_));
INVX1 INVX1_1246 ( .A(u2_remHi_407_), .Y(u2__abc_52138_new_n6198_));
INVX1 INVX1_1247 ( .A(u2_remHi_406_), .Y(u2__abc_52138_new_n6201_));
INVX1 INVX1_1248 ( .A(u2_o_406_), .Y(u2__abc_52138_new_n6203_));
INVX1 INVX1_1249 ( .A(u2_remHi_412_), .Y(u2__abc_52138_new_n6208_));
INVX1 INVX1_125 ( .A(\a[20] ), .Y(_abc_65734_new_n1218_));
INVX1 INVX1_1250 ( .A(u2_o_412_), .Y(u2__abc_52138_new_n6210_));
INVX1 INVX1_1251 ( .A(u2_remHi_413_), .Y(u2__abc_52138_new_n6213_));
INVX1 INVX1_1252 ( .A(u2_o_413_), .Y(u2__abc_52138_new_n6215_));
INVX1 INVX1_1253 ( .A(u2_o_411_), .Y(u2__abc_52138_new_n6219_));
INVX1 INVX1_1254 ( .A(u2_remHi_411_), .Y(u2__abc_52138_new_n6221_));
INVX1 INVX1_1255 ( .A(u2_remHi_410_), .Y(u2__abc_52138_new_n6224_));
INVX1 INVX1_1256 ( .A(u2_o_410_), .Y(u2__abc_52138_new_n6226_));
INVX1 INVX1_1257 ( .A(u2_remHi_398_), .Y(u2__abc_52138_new_n6232_));
INVX1 INVX1_1258 ( .A(u2_o_398_), .Y(u2__abc_52138_new_n6234_));
INVX1 INVX1_1259 ( .A(u2_o_399_), .Y(u2__abc_52138_new_n6237_));
INVX1 INVX1_126 ( .A(\a[22] ), .Y(_abc_65734_new_n1223_));
INVX1 INVX1_1260 ( .A(u2_remHi_399_), .Y(u2__abc_52138_new_n6239_));
INVX1 INVX1_1261 ( .A(u2_remHi_400_), .Y(u2__abc_52138_new_n6243_));
INVX1 INVX1_1262 ( .A(u2_o_400_), .Y(u2__abc_52138_new_n6245_));
INVX1 INVX1_1263 ( .A(u2_o_401_), .Y(u2__abc_52138_new_n6248_));
INVX1 INVX1_1264 ( .A(u2_remHi_401_), .Y(u2__abc_52138_new_n6250_));
INVX1 INVX1_1265 ( .A(u2_remHi_404_), .Y(u2__abc_52138_new_n6255_));
INVX1 INVX1_1266 ( .A(u2_o_404_), .Y(u2__abc_52138_new_n6257_));
INVX1 INVX1_1267 ( .A(u2_remHi_405_), .Y(u2__abc_52138_new_n6260_));
INVX1 INVX1_1268 ( .A(u2_o_405_), .Y(u2__abc_52138_new_n6262_));
INVX1 INVX1_1269 ( .A(u2_o_403_), .Y(u2__abc_52138_new_n6266_));
INVX1 INVX1_127 ( .A(\a[24] ), .Y(_abc_65734_new_n1228_));
INVX1 INVX1_1270 ( .A(u2_remHi_403_), .Y(u2__abc_52138_new_n6268_));
INVX1 INVX1_1271 ( .A(u2_remHi_402_), .Y(u2__abc_52138_new_n6271_));
INVX1 INVX1_1272 ( .A(u2_o_402_), .Y(u2__abc_52138_new_n6273_));
INVX1 INVX1_1273 ( .A(u2_remHi_392_), .Y(u2__abc_52138_new_n6280_));
INVX1 INVX1_1274 ( .A(u2_o_392_), .Y(u2__abc_52138_new_n6282_));
INVX1 INVX1_1275 ( .A(u2_o_393_), .Y(u2__abc_52138_new_n6285_));
INVX1 INVX1_1276 ( .A(u2__abc_52138_new_n6286_), .Y(u2__abc_52138_new_n6287_));
INVX1 INVX1_1277 ( .A(u2__abc_52138_new_n6289_), .Y(u2__abc_52138_new_n6290_));
INVX1 INVX1_1278 ( .A(u2_remHi_390_), .Y(u2__abc_52138_new_n6292_));
INVX1 INVX1_1279 ( .A(u2__abc_52138_new_n6294_), .Y(u2__abc_52138_new_n6295_));
INVX1 INVX1_128 ( .A(\a[26] ), .Y(_abc_65734_new_n1233_));
INVX1 INVX1_1280 ( .A(u2_remHi_391_), .Y(u2__abc_52138_new_n6297_));
INVX1 INVX1_1281 ( .A(u2__abc_52138_new_n6298_), .Y(u2__abc_52138_new_n6299_));
INVX1 INVX1_1282 ( .A(u2_remHi_396_), .Y(u2__abc_52138_new_n6304_));
INVX1 INVX1_1283 ( .A(u2_o_396_), .Y(u2__abc_52138_new_n6306_));
INVX1 INVX1_1284 ( .A(u2_remHi_397_), .Y(u2__abc_52138_new_n6309_));
INVX1 INVX1_1285 ( .A(u2_o_397_), .Y(u2__abc_52138_new_n6311_));
INVX1 INVX1_1286 ( .A(u2_o_395_), .Y(u2__abc_52138_new_n6315_));
INVX1 INVX1_1287 ( .A(u2_remHi_395_), .Y(u2__abc_52138_new_n6317_));
INVX1 INVX1_1288 ( .A(u2_remHi_394_), .Y(u2__abc_52138_new_n6320_));
INVX1 INVX1_1289 ( .A(u2__abc_52138_new_n6321_), .Y(u2__abc_52138_new_n6322_));
INVX1 INVX1_129 ( .A(\a[28] ), .Y(_abc_65734_new_n1238_));
INVX1 INVX1_1290 ( .A(u2__abc_52138_new_n6327_), .Y(u2__abc_52138_new_n6328_));
INVX1 INVX1_1291 ( .A(u2__abc_52138_new_n6329_), .Y(u2__abc_52138_new_n6330_));
INVX1 INVX1_1292 ( .A(u2__abc_52138_new_n6135_), .Y(u2__abc_52138_new_n6333_));
INVX1 INVX1_1293 ( .A(u2__abc_52138_new_n6174_), .Y(u2__abc_52138_new_n6334_));
INVX1 INVX1_1294 ( .A(u2__abc_52138_new_n6168_), .Y(u2__abc_52138_new_n6336_));
INVX1 INVX1_1295 ( .A(u2__abc_52138_new_n6150_), .Y(u2__abc_52138_new_n6339_));
INVX1 INVX1_1296 ( .A(u2__abc_52138_new_n6314_), .Y(u2__abc_52138_new_n6345_));
INVX1 INVX1_1297 ( .A(u2__abc_52138_new_n6316_), .Y(u2__abc_52138_new_n6346_));
INVX1 INVX1_1298 ( .A(u2__abc_52138_new_n6300_), .Y(u2__abc_52138_new_n6350_));
INVX1 INVX1_1299 ( .A(u2_remHi_393_), .Y(u2__abc_52138_new_n6352_));
INVX1 INVX1_13 ( .A(sqrto_87_), .Y(_abc_65734_new_n863_));
INVX1 INVX1_130 ( .A(\a[30] ), .Y(_abc_65734_new_n1243_));
INVX1 INVX1_1300 ( .A(u2__abc_52138_new_n6199_), .Y(u2__abc_52138_new_n6358_));
INVX1 INVX1_1301 ( .A(u2__abc_52138_new_n6193_), .Y(u2__abc_52138_new_n6360_));
INVX1 INVX1_1302 ( .A(u2__abc_52138_new_n6218_), .Y(u2__abc_52138_new_n6364_));
INVX1 INVX1_1303 ( .A(u2__abc_52138_new_n6220_), .Y(u2__abc_52138_new_n6365_));
INVX1 INVX1_1304 ( .A(u2__abc_52138_new_n6227_), .Y(u2__abc_52138_new_n6366_));
INVX1 INVX1_1305 ( .A(u2__abc_52138_new_n6214_), .Y(u2__abc_52138_new_n6368_));
INVX1 INVX1_1306 ( .A(u2__abc_52138_new_n6369_), .Y(u2__abc_52138_new_n6370_));
INVX1 INVX1_1307 ( .A(u2__abc_52138_new_n6240_), .Y(u2__abc_52138_new_n6373_));
INVX1 INVX1_1308 ( .A(u2__abc_52138_new_n6251_), .Y(u2__abc_52138_new_n6375_));
INVX1 INVX1_1309 ( .A(u2__abc_52138_new_n6269_), .Y(u2__abc_52138_new_n6378_));
INVX1 INVX1_131 ( .A(\a[32] ), .Y(_abc_65734_new_n1248_));
INVX1 INVX1_1310 ( .A(u2__abc_52138_new_n6261_), .Y(u2__abc_52138_new_n6380_));
INVX1 INVX1_1311 ( .A(u2__abc_52138_new_n6107_), .Y(u2__abc_52138_new_n6387_));
INVX1 INVX1_1312 ( .A(u2__abc_52138_new_n6121_), .Y(u2__abc_52138_new_n6388_));
INVX1 INVX1_1313 ( .A(u2__abc_52138_new_n6128_), .Y(u2__abc_52138_new_n6389_));
INVX1 INVX1_1314 ( .A(u2__abc_52138_new_n6097_), .Y(u2__abc_52138_new_n6393_));
INVX1 INVX1_1315 ( .A(u2__abc_52138_new_n6104_), .Y(u2__abc_52138_new_n6394_));
INVX1 INVX1_1316 ( .A(u2__abc_52138_new_n6046_), .Y(u2__abc_52138_new_n6400_));
INVX1 INVX1_1317 ( .A(u2__abc_52138_new_n6055_), .Y(u2__abc_52138_new_n6401_));
INVX1 INVX1_1318 ( .A(u2__abc_52138_new_n6071_), .Y(u2__abc_52138_new_n6406_));
INVX1 INVX1_1319 ( .A(u2__abc_52138_new_n6078_), .Y(u2__abc_52138_new_n6407_));
INVX1 INVX1_132 ( .A(\a[34] ), .Y(_abc_65734_new_n1253_));
INVX1 INVX1_1320 ( .A(u2__abc_52138_new_n5984_), .Y(u2__abc_52138_new_n6413_));
INVX1 INVX1_1321 ( .A(u2_o_439_), .Y(u2__abc_52138_new_n6414_));
INVX1 INVX1_1322 ( .A(u2_remHi_439_), .Y(u2__abc_52138_new_n6415_));
INVX1 INVX1_1323 ( .A(u2__abc_52138_new_n5952_), .Y(u2__abc_52138_new_n6424_));
INVX1 INVX1_1324 ( .A(u2__abc_52138_new_n6018_), .Y(u2__abc_52138_new_n6427_));
INVX1 INVX1_1325 ( .A(u2__abc_52138_new_n6001_), .Y(u2__abc_52138_new_n6431_));
INVX1 INVX1_1326 ( .A(u2__abc_52138_new_n5993_), .Y(u2__abc_52138_new_n6433_));
INVX1 INVX1_1327 ( .A(u2_o_449_), .Y(u2__abc_52138_new_n6446_));
INVX1 INVX1_1328 ( .A(u2_remHi_449_), .Y(u2__abc_52138_new_n6447_));
INVX1 INVX1_1329 ( .A(sqrto_4_), .Y(u2__abc_52138_new_n6458_));
INVX1 INVX1_133 ( .A(\a[36] ), .Y(_abc_65734_new_n1258_));
INVX1 INVX1_1330 ( .A(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n6499_));
INVX1 INVX1_1331 ( .A(u2_remHi_0_), .Y(u2__abc_52138_new_n6502_));
INVX1 INVX1_1332 ( .A(u2_state_2_), .Y(u2__abc_52138_new_n6503_));
INVX1 INVX1_1333 ( .A(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n6505_));
INVX1 INVX1_1334 ( .A(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6510_));
INVX1 INVX1_1335 ( .A(u2_remHi_1_), .Y(u2__abc_52138_new_n6515_));
INVX1 INVX1_1336 ( .A(u2__abc_52138_new_n6450_), .Y(u2__abc_52138_new_n6538_));
INVX1 INVX1_1337 ( .A(u2__abc_52138_new_n6540_), .Y(u2__abc_52138_new_n6541_));
INVX1 INVX1_1338 ( .A(u2__abc_52138_new_n6542_), .Y(u2__abc_52138_new_n6550_));
INVX1 INVX1_1339 ( .A(u2__abc_52138_new_n6459_), .Y(u2__abc_52138_new_n6578_));
INVX1 INVX1_134 ( .A(\a[38] ), .Y(_abc_65734_new_n1263_));
INVX1 INVX1_1340 ( .A(u2__abc_52138_new_n3057_), .Y(u2__abc_52138_new_n6579_));
INVX1 INVX1_1341 ( .A(u2_remHi_8_), .Y(u2__abc_52138_new_n6586_));
INVX1 INVX1_1342 ( .A(u2__abc_52138_new_n3041_), .Y(u2__abc_52138_new_n6600_));
INVX1 INVX1_1343 ( .A(u2__abc_52138_new_n3046_), .Y(u2__abc_52138_new_n6601_));
INVX1 INVX1_1344 ( .A(u2__abc_52138_new_n6603_), .Y(u2__abc_52138_new_n6604_));
INVX1 INVX1_1345 ( .A(u2__abc_52138_new_n6606_), .Y(u2__abc_52138_new_n6607_));
INVX1 INVX1_1346 ( .A(u2__abc_52138_new_n6628_), .Y(u2__abc_52138_new_n6643_));
INVX1 INVX1_1347 ( .A(sqrto_12_), .Y(u2__abc_52138_new_n6654_));
INVX1 INVX1_1348 ( .A(u2__abc_52138_new_n3171_), .Y(u2__abc_52138_new_n6664_));
INVX1 INVX1_1349 ( .A(u2__abc_52138_new_n6673_), .Y(u2__abc_52138_new_n6674_));
INVX1 INVX1_135 ( .A(\a[40] ), .Y(_abc_65734_new_n1268_));
INVX1 INVX1_1350 ( .A(u2__abc_52138_new_n3160_), .Y(u2__abc_52138_new_n6691_));
INVX1 INVX1_1351 ( .A(u2__abc_52138_new_n3176_), .Y(u2__abc_52138_new_n6692_));
INVX1 INVX1_1352 ( .A(u2_remHi_19_), .Y(u2__abc_52138_new_n6706_));
INVX1 INVX1_1353 ( .A(u2__abc_52138_new_n3165_), .Y(u2__abc_52138_new_n6713_));
INVX1 INVX1_1354 ( .A(sqrto_20_), .Y(u2__abc_52138_new_n6733_));
INVX1 INVX1_1355 ( .A(u2__abc_52138_new_n6734_), .Y(u2__abc_52138_new_n6760_));
INVX1 INVX1_1356 ( .A(u2__abc_52138_new_n3132_), .Y(u2__abc_52138_new_n6765_));
INVX1 INVX1_1357 ( .A(u2__abc_52138_new_n6801_), .Y(u2__abc_52138_new_n6802_));
INVX1 INVX1_1358 ( .A(u2__abc_52138_new_n6803_), .Y(u2__abc_52138_new_n6804_));
INVX1 INVX1_1359 ( .A(u2__abc_52138_new_n6805_), .Y(u2__abc_52138_new_n6806_));
INVX1 INVX1_136 ( .A(\a[42] ), .Y(_abc_65734_new_n1273_));
INVX1 INVX1_1360 ( .A(u2__abc_52138_new_n6808_), .Y(u2__abc_52138_new_n6809_));
INVX1 INVX1_1361 ( .A(u2_remHi_32_), .Y(u2__abc_52138_new_n6848_));
INVX1 INVX1_1362 ( .A(u2__abc_52138_new_n6844_), .Y(u2__abc_52138_new_n6853_));
INVX1 INVX1_1363 ( .A(u2__abc_52138_new_n6854_), .Y(u2__abc_52138_new_n6862_));
INVX1 INVX1_1364 ( .A(u2__abc_52138_new_n6887_), .Y(u2__abc_52138_new_n6888_));
INVX1 INVX1_1365 ( .A(u2__abc_52138_new_n3402_), .Y(u2__abc_52138_new_n6904_));
INVX1 INVX1_1366 ( .A(u2__abc_52138_new_n3350_), .Y(u2__abc_52138_new_n6923_));
INVX1 INVX1_1367 ( .A(u2__abc_52138_new_n6931_), .Y(u2__abc_52138_new_n6932_));
INVX1 INVX1_1368 ( .A(u2__abc_52138_new_n3352_), .Y(u2__abc_52138_new_n6947_));
INVX1 INVX1_1369 ( .A(u2__abc_52138_new_n3347_), .Y(u2__abc_52138_new_n6966_));
INVX1 INVX1_137 ( .A(\a[44] ), .Y(_abc_65734_new_n1278_));
INVX1 INVX1_1370 ( .A(u2__abc_52138_new_n3372_), .Y(u2__abc_52138_new_n6988_));
INVX1 INVX1_1371 ( .A(u2__abc_52138_new_n3359_), .Y(u2__abc_52138_new_n6998_));
INVX1 INVX1_1372 ( .A(u2__abc_52138_new_n7012_), .Y(u2__abc_52138_new_n7014_));
INVX1 INVX1_1373 ( .A(u2__abc_52138_new_n3301_), .Y(u2__abc_52138_new_n7030_));
INVX1 INVX1_1374 ( .A(u2__abc_52138_new_n7053_), .Y(u2__abc_52138_new_n7054_));
INVX1 INVX1_1375 ( .A(u2__abc_52138_new_n3325_), .Y(u2__abc_52138_new_n7073_));
INVX1 INVX1_1376 ( .A(u2__abc_52138_new_n7074_), .Y(u2__abc_52138_new_n7075_));
INVX1 INVX1_1377 ( .A(u2__abc_52138_new_n7055_), .Y(u2__abc_52138_new_n7094_));
INVX1 INVX1_1378 ( .A(u2__abc_52138_new_n7110_), .Y(u2__abc_52138_new_n7117_));
INVX1 INVX1_1379 ( .A(u2__abc_52138_new_n3283_), .Y(u2__abc_52138_new_n7135_));
INVX1 INVX1_138 ( .A(\a[46] ), .Y(_abc_65734_new_n1283_));
INVX1 INVX1_1380 ( .A(u2__abc_52138_new_n7140_), .Y(u2__abc_52138_new_n7141_));
INVX1 INVX1_1381 ( .A(u2__abc_52138_new_n7185_), .Y(u2__abc_52138_new_n7186_));
INVX1 INVX1_1382 ( .A(u2__abc_52138_new_n3849_), .Y(u2__abc_52138_new_n7212_));
INVX1 INVX1_1383 ( .A(u2__abc_52138_new_n7203_), .Y(u2__abc_52138_new_n7223_));
INVX1 INVX1_1384 ( .A(u2__abc_52138_new_n3844_), .Y(u2__abc_52138_new_n7224_));
INVX1 INVX1_1385 ( .A(sqrto_68_), .Y(u2__abc_52138_new_n7264_));
INVX1 INVX1_1386 ( .A(u2__abc_52138_new_n7268_), .Y(u2__abc_52138_new_n7269_));
INVX1 INVX1_1387 ( .A(u2__abc_52138_new_n7270_), .Y(u2__abc_52138_new_n7271_));
INVX1 INVX1_1388 ( .A(u2__abc_52138_new_n7289_), .Y(u2__abc_52138_new_n7311_));
INVX1 INVX1_1389 ( .A(u2__abc_52138_new_n7315_), .Y(u2__abc_52138_new_n7316_));
INVX1 INVX1_139 ( .A(\a[48] ), .Y(_abc_65734_new_n1288_));
INVX1 INVX1_1390 ( .A(u2__abc_52138_new_n7325_), .Y(u2__abc_52138_new_n7326_));
INVX1 INVX1_1391 ( .A(u2__abc_52138_new_n3822_), .Y(u2__abc_52138_new_n7357_));
INVX1 INVX1_1392 ( .A(u2__abc_52138_new_n3747_), .Y(u2__abc_52138_new_n7371_));
INVX1 INVX1_1393 ( .A(u2__abc_52138_new_n7380_), .Y(u2__abc_52138_new_n7381_));
INVX1 INVX1_1394 ( .A(u2__abc_52138_new_n3781_), .Y(u2__abc_52138_new_n7399_));
INVX1 INVX1_1395 ( .A(u2__abc_52138_new_n7407_), .Y(u2__abc_52138_new_n7408_));
INVX1 INVX1_1396 ( .A(u2__abc_52138_new_n7452_), .Y(u2__abc_52138_new_n7453_));
INVX1 INVX1_1397 ( .A(u2__abc_52138_new_n7463_), .Y(u2__abc_52138_new_n7464_));
INVX1 INVX1_1398 ( .A(u2__abc_52138_new_n3717_), .Y(u2__abc_52138_new_n7472_));
INVX1 INVX1_1399 ( .A(u2__abc_52138_new_n7474_), .Y(u2__abc_52138_new_n7475_));
INVX1 INVX1_14 ( .A(sqrto_88_), .Y(_abc_65734_new_n866_));
INVX1 INVX1_140 ( .A(\a[50] ), .Y(_abc_65734_new_n1293_));
INVX1 INVX1_1400 ( .A(u2__abc_52138_new_n7494_), .Y(u2__abc_52138_new_n7495_));
INVX1 INVX1_1401 ( .A(u2__abc_52138_new_n3692_), .Y(u2__abc_52138_new_n7522_));
INVX1 INVX1_1402 ( .A(u2__abc_52138_new_n3662_), .Y(u2__abc_52138_new_n7543_));
INVX1 INVX1_1403 ( .A(u2__abc_52138_new_n3685_), .Y(u2__abc_52138_new_n7579_));
INVX1 INVX1_1404 ( .A(u2__abc_52138_new_n7581_), .Y(u2__abc_52138_new_n7582_));
INVX1 INVX1_1405 ( .A(u2__abc_52138_new_n7583_), .Y(u2__abc_52138_new_n7584_));
INVX1 INVX1_1406 ( .A(u2__abc_52138_new_n7587_), .Y(u2__abc_52138_new_n7588_));
INVX1 INVX1_1407 ( .A(u2__abc_52138_new_n3674_), .Y(u2__abc_52138_new_n7616_));
INVX1 INVX1_1408 ( .A(u2__abc_52138_new_n7629_), .Y(u2__abc_52138_new_n7630_));
INVX1 INVX1_1409 ( .A(u2__abc_52138_new_n7632_), .Y(u2__abc_52138_new_n7633_));
INVX1 INVX1_141 ( .A(\a[52] ), .Y(_abc_65734_new_n1298_));
INVX1 INVX1_1410 ( .A(u2__abc_52138_new_n3627_), .Y(u2__abc_52138_new_n7703_));
INVX1 INVX1_1411 ( .A(u2__abc_52138_new_n7695_), .Y(u2__abc_52138_new_n7705_));
INVX1 INVX1_1412 ( .A(u2__abc_52138_new_n7721_), .Y(u2__abc_52138_new_n7729_));
INVX1 INVX1_1413 ( .A(u2__abc_52138_new_n7738_), .Y(u2__abc_52138_new_n7757_));
INVX1 INVX1_1414 ( .A(u2__abc_52138_new_n3587_), .Y(u2__abc_52138_new_n7771_));
INVX1 INVX1_1415 ( .A(rst), .Y(u2__abc_52138_new_n7779_));
INVX1 INVX1_1416 ( .A(u2__abc_52138_new_n3514_), .Y(u2__abc_52138_new_n7819_));
INVX1 INVX1_1417 ( .A(u2__abc_52138_new_n3520_), .Y(u2__abc_52138_new_n7828_));
INVX1 INVX1_1418 ( .A(u2__abc_52138_new_n7829_), .Y(u2__abc_52138_new_n7830_));
INVX1 INVX1_1419 ( .A(u2__abc_52138_new_n7852_), .Y(u2__abc_52138_new_n7853_));
INVX1 INVX1_142 ( .A(\a[54] ), .Y(_abc_65734_new_n1303_));
INVX1 INVX1_1420 ( .A(u2__abc_52138_new_n3528_), .Y(u2__abc_52138_new_n7890_));
INVX1 INVX1_1421 ( .A(u2_remHi_128_), .Y(u2__abc_52138_new_n7905_));
INVX1 INVX1_1422 ( .A(u2__abc_52138_new_n7918_), .Y(u2__abc_52138_new_n7919_));
INVX1 INVX1_1423 ( .A(u2__abc_52138_new_n7944_), .Y(u2__abc_52138_new_n7945_));
INVX1 INVX1_1424 ( .A(u2__abc_52138_new_n4681_), .Y(u2__abc_52138_new_n7981_));
INVX1 INVX1_1425 ( .A(u2__abc_52138_new_n4734_), .Y(u2__abc_52138_new_n7984_));
INVX1 INVX1_1426 ( .A(u2__abc_52138_new_n7989_), .Y(u2__abc_52138_new_n7990_));
INVX1 INVX1_1427 ( .A(u2__abc_52138_new_n4683_), .Y(u2__abc_52138_new_n8007_));
INVX1 INVX1_1428 ( .A(u2__abc_52138_new_n4678_), .Y(u2__abc_52138_new_n8030_));
INVX1 INVX1_1429 ( .A(u2__abc_52138_new_n7987_), .Y(u2__abc_52138_new_n8072_));
INVX1 INVX1_143 ( .A(\a[56] ), .Y(_abc_65734_new_n1308_));
INVX1 INVX1_1430 ( .A(u2__abc_52138_new_n8082_), .Y(u2__abc_52138_new_n8083_));
INVX1 INVX1_1431 ( .A(u2__abc_52138_new_n4634_), .Y(u2__abc_52138_new_n8132_));
INVX1 INVX1_1432 ( .A(u2__abc_52138_new_n4593_), .Y(u2__abc_52138_new_n8162_));
INVX1 INVX1_1433 ( .A(u2__abc_52138_new_n8172_), .Y(u2__abc_52138_new_n8189_));
INVX1 INVX1_1434 ( .A(u2__abc_52138_new_n8211_), .Y(u2__abc_52138_new_n8212_));
INVX1 INVX1_1435 ( .A(u2__abc_52138_new_n4610_), .Y(u2__abc_52138_new_n8229_));
INVX1 INVX1_1436 ( .A(u2_remHi_159_), .Y(u2__abc_52138_new_n8243_));
INVX1 INVX1_1437 ( .A(u2__abc_52138_new_n8256_), .Y(u2__abc_52138_new_n8257_));
INVX1 INVX1_1438 ( .A(u2__abc_52138_new_n8258_), .Y(u2__abc_52138_new_n8259_));
INVX1 INVX1_1439 ( .A(u2__abc_52138_new_n8303_), .Y(u2__abc_52138_new_n8304_));
INVX1 INVX1_144 ( .A(\a[58] ), .Y(_abc_65734_new_n1313_));
INVX1 INVX1_1440 ( .A(u2__abc_52138_new_n4563_), .Y(u2__abc_52138_new_n8312_));
INVX1 INVX1_1441 ( .A(u2__abc_52138_new_n8321_), .Y(u2__abc_52138_new_n8322_));
INVX1 INVX1_1442 ( .A(u2__abc_52138_new_n4549_), .Y(u2__abc_52138_new_n8331_));
INVX1 INVX1_1443 ( .A(u2__abc_52138_new_n8342_), .Y(u2__abc_52138_new_n8343_));
INVX1 INVX1_1444 ( .A(u2__abc_52138_new_n8344_), .Y(u2__abc_52138_new_n8345_));
INVX1 INVX1_1445 ( .A(u2__abc_52138_new_n8346_), .Y(u2__abc_52138_new_n8347_));
INVX1 INVX1_1446 ( .A(u2__abc_52138_new_n4513_), .Y(u2__abc_52138_new_n8363_));
INVX1 INVX1_1447 ( .A(u2__abc_52138_new_n8384_), .Y(u2__abc_52138_new_n8385_));
INVX1 INVX1_1448 ( .A(u2__abc_52138_new_n4511_), .Y(u2__abc_52138_new_n8418_));
INVX1 INVX1_1449 ( .A(u2__abc_52138_new_n4488_), .Y(u2__abc_52138_new_n8422_));
INVX1 INVX1_145 ( .A(\a[60] ), .Y(_abc_65734_new_n1318_));
INVX1 INVX1_1450 ( .A(u2__abc_52138_new_n4479_), .Y(u2__abc_52138_new_n8424_));
INVX1 INVX1_1451 ( .A(u2__abc_52138_new_n4484_), .Y(u2__abc_52138_new_n8425_));
INVX1 INVX1_1452 ( .A(u2__abc_52138_new_n4456_), .Y(u2__abc_52138_new_n8448_));
INVX1 INVX1_1453 ( .A(u2__abc_52138_new_n4472_), .Y(u2__abc_52138_new_n8450_));
INVX1 INVX1_1454 ( .A(u2__abc_52138_new_n8451_), .Y(u2__abc_52138_new_n8452_));
INVX1 INVX1_1455 ( .A(u2__abc_52138_new_n8473_), .Y(u2__abc_52138_new_n8474_));
INVX1 INVX1_1456 ( .A(u2__abc_52138_new_n8475_), .Y(u2__abc_52138_new_n8476_));
INVX1 INVX1_1457 ( .A(u2__abc_52138_new_n8515_), .Y(u2__abc_52138_new_n8523_));
INVX1 INVX1_1458 ( .A(u2__abc_52138_new_n8532_), .Y(u2__abc_52138_new_n8533_));
INVX1 INVX1_1459 ( .A(u2__abc_52138_new_n8535_), .Y(u2__abc_52138_new_n8543_));
INVX1 INVX1_146 ( .A(\a[62] ), .Y(_abc_65734_new_n1323_));
INVX1 INVX1_1460 ( .A(u2__abc_52138_new_n8554_), .Y(u2__abc_52138_new_n8555_));
INVX1 INVX1_1461 ( .A(u2__abc_52138_new_n8573_), .Y(u2__abc_52138_new_n8594_));
INVX1 INVX1_1462 ( .A(u2__abc_52138_new_n4406_), .Y(u2__abc_52138_new_n8596_));
INVX1 INVX1_1463 ( .A(u2__abc_52138_new_n8603_), .Y(u2__abc_52138_new_n8604_));
INVX1 INVX1_1464 ( .A(u2__abc_52138_new_n8605_), .Y(u2__abc_52138_new_n8606_));
INVX1 INVX1_1465 ( .A(u2__abc_52138_new_n8623_), .Y(u2__abc_52138_new_n8624_));
INVX1 INVX1_1466 ( .A(u2__abc_52138_new_n4346_), .Y(u2__abc_52138_new_n8654_));
INVX1 INVX1_1467 ( .A(u2__abc_52138_new_n4309_), .Y(u2__abc_52138_new_n8685_));
INVX1 INVX1_1468 ( .A(u2__abc_52138_new_n8692_), .Y(u2__abc_52138_new_n8709_));
INVX1 INVX1_1469 ( .A(u2__abc_52138_new_n8731_), .Y(u2__abc_52138_new_n8732_));
INVX1 INVX1_147 ( .A(\a[64] ), .Y(_abc_65734_new_n1328_));
INVX1 INVX1_1470 ( .A(u2__abc_52138_new_n4324_), .Y(u2__abc_52138_new_n8749_));
INVX1 INVX1_1471 ( .A(u2__abc_52138_new_n4256_), .Y(u2__abc_52138_new_n8767_));
INVX1 INVX1_1472 ( .A(u2__abc_52138_new_n8785_), .Y(u2__abc_52138_new_n8793_));
INVX1 INVX1_1473 ( .A(u2__abc_52138_new_n4281_), .Y(u2__abc_52138_new_n8852_));
INVX1 INVX1_1474 ( .A(u2__abc_52138_new_n8858_), .Y(u2__abc_52138_new_n8866_));
INVX1 INVX1_1475 ( .A(u2__abc_52138_new_n8875_), .Y(u2__abc_52138_new_n8876_));
INVX1 INVX1_1476 ( .A(u2__abc_52138_new_n8877_), .Y(u2__abc_52138_new_n8885_));
INVX1 INVX1_1477 ( .A(u2__abc_52138_new_n4237_), .Y(u2__abc_52138_new_n8894_));
INVX1 INVX1_1478 ( .A(u2__abc_52138_new_n8898_), .Y(u2__abc_52138_new_n8899_));
INVX1 INVX1_1479 ( .A(u2__abc_52138_new_n4218_), .Y(u2__abc_52138_new_n8926_));
INVX1 INVX1_148 ( .A(\a[66] ), .Y(_abc_65734_new_n1333_));
INVX1 INVX1_1480 ( .A(u2__abc_52138_new_n4166_), .Y(u2__abc_52138_new_n8935_));
INVX1 INVX1_1481 ( .A(u2__abc_52138_new_n8944_), .Y(u2__abc_52138_new_n8945_));
INVX1 INVX1_1482 ( .A(u2__abc_52138_new_n8946_), .Y(u2__abc_52138_new_n8947_));
INVX1 INVX1_1483 ( .A(u2__abc_52138_new_n8983_), .Y(u2__abc_52138_new_n8984_));
INVX1 INVX1_1484 ( .A(u2__abc_52138_new_n4183_), .Y(u2__abc_52138_new_n9001_));
INVX1 INVX1_1485 ( .A(u2__abc_52138_new_n4170_), .Y(u2__abc_52138_new_n9020_));
INVX1 INVX1_1486 ( .A(u2__abc_52138_new_n9101_), .Y(u2__abc_52138_new_n9102_));
INVX1 INVX1_1487 ( .A(u2__abc_52138_new_n9107_), .Y(u2__abc_52138_new_n9115_));
INVX1 INVX1_1488 ( .A(u2__abc_52138_new_n9124_), .Y(u2__abc_52138_new_n9125_));
INVX1 INVX1_1489 ( .A(u2__abc_52138_new_n9126_), .Y(u2__abc_52138_new_n9134_));
INVX1 INVX1_149 ( .A(\a[68] ), .Y(_abc_65734_new_n1338_));
INVX1 INVX1_1490 ( .A(u2__abc_52138_new_n4094_), .Y(u2__abc_52138_new_n9143_));
INVX1 INVX1_1491 ( .A(u2__abc_52138_new_n9145_), .Y(u2__abc_52138_new_n9146_));
INVX1 INVX1_1492 ( .A(u2__abc_52138_new_n4078_), .Y(u2__abc_52138_new_n9163_));
INVX1 INVX1_1493 ( .A(u2__abc_52138_new_n4075_), .Y(u2__abc_52138_new_n9173_));
INVX1 INVX1_1494 ( .A(u2__abc_52138_new_n4086_), .Y(u2__abc_52138_new_n9182_));
INVX1 INVX1_1495 ( .A(u2__abc_52138_new_n4018_), .Y(u2__abc_52138_new_n9205_));
INVX1 INVX1_1496 ( .A(u2__abc_52138_new_n9206_), .Y(u2__abc_52138_new_n9207_));
INVX1 INVX1_1497 ( .A(u2__abc_52138_new_n4046_), .Y(u2__abc_52138_new_n9226_));
INVX1 INVX1_1498 ( .A(u2__abc_52138_new_n9230_), .Y(u2__abc_52138_new_n9231_));
INVX1 INVX1_1499 ( .A(u2__abc_52138_new_n9265_), .Y(u2__abc_52138_new_n9287_));
INVX1 INVX1_15 ( .A(sqrto_89_), .Y(_abc_65734_new_n869_));
INVX1 INVX1_150 ( .A(\a[70] ), .Y(_abc_65734_new_n1343_));
INVX1 INVX1_1500 ( .A(u2__abc_52138_new_n9278_), .Y(u2__abc_52138_new_n9288_));
INVX1 INVX1_1501 ( .A(u2__abc_52138_new_n5698_), .Y(u2__abc_52138_new_n9306_));
INVX1 INVX1_1502 ( .A(u2__abc_52138_new_n9298_), .Y(u2__abc_52138_new_n9307_));
INVX1 INVX1_1503 ( .A(u2__abc_52138_new_n5708_), .Y(u2__abc_52138_new_n9316_));
INVX1 INVX1_1504 ( .A(u2__abc_52138_new_n9317_), .Y(u2__abc_52138_new_n9318_));
INVX1 INVX1_1505 ( .A(u2__abc_52138_new_n9319_), .Y(u2__abc_52138_new_n9320_));
INVX1 INVX1_1506 ( .A(u2__abc_52138_new_n9322_), .Y(u2__abc_52138_new_n9323_));
INVX1 INVX1_1507 ( .A(u2__abc_52138_new_n5728_), .Y(u2__abc_52138_new_n9340_));
INVX1 INVX1_1508 ( .A(u2__abc_52138_new_n9341_), .Y(u2__abc_52138_new_n9342_));
INVX1 INVX1_1509 ( .A(u2__abc_52138_new_n9351_), .Y(u2__abc_52138_new_n9352_));
INVX1 INVX1_151 ( .A(\a[72] ), .Y(_abc_65734_new_n1348_));
INVX1 INVX1_1510 ( .A(u2__abc_52138_new_n5677_), .Y(u2__abc_52138_new_n9372_));
INVX1 INVX1_1511 ( .A(u2__abc_52138_new_n9364_), .Y(u2__abc_52138_new_n9373_));
INVX1 INVX1_1512 ( .A(u2__abc_52138_new_n5652_), .Y(u2__abc_52138_new_n9418_));
INVX1 INVX1_1513 ( .A(u2__abc_52138_new_n5659_), .Y(u2__abc_52138_new_n9420_));
INVX1 INVX1_1514 ( .A(u2__abc_52138_new_n9421_), .Y(u2__abc_52138_new_n9422_));
INVX1 INVX1_1515 ( .A(u2__abc_52138_new_n5643_), .Y(u2__abc_52138_new_n9430_));
INVX1 INVX1_1516 ( .A(u2__abc_52138_new_n9446_), .Y(u2__abc_52138_new_n9447_));
INVX1 INVX1_1517 ( .A(u2__abc_52138_new_n9448_), .Y(u2__abc_52138_new_n9449_));
INVX1 INVX1_1518 ( .A(u2__abc_52138_new_n9466_), .Y(u2__abc_52138_new_n9467_));
INVX1 INVX1_1519 ( .A(u2_remHi_274_), .Y(u2__abc_52138_new_n9471_));
INVX1 INVX1_152 ( .A(\a[74] ), .Y(_abc_65734_new_n1353_));
INVX1 INVX1_1520 ( .A(u2__abc_52138_new_n5596_), .Y(u2__abc_52138_new_n9476_));
INVX1 INVX1_1521 ( .A(u2__abc_52138_new_n5617_), .Y(u2__abc_52138_new_n9485_));
INVX1 INVX1_1522 ( .A(u2__abc_52138_new_n9488_), .Y(u2__abc_52138_new_n9489_));
INVX1 INVX1_1523 ( .A(u2__abc_52138_new_n9491_), .Y(u2__abc_52138_new_n9492_));
INVX1 INVX1_1524 ( .A(u2__abc_52138_new_n5631_), .Y(u2__abc_52138_new_n9508_));
INVX1 INVX1_1525 ( .A(u2__abc_52138_new_n9510_), .Y(u2__abc_52138_new_n9511_));
INVX1 INVX1_1526 ( .A(u2__abc_52138_new_n5619_), .Y(u2__abc_52138_new_n9519_));
INVX1 INVX1_1527 ( .A(u2__abc_52138_new_n9533_), .Y(u2__abc_52138_new_n9534_));
INVX1 INVX1_1528 ( .A(u2__abc_52138_new_n9551_), .Y(u2__abc_52138_new_n9552_));
INVX1 INVX1_1529 ( .A(u2__abc_52138_new_n5549_), .Y(u2__abc_52138_new_n9560_));
INVX1 INVX1_153 ( .A(\a[76] ), .Y(_abc_65734_new_n1358_));
INVX1 INVX1_1530 ( .A(u2__abc_52138_new_n9570_), .Y(u2__abc_52138_new_n9571_));
INVX1 INVX1_1531 ( .A(u2__abc_52138_new_n9573_), .Y(u2__abc_52138_new_n9574_));
INVX1 INVX1_1532 ( .A(u2__abc_52138_new_n9575_), .Y(u2__abc_52138_new_n9576_));
INVX1 INVX1_1533 ( .A(u2__abc_52138_new_n5583_), .Y(u2__abc_52138_new_n9584_));
INVX1 INVX1_1534 ( .A(u2__abc_52138_new_n5590_), .Y(u2__abc_52138_new_n9594_));
INVX1 INVX1_1535 ( .A(u2__abc_52138_new_n9595_), .Y(u2__abc_52138_new_n9596_));
INVX1 INVX1_1536 ( .A(u2__abc_52138_new_n9621_), .Y(u2__abc_52138_new_n9622_));
INVX1 INVX1_1537 ( .A(u2__abc_52138_new_n9623_), .Y(u2__abc_52138_new_n9624_));
INVX1 INVX1_1538 ( .A(u2__abc_52138_new_n9641_), .Y(u2__abc_52138_new_n9642_));
INVX1 INVX1_1539 ( .A(u2_remHi_290_), .Y(u2__abc_52138_new_n9646_));
INVX1 INVX1_154 ( .A(\a[78] ), .Y(_abc_65734_new_n1363_));
INVX1 INVX1_1540 ( .A(u2__abc_52138_new_n5503_), .Y(u2__abc_52138_new_n9651_));
INVX1 INVX1_1541 ( .A(u2__abc_52138_new_n9662_), .Y(u2__abc_52138_new_n9663_));
INVX1 INVX1_1542 ( .A(u2__abc_52138_new_n9664_), .Y(u2__abc_52138_new_n9665_));
INVX1 INVX1_1543 ( .A(u2__abc_52138_new_n9667_), .Y(u2__abc_52138_new_n9668_));
INVX1 INVX1_1544 ( .A(u2__abc_52138_new_n5538_), .Y(u2__abc_52138_new_n9684_));
INVX1 INVX1_1545 ( .A(u2__abc_52138_new_n9686_), .Y(u2__abc_52138_new_n9687_));
INVX1 INVX1_1546 ( .A(u2__abc_52138_new_n5526_), .Y(u2__abc_52138_new_n9695_));
INVX1 INVX1_1547 ( .A(u2__abc_52138_new_n5458_), .Y(u2__abc_52138_new_n9716_));
INVX1 INVX1_1548 ( .A(u2__abc_52138_new_n9708_), .Y(u2__abc_52138_new_n9717_));
INVX1 INVX1_1549 ( .A(u2__abc_52138_new_n9747_), .Y(u2__abc_52138_new_n9748_));
INVX1 INVX1_155 ( .A(\a[80] ), .Y(_abc_65734_new_n1368_));
INVX1 INVX1_1550 ( .A(u2__abc_52138_new_n9749_), .Y(u2__abc_52138_new_n9750_));
INVX1 INVX1_1551 ( .A(u2__abc_52138_new_n5495_), .Y(u2__abc_52138_new_n9766_));
INVX1 INVX1_1552 ( .A(u2__abc_52138_new_n5497_), .Y(u2__abc_52138_new_n9768_));
INVX1 INVX1_1553 ( .A(u2__abc_52138_new_n9769_), .Y(u2__abc_52138_new_n9770_));
INVX1 INVX1_1554 ( .A(u2__abc_52138_new_n5410_), .Y(u2__abc_52138_new_n9802_));
INVX1 INVX1_1555 ( .A(u2__abc_52138_new_n9794_), .Y(u2__abc_52138_new_n9803_));
INVX1 INVX1_1556 ( .A(u2__abc_52138_new_n5429_), .Y(u2__abc_52138_new_n9830_));
INVX1 INVX1_1557 ( .A(u2__abc_52138_new_n9832_), .Y(u2__abc_52138_new_n9833_));
INVX1 INVX1_1558 ( .A(u2__abc_52138_new_n9835_), .Y(u2__abc_52138_new_n9836_));
INVX1 INVX1_1559 ( .A(u2__abc_52138_new_n9844_), .Y(u2__abc_52138_new_n9845_));
INVX1 INVX1_156 ( .A(\a[82] ), .Y(_abc_65734_new_n1373_));
INVX1 INVX1_1560 ( .A(u2_remHi_310_), .Y(u2__abc_52138_new_n9858_));
INVX1 INVX1_1561 ( .A(u2__abc_52138_new_n9877_), .Y(u2__abc_52138_new_n9878_));
INVX1 INVX1_1562 ( .A(u2__abc_52138_new_n5381_), .Y(u2__abc_52138_new_n9894_));
INVX1 INVX1_1563 ( .A(u2__abc_52138_new_n9896_), .Y(u2__abc_52138_new_n9897_));
INVX1 INVX1_1564 ( .A(u2__abc_52138_new_n5369_), .Y(u2__abc_52138_new_n9905_));
INVX1 INVX1_1565 ( .A(u2__abc_52138_new_n9916_), .Y(u2__abc_52138_new_n9917_));
INVX1 INVX1_1566 ( .A(u2__abc_52138_new_n9920_), .Y(u2__abc_52138_new_n9921_));
INVX1 INVX1_1567 ( .A(u2__abc_52138_new_n5400_), .Y(u2__abc_52138_new_n9937_));
INVX1 INVX1_1568 ( .A(u2__abc_52138_new_n9939_), .Y(u2__abc_52138_new_n9940_));
INVX1 INVX1_1569 ( .A(u2__abc_52138_new_n5388_), .Y(u2__abc_52138_new_n9948_));
INVX1 INVX1_157 ( .A(\a[84] ), .Y(_abc_65734_new_n1378_));
INVX1 INVX1_1570 ( .A(u2__abc_52138_new_n9792_), .Y(u2__abc_52138_new_n9959_));
INVX1 INVX1_1571 ( .A(u2__abc_52138_new_n9967_), .Y(u2__abc_52138_new_n9968_));
INVX1 INVX1_1572 ( .A(u2__abc_52138_new_n5344_), .Y(u2__abc_52138_new_n9976_));
INVX1 INVX1_1573 ( .A(u2__abc_52138_new_n9986_), .Y(u2__abc_52138_new_n9987_));
INVX1 INVX1_1574 ( .A(u2_remHi_322_), .Y(u2__abc_52138_new_n9992_));
INVX1 INVX1_1575 ( .A(u2__abc_52138_new_n10007_), .Y(u2__abc_52138_new_n10008_));
INVX1 INVX1_1576 ( .A(u2__abc_52138_new_n10010_), .Y(u2__abc_52138_new_n10011_));
INVX1 INVX1_1577 ( .A(u2__abc_52138_new_n10028_), .Y(u2__abc_52138_new_n10029_));
INVX1 INVX1_1578 ( .A(u2__abc_52138_new_n5324_), .Y(u2__abc_52138_new_n10037_));
INVX1 INVX1_1579 ( .A(u2__abc_52138_new_n5277_), .Y(u2__abc_52138_new_n10060_));
INVX1 INVX1_158 ( .A(\a[86] ), .Y(_abc_65734_new_n1383_));
INVX1 INVX1_1580 ( .A(u2__abc_52138_new_n10052_), .Y(u2__abc_52138_new_n10061_));
INVX1 INVX1_1581 ( .A(u2__abc_52138_new_n10091_), .Y(u2__abc_52138_new_n10092_));
INVX1 INVX1_1582 ( .A(u2__abc_52138_new_n10093_), .Y(u2__abc_52138_new_n10094_));
INVX1 INVX1_1583 ( .A(u2__abc_52138_new_n5309_), .Y(u2__abc_52138_new_n10102_));
INVX1 INVX1_1584 ( .A(u2__abc_52138_new_n5316_), .Y(u2__abc_52138_new_n10112_));
INVX1 INVX1_1585 ( .A(u2__abc_52138_new_n10113_), .Y(u2__abc_52138_new_n10114_));
INVX1 INVX1_1586 ( .A(u2__abc_52138_new_n10050_), .Y(u2__abc_52138_new_n10131_));
INVX1 INVX1_1587 ( .A(u2__abc_52138_new_n10138_), .Y(u2__abc_52138_new_n10139_));
INVX1 INVX1_1588 ( .A(u2__abc_52138_new_n10156_), .Y(u2__abc_52138_new_n10157_));
INVX1 INVX1_1589 ( .A(u2__abc_52138_new_n5230_), .Y(u2__abc_52138_new_n10165_));
INVX1 INVX1_159 ( .A(\a[88] ), .Y(_abc_65734_new_n1388_));
INVX1 INVX1_1590 ( .A(u2__abc_52138_new_n10137_), .Y(u2__abc_52138_new_n10174_));
INVX1 INVX1_1591 ( .A(u2__abc_52138_new_n10176_), .Y(u2__abc_52138_new_n10177_));
INVX1 INVX1_1592 ( .A(u2__abc_52138_new_n10178_), .Y(u2__abc_52138_new_n10179_));
INVX1 INVX1_1593 ( .A(u2__abc_52138_new_n10181_), .Y(u2__abc_52138_new_n10182_));
INVX1 INVX1_1594 ( .A(u2__abc_52138_new_n10199_), .Y(u2__abc_52138_new_n10200_));
INVX1 INVX1_1595 ( .A(u2__abc_52138_new_n5255_), .Y(u2__abc_52138_new_n10218_));
INVX1 INVX1_1596 ( .A(u2__abc_52138_new_n10222_), .Y(u2__abc_52138_new_n10223_));
INVX1 INVX1_1597 ( .A(u2__abc_52138_new_n10224_), .Y(u2__abc_52138_new_n10225_));
INVX1 INVX1_1598 ( .A(u2__abc_52138_new_n5196_), .Y(u2__abc_52138_new_n10233_));
INVX1 INVX1_1599 ( .A(u2__abc_52138_new_n5203_), .Y(u2__abc_52138_new_n10243_));
INVX1 INVX1_16 ( .A(sqrto_90_), .Y(_abc_65734_new_n872_));
INVX1 INVX1_160 ( .A(\a[90] ), .Y(_abc_65734_new_n1393_));
INVX1 INVX1_1600 ( .A(u2__abc_52138_new_n10244_), .Y(u2__abc_52138_new_n10245_));
INVX1 INVX1_1601 ( .A(u2__abc_52138_new_n5184_), .Y(u2__abc_52138_new_n10263_));
INVX1 INVX1_1602 ( .A(u2__abc_52138_new_n10265_), .Y(u2__abc_52138_new_n10266_));
INVX1 INVX1_1603 ( .A(u2__abc_52138_new_n10268_), .Y(u2__abc_52138_new_n10269_));
INVX1 INVX1_1604 ( .A(u2__abc_52138_new_n10314_), .Y(u2__abc_52138_new_n10315_));
INVX1 INVX1_1605 ( .A(u2__abc_52138_new_n10332_), .Y(u2__abc_52138_new_n10333_));
INVX1 INVX1_1606 ( .A(u2__abc_52138_new_n5135_), .Y(u2__abc_52138_new_n10341_));
INVX1 INVX1_1607 ( .A(u2__abc_52138_new_n10351_), .Y(u2__abc_52138_new_n10352_));
INVX1 INVX1_1608 ( .A(u2__abc_52138_new_n10354_), .Y(u2__abc_52138_new_n10355_));
INVX1 INVX1_1609 ( .A(u2__abc_52138_new_n10356_), .Y(u2__abc_52138_new_n10357_));
INVX1 INVX1_161 ( .A(\a[92] ), .Y(_abc_65734_new_n1398_));
INVX1 INVX1_1610 ( .A(u2__abc_52138_new_n5169_), .Y(u2__abc_52138_new_n10365_));
INVX1 INVX1_1611 ( .A(u2__abc_52138_new_n5176_), .Y(u2__abc_52138_new_n10375_));
INVX1 INVX1_1612 ( .A(u2__abc_52138_new_n10376_), .Y(u2__abc_52138_new_n10377_));
INVX1 INVX1_1613 ( .A(u2__abc_52138_new_n5158_), .Y(u2__abc_52138_new_n10385_));
INVX1 INVX1_1614 ( .A(u2__abc_52138_new_n10397_), .Y(u2__abc_52138_new_n10398_));
INVX1 INVX1_1615 ( .A(u2__abc_52138_new_n10400_), .Y(u2__abc_52138_new_n10401_));
INVX1 INVX1_1616 ( .A(u2__abc_52138_new_n10419_), .Y(u2__abc_52138_new_n10420_));
INVX1 INVX1_1617 ( .A(u2_remHi_362_), .Y(u2__abc_52138_new_n10425_));
INVX1 INVX1_1618 ( .A(u2__abc_52138_new_n10444_), .Y(u2__abc_52138_new_n10445_));
INVX1 INVX1_1619 ( .A(u2__abc_52138_new_n10462_), .Y(u2__abc_52138_new_n10463_));
INVX1 INVX1_162 ( .A(\a[94] ), .Y(_abc_65734_new_n1403_));
INVX1 INVX1_1620 ( .A(u2__abc_52138_new_n5115_), .Y(u2__abc_52138_new_n10471_));
INVX1 INVX1_1621 ( .A(u2__abc_52138_new_n10486_), .Y(u2__abc_52138_new_n10487_));
INVX1 INVX1_1622 ( .A(u2__abc_52138_new_n10488_), .Y(u2__abc_52138_new_n10489_));
INVX1 INVX1_1623 ( .A(u2__abc_52138_new_n10506_), .Y(u2__abc_52138_new_n10507_));
INVX1 INVX1_1624 ( .A(u2__abc_52138_new_n5046_), .Y(u2__abc_52138_new_n10515_));
INVX1 INVX1_1625 ( .A(u2__abc_52138_new_n10537_), .Y(u2__abc_52138_new_n10545_));
INVX1 INVX1_1626 ( .A(u2__abc_52138_new_n5088_), .Y(u2__abc_52138_new_n10564_));
INVX1 INVX1_1627 ( .A(u2__abc_52138_new_n5029_), .Y(u2__abc_52138_new_n10585_));
INVX1 INVX1_1628 ( .A(u2__abc_52138_new_n5021_), .Y(u2__abc_52138_new_n10586_));
INVX1 INVX1_1629 ( .A(u2_remHi_378_), .Y(u2__abc_52138_new_n10593_));
INVX1 INVX1_163 ( .A(\a[96] ), .Y(_abc_65734_new_n1408_));
INVX1 INVX1_1630 ( .A(u2__abc_52138_new_n5041_), .Y(u2__abc_52138_new_n10598_));
INVX1 INVX1_1631 ( .A(u2__abc_52138_new_n10609_), .Y(u2__abc_52138_new_n10610_));
INVX1 INVX1_1632 ( .A(u2__abc_52138_new_n5012_), .Y(u2__abc_52138_new_n10626_));
INVX1 INVX1_1633 ( .A(u2__abc_52138_new_n10628_), .Y(u2__abc_52138_new_n10629_));
INVX1 INVX1_1634 ( .A(u2__abc_52138_new_n5000_), .Y(u2__abc_52138_new_n10637_));
INVX1 INVX1_1635 ( .A(u2__abc_52138_new_n5736_), .Y(u2__abc_52138_new_n10646_));
INVX1 INVX1_1636 ( .A(u2__abc_52138_new_n5367_), .Y(u2__abc_52138_new_n10648_));
INVX1 INVX1_1637 ( .A(u2__abc_52138_new_n10587_), .Y(u2__abc_52138_new_n10651_));
INVX1 INVX1_1638 ( .A(u2__abc_52138_new_n10660_), .Y(u2__abc_52138_new_n10661_));
INVX1 INVX1_1639 ( .A(u2__abc_52138_new_n10662_), .Y(u2__abc_52138_new_n10663_));
INVX1 INVX1_164 ( .A(\a[98] ), .Y(_abc_65734_new_n1413_));
INVX1 INVX1_1640 ( .A(u2__abc_52138_new_n6172_), .Y(u2__abc_52138_new_n10679_));
INVX1 INVX1_1641 ( .A(u2__abc_52138_new_n10681_), .Y(u2__abc_52138_new_n10682_));
INVX1 INVX1_1642 ( .A(u2__abc_52138_new_n6161_), .Y(u2__abc_52138_new_n10690_));
INVX1 INVX1_1643 ( .A(u2__abc_52138_new_n10700_), .Y(u2__abc_52138_new_n10701_));
INVX1 INVX1_1644 ( .A(u2__abc_52138_new_n10702_), .Y(u2__abc_52138_new_n10703_));
INVX1 INVX1_1645 ( .A(u2__abc_52138_new_n10705_), .Y(u2__abc_52138_new_n10706_));
INVX1 INVX1_1646 ( .A(u2__abc_52138_new_n6140_), .Y(u2__abc_52138_new_n10722_));
INVX1 INVX1_1647 ( .A(u2__abc_52138_new_n6148_), .Y(u2__abc_52138_new_n10723_));
INVX1 INVX1_1648 ( .A(u2__abc_52138_new_n6137_), .Y(u2__abc_52138_new_n10735_));
INVX1 INVX1_1649 ( .A(u2__abc_52138_new_n6142_), .Y(u2__abc_52138_new_n10745_));
INVX1 INVX1_165 ( .A(\a[100] ), .Y(_abc_65734_new_n1418_));
INVX1 INVX1_1650 ( .A(u2__abc_52138_new_n10748_), .Y(u2__abc_52138_new_n10749_));
INVX1 INVX1_1651 ( .A(u2__abc_52138_new_n10760_), .Y(u2__abc_52138_new_n10762_));
INVX1 INVX1_1652 ( .A(u2__abc_52138_new_n6281_), .Y(u2__abc_52138_new_n10788_));
INVX1 INVX1_1653 ( .A(u2__abc_52138_new_n10789_), .Y(u2__abc_52138_new_n10790_));
INVX1 INVX1_1654 ( .A(u2__abc_52138_new_n10792_), .Y(u2__abc_52138_new_n10793_));
INVX1 INVX1_1655 ( .A(u2__abc_52138_new_n10794_), .Y(u2__abc_52138_new_n10795_));
INVX1 INVX1_1656 ( .A(u2__abc_52138_new_n10812_), .Y(u2__abc_52138_new_n10813_));
INVX1 INVX1_1657 ( .A(u2__abc_52138_new_n10835_), .Y(u2__abc_52138_new_n10836_));
INVX1 INVX1_1658 ( .A(u2__abc_52138_new_n6233_), .Y(u2__abc_52138_new_n10844_));
INVX1 INVX1_1659 ( .A(u2__abc_52138_new_n10853_), .Y(u2__abc_52138_new_n10854_));
INVX1 INVX1_166 ( .A(\a[102] ), .Y(_abc_65734_new_n1423_));
INVX1 INVX1_1660 ( .A(u2__abc_52138_new_n6254_), .Y(u2__abc_52138_new_n10872_));
INVX1 INVX1_1661 ( .A(u2__abc_52138_new_n6253_), .Y(u2__abc_52138_new_n10873_));
INVX1 INVX1_1662 ( .A(u2__abc_52138_new_n6244_), .Y(u2__abc_52138_new_n10874_));
INVX1 INVX1_1663 ( .A(u2__abc_52138_new_n10878_), .Y(u2__abc_52138_new_n10879_));
INVX1 INVX1_1664 ( .A(u2__abc_52138_new_n6267_), .Y(u2__abc_52138_new_n10895_));
INVX1 INVX1_1665 ( .A(u2__abc_52138_new_n10897_), .Y(u2__abc_52138_new_n10898_));
INVX1 INVX1_1666 ( .A(u2__abc_52138_new_n6256_), .Y(u2__abc_52138_new_n10906_));
INVX1 INVX1_1667 ( .A(u2__abc_52138_new_n6277_), .Y(u2__abc_52138_new_n10915_));
INVX1 INVX1_1668 ( .A(u2__abc_52138_new_n10922_), .Y(u2__abc_52138_new_n10923_));
INVX1 INVX1_1669 ( .A(u2__abc_52138_new_n6197_), .Y(u2__abc_52138_new_n10939_));
INVX1 INVX1_167 ( .A(\a[104] ), .Y(_abc_65734_new_n1428_));
INVX1 INVX1_1670 ( .A(u2__abc_52138_new_n10941_), .Y(u2__abc_52138_new_n10942_));
INVX1 INVX1_1671 ( .A(u2__abc_52138_new_n6186_), .Y(u2__abc_52138_new_n10950_));
INVX1 INVX1_1672 ( .A(u2__abc_52138_new_n10960_), .Y(u2__abc_52138_new_n10961_));
INVX1 INVX1_1673 ( .A(u2__abc_52138_new_n10963_), .Y(u2__abc_52138_new_n10964_));
INVX1 INVX1_1674 ( .A(u2__abc_52138_new_n10965_), .Y(u2__abc_52138_new_n10966_));
INVX1 INVX1_1675 ( .A(u2__abc_52138_new_n6225_), .Y(u2__abc_52138_new_n10974_));
INVX1 INVX1_1676 ( .A(u2__abc_52138_new_n10984_), .Y(u2__abc_52138_new_n10985_));
INVX1 INVX1_1677 ( .A(u2__abc_52138_new_n6209_), .Y(u2__abc_52138_new_n10993_));
INVX1 INVX1_1678 ( .A(u2__abc_52138_new_n11012_), .Y(u2__abc_52138_new_n11013_));
INVX1 INVX1_1679 ( .A(u2__abc_52138_new_n6123_), .Y(u2__abc_52138_new_n11029_));
INVX1 INVX1_168 ( .A(\a[106] ), .Y(_abc_65734_new_n1433_));
INVX1 INVX1_1680 ( .A(u2__abc_52138_new_n6117_), .Y(u2__abc_52138_new_n11041_));
INVX1 INVX1_1681 ( .A(u2__abc_52138_new_n11051_), .Y(u2__abc_52138_new_n11052_));
INVX1 INVX1_1682 ( .A(u2__abc_52138_new_n11054_), .Y(u2__abc_52138_new_n11055_));
INVX1 INVX1_1683 ( .A(u2__abc_52138_new_n11056_), .Y(u2__abc_52138_new_n11057_));
INVX1 INVX1_1684 ( .A(u2__abc_52138_new_n6102_), .Y(u2__abc_52138_new_n11065_));
INVX1 INVX1_1685 ( .A(u2__abc_52138_new_n6093_), .Y(u2__abc_52138_new_n11085_));
INVX1 INVX1_1686 ( .A(u2__abc_52138_new_n11053_), .Y(u2__abc_52138_new_n11094_));
INVX1 INVX1_1687 ( .A(u2__abc_52138_new_n11099_), .Y(u2__abc_52138_new_n11100_));
INVX1 INVX1_1688 ( .A(u2__abc_52138_new_n6048_), .Y(u2__abc_52138_new_n11108_));
INVX1 INVX1_1689 ( .A(u2__abc_52138_new_n6053_), .Y(u2__abc_52138_new_n11117_));
INVX1 INVX1_169 ( .A(\a[108] ), .Y(_abc_65734_new_n1438_));
INVX1 INVX1_1690 ( .A(u2__abc_52138_new_n6045_), .Y(u2__abc_52138_new_n11128_));
INVX1 INVX1_1691 ( .A(u2__abc_52138_new_n11141_), .Y(u2__abc_52138_new_n11142_));
INVX1 INVX1_1692 ( .A(u2__abc_52138_new_n11158_), .Y(u2__abc_52138_new_n11159_));
INVX1 INVX1_1693 ( .A(u2__abc_52138_new_n6067_), .Y(u2__abc_52138_new_n11170_));
INVX1 INVX1_1694 ( .A(u2__abc_52138_new_n11011_), .Y(u2__abc_52138_new_n11179_));
INVX1 INVX1_1695 ( .A(u2__abc_52138_new_n6011_), .Y(u2__abc_52138_new_n11193_));
INVX1 INVX1_1696 ( .A(u2__abc_52138_new_n11185_), .Y(u2__abc_52138_new_n11194_));
INVX1 INVX1_1697 ( .A(u2__abc_52138_new_n11203_), .Y(u2__abc_52138_new_n11204_));
INVX1 INVX1_1698 ( .A(u2__abc_52138_new_n11206_), .Y(u2__abc_52138_new_n11207_));
INVX1 INVX1_1699 ( .A(u2__abc_52138_new_n6027_), .Y(u2__abc_52138_new_n11223_));
INVX1 INVX1_17 ( .A(sqrto_91_), .Y(_abc_65734_new_n875_));
INVX1 INVX1_170 ( .A(\a[110] ), .Y(_abc_65734_new_n1443_));
INVX1 INVX1_1700 ( .A(u2__abc_52138_new_n11225_), .Y(u2__abc_52138_new_n11226_));
INVX1 INVX1_1701 ( .A(u2__abc_52138_new_n6004_), .Y(u2__abc_52138_new_n11234_));
INVX1 INVX1_1702 ( .A(u2__abc_52138_new_n11236_), .Y(u2__abc_52138_new_n11237_));
INVX1 INVX1_1703 ( .A(u2__abc_52138_new_n5978_), .Y(u2__abc_52138_new_n11286_));
INVX1 INVX1_1704 ( .A(u2__abc_52138_new_n5973_), .Y(u2__abc_52138_new_n11287_));
INVX1 INVX1_1705 ( .A(u2__abc_52138_new_n5975_), .Y(u2__abc_52138_new_n11300_));
INVX1 INVX1_1706 ( .A(u2__abc_52138_new_n5982_), .Y(u2__abc_52138_new_n11309_));
INVX1 INVX1_1707 ( .A(u2__abc_52138_new_n11314_), .Y(u2__abc_52138_new_n11315_));
INVX1 INVX1_1708 ( .A(u2__abc_52138_new_n5956_), .Y(u2__abc_52138_new_n11331_));
INVX1 INVX1_1709 ( .A(u2__abc_52138_new_n11332_), .Y(u2__abc_52138_new_n11333_));
INVX1 INVX1_171 ( .A(fracta_112_), .Y(_abc_65734_new_n1448_));
INVX1 INVX1_1710 ( .A(u2__abc_52138_new_n11334_), .Y(u2__abc_52138_new_n11335_));
INVX1 INVX1_1711 ( .A(u2__abc_52138_new_n5945_), .Y(u2__abc_52138_new_n11343_));
INVX1 INVX1_1712 ( .A(u2__abc_52138_new_n5966_), .Y(u2__abc_52138_new_n11353_));
INVX1 INVX1_1713 ( .A(u2__abc_52138_new_n11360_), .Y(u2__abc_52138_new_n11361_));
INVX1 INVX1_1714 ( .A(u2__abc_52138_new_n3009_), .Y(u2__abc_52138_new_n11369_));
INVX1 INVX1_1715 ( .A(u2_cnt_0_), .Y(u2__abc_52138_new_n11377_));
INVX1 INVX1_1716 ( .A(u2_cnt_2_), .Y(u2__abc_52138_new_n11386_));
INVX1 INVX1_1717 ( .A(u2__abc_52138_new_n11392_), .Y(u2__abc_52138_new_n11393_));
INVX1 INVX1_1718 ( .A(u2__abc_52138_new_n2965_), .Y(u2__abc_52138_new_n11394_));
INVX1 INVX1_1719 ( .A(u2__abc_52138_new_n11401_), .Y(u2__abc_52138_new_n11402_));
INVX1 INVX1_172 ( .A(\a[113] ), .Y(_abc_65734_new_n1456_));
INVX1 INVX1_1720 ( .A(u2_cnt_6_), .Y(u2__abc_52138_new_n11406_));
INVX1 INVX1_1721 ( .A(u2_remLo_32_), .Y(u2__abc_52138_new_n11507_));
INVX1 INVX1_1722 ( .A(u2_remLo_33_), .Y(u2__abc_52138_new_n11512_));
INVX1 INVX1_1723 ( .A(u2__abc_52138_new_n11514_), .Y(u2__abc_52138_new_n11515_));
INVX1 INVX1_1724 ( .A(u2_remLo_35_), .Y(u2__abc_52138_new_n11521_));
INVX1 INVX1_1725 ( .A(u2_remLo_36_), .Y(u2__abc_52138_new_n11524_));
INVX1 INVX1_1726 ( .A(u2__abc_52138_new_n11526_), .Y(u2__abc_52138_new_n11527_));
INVX1 INVX1_1727 ( .A(u2_remLo_37_), .Y(u2__abc_52138_new_n11530_));
INVX1 INVX1_1728 ( .A(u2_remLo_38_), .Y(u2__abc_52138_new_n11533_));
INVX1 INVX1_1729 ( .A(u2_remLo_39_), .Y(u2__abc_52138_new_n11536_));
INVX1 INVX1_173 ( .A(\a[114] ), .Y(_abc_65734_new_n1458_));
INVX1 INVX1_1730 ( .A(u2_remLo_40_), .Y(u2__abc_52138_new_n11539_));
INVX1 INVX1_1731 ( .A(u2_remLo_41_), .Y(u2__abc_52138_new_n11542_));
INVX1 INVX1_1732 ( .A(u2_remLo_42_), .Y(u2__abc_52138_new_n11545_));
INVX1 INVX1_1733 ( .A(u2_remLo_43_), .Y(u2__abc_52138_new_n11548_));
INVX1 INVX1_1734 ( .A(u2_remLo_44_), .Y(u2__abc_52138_new_n11551_));
INVX1 INVX1_1735 ( .A(u2_remLo_45_), .Y(u2__abc_52138_new_n11554_));
INVX1 INVX1_1736 ( .A(u2_remLo_47_), .Y(u2__abc_52138_new_n11560_));
INVX1 INVX1_1737 ( .A(u2_remLo_48_), .Y(u2__abc_52138_new_n11563_));
INVX1 INVX1_1738 ( .A(u2__abc_52138_new_n11565_), .Y(u2__abc_52138_new_n11566_));
INVX1 INVX1_1739 ( .A(u2_remLo_49_), .Y(u2__abc_52138_new_n11569_));
INVX1 INVX1_174 ( .A(\a[115] ), .Y(_abc_65734_new_n1463_));
INVX1 INVX1_1740 ( .A(u2_remLo_50_), .Y(u2__abc_52138_new_n11572_));
INVX1 INVX1_1741 ( .A(u2_remLo_51_), .Y(u2__abc_52138_new_n11575_));
INVX1 INVX1_1742 ( .A(u2_remLo_52_), .Y(u2__abc_52138_new_n11578_));
INVX1 INVX1_1743 ( .A(u2_remLo_53_), .Y(u2__abc_52138_new_n11581_));
INVX1 INVX1_1744 ( .A(u2_remLo_54_), .Y(u2__abc_52138_new_n11584_));
INVX1 INVX1_1745 ( .A(u2_remLo_55_), .Y(u2__abc_52138_new_n11587_));
INVX1 INVX1_1746 ( .A(u2_remLo_56_), .Y(u2__abc_52138_new_n11590_));
INVX1 INVX1_1747 ( .A(u2_remLo_57_), .Y(u2__abc_52138_new_n11593_));
INVX1 INVX1_1748 ( .A(u2_remLo_58_), .Y(u2__abc_52138_new_n11596_));
INVX1 INVX1_1749 ( .A(u2_remLo_59_), .Y(u2__abc_52138_new_n11599_));
INVX1 INVX1_175 ( .A(\a[116] ), .Y(_abc_65734_new_n1473_));
INVX1 INVX1_1750 ( .A(u2_remLo_60_), .Y(u2__abc_52138_new_n11602_));
INVX1 INVX1_1751 ( .A(u2_remLo_62_), .Y(u2__abc_52138_new_n11608_));
INVX1 INVX1_1752 ( .A(u2_remLo_63_), .Y(u2__abc_52138_new_n11611_));
INVX1 INVX1_1753 ( .A(u2_remLo_64_), .Y(u2__abc_52138_new_n11614_));
INVX1 INVX1_1754 ( .A(u2_remLo_66_), .Y(u2__abc_52138_new_n11620_));
INVX1 INVX1_1755 ( .A(u2_remLo_67_), .Y(u2__abc_52138_new_n11623_));
INVX1 INVX1_1756 ( .A(u2__abc_52138_new_n11625_), .Y(u2__abc_52138_new_n11626_));
INVX1 INVX1_1757 ( .A(u2_remLo_68_), .Y(u2__abc_52138_new_n11629_));
INVX1 INVX1_1758 ( .A(u2_remLo_69_), .Y(u2__abc_52138_new_n11632_));
INVX1 INVX1_1759 ( .A(u2_remLo_70_), .Y(u2__abc_52138_new_n11635_));
INVX1 INVX1_176 ( .A(\a[117] ), .Y(_abc_65734_new_n1481_));
INVX1 INVX1_1760 ( .A(u2_remLo_71_), .Y(u2__abc_52138_new_n11638_));
INVX1 INVX1_1761 ( .A(u2_remLo_72_), .Y(u2__abc_52138_new_n11641_));
INVX1 INVX1_1762 ( .A(u2_remLo_73_), .Y(u2__abc_52138_new_n11644_));
INVX1 INVX1_1763 ( .A(u2_remLo_75_), .Y(u2__abc_52138_new_n11650_));
INVX1 INVX1_1764 ( .A(u2_remLo_76_), .Y(u2__abc_52138_new_n11653_));
INVX1 INVX1_1765 ( .A(u2__abc_52138_new_n11655_), .Y(u2__abc_52138_new_n11656_));
INVX1 INVX1_1766 ( .A(u2_remLo_77_), .Y(u2__abc_52138_new_n11659_));
INVX1 INVX1_1767 ( .A(u2_remLo_78_), .Y(u2__abc_52138_new_n11662_));
INVX1 INVX1_1768 ( .A(u2_remLo_79_), .Y(u2__abc_52138_new_n11665_));
INVX1 INVX1_1769 ( .A(u2_remLo_81_), .Y(u2__abc_52138_new_n11671_));
INVX1 INVX1_177 ( .A(_abc_65734_new_n1483_), .Y(_abc_65734_new_n1484_));
INVX1 INVX1_1770 ( .A(u2_remLo_82_), .Y(u2__abc_52138_new_n11674_));
INVX1 INVX1_1771 ( .A(u2_remLo_83_), .Y(u2__abc_52138_new_n11677_));
INVX1 INVX1_1772 ( .A(u2_remLo_84_), .Y(u2__abc_52138_new_n11680_));
INVX1 INVX1_1773 ( .A(u2_remLo_85_), .Y(u2__abc_52138_new_n11683_));
INVX1 INVX1_1774 ( .A(u2_remLo_86_), .Y(u2__abc_52138_new_n11686_));
INVX1 INVX1_1775 ( .A(u2_remLo_87_), .Y(u2__abc_52138_new_n11689_));
INVX1 INVX1_1776 ( .A(u2_remLo_88_), .Y(u2__abc_52138_new_n11692_));
INVX1 INVX1_1777 ( .A(u2_remLo_89_), .Y(u2__abc_52138_new_n11695_));
INVX1 INVX1_1778 ( .A(u2_remLo_90_), .Y(u2__abc_52138_new_n11698_));
INVX1 INVX1_1779 ( .A(u2_remLo_91_), .Y(u2__abc_52138_new_n11701_));
INVX1 INVX1_178 ( .A(\a[118] ), .Y(_abc_65734_new_n1493_));
INVX1 INVX1_1780 ( .A(u2_remLo_92_), .Y(u2__abc_52138_new_n11704_));
INVX1 INVX1_1781 ( .A(u2_remLo_93_), .Y(u2__abc_52138_new_n11707_));
INVX1 INVX1_1782 ( .A(u2_remLo_94_), .Y(u2__abc_52138_new_n11710_));
INVX1 INVX1_1783 ( .A(u2_remLo_95_), .Y(u2__abc_52138_new_n11713_));
INVX1 INVX1_1784 ( .A(u2_remLo_96_), .Y(u2__abc_52138_new_n11716_));
INVX1 INVX1_1785 ( .A(u2_remLo_98_), .Y(u2__abc_52138_new_n11724_));
INVX1 INVX1_1786 ( .A(u2_remLo_99_), .Y(u2__abc_52138_new_n11728_));
INVX1 INVX1_1787 ( .A(u2__abc_52138_new_n11730_), .Y(u2__abc_52138_new_n11731_));
INVX1 INVX1_1788 ( .A(u2_remLo_100_), .Y(u2__abc_52138_new_n11734_));
INVX1 INVX1_1789 ( .A(u2_remLo_101_), .Y(u2__abc_52138_new_n11737_));
INVX1 INVX1_179 ( .A(\a[119] ), .Y(_abc_65734_new_n1500_));
INVX1 INVX1_1790 ( .A(u2_remLo_102_), .Y(u2__abc_52138_new_n11740_));
INVX1 INVX1_1791 ( .A(u2_remLo_103_), .Y(u2__abc_52138_new_n11743_));
INVX1 INVX1_1792 ( .A(u2_remLo_104_), .Y(u2__abc_52138_new_n11746_));
INVX1 INVX1_1793 ( .A(u2_remLo_105_), .Y(u2__abc_52138_new_n11749_));
INVX1 INVX1_1794 ( .A(u2_remLo_106_), .Y(u2__abc_52138_new_n11752_));
INVX1 INVX1_1795 ( .A(u2_remLo_107_), .Y(u2__abc_52138_new_n11755_));
INVX1 INVX1_1796 ( .A(u2_remLo_108_), .Y(u2__abc_52138_new_n11758_));
INVX1 INVX1_1797 ( .A(u2_remLo_109_), .Y(u2__abc_52138_new_n11761_));
INVX1 INVX1_1798 ( .A(u2_remLo_111_), .Y(u2__abc_52138_new_n11767_));
INVX1 INVX1_1799 ( .A(u2_remLo_112_), .Y(u2__abc_52138_new_n11770_));
INVX1 INVX1_18 ( .A(sqrto_92_), .Y(_abc_65734_new_n878_));
INVX1 INVX1_180 ( .A(\a[120] ), .Y(_abc_65734_new_n1510_));
INVX1 INVX1_1800 ( .A(u2_remLo_113_), .Y(u2__abc_52138_new_n11773_));
INVX1 INVX1_1801 ( .A(u2_remLo_115_), .Y(u2__abc_52138_new_n11779_));
INVX1 INVX1_1802 ( .A(u2_remLo_116_), .Y(u2__abc_52138_new_n11782_));
INVX1 INVX1_1803 ( .A(u2__abc_52138_new_n11784_), .Y(u2__abc_52138_new_n11785_));
INVX1 INVX1_1804 ( .A(u2_remLo_117_), .Y(u2__abc_52138_new_n11788_));
INVX1 INVX1_1805 ( .A(u2_remLo_118_), .Y(u2__abc_52138_new_n11791_));
INVX1 INVX1_1806 ( .A(u2_remLo_119_), .Y(u2__abc_52138_new_n11794_));
INVX1 INVX1_1807 ( .A(u2_remLo_120_), .Y(u2__abc_52138_new_n11797_));
INVX1 INVX1_1808 ( .A(u2_remLo_121_), .Y(u2__abc_52138_new_n11800_));
INVX1 INVX1_1809 ( .A(u2_remLo_122_), .Y(u2__abc_52138_new_n11803_));
INVX1 INVX1_181 ( .A(\a[121] ), .Y(_abc_65734_new_n1523_));
INVX1 INVX1_1810 ( .A(u2_remLo_123_), .Y(u2__abc_52138_new_n11806_));
INVX1 INVX1_1811 ( .A(u2_remLo_124_), .Y(u2__abc_52138_new_n11809_));
INVX1 INVX1_1812 ( .A(u2_remLo_125_), .Y(u2__abc_52138_new_n11812_));
INVX1 INVX1_1813 ( .A(u2_remLo_126_), .Y(u2__abc_52138_new_n11815_));
INVX1 INVX1_1814 ( .A(u2_remLo_127_), .Y(u2__abc_52138_new_n11818_));
INVX1 INVX1_1815 ( .A(u2_remLo_128_), .Y(u2__abc_52138_new_n11821_));
INVX1 INVX1_1816 ( .A(u2_remLo_130_), .Y(u2__abc_52138_new_n11827_));
INVX1 INVX1_1817 ( .A(u2_remLo_131_), .Y(u2__abc_52138_new_n11830_));
INVX1 INVX1_1818 ( .A(u2__abc_52138_new_n11832_), .Y(u2__abc_52138_new_n11833_));
INVX1 INVX1_1819 ( .A(u2_remLo_132_), .Y(u2__abc_52138_new_n11836_));
INVX1 INVX1_182 ( .A(\a[122] ), .Y(_abc_65734_new_n1533_));
INVX1 INVX1_1820 ( .A(u2_remLo_133_), .Y(u2__abc_52138_new_n11839_));
INVX1 INVX1_1821 ( .A(u2_remLo_134_), .Y(u2__abc_52138_new_n11843_));
INVX1 INVX1_1822 ( .A(u2_remLo_135_), .Y(u2__abc_52138_new_n11846_));
INVX1 INVX1_1823 ( .A(u2_remLo_136_), .Y(u2__abc_52138_new_n11849_));
INVX1 INVX1_1824 ( .A(u2_remLo_137_), .Y(u2__abc_52138_new_n11852_));
INVX1 INVX1_1825 ( .A(u2_remLo_138_), .Y(u2__abc_52138_new_n11855_));
INVX1 INVX1_1826 ( .A(u2_remLo_139_), .Y(u2__abc_52138_new_n11858_));
INVX1 INVX1_1827 ( .A(u2_remLo_140_), .Y(u2__abc_52138_new_n11861_));
INVX1 INVX1_1828 ( .A(u2_remLo_141_), .Y(u2__abc_52138_new_n11864_));
INVX1 INVX1_1829 ( .A(u2_remLo_143_), .Y(u2__abc_52138_new_n11870_));
INVX1 INVX1_183 ( .A(_abc_65734_new_n1534_), .Y(_abc_65734_new_n1535_));
INVX1 INVX1_1830 ( .A(u2_remLo_144_), .Y(u2__abc_52138_new_n11873_));
INVX1 INVX1_1831 ( .A(u2_remLo_145_), .Y(u2__abc_52138_new_n11876_));
INVX1 INVX1_1832 ( .A(u2_remLo_146_), .Y(u2__abc_52138_new_n11879_));
INVX1 INVX1_1833 ( .A(u2_remLo_147_), .Y(u2__abc_52138_new_n11882_));
INVX1 INVX1_1834 ( .A(u2_remLo_148_), .Y(u2__abc_52138_new_n11885_));
INVX1 INVX1_1835 ( .A(u2_remLo_149_), .Y(u2__abc_52138_new_n11888_));
INVX1 INVX1_1836 ( .A(u2_remLo_150_), .Y(u2__abc_52138_new_n11891_));
INVX1 INVX1_1837 ( .A(u2_remLo_151_), .Y(u2__abc_52138_new_n11894_));
INVX1 INVX1_1838 ( .A(u2_remLo_152_), .Y(u2__abc_52138_new_n11897_));
INVX1 INVX1_1839 ( .A(u2_remLo_153_), .Y(u2__abc_52138_new_n11900_));
INVX1 INVX1_184 ( .A(\a[123] ), .Y(_abc_65734_new_n1545_));
INVX1 INVX1_1840 ( .A(u2_remLo_154_), .Y(u2__abc_52138_new_n11903_));
INVX1 INVX1_1841 ( .A(u2_remLo_155_), .Y(u2__abc_52138_new_n11906_));
INVX1 INVX1_1842 ( .A(u2_remLo_156_), .Y(u2__abc_52138_new_n11909_));
INVX1 INVX1_1843 ( .A(u2_remLo_157_), .Y(u2__abc_52138_new_n11912_));
INVX1 INVX1_1844 ( .A(u2_remLo_158_), .Y(u2__abc_52138_new_n11915_));
INVX1 INVX1_1845 ( .A(u2_remLo_159_), .Y(u2__abc_52138_new_n11918_));
INVX1 INVX1_1846 ( .A(u2_remLo_162_), .Y(u2__abc_52138_new_n11927_));
INVX1 INVX1_1847 ( .A(u2_remLo_163_), .Y(u2__abc_52138_new_n11930_));
INVX1 INVX1_1848 ( .A(u2__abc_52138_new_n11932_), .Y(u2__abc_52138_new_n11933_));
INVX1 INVX1_1849 ( .A(u2_remLo_164_), .Y(u2__abc_52138_new_n11936_));
INVX1 INVX1_185 ( .A(\a[124] ), .Y(_abc_65734_new_n1555_));
INVX1 INVX1_1850 ( .A(u2_remLo_165_), .Y(u2__abc_52138_new_n11939_));
INVX1 INVX1_1851 ( .A(u2_remLo_166_), .Y(u2__abc_52138_new_n11942_));
INVX1 INVX1_1852 ( .A(u2_remLo_167_), .Y(u2__abc_52138_new_n11945_));
INVX1 INVX1_1853 ( .A(u2_remLo_168_), .Y(u2__abc_52138_new_n11948_));
INVX1 INVX1_1854 ( .A(u2_remLo_169_), .Y(u2__abc_52138_new_n11951_));
INVX1 INVX1_1855 ( .A(u2_remLo_170_), .Y(u2__abc_52138_new_n11954_));
INVX1 INVX1_1856 ( .A(u2_remLo_171_), .Y(u2__abc_52138_new_n11957_));
INVX1 INVX1_1857 ( .A(u2_remLo_172_), .Y(u2__abc_52138_new_n11960_));
INVX1 INVX1_1858 ( .A(u2_remLo_173_), .Y(u2__abc_52138_new_n11963_));
INVX1 INVX1_1859 ( .A(u2_remLo_174_), .Y(u2__abc_52138_new_n11966_));
INVX1 INVX1_186 ( .A(_abc_65734_new_n1550_), .Y(_abc_65734_new_n1558_));
INVX1 INVX1_1860 ( .A(u2_remLo_175_), .Y(u2__abc_52138_new_n11970_));
INVX1 INVX1_1861 ( .A(u2_remLo_176_), .Y(u2__abc_52138_new_n11973_));
INVX1 INVX1_1862 ( .A(u2_remLo_177_), .Y(u2__abc_52138_new_n11976_));
INVX1 INVX1_1863 ( .A(u2_remLo_178_), .Y(u2__abc_52138_new_n11979_));
INVX1 INVX1_1864 ( .A(u2_remLo_179_), .Y(u2__abc_52138_new_n11982_));
INVX1 INVX1_1865 ( .A(u2_remLo_180_), .Y(u2__abc_52138_new_n11985_));
INVX1 INVX1_1866 ( .A(u2_remLo_181_), .Y(u2__abc_52138_new_n11988_));
INVX1 INVX1_1867 ( .A(u2_remLo_182_), .Y(u2__abc_52138_new_n11991_));
INVX1 INVX1_1868 ( .A(u2_remLo_183_), .Y(u2__abc_52138_new_n11994_));
INVX1 INVX1_1869 ( .A(u2_remLo_184_), .Y(u2__abc_52138_new_n11997_));
INVX1 INVX1_187 ( .A(\a[125] ), .Y(_abc_65734_new_n1563_));
INVX1 INVX1_1870 ( .A(u2_remLo_185_), .Y(u2__abc_52138_new_n12000_));
INVX1 INVX1_1871 ( .A(u2_remLo_186_), .Y(u2__abc_52138_new_n12003_));
INVX1 INVX1_1872 ( .A(u2_remLo_187_), .Y(u2__abc_52138_new_n12006_));
INVX1 INVX1_1873 ( .A(u2_remLo_188_), .Y(u2__abc_52138_new_n12009_));
INVX1 INVX1_1874 ( .A(u2_remLo_189_), .Y(u2__abc_52138_new_n12012_));
INVX1 INVX1_1875 ( .A(u2_remLo_190_), .Y(u2__abc_52138_new_n12015_));
INVX1 INVX1_1876 ( .A(u2_remLo_191_), .Y(u2__abc_52138_new_n12018_));
INVX1 INVX1_1877 ( .A(u2_remLo_192_), .Y(u2__abc_52138_new_n12021_));
INVX1 INVX1_1878 ( .A(u2_remLo_194_), .Y(u2__abc_52138_new_n12027_));
INVX1 INVX1_1879 ( .A(u2_remLo_195_), .Y(u2__abc_52138_new_n12030_));
INVX1 INVX1_188 ( .A(_abc_65734_new_n1567_), .Y(_abc_65734_new_n1571_));
INVX1 INVX1_1880 ( .A(u2__abc_52138_new_n12032_), .Y(u2__abc_52138_new_n12033_));
INVX1 INVX1_1881 ( .A(u2_remLo_196_), .Y(u2__abc_52138_new_n12036_));
INVX1 INVX1_1882 ( .A(u2_remLo_197_), .Y(u2__abc_52138_new_n12039_));
INVX1 INVX1_1883 ( .A(u2_remLo_198_), .Y(u2__abc_52138_new_n12042_));
INVX1 INVX1_1884 ( .A(u2_remLo_199_), .Y(u2__abc_52138_new_n12045_));
INVX1 INVX1_1885 ( .A(u2_remLo_200_), .Y(u2__abc_52138_new_n12048_));
INVX1 INVX1_1886 ( .A(u2_remLo_201_), .Y(u2__abc_52138_new_n12051_));
INVX1 INVX1_1887 ( .A(u2_remLo_203_), .Y(u2__abc_52138_new_n12057_));
INVX1 INVX1_1888 ( .A(u2_remLo_204_), .Y(u2__abc_52138_new_n12060_));
INVX1 INVX1_1889 ( .A(u2__abc_52138_new_n12062_), .Y(u2__abc_52138_new_n12063_));
INVX1 INVX1_189 ( .A(\a[112] ), .Y(u1__abc_51895_new_n144_));
INVX1 INVX1_1890 ( .A(u2_remLo_205_), .Y(u2__abc_52138_new_n12066_));
INVX1 INVX1_1891 ( .A(u2_remLo_206_), .Y(u2__abc_52138_new_n12069_));
INVX1 INVX1_1892 ( .A(u2_remLo_207_), .Y(u2__abc_52138_new_n12073_));
INVX1 INVX1_1893 ( .A(u2_remLo_208_), .Y(u2__abc_52138_new_n12076_));
INVX1 INVX1_1894 ( .A(u2_remLo_209_), .Y(u2__abc_52138_new_n12079_));
INVX1 INVX1_1895 ( .A(u2_remLo_210_), .Y(u2__abc_52138_new_n12082_));
INVX1 INVX1_1896 ( .A(u2_remLo_211_), .Y(u2__abc_52138_new_n12085_));
INVX1 INVX1_1897 ( .A(u2_remLo_212_), .Y(u2__abc_52138_new_n12088_));
INVX1 INVX1_1898 ( .A(u2_remLo_213_), .Y(u2__abc_52138_new_n12091_));
INVX1 INVX1_1899 ( .A(u2_remLo_214_), .Y(u2__abc_52138_new_n12094_));
INVX1 INVX1_19 ( .A(sqrto_93_), .Y(_abc_65734_new_n881_));
INVX1 INVX1_190 ( .A(u1_xinf), .Y(u1__abc_51895_new_n278_));
INVX1 INVX1_1900 ( .A(u2_remLo_215_), .Y(u2__abc_52138_new_n12097_));
INVX1 INVX1_1901 ( .A(u2_remLo_216_), .Y(u2__abc_52138_new_n12100_));
INVX1 INVX1_1902 ( .A(u2_remLo_217_), .Y(u2__abc_52138_new_n12103_));
INVX1 INVX1_1903 ( .A(u2_remLo_218_), .Y(u2__abc_52138_new_n12106_));
INVX1 INVX1_1904 ( .A(u2_remLo_219_), .Y(u2__abc_52138_new_n12109_));
INVX1 INVX1_1905 ( .A(u2_remLo_220_), .Y(u2__abc_52138_new_n12112_));
INVX1 INVX1_1906 ( .A(u2_remLo_221_), .Y(u2__abc_52138_new_n12115_));
INVX1 INVX1_1907 ( .A(u2_remLo_222_), .Y(u2__abc_52138_new_n12118_));
INVX1 INVX1_1908 ( .A(u2_remLo_223_), .Y(u2__abc_52138_new_n12121_));
INVX1 INVX1_1909 ( .A(u2_remLo_224_), .Y(u2__abc_52138_new_n12124_));
INVX1 INVX1_191 ( .A(ld), .Y(u2__abc_52138_new_n2962_));
INVX1 INVX1_1910 ( .A(u2_remLo_227_), .Y(u2__abc_52138_new_n12133_));
INVX1 INVX1_1911 ( .A(u2__abc_52138_new_n12135_), .Y(u2__abc_52138_new_n12136_));
INVX1 INVX1_1912 ( .A(u2_remLo_228_), .Y(u2__abc_52138_new_n12139_));
INVX1 INVX1_1913 ( .A(u2__abc_52138_new_n12141_), .Y(u2__abc_52138_new_n12142_));
INVX1 INVX1_1914 ( .A(u2_remLo_229_), .Y(u2__abc_52138_new_n12145_));
INVX1 INVX1_1915 ( .A(u2_remLo_230_), .Y(u2__abc_52138_new_n12148_));
INVX1 INVX1_1916 ( .A(u2_remLo_231_), .Y(u2__abc_52138_new_n12151_));
INVX1 INVX1_1917 ( .A(u2_remLo_232_), .Y(u2__abc_52138_new_n12154_));
INVX1 INVX1_1918 ( .A(u2_remLo_233_), .Y(u2__abc_52138_new_n12157_));
INVX1 INVX1_1919 ( .A(u2_remLo_234_), .Y(u2__abc_52138_new_n12160_));
INVX1 INVX1_192 ( .A(u2_state_0_), .Y(u2__abc_52138_new_n2963_));
INVX1 INVX1_1920 ( .A(u2_remLo_235_), .Y(u2__abc_52138_new_n12164_));
INVX1 INVX1_1921 ( .A(u2_remLo_236_), .Y(u2__abc_52138_new_n12167_));
INVX1 INVX1_1922 ( .A(u2_remLo_237_), .Y(u2__abc_52138_new_n12170_));
INVX1 INVX1_1923 ( .A(u2_remLo_238_), .Y(u2__abc_52138_new_n12173_));
INVX1 INVX1_1924 ( .A(u2_remLo_239_), .Y(u2__abc_52138_new_n12176_));
INVX1 INVX1_1925 ( .A(u2_remLo_241_), .Y(u2__abc_52138_new_n12182_));
INVX1 INVX1_1926 ( .A(u2_remLo_242_), .Y(u2__abc_52138_new_n12185_));
INVX1 INVX1_1927 ( .A(u2_remLo_243_), .Y(u2__abc_52138_new_n12188_));
INVX1 INVX1_1928 ( .A(u2_remLo_244_), .Y(u2__abc_52138_new_n12191_));
INVX1 INVX1_1929 ( .A(u2_remLo_245_), .Y(u2__abc_52138_new_n12194_));
INVX1 INVX1_193 ( .A(ce), .Y(u2__abc_52138_new_n2966_));
INVX1 INVX1_1930 ( .A(u2_remLo_246_), .Y(u2__abc_52138_new_n12197_));
INVX1 INVX1_1931 ( .A(u2_remLo_247_), .Y(u2__abc_52138_new_n12200_));
INVX1 INVX1_1932 ( .A(u2_remLo_248_), .Y(u2__abc_52138_new_n12203_));
INVX1 INVX1_1933 ( .A(u2_remLo_249_), .Y(u2__abc_52138_new_n12206_));
INVX1 INVX1_1934 ( .A(u2_remLo_250_), .Y(u2__abc_52138_new_n12209_));
INVX1 INVX1_1935 ( .A(u2_remLo_251_), .Y(u2__abc_52138_new_n12212_));
INVX1 INVX1_1936 ( .A(u2_remLo_252_), .Y(u2__abc_52138_new_n12215_));
INVX1 INVX1_1937 ( .A(u2_remLo_253_), .Y(u2__abc_52138_new_n12218_));
INVX1 INVX1_1938 ( .A(u2_remLo_254_), .Y(u2__abc_52138_new_n12221_));
INVX1 INVX1_1939 ( .A(u2_remLo_255_), .Y(u2__abc_52138_new_n12224_));
INVX1 INVX1_194 ( .A(u2_cnt_4_), .Y(u2__abc_52138_new_n2967_));
INVX1 INVX1_1940 ( .A(u2_remLo_256_), .Y(u2__abc_52138_new_n12227_));
INVX1 INVX1_1941 ( .A(u2__abc_52138_new_n3207_), .Y(u2__abc_52138_new_n12844_));
INVX1 INVX1_1942 ( .A(u2__abc_52138_new_n3208_), .Y(u2__abc_52138_new_n12845_));
INVX1 INVX1_1943 ( .A(u2__abc_52138_new_n3232_), .Y(u2__abc_52138_new_n12851_));
INVX1 INVX1_1944 ( .A(u2__abc_52138_new_n3395_), .Y(u2__abc_52138_new_n12858_));
INVX1 INVX1_1945 ( .A(u2__abc_52138_new_n3483_), .Y(u2__abc_52138_new_n12876_));
INVX1 INVX1_1946 ( .A(u2__abc_52138_new_n3827_), .Y(u2__abc_52138_new_n12904_));
INVX1 INVX1_1947 ( .A(u2__abc_52138_new_n3904_), .Y(u2__abc_52138_new_n12906_));
INVX1 INVX1_1948 ( .A(u2__abc_52138_new_n3953_), .Y(u2__abc_52138_new_n12931_));
INVX1 INVX1_1949 ( .A(u2__abc_52138_new_n4720_), .Y(u2__abc_52138_new_n12955_));
INVX1 INVX1_195 ( .A(u2__abc_52138_new_n2969_), .Y(u2__abc_52138_new_n2970_));
INVX1 INVX1_1950 ( .A(u2__abc_52138_new_n4812_), .Y(u2__abc_52138_new_n12973_));
INVX1 INVX1_1951 ( .A(u2__abc_52138_new_n4832_), .Y(u2__abc_52138_new_n12982_));
INVX1 INVX1_1952 ( .A(u2__abc_52138_new_n4886_), .Y(u2__abc_52138_new_n12997_));
INVX1 INVX1_1953 ( .A(u2__abc_52138_new_n4919_), .Y(u2__abc_52138_new_n13008_));
INVX1 INVX1_1954 ( .A(u2__abc_52138_new_n4925_), .Y(u2__abc_52138_new_n13012_));
INVX1 INVX1_1955 ( .A(u2__abc_52138_new_n6332_), .Y(u2__abc_52138_new_n13040_));
INVX1 INVX1_1956 ( .A(u2__abc_52138_new_n6440_), .Y(u2__abc_52138_new_n13041_));
INVX1 INVX1_1957 ( .A(u2__abc_52138_new_n13067_), .Y(u2__abc_52138_new_n13068_));
INVX1 INVX1_1958 ( .A(u2__abc_52138_new_n13098_), .Y(u2__abc_52138_new_n13099_));
INVX1 INVX1_1959 ( .A(u2__abc_52138_new_n13129_), .Y(u2__abc_52138_new_n13130_));
INVX1 INVX1_196 ( .A(u2__abc_52138_new_n2972_), .Y(u2__abc_52138_new_n2973_));
INVX1 INVX1_1960 ( .A(u2__abc_52138_new_n13160_), .Y(u2__abc_52138_new_n13161_));
INVX1 INVX1_1961 ( .A(u2__abc_52138_new_n13191_), .Y(u2__abc_52138_new_n13192_));
INVX1 INVX1_1962 ( .A(u2__abc_52138_new_n13222_), .Y(u2__abc_52138_new_n13223_));
INVX1 INVX1_1963 ( .A(u2__abc_52138_new_n13253_), .Y(u2__abc_52138_new_n13254_));
INVX1 INVX1_1964 ( .A(u2__abc_52138_new_n13284_), .Y(u2__abc_52138_new_n13285_));
INVX1 INVX1_1965 ( .A(sqrto_34_), .Y(u2__abc_52138_new_n13310_));
INVX1 INVX1_1966 ( .A(u2__abc_52138_new_n13316_), .Y(u2__abc_52138_new_n13317_));
INVX1 INVX1_1967 ( .A(u2__abc_52138_new_n13347_), .Y(u2__abc_52138_new_n13348_));
INVX1 INVX1_1968 ( .A(u2__abc_52138_new_n13378_), .Y(u2__abc_52138_new_n13379_));
INVX1 INVX1_1969 ( .A(u2__abc_52138_new_n13409_), .Y(u2__abc_52138_new_n13410_));
INVX1 INVX1_197 ( .A(u2_cnt_1_), .Y(u2__abc_52138_new_n2974_));
INVX1 INVX1_1970 ( .A(u2__abc_52138_new_n13440_), .Y(u2__abc_52138_new_n13441_));
INVX1 INVX1_1971 ( .A(u2__abc_52138_new_n13471_), .Y(u2__abc_52138_new_n13472_));
INVX1 INVX1_1972 ( .A(u2__abc_52138_new_n13502_), .Y(u2__abc_52138_new_n13503_));
INVX1 INVX1_1973 ( .A(u2__abc_52138_new_n13533_), .Y(u2__abc_52138_new_n13534_));
INVX1 INVX1_1974 ( .A(u2__abc_52138_new_n13564_), .Y(u2__abc_52138_new_n13565_));
INVX1 INVX1_1975 ( .A(u2__abc_52138_new_n13595_), .Y(u2__abc_52138_new_n13596_));
INVX1 INVX1_1976 ( .A(u2__abc_52138_new_n13626_), .Y(u2__abc_52138_new_n13627_));
INVX1 INVX1_1977 ( .A(u2__abc_52138_new_n13657_), .Y(u2__abc_52138_new_n13658_));
INVX1 INVX1_1978 ( .A(u2__abc_52138_new_n13688_), .Y(u2__abc_52138_new_n13689_));
INVX1 INVX1_1979 ( .A(u2__abc_52138_new_n13719_), .Y(u2__abc_52138_new_n13720_));
INVX1 INVX1_198 ( .A(u2__abc_52138_new_n2975_), .Y(u2__abc_52138_new_n2976_));
INVX1 INVX1_1980 ( .A(u2__abc_52138_new_n13750_), .Y(u2__abc_52138_new_n13751_));
INVX1 INVX1_1981 ( .A(u2__abc_52138_new_n13781_), .Y(u2__abc_52138_new_n13782_));
INVX1 INVX1_1982 ( .A(u2__abc_52138_new_n13812_), .Y(u2__abc_52138_new_n13813_));
INVX1 INVX1_1983 ( .A(u2__abc_52138_new_n13843_), .Y(u2__abc_52138_new_n13844_));
INVX1 INVX1_1984 ( .A(u2__abc_52138_new_n13874_), .Y(u2__abc_52138_new_n13875_));
INVX1 INVX1_1985 ( .A(u2__abc_52138_new_n13905_), .Y(u2__abc_52138_new_n13906_));
INVX1 INVX1_1986 ( .A(u2__abc_52138_new_n13936_), .Y(u2__abc_52138_new_n13937_));
INVX1 INVX1_1987 ( .A(sqrto_118_), .Y(u2__abc_52138_new_n13962_));
INVX1 INVX1_1988 ( .A(u2__abc_52138_new_n13968_), .Y(u2__abc_52138_new_n13969_));
INVX1 INVX1_1989 ( .A(u2__abc_52138_new_n13999_), .Y(u2__abc_52138_new_n14000_));
INVX1 INVX1_199 ( .A(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n2986_));
INVX1 INVX1_1990 ( .A(u2__abc_52138_new_n14030_), .Y(u2__abc_52138_new_n14031_));
INVX1 INVX1_1991 ( .A(sqrto_130_), .Y(u2__abc_52138_new_n14056_));
INVX1 INVX1_1992 ( .A(u2__abc_52138_new_n14062_), .Y(u2__abc_52138_new_n14063_));
INVX1 INVX1_1993 ( .A(u2__abc_52138_new_n14093_), .Y(u2__abc_52138_new_n14094_));
INVX1 INVX1_1994 ( .A(u2__abc_52138_new_n14124_), .Y(u2__abc_52138_new_n14125_));
INVX1 INVX1_1995 ( .A(u2__abc_52138_new_n14155_), .Y(u2__abc_52138_new_n14156_));
INVX1 INVX1_1996 ( .A(u2__abc_52138_new_n14186_), .Y(u2__abc_52138_new_n14187_));
INVX1 INVX1_1997 ( .A(u2__abc_52138_new_n14217_), .Y(u2__abc_52138_new_n14218_));
INVX1 INVX1_1998 ( .A(u2__abc_52138_new_n14248_), .Y(u2__abc_52138_new_n14249_));
INVX1 INVX1_1999 ( .A(u2__abc_52138_new_n14279_), .Y(u2__abc_52138_new_n14280_));
INVX1 INVX1_2 ( .A(sqrto_76_), .Y(_abc_65734_new_n830_));
INVX1 INVX1_20 ( .A(sqrto_94_), .Y(_abc_65734_new_n884_));
INVX1 INVX1_200 ( .A(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n2991_));
INVX1 INVX1_2000 ( .A(u2__abc_52138_new_n14310_), .Y(u2__abc_52138_new_n14311_));
INVX1 INVX1_2001 ( .A(u2__abc_52138_new_n14341_), .Y(u2__abc_52138_new_n14342_));
INVX1 INVX1_2002 ( .A(u2__abc_52138_new_n14372_), .Y(u2__abc_52138_new_n14373_));
INVX1 INVX1_2003 ( .A(u2__abc_52138_new_n14403_), .Y(u2__abc_52138_new_n14404_));
INVX1 INVX1_2004 ( .A(u2__abc_52138_new_n14434_), .Y(u2__abc_52138_new_n14435_));
INVX1 INVX1_2005 ( .A(u2__abc_52138_new_n14465_), .Y(u2__abc_52138_new_n14466_));
INVX1 INVX1_2006 ( .A(u2__abc_52138_new_n14496_), .Y(u2__abc_52138_new_n14497_));
INVX1 INVX1_2007 ( .A(u2__abc_52138_new_n14527_), .Y(u2__abc_52138_new_n14528_));
INVX1 INVX1_2008 ( .A(u2__abc_52138_new_n14558_), .Y(u2__abc_52138_new_n14559_));
INVX1 INVX1_2009 ( .A(u2__abc_52138_new_n14589_), .Y(u2__abc_52138_new_n14590_));
INVX1 INVX1_201 ( .A(u2_remHiShift_0_), .Y(u2__abc_52138_new_n2996_));
INVX1 INVX1_2010 ( .A(sqrto_202_), .Y(u2__abc_52138_new_n14615_));
INVX1 INVX1_2011 ( .A(u2__abc_52138_new_n14621_), .Y(u2__abc_52138_new_n14622_));
INVX1 INVX1_2012 ( .A(u2__abc_52138_new_n14652_), .Y(u2__abc_52138_new_n14653_));
INVX1 INVX1_2013 ( .A(u2__abc_52138_new_n14683_), .Y(u2__abc_52138_new_n14684_));
INVX1 INVX1_2014 ( .A(u2__abc_52138_new_n14714_), .Y(u2__abc_52138_new_n14715_));
INVX1 INVX1_2015 ( .A(u2__abc_52138_new_n14745_), .Y(u2__abc_52138_new_n14746_));
INVX1 INVX1_2016 ( .A(u2__abc_52138_new_n14776_), .Y(u2__abc_52138_new_n14777_));
INVX1 INVX1_2017 ( .A(u2__abc_52138_new_n14807_), .Y(u2__abc_52138_new_n14808_));
INVX1 INVX1_2018 ( .A(u2__abc_52138_new_n14838_), .Y(u2__abc_52138_new_n14839_));
INVX1 INVX1_2019 ( .A(u2__abc_52138_new_n14869_), .Y(u2__abc_52138_new_n14870_));
INVX1 INVX1_202 ( .A(u2_o_448_), .Y(u2__abc_52138_new_n2997_));
INVX1 INVX1_2020 ( .A(u2__abc_52138_new_n14900_), .Y(u2__abc_52138_new_n14901_));
INVX1 INVX1_2021 ( .A(u2__abc_52138_new_n14931_), .Y(u2__abc_52138_new_n14932_));
INVX1 INVX1_2022 ( .A(u2__abc_52138_new_n14962_), .Y(u2__abc_52138_new_n14963_));
INVX1 INVX1_2023 ( .A(u2__abc_52138_new_n14993_), .Y(u2__abc_52138_new_n14994_));
INVX1 INVX1_2024 ( .A(u2__abc_52138_new_n15024_), .Y(u2__abc_52138_new_n15025_));
INVX1 INVX1_2025 ( .A(u2__abc_52138_new_n15055_), .Y(u2__abc_52138_new_n15056_));
INVX1 INVX1_2026 ( .A(u2__abc_52138_new_n15086_), .Y(u2__abc_52138_new_n15087_));
INVX1 INVX1_2027 ( .A(u2__abc_52138_new_n15117_), .Y(u2__abc_52138_new_n15118_));
INVX1 INVX1_2028 ( .A(u2__abc_52138_new_n15148_), .Y(u2__abc_52138_new_n15149_));
INVX1 INVX1_2029 ( .A(u2__abc_52138_new_n15179_), .Y(u2__abc_52138_new_n15180_));
INVX1 INVX1_203 ( .A(u2_remHi_448_), .Y(u2__abc_52138_new_n2999_));
INVX1 INVX1_2030 ( .A(u2__abc_52138_new_n15210_), .Y(u2__abc_52138_new_n15211_));
INVX1 INVX1_2031 ( .A(u2__abc_52138_new_n15241_), .Y(u2__abc_52138_new_n15242_));
INVX1 INVX1_2032 ( .A(u2__abc_52138_new_n15272_), .Y(u2__abc_52138_new_n15273_));
INVX1 INVX1_2033 ( .A(u2__abc_52138_new_n15303_), .Y(u2__abc_52138_new_n15304_));
INVX1 INVX1_2034 ( .A(u2__abc_52138_new_n15334_), .Y(u2__abc_52138_new_n15335_));
INVX1 INVX1_2035 ( .A(u2__abc_52138_new_n15365_), .Y(u2__abc_52138_new_n15366_));
INVX1 INVX1_2036 ( .A(u2__abc_52138_new_n15396_), .Y(u2__abc_52138_new_n15397_));
INVX1 INVX1_2037 ( .A(u2__abc_52138_new_n15427_), .Y(u2__abc_52138_new_n15428_));
INVX1 INVX1_2038 ( .A(u2__abc_52138_new_n15458_), .Y(u2__abc_52138_new_n15459_));
INVX1 INVX1_2039 ( .A(u2_o_314_), .Y(u2__abc_52138_new_n15484_));
INVX1 INVX1_204 ( .A(u2_remHi_447_), .Y(u2__abc_52138_new_n3003_));
INVX1 INVX1_2040 ( .A(u2__abc_52138_new_n15490_), .Y(u2__abc_52138_new_n15491_));
INVX1 INVX1_2041 ( .A(u2__abc_52138_new_n15521_), .Y(u2__abc_52138_new_n15522_));
INVX1 INVX1_2042 ( .A(u2__abc_52138_new_n15552_), .Y(u2__abc_52138_new_n15553_));
INVX1 INVX1_2043 ( .A(u2__abc_52138_new_n15583_), .Y(u2__abc_52138_new_n15584_));
INVX1 INVX1_2044 ( .A(u2__abc_52138_new_n15614_), .Y(u2__abc_52138_new_n15615_));
INVX1 INVX1_2045 ( .A(u2_o_334_), .Y(u2__abc_52138_new_n15640_));
INVX1 INVX1_2046 ( .A(u2__abc_52138_new_n15646_), .Y(u2__abc_52138_new_n15647_));
INVX1 INVX1_2047 ( .A(u2_o_338_), .Y(u2__abc_52138_new_n15672_));
INVX1 INVX1_2048 ( .A(u2__abc_52138_new_n15678_), .Y(u2__abc_52138_new_n15679_));
INVX1 INVX1_2049 ( .A(u2__abc_52138_new_n15709_), .Y(u2__abc_52138_new_n15710_));
INVX1 INVX1_205 ( .A(u2_o_447_), .Y(u2__abc_52138_new_n3005_));
INVX1 INVX1_2050 ( .A(u2__abc_52138_new_n15740_), .Y(u2__abc_52138_new_n15741_));
INVX1 INVX1_2051 ( .A(u2__abc_52138_new_n15771_), .Y(u2__abc_52138_new_n15772_));
INVX1 INVX1_2052 ( .A(u2__abc_52138_new_n15802_), .Y(u2__abc_52138_new_n15803_));
INVX1 INVX1_2053 ( .A(u2__abc_52138_new_n15833_), .Y(u2__abc_52138_new_n15834_));
INVX1 INVX1_2054 ( .A(u2__abc_52138_new_n15864_), .Y(u2__abc_52138_new_n15865_));
INVX1 INVX1_2055 ( .A(u2__abc_52138_new_n15895_), .Y(u2__abc_52138_new_n15896_));
INVX1 INVX1_2056 ( .A(u2_o_369_), .Y(u2__abc_52138_new_n15913_));
INVX1 INVX1_2057 ( .A(u2__abc_52138_new_n15927_), .Y(u2__abc_52138_new_n15928_));
INVX1 INVX1_2058 ( .A(u2__abc_52138_new_n15958_), .Y(u2__abc_52138_new_n15959_));
INVX1 INVX1_2059 ( .A(u2__abc_52138_new_n15989_), .Y(u2__abc_52138_new_n15990_));
INVX1 INVX1_206 ( .A(u2_remHi_446_), .Y(u2__abc_52138_new_n3008_));
INVX1 INVX1_2060 ( .A(u2__abc_52138_new_n16020_), .Y(u2__abc_52138_new_n16021_));
INVX1 INVX1_2061 ( .A(u2__abc_52138_new_n16051_), .Y(u2__abc_52138_new_n16052_));
INVX1 INVX1_2062 ( .A(u2_o_390_), .Y(u2__abc_52138_new_n16077_));
INVX1 INVX1_2063 ( .A(u2__abc_52138_new_n16083_), .Y(u2__abc_52138_new_n16084_));
INVX1 INVX1_2064 ( .A(u2_o_391_), .Y(u2__abc_52138_new_n16086_));
INVX1 INVX1_2065 ( .A(u2_o_394_), .Y(u2__abc_52138_new_n16110_));
INVX1 INVX1_2066 ( .A(u2__abc_52138_new_n16116_), .Y(u2__abc_52138_new_n16117_));
INVX1 INVX1_2067 ( .A(u2__abc_52138_new_n16147_), .Y(u2__abc_52138_new_n16148_));
INVX1 INVX1_2068 ( .A(u2__abc_52138_new_n16178_), .Y(u2__abc_52138_new_n16179_));
INVX1 INVX1_2069 ( .A(u2__abc_52138_new_n16209_), .Y(u2__abc_52138_new_n16210_));
INVX1 INVX1_207 ( .A(u2_o_446_), .Y(u2__abc_52138_new_n3010_));
INVX1 INVX1_2070 ( .A(u2__abc_52138_new_n16240_), .Y(u2__abc_52138_new_n16241_));
INVX1 INVX1_2071 ( .A(u2__abc_52138_new_n16271_), .Y(u2__abc_52138_new_n16272_));
INVX1 INVX1_2072 ( .A(u2__abc_52138_new_n16302_), .Y(u2__abc_52138_new_n16303_));
INVX1 INVX1_2073 ( .A(u2__abc_52138_new_n16333_), .Y(u2__abc_52138_new_n16334_));
INVX1 INVX1_2074 ( .A(u2__abc_52138_new_n16364_), .Y(u2__abc_52138_new_n16365_));
INVX1 INVX1_2075 ( .A(u2__abc_52138_new_n16395_), .Y(u2__abc_52138_new_n16396_));
INVX1 INVX1_2076 ( .A(u2__abc_52138_new_n16426_), .Y(u2__abc_52138_new_n16427_));
INVX1 INVX1_2077 ( .A(u2__abc_52138_new_n16457_), .Y(u2__abc_52138_new_n16458_));
INVX1 INVX1_2078 ( .A(u2__abc_52138_new_n16488_), .Y(u2__abc_52138_new_n16489_));
INVX1 INVX1_2079 ( .A(u2__abc_52138_new_n16519_), .Y(u2__abc_52138_new_n16520_));
INVX1 INVX1_208 ( .A(u2__abc_52138_new_n3014_), .Y(u2__abc_52138_new_n3015_));
INVX1 INVX1_209 ( .A(u2_remHi_13_), .Y(u2__abc_52138_new_n3017_));
INVX1 INVX1_21 ( .A(sqrto_95_), .Y(_abc_65734_new_n887_));
INVX1 INVX1_210 ( .A(sqrto_13_), .Y(u2__abc_52138_new_n3019_));
INVX1 INVX1_211 ( .A(sqrto_11_), .Y(u2__abc_52138_new_n3022_));
INVX1 INVX1_212 ( .A(u2_remHi_11_), .Y(u2__abc_52138_new_n3024_));
INVX1 INVX1_213 ( .A(sqrto_10_), .Y(u2__abc_52138_new_n3027_));
INVX1 INVX1_214 ( .A(u2_remHi_10_), .Y(u2__abc_52138_new_n3029_));
INVX1 INVX1_215 ( .A(sqrto_9_), .Y(u2__abc_52138_new_n3035_));
INVX1 INVX1_216 ( .A(u2_remHi_9_), .Y(u2__abc_52138_new_n3037_));
INVX1 INVX1_217 ( .A(sqrto_7_), .Y(u2__abc_52138_new_n3040_));
INVX1 INVX1_218 ( .A(u2_remHi_7_), .Y(u2__abc_52138_new_n3042_));
INVX1 INVX1_219 ( .A(sqrto_6_), .Y(u2__abc_52138_new_n3045_));
INVX1 INVX1_22 ( .A(sqrto_96_), .Y(_abc_65734_new_n890_));
INVX1 INVX1_220 ( .A(u2_remHi_6_), .Y(u2__abc_52138_new_n3047_));
INVX1 INVX1_221 ( .A(u2_remHi_5_), .Y(u2__abc_52138_new_n3054_));
INVX1 INVX1_222 ( .A(sqrto_5_), .Y(u2__abc_52138_new_n3056_));
INVX1 INVX1_223 ( .A(sqrto_2_), .Y(u2__abc_52138_new_n3060_));
INVX1 INVX1_224 ( .A(u2_remHi_2_), .Y(u2__abc_52138_new_n3062_));
INVX1 INVX1_225 ( .A(u2_root_0_), .Y(u2__abc_52138_new_n3069_));
INVX1 INVX1_226 ( .A(u2__abc_52138_new_n3070_), .Y(u2__abc_52138_new_n3071_));
INVX1 INVX1_227 ( .A(sqrto_0_), .Y(u2__abc_52138_new_n3072_));
INVX1 INVX1_228 ( .A(sqrto_1_), .Y(u2__abc_52138_new_n3074_));
INVX1 INVX1_229 ( .A(sqrto_3_), .Y(u2__abc_52138_new_n3079_));
INVX1 INVX1_23 ( .A(sqrto_97_), .Y(_abc_65734_new_n893_));
INVX1 INVX1_230 ( .A(u2_remHi_3_), .Y(u2__abc_52138_new_n3081_));
INVX1 INVX1_231 ( .A(u2__abc_52138_new_n3082_), .Y(u2__abc_52138_new_n3083_));
INVX1 INVX1_232 ( .A(u2__abc_52138_new_n3063_), .Y(u2__abc_52138_new_n3084_));
INVX1 INVX1_233 ( .A(u2_remHi_4_), .Y(u2__abc_52138_new_n3086_));
INVX1 INVX1_234 ( .A(u2__abc_52138_new_n3087_), .Y(u2__abc_52138_new_n3088_));
INVX1 INVX1_235 ( .A(u2__abc_52138_new_n3055_), .Y(u2__abc_52138_new_n3089_));
INVX1 INVX1_236 ( .A(u2__abc_52138_new_n3043_), .Y(u2__abc_52138_new_n3093_));
INVX1 INVX1_237 ( .A(u2__abc_52138_new_n3048_), .Y(u2__abc_52138_new_n3094_));
INVX1 INVX1_238 ( .A(sqrto_8_), .Y(u2__abc_52138_new_n3096_));
INVX1 INVX1_239 ( .A(u2_remHi_12_), .Y(u2__abc_52138_new_n3101_));
INVX1 INVX1_24 ( .A(sqrto_98_), .Y(_abc_65734_new_n896_));
INVX1 INVX1_240 ( .A(u2__abc_52138_new_n3102_), .Y(u2__abc_52138_new_n3103_));
INVX1 INVX1_241 ( .A(u2__abc_52138_new_n3018_), .Y(u2__abc_52138_new_n3104_));
INVX1 INVX1_242 ( .A(u2__abc_52138_new_n3025_), .Y(u2__abc_52138_new_n3106_));
INVX1 INVX1_243 ( .A(u2__abc_52138_new_n3030_), .Y(u2__abc_52138_new_n3107_));
INVX1 INVX1_244 ( .A(sqrto_24_), .Y(u2__abc_52138_new_n3112_));
INVX1 INVX1_245 ( .A(u2_remHi_24_), .Y(u2__abc_52138_new_n3114_));
INVX1 INVX1_246 ( .A(sqrto_25_), .Y(u2__abc_52138_new_n3117_));
INVX1 INVX1_247 ( .A(u2_remHi_25_), .Y(u2__abc_52138_new_n3119_));
INVX1 INVX1_248 ( .A(sqrto_23_), .Y(u2__abc_52138_new_n3123_));
INVX1 INVX1_249 ( .A(u2_remHi_23_), .Y(u2__abc_52138_new_n3125_));
INVX1 INVX1_25 ( .A(sqrto_99_), .Y(_abc_65734_new_n899_));
INVX1 INVX1_250 ( .A(sqrto_22_), .Y(u2__abc_52138_new_n3128_));
INVX1 INVX1_251 ( .A(u2_remHi_22_), .Y(u2__abc_52138_new_n3130_));
INVX1 INVX1_252 ( .A(sqrto_28_), .Y(u2__abc_52138_new_n3135_));
INVX1 INVX1_253 ( .A(u2_remHi_28_), .Y(u2__abc_52138_new_n3137_));
INVX1 INVX1_254 ( .A(u2_remHi_29_), .Y(u2__abc_52138_new_n3140_));
INVX1 INVX1_255 ( .A(sqrto_29_), .Y(u2__abc_52138_new_n3142_));
INVX1 INVX1_256 ( .A(sqrto_27_), .Y(u2__abc_52138_new_n3146_));
INVX1 INVX1_257 ( .A(u2_remHi_27_), .Y(u2__abc_52138_new_n3148_));
INVX1 INVX1_258 ( .A(sqrto_26_), .Y(u2__abc_52138_new_n3151_));
INVX1 INVX1_259 ( .A(u2_remHi_26_), .Y(u2__abc_52138_new_n3153_));
INVX1 INVX1_26 ( .A(sqrto_100_), .Y(_abc_65734_new_n902_));
INVX1 INVX1_260 ( .A(sqrto_16_), .Y(u2__abc_52138_new_n3159_));
INVX1 INVX1_261 ( .A(u2_remHi_16_), .Y(u2__abc_52138_new_n3161_));
INVX1 INVX1_262 ( .A(sqrto_17_), .Y(u2__abc_52138_new_n3164_));
INVX1 INVX1_263 ( .A(u2_remHi_17_), .Y(u2__abc_52138_new_n3166_));
INVX1 INVX1_264 ( .A(sqrto_14_), .Y(u2__abc_52138_new_n3170_));
INVX1 INVX1_265 ( .A(u2_remHi_14_), .Y(u2__abc_52138_new_n3172_));
INVX1 INVX1_266 ( .A(sqrto_15_), .Y(u2__abc_52138_new_n3175_));
INVX1 INVX1_267 ( .A(u2_remHi_15_), .Y(u2__abc_52138_new_n3177_));
INVX1 INVX1_268 ( .A(sqrto_21_), .Y(u2__abc_52138_new_n3183_));
INVX1 INVX1_269 ( .A(u2_remHi_21_), .Y(u2__abc_52138_new_n3185_));
INVX1 INVX1_27 ( .A(sqrto_101_), .Y(_abc_65734_new_n905_));
INVX1 INVX1_270 ( .A(sqrto_18_), .Y(u2__abc_52138_new_n3189_));
INVX1 INVX1_271 ( .A(u2_remHi_18_), .Y(u2__abc_52138_new_n3191_));
INVX1 INVX1_272 ( .A(u2__abc_52138_new_n3173_), .Y(u2__abc_52138_new_n3199_));
INVX1 INVX1_273 ( .A(u2__abc_52138_new_n3178_), .Y(u2__abc_52138_new_n3200_));
INVX1 INVX1_274 ( .A(u2__abc_52138_new_n3162_), .Y(u2__abc_52138_new_n3202_));
INVX1 INVX1_275 ( .A(u2__abc_52138_new_n3167_), .Y(u2__abc_52138_new_n3203_));
INVX1 INVX1_276 ( .A(sqrto_19_), .Y(u2__abc_52138_new_n3206_));
INVX1 INVX1_277 ( .A(u2__abc_52138_new_n3192_), .Y(u2__abc_52138_new_n3209_));
INVX1 INVX1_278 ( .A(u2_remHi_20_), .Y(u2__abc_52138_new_n3211_));
INVX1 INVX1_279 ( .A(u2__abc_52138_new_n3214_), .Y(u2__abc_52138_new_n3215_));
INVX1 INVX1_28 ( .A(sqrto_102_), .Y(_abc_65734_new_n908_));
INVX1 INVX1_280 ( .A(u2__abc_52138_new_n3126_), .Y(u2__abc_52138_new_n3222_));
INVX1 INVX1_281 ( .A(u2__abc_52138_new_n3131_), .Y(u2__abc_52138_new_n3223_));
INVX1 INVX1_282 ( .A(u2__abc_52138_new_n3226_), .Y(u2__abc_52138_new_n3227_));
INVX1 INVX1_283 ( .A(u2__abc_52138_new_n3138_), .Y(u2__abc_52138_new_n3230_));
INVX1 INVX1_284 ( .A(u2__abc_52138_new_n3149_), .Y(u2__abc_52138_new_n3233_));
INVX1 INVX1_285 ( .A(u2__abc_52138_new_n3154_), .Y(u2__abc_52138_new_n3234_));
INVX1 INVX1_286 ( .A(sqrto_56_), .Y(u2__abc_52138_new_n3240_));
INVX1 INVX1_287 ( .A(u2_remHi_56_), .Y(u2__abc_52138_new_n3242_));
INVX1 INVX1_288 ( .A(sqrto_57_), .Y(u2__abc_52138_new_n3245_));
INVX1 INVX1_289 ( .A(u2_remHi_57_), .Y(u2__abc_52138_new_n3247_));
INVX1 INVX1_29 ( .A(sqrto_103_), .Y(_abc_65734_new_n911_));
INVX1 INVX1_290 ( .A(sqrto_54_), .Y(u2__abc_52138_new_n3251_));
INVX1 INVX1_291 ( .A(u2_remHi_54_), .Y(u2__abc_52138_new_n3253_));
INVX1 INVX1_292 ( .A(sqrto_55_), .Y(u2__abc_52138_new_n3256_));
INVX1 INVX1_293 ( .A(u2_remHi_55_), .Y(u2__abc_52138_new_n3258_));
INVX1 INVX1_294 ( .A(sqrto_60_), .Y(u2__abc_52138_new_n3263_));
INVX1 INVX1_295 ( .A(u2_remHi_60_), .Y(u2__abc_52138_new_n3265_));
INVX1 INVX1_296 ( .A(u2_remHi_61_), .Y(u2__abc_52138_new_n3268_));
INVX1 INVX1_297 ( .A(sqrto_61_), .Y(u2__abc_52138_new_n3270_));
INVX1 INVX1_298 ( .A(sqrto_59_), .Y(u2__abc_52138_new_n3274_));
INVX1 INVX1_299 ( .A(u2_remHi_59_), .Y(u2__abc_52138_new_n3276_));
INVX1 INVX1_3 ( .A(sqrto_77_), .Y(_abc_65734_new_n833_));
INVX1 INVX1_30 ( .A(sqrto_104_), .Y(_abc_65734_new_n914_));
INVX1 INVX1_300 ( .A(sqrto_58_), .Y(u2__abc_52138_new_n3279_));
INVX1 INVX1_301 ( .A(u2_remHi_58_), .Y(u2__abc_52138_new_n3281_));
INVX1 INVX1_302 ( .A(u2_remHi_48_), .Y(u2__abc_52138_new_n3287_));
INVX1 INVX1_303 ( .A(sqrto_48_), .Y(u2__abc_52138_new_n3289_));
INVX1 INVX1_304 ( .A(u2_remHi_49_), .Y(u2__abc_52138_new_n3292_));
INVX1 INVX1_305 ( .A(sqrto_49_), .Y(u2__abc_52138_new_n3294_));
INVX1 INVX1_306 ( .A(u2_remHi_47_), .Y(u2__abc_52138_new_n3298_));
INVX1 INVX1_307 ( .A(sqrto_47_), .Y(u2__abc_52138_new_n3300_));
INVX1 INVX1_308 ( .A(sqrto_46_), .Y(u2__abc_52138_new_n3303_));
INVX1 INVX1_309 ( .A(u2_remHi_46_), .Y(u2__abc_52138_new_n3305_));
INVX1 INVX1_31 ( .A(sqrto_105_), .Y(_abc_65734_new_n917_));
INVX1 INVX1_310 ( .A(u2__abc_52138_new_n3307_), .Y(u2__abc_52138_new_n3308_));
INVX1 INVX1_311 ( .A(sqrto_52_), .Y(u2__abc_52138_new_n3311_));
INVX1 INVX1_312 ( .A(u2_remHi_52_), .Y(u2__abc_52138_new_n3313_));
INVX1 INVX1_313 ( .A(sqrto_53_), .Y(u2__abc_52138_new_n3316_));
INVX1 INVX1_314 ( .A(u2_remHi_53_), .Y(u2__abc_52138_new_n3318_));
INVX1 INVX1_315 ( .A(sqrto_51_), .Y(u2__abc_52138_new_n3322_));
INVX1 INVX1_316 ( .A(u2_remHi_51_), .Y(u2__abc_52138_new_n3324_));
INVX1 INVX1_317 ( .A(sqrto_50_), .Y(u2__abc_52138_new_n3327_));
INVX1 INVX1_318 ( .A(u2_remHi_50_), .Y(u2__abc_52138_new_n3329_));
INVX1 INVX1_319 ( .A(sqrto_40_), .Y(u2__abc_52138_new_n3335_));
INVX1 INVX1_32 ( .A(sqrto_106_), .Y(_abc_65734_new_n920_));
INVX1 INVX1_320 ( .A(u2_remHi_40_), .Y(u2__abc_52138_new_n3337_));
INVX1 INVX1_321 ( .A(sqrto_41_), .Y(u2__abc_52138_new_n3340_));
INVX1 INVX1_322 ( .A(u2_remHi_41_), .Y(u2__abc_52138_new_n3342_));
INVX1 INVX1_323 ( .A(sqrto_38_), .Y(u2__abc_52138_new_n3346_));
INVX1 INVX1_324 ( .A(u2_remHi_38_), .Y(u2__abc_52138_new_n3348_));
INVX1 INVX1_325 ( .A(sqrto_39_), .Y(u2__abc_52138_new_n3351_));
INVX1 INVX1_326 ( .A(u2_remHi_39_), .Y(u2__abc_52138_new_n3353_));
INVX1 INVX1_327 ( .A(sqrto_44_), .Y(u2__abc_52138_new_n3358_));
INVX1 INVX1_328 ( .A(u2_remHi_44_), .Y(u2__abc_52138_new_n3360_));
INVX1 INVX1_329 ( .A(sqrto_45_), .Y(u2__abc_52138_new_n3363_));
INVX1 INVX1_33 ( .A(sqrto_107_), .Y(_abc_65734_new_n923_));
INVX1 INVX1_330 ( .A(u2_remHi_45_), .Y(u2__abc_52138_new_n3365_));
INVX1 INVX1_331 ( .A(sqrto_43_), .Y(u2__abc_52138_new_n3369_));
INVX1 INVX1_332 ( .A(u2_remHi_43_), .Y(u2__abc_52138_new_n3371_));
INVX1 INVX1_333 ( .A(sqrto_42_), .Y(u2__abc_52138_new_n3374_));
INVX1 INVX1_334 ( .A(u2_remHi_42_), .Y(u2__abc_52138_new_n3376_));
INVX1 INVX1_335 ( .A(sqrto_33_), .Y(u2__abc_52138_new_n3383_));
INVX1 INVX1_336 ( .A(u2_remHi_33_), .Y(u2__abc_52138_new_n3385_));
INVX1 INVX1_337 ( .A(sqrto_30_), .Y(u2__abc_52138_new_n3389_));
INVX1 INVX1_338 ( .A(u2_remHi_30_), .Y(u2__abc_52138_new_n3391_));
INVX1 INVX1_339 ( .A(sqrto_31_), .Y(u2__abc_52138_new_n3394_));
INVX1 INVX1_34 ( .A(sqrto_108_), .Y(_abc_65734_new_n926_));
INVX1 INVX1_340 ( .A(u2_remHi_31_), .Y(u2__abc_52138_new_n3396_));
INVX1 INVX1_341 ( .A(sqrto_36_), .Y(u2__abc_52138_new_n3401_));
INVX1 INVX1_342 ( .A(u2_remHi_36_), .Y(u2__abc_52138_new_n3403_));
INVX1 INVX1_343 ( .A(sqrto_37_), .Y(u2__abc_52138_new_n3406_));
INVX1 INVX1_344 ( .A(u2_remHi_37_), .Y(u2__abc_52138_new_n3408_));
INVX1 INVX1_345 ( .A(sqrto_35_), .Y(u2__abc_52138_new_n3412_));
INVX1 INVX1_346 ( .A(u2_remHi_35_), .Y(u2__abc_52138_new_n3414_));
INVX1 INVX1_347 ( .A(u2__abc_52138_new_n3392_), .Y(u2__abc_52138_new_n3434_));
INVX1 INVX1_348 ( .A(u2__abc_52138_new_n3397_), .Y(u2__abc_52138_new_n3435_));
INVX1 INVX1_349 ( .A(sqrto_32_), .Y(u2__abc_52138_new_n3437_));
INVX1 INVX1_35 ( .A(sqrto_109_), .Y(_abc_65734_new_n929_));
INVX1 INVX1_350 ( .A(u2__abc_52138_new_n3386_), .Y(u2__abc_52138_new_n3439_));
INVX1 INVX1_351 ( .A(u2__abc_52138_new_n3415_), .Y(u2__abc_52138_new_n3442_));
INVX1 INVX1_352 ( .A(u2_remHi_34_), .Y(u2__abc_52138_new_n3443_));
INVX1 INVX1_353 ( .A(u2__abc_52138_new_n3444_), .Y(u2__abc_52138_new_n3445_));
INVX1 INVX1_354 ( .A(u2__abc_52138_new_n3404_), .Y(u2__abc_52138_new_n3447_));
INVX1 INVX1_355 ( .A(u2__abc_52138_new_n3409_), .Y(u2__abc_52138_new_n3448_));
INVX1 INVX1_356 ( .A(u2__abc_52138_new_n3349_), .Y(u2__abc_52138_new_n3453_));
INVX1 INVX1_357 ( .A(u2__abc_52138_new_n3354_), .Y(u2__abc_52138_new_n3454_));
INVX1 INVX1_358 ( .A(u2__abc_52138_new_n3457_), .Y(u2__abc_52138_new_n3458_));
INVX1 INVX1_359 ( .A(u2__abc_52138_new_n3370_), .Y(u2__abc_52138_new_n3460_));
INVX1 INVX1_36 ( .A(sqrto_110_), .Y(_abc_65734_new_n932_));
INVX1 INVX1_360 ( .A(u2__abc_52138_new_n3364_), .Y(u2__abc_52138_new_n3463_));
INVX1 INVX1_361 ( .A(u2__abc_52138_new_n3464_), .Y(u2__abc_52138_new_n3465_));
INVX1 INVX1_362 ( .A(u2__abc_52138_new_n3299_), .Y(u2__abc_52138_new_n3469_));
INVX1 INVX1_363 ( .A(u2__abc_52138_new_n3306_), .Y(u2__abc_52138_new_n3470_));
INVX1 INVX1_364 ( .A(u2__abc_52138_new_n3474_), .Y(u2__abc_52138_new_n3475_));
INVX1 INVX1_365 ( .A(u2__abc_52138_new_n3479_), .Y(u2__abc_52138_new_n3480_));
INVX1 INVX1_366 ( .A(u2__abc_52138_new_n3314_), .Y(u2__abc_52138_new_n3481_));
INVX1 INVX1_367 ( .A(u2__abc_52138_new_n3319_), .Y(u2__abc_52138_new_n3482_));
INVX1 INVX1_368 ( .A(u2__abc_52138_new_n3285_), .Y(u2__abc_52138_new_n3486_));
INVX1 INVX1_369 ( .A(u2__abc_52138_new_n3254_), .Y(u2__abc_52138_new_n3488_));
INVX1 INVX1_37 ( .A(sqrto_111_), .Y(_abc_65734_new_n935_));
INVX1 INVX1_370 ( .A(u2__abc_52138_new_n3259_), .Y(u2__abc_52138_new_n3489_));
INVX1 INVX1_371 ( .A(u2__abc_52138_new_n3491_), .Y(u2__abc_52138_new_n3492_));
INVX1 INVX1_372 ( .A(u2__abc_52138_new_n3275_), .Y(u2__abc_52138_new_n3494_));
INVX1 INVX1_373 ( .A(u2_remHi_118_), .Y(u2__abc_52138_new_n3503_));
INVX1 INVX1_374 ( .A(u2__abc_52138_new_n3504_), .Y(u2__abc_52138_new_n3505_));
INVX1 INVX1_375 ( .A(u2_remHi_119_), .Y(u2__abc_52138_new_n3508_));
INVX1 INVX1_376 ( .A(u2__abc_52138_new_n3509_), .Y(u2__abc_52138_new_n3510_));
INVX1 INVX1_377 ( .A(sqrto_119_), .Y(u2__abc_52138_new_n3511_));
INVX1 INVX1_378 ( .A(u2__abc_52138_new_n3512_), .Y(u2__abc_52138_new_n3513_));
INVX1 INVX1_379 ( .A(sqrto_120_), .Y(u2__abc_52138_new_n3516_));
INVX1 INVX1_38 ( .A(sqrto_112_), .Y(_abc_65734_new_n938_));
INVX1 INVX1_380 ( .A(u2_remHi_120_), .Y(u2__abc_52138_new_n3518_));
INVX1 INVX1_381 ( .A(sqrto_121_), .Y(u2__abc_52138_new_n3521_));
INVX1 INVX1_382 ( .A(u2_remHi_121_), .Y(u2__abc_52138_new_n3523_));
INVX1 INVX1_383 ( .A(sqrto_124_), .Y(u2__abc_52138_new_n3527_));
INVX1 INVX1_384 ( .A(u2_remHi_124_), .Y(u2__abc_52138_new_n3529_));
INVX1 INVX1_385 ( .A(u2_remHi_125_), .Y(u2__abc_52138_new_n3532_));
INVX1 INVX1_386 ( .A(sqrto_125_), .Y(u2__abc_52138_new_n3534_));
INVX1 INVX1_387 ( .A(sqrto_123_), .Y(u2__abc_52138_new_n3538_));
INVX1 INVX1_388 ( .A(u2_remHi_123_), .Y(u2__abc_52138_new_n3540_));
INVX1 INVX1_389 ( .A(u2_remHi_122_), .Y(u2__abc_52138_new_n3542_));
INVX1 INVX1_39 ( .A(sqrto_113_), .Y(_abc_65734_new_n941_));
INVX1 INVX1_390 ( .A(sqrto_122_), .Y(u2__abc_52138_new_n3544_));
INVX1 INVX1_391 ( .A(sqrto_110_), .Y(u2__abc_52138_new_n3550_));
INVX1 INVX1_392 ( .A(u2_remHi_110_), .Y(u2__abc_52138_new_n3552_));
INVX1 INVX1_393 ( .A(sqrto_111_), .Y(u2__abc_52138_new_n3555_));
INVX1 INVX1_394 ( .A(u2_remHi_111_), .Y(u2__abc_52138_new_n3557_));
INVX1 INVX1_395 ( .A(sqrto_112_), .Y(u2__abc_52138_new_n3561_));
INVX1 INVX1_396 ( .A(u2_remHi_112_), .Y(u2__abc_52138_new_n3563_));
INVX1 INVX1_397 ( .A(sqrto_113_), .Y(u2__abc_52138_new_n3566_));
INVX1 INVX1_398 ( .A(u2_remHi_113_), .Y(u2__abc_52138_new_n3568_));
INVX1 INVX1_399 ( .A(u2_remHi_116_), .Y(u2__abc_52138_new_n3573_));
INVX1 INVX1_4 ( .A(sqrto_78_), .Y(_abc_65734_new_n836_));
INVX1 INVX1_40 ( .A(sqrto_114_), .Y(_abc_65734_new_n944_));
INVX1 INVX1_400 ( .A(sqrto_116_), .Y(u2__abc_52138_new_n3575_));
INVX1 INVX1_401 ( .A(sqrto_117_), .Y(u2__abc_52138_new_n3578_));
INVX1 INVX1_402 ( .A(u2_remHi_117_), .Y(u2__abc_52138_new_n3580_));
INVX1 INVX1_403 ( .A(sqrto_115_), .Y(u2__abc_52138_new_n3583_));
INVX1 INVX1_404 ( .A(u2_remHi_115_), .Y(u2__abc_52138_new_n3585_));
INVX1 INVX1_405 ( .A(sqrto_114_), .Y(u2__abc_52138_new_n3588_));
INVX1 INVX1_406 ( .A(u2_remHi_114_), .Y(u2__abc_52138_new_n3590_));
INVX1 INVX1_407 ( .A(sqrto_104_), .Y(u2__abc_52138_new_n3597_));
INVX1 INVX1_408 ( .A(u2_remHi_104_), .Y(u2__abc_52138_new_n3599_));
INVX1 INVX1_409 ( .A(sqrto_105_), .Y(u2__abc_52138_new_n3602_));
INVX1 INVX1_41 ( .A(sqrto_115_), .Y(_abc_65734_new_n947_));
INVX1 INVX1_410 ( .A(u2_remHi_105_), .Y(u2__abc_52138_new_n3604_));
INVX1 INVX1_411 ( .A(sqrto_103_), .Y(u2__abc_52138_new_n3608_));
INVX1 INVX1_412 ( .A(u2_remHi_103_), .Y(u2__abc_52138_new_n3610_));
INVX1 INVX1_413 ( .A(u2_remHi_102_), .Y(u2__abc_52138_new_n3612_));
INVX1 INVX1_414 ( .A(sqrto_102_), .Y(u2__abc_52138_new_n3614_));
INVX1 INVX1_415 ( .A(sqrto_108_), .Y(u2__abc_52138_new_n3619_));
INVX1 INVX1_416 ( .A(u2_remHi_108_), .Y(u2__abc_52138_new_n3621_));
INVX1 INVX1_417 ( .A(sqrto_109_), .Y(u2__abc_52138_new_n3624_));
INVX1 INVX1_418 ( .A(u2_remHi_109_), .Y(u2__abc_52138_new_n3626_));
INVX1 INVX1_419 ( .A(sqrto_107_), .Y(u2__abc_52138_new_n3630_));
INVX1 INVX1_42 ( .A(sqrto_116_), .Y(_abc_65734_new_n950_));
INVX1 INVX1_420 ( .A(u2_remHi_107_), .Y(u2__abc_52138_new_n3632_));
INVX1 INVX1_421 ( .A(u2_remHi_106_), .Y(u2__abc_52138_new_n3634_));
INVX1 INVX1_422 ( .A(sqrto_106_), .Y(u2__abc_52138_new_n3636_));
INVX1 INVX1_423 ( .A(u2_remHi_96_), .Y(u2__abc_52138_new_n3642_));
INVX1 INVX1_424 ( .A(sqrto_96_), .Y(u2__abc_52138_new_n3644_));
INVX1 INVX1_425 ( .A(u2_remHi_97_), .Y(u2__abc_52138_new_n3647_));
INVX1 INVX1_426 ( .A(sqrto_97_), .Y(u2__abc_52138_new_n3649_));
INVX1 INVX1_427 ( .A(sqrto_95_), .Y(u2__abc_52138_new_n3653_));
INVX1 INVX1_428 ( .A(u2_remHi_95_), .Y(u2__abc_52138_new_n3655_));
INVX1 INVX1_429 ( .A(sqrto_94_), .Y(u2__abc_52138_new_n3658_));
INVX1 INVX1_43 ( .A(sqrto_117_), .Y(_abc_65734_new_n953_));
INVX1 INVX1_430 ( .A(u2_remHi_94_), .Y(u2__abc_52138_new_n3660_));
INVX1 INVX1_431 ( .A(sqrto_100_), .Y(u2__abc_52138_new_n3665_));
INVX1 INVX1_432 ( .A(u2_remHi_100_), .Y(u2__abc_52138_new_n3667_));
INVX1 INVX1_433 ( .A(sqrto_101_), .Y(u2__abc_52138_new_n3670_));
INVX1 INVX1_434 ( .A(u2_remHi_101_), .Y(u2__abc_52138_new_n3672_));
INVX1 INVX1_435 ( .A(sqrto_99_), .Y(u2__abc_52138_new_n3676_));
INVX1 INVX1_436 ( .A(u2_remHi_99_), .Y(u2__abc_52138_new_n3678_));
INVX1 INVX1_437 ( .A(sqrto_98_), .Y(u2__abc_52138_new_n3681_));
INVX1 INVX1_438 ( .A(u2_remHi_98_), .Y(u2__abc_52138_new_n3683_));
INVX1 INVX1_439 ( .A(sqrto_92_), .Y(u2__abc_52138_new_n3691_));
INVX1 INVX1_44 ( .A(sqrto_118_), .Y(_abc_65734_new_n956_));
INVX1 INVX1_440 ( .A(u2_remHi_92_), .Y(u2__abc_52138_new_n3693_));
INVX1 INVX1_441 ( .A(sqrto_93_), .Y(u2__abc_52138_new_n3696_));
INVX1 INVX1_442 ( .A(u2_remHi_93_), .Y(u2__abc_52138_new_n3698_));
INVX1 INVX1_443 ( .A(sqrto_91_), .Y(u2__abc_52138_new_n3702_));
INVX1 INVX1_444 ( .A(u2_remHi_91_), .Y(u2__abc_52138_new_n3704_));
INVX1 INVX1_445 ( .A(u2_remHi_90_), .Y(u2__abc_52138_new_n3706_));
INVX1 INVX1_446 ( .A(sqrto_90_), .Y(u2__abc_52138_new_n3708_));
INVX1 INVX1_447 ( .A(sqrto_88_), .Y(u2__abc_52138_new_n3713_));
INVX1 INVX1_448 ( .A(u2_remHi_88_), .Y(u2__abc_52138_new_n3715_));
INVX1 INVX1_449 ( .A(sqrto_89_), .Y(u2__abc_52138_new_n3718_));
INVX1 INVX1_45 ( .A(sqrto_119_), .Y(_abc_65734_new_n959_));
INVX1 INVX1_450 ( .A(u2_remHi_89_), .Y(u2__abc_52138_new_n3720_));
INVX1 INVX1_451 ( .A(u2_remHi_87_), .Y(u2__abc_52138_new_n3724_));
INVX1 INVX1_452 ( .A(u2__abc_52138_new_n3725_), .Y(u2__abc_52138_new_n3726_));
INVX1 INVX1_453 ( .A(sqrto_87_), .Y(u2__abc_52138_new_n3727_));
INVX1 INVX1_454 ( .A(u2__abc_52138_new_n3728_), .Y(u2__abc_52138_new_n3729_));
INVX1 INVX1_455 ( .A(u2_remHi_86_), .Y(u2__abc_52138_new_n3730_));
INVX1 INVX1_456 ( .A(sqrto_86_), .Y(u2__abc_52138_new_n3732_));
INVX1 INVX1_457 ( .A(sqrto_78_), .Y(u2__abc_52138_new_n3738_));
INVX1 INVX1_458 ( .A(u2_remHi_78_), .Y(u2__abc_52138_new_n3740_));
INVX1 INVX1_459 ( .A(sqrto_79_), .Y(u2__abc_52138_new_n3743_));
INVX1 INVX1_46 ( .A(sqrto_120_), .Y(_abc_65734_new_n962_));
INVX1 INVX1_460 ( .A(u2_remHi_79_), .Y(u2__abc_52138_new_n3745_));
INVX1 INVX1_461 ( .A(sqrto_80_), .Y(u2__abc_52138_new_n3749_));
INVX1 INVX1_462 ( .A(u2_remHi_80_), .Y(u2__abc_52138_new_n3751_));
INVX1 INVX1_463 ( .A(sqrto_81_), .Y(u2__abc_52138_new_n3754_));
INVX1 INVX1_464 ( .A(u2_remHi_81_), .Y(u2__abc_52138_new_n3756_));
INVX1 INVX1_465 ( .A(sqrto_84_), .Y(u2__abc_52138_new_n3761_));
INVX1 INVX1_466 ( .A(u2_remHi_84_), .Y(u2__abc_52138_new_n3763_));
INVX1 INVX1_467 ( .A(sqrto_85_), .Y(u2__abc_52138_new_n3766_));
INVX1 INVX1_468 ( .A(u2_remHi_85_), .Y(u2__abc_52138_new_n3768_));
INVX1 INVX1_469 ( .A(sqrto_83_), .Y(u2__abc_52138_new_n3772_));
INVX1 INVX1_47 ( .A(sqrto_121_), .Y(_abc_65734_new_n965_));
INVX1 INVX1_470 ( .A(u2_remHi_83_), .Y(u2__abc_52138_new_n3774_));
INVX1 INVX1_471 ( .A(sqrto_82_), .Y(u2__abc_52138_new_n3777_));
INVX1 INVX1_472 ( .A(u2_remHi_82_), .Y(u2__abc_52138_new_n3779_));
INVX1 INVX1_473 ( .A(u2_remHi_70_), .Y(u2__abc_52138_new_n3786_));
INVX1 INVX1_474 ( .A(sqrto_70_), .Y(u2__abc_52138_new_n3788_));
INVX1 INVX1_475 ( .A(u2_remHi_71_), .Y(u2__abc_52138_new_n3791_));
INVX1 INVX1_476 ( .A(sqrto_71_), .Y(u2__abc_52138_new_n3793_));
INVX1 INVX1_477 ( .A(sqrto_72_), .Y(u2__abc_52138_new_n3797_));
INVX1 INVX1_478 ( .A(u2_remHi_72_), .Y(u2__abc_52138_new_n3799_));
INVX1 INVX1_479 ( .A(sqrto_73_), .Y(u2__abc_52138_new_n3802_));
INVX1 INVX1_48 ( .A(sqrto_122_), .Y(_abc_65734_new_n968_));
INVX1 INVX1_480 ( .A(u2_remHi_73_), .Y(u2__abc_52138_new_n3804_));
INVX1 INVX1_481 ( .A(u2_remHi_76_), .Y(u2__abc_52138_new_n3808_));
INVX1 INVX1_482 ( .A(sqrto_76_), .Y(u2__abc_52138_new_n3810_));
INVX1 INVX1_483 ( .A(u2_remHi_77_), .Y(u2__abc_52138_new_n3813_));
INVX1 INVX1_484 ( .A(sqrto_77_), .Y(u2__abc_52138_new_n3815_));
INVX1 INVX1_485 ( .A(u2_remHi_75_), .Y(u2__abc_52138_new_n3819_));
INVX1 INVX1_486 ( .A(sqrto_75_), .Y(u2__abc_52138_new_n3821_));
INVX1 INVX1_487 ( .A(u2_remHi_74_), .Y(u2__abc_52138_new_n3824_));
INVX1 INVX1_488 ( .A(sqrto_74_), .Y(u2__abc_52138_new_n3826_));
INVX1 INVX1_489 ( .A(sqrto_62_), .Y(u2__abc_52138_new_n3832_));
INVX1 INVX1_49 ( .A(sqrto_123_), .Y(_abc_65734_new_n971_));
INVX1 INVX1_490 ( .A(u2_remHi_62_), .Y(u2__abc_52138_new_n3834_));
INVX1 INVX1_491 ( .A(sqrto_63_), .Y(u2__abc_52138_new_n3837_));
INVX1 INVX1_492 ( .A(u2_remHi_63_), .Y(u2__abc_52138_new_n3839_));
INVX1 INVX1_493 ( .A(sqrto_64_), .Y(u2__abc_52138_new_n3843_));
INVX1 INVX1_494 ( .A(u2_remHi_64_), .Y(u2__abc_52138_new_n3845_));
INVX1 INVX1_495 ( .A(sqrto_65_), .Y(u2__abc_52138_new_n3848_));
INVX1 INVX1_496 ( .A(u2_remHi_65_), .Y(u2__abc_52138_new_n3850_));
INVX1 INVX1_497 ( .A(sqrto_69_), .Y(u2__abc_52138_new_n3856_));
INVX1 INVX1_498 ( .A(u2_remHi_69_), .Y(u2__abc_52138_new_n3858_));
INVX1 INVX1_499 ( .A(sqrto_66_), .Y(u2__abc_52138_new_n3862_));
INVX1 INVX1_5 ( .A(sqrto_79_), .Y(_abc_65734_new_n839_));
INVX1 INVX1_50 ( .A(sqrto_124_), .Y(_abc_65734_new_n974_));
INVX1 INVX1_500 ( .A(u2_remHi_66_), .Y(u2__abc_52138_new_n3864_));
INVX1 INVX1_501 ( .A(u2__abc_52138_new_n3835_), .Y(u2__abc_52138_new_n3874_));
INVX1 INVX1_502 ( .A(u2__abc_52138_new_n3840_), .Y(u2__abc_52138_new_n3875_));
INVX1 INVX1_503 ( .A(u2__abc_52138_new_n3846_), .Y(u2__abc_52138_new_n3877_));
INVX1 INVX1_504 ( .A(u2__abc_52138_new_n3851_), .Y(u2__abc_52138_new_n3878_));
INVX1 INVX1_505 ( .A(sqrto_67_), .Y(u2__abc_52138_new_n3881_));
INVX1 INVX1_506 ( .A(u2_remHi_67_), .Y(u2__abc_52138_new_n3883_));
INVX1 INVX1_507 ( .A(u2__abc_52138_new_n3884_), .Y(u2__abc_52138_new_n3885_));
INVX1 INVX1_508 ( .A(u2__abc_52138_new_n3865_), .Y(u2__abc_52138_new_n3886_));
INVX1 INVX1_509 ( .A(u2_remHi_68_), .Y(u2__abc_52138_new_n3888_));
INVX1 INVX1_51 ( .A(sqrto_125_), .Y(_abc_65734_new_n977_));
INVX1 INVX1_510 ( .A(u2__abc_52138_new_n3891_), .Y(u2__abc_52138_new_n3892_));
INVX1 INVX1_511 ( .A(u2__abc_52138_new_n3792_), .Y(u2__abc_52138_new_n3895_));
INVX1 INVX1_512 ( .A(u2__abc_52138_new_n3800_), .Y(u2__abc_52138_new_n3897_));
INVX1 INVX1_513 ( .A(u2__abc_52138_new_n3805_), .Y(u2__abc_52138_new_n3898_));
INVX1 INVX1_514 ( .A(u2__abc_52138_new_n3820_), .Y(u2__abc_52138_new_n3901_));
INVX1 INVX1_515 ( .A(u2__abc_52138_new_n3741_), .Y(u2__abc_52138_new_n3908_));
INVX1 INVX1_516 ( .A(u2__abc_52138_new_n3746_), .Y(u2__abc_52138_new_n3909_));
INVX1 INVX1_517 ( .A(u2__abc_52138_new_n3752_), .Y(u2__abc_52138_new_n3911_));
INVX1 INVX1_518 ( .A(u2__abc_52138_new_n3757_), .Y(u2__abc_52138_new_n3912_));
INVX1 INVX1_519 ( .A(u2__abc_52138_new_n3919_), .Y(u2__abc_52138_new_n3920_));
INVX1 INVX1_52 ( .A(sqrto_126_), .Y(_abc_65734_new_n980_));
INVX1 INVX1_520 ( .A(u2__abc_52138_new_n3925_), .Y(u2__abc_52138_new_n3926_));
INVX1 INVX1_521 ( .A(u2__abc_52138_new_n3697_), .Y(u2__abc_52138_new_n3932_));
INVX1 INVX1_522 ( .A(u2__abc_52138_new_n3933_), .Y(u2__abc_52138_new_n3934_));
INVX1 INVX1_523 ( .A(u2__abc_52138_new_n3656_), .Y(u2__abc_52138_new_n3939_));
INVX1 INVX1_524 ( .A(u2__abc_52138_new_n3661_), .Y(u2__abc_52138_new_n3940_));
INVX1 INVX1_525 ( .A(u2__abc_52138_new_n3944_), .Y(u2__abc_52138_new_n3945_));
INVX1 INVX1_526 ( .A(u2__abc_52138_new_n3679_), .Y(u2__abc_52138_new_n3948_));
INVX1 INVX1_527 ( .A(u2__abc_52138_new_n3684_), .Y(u2__abc_52138_new_n3949_));
INVX1 INVX1_528 ( .A(u2__abc_52138_new_n3603_), .Y(u2__abc_52138_new_n3958_));
INVX1 INVX1_529 ( .A(u2__abc_52138_new_n3959_), .Y(u2__abc_52138_new_n3960_));
INVX1 INVX1_53 ( .A(sqrto_127_), .Y(_abc_65734_new_n983_));
INVX1 INVX1_530 ( .A(u2__abc_52138_new_n3625_), .Y(u2__abc_52138_new_n3966_));
INVX1 INVX1_531 ( .A(u2__abc_52138_new_n3553_), .Y(u2__abc_52138_new_n3972_));
INVX1 INVX1_532 ( .A(u2__abc_52138_new_n3558_), .Y(u2__abc_52138_new_n3973_));
INVX1 INVX1_533 ( .A(u2__abc_52138_new_n3567_), .Y(u2__abc_52138_new_n3975_));
INVX1 INVX1_534 ( .A(u2__abc_52138_new_n3976_), .Y(u2__abc_52138_new_n3977_));
INVX1 INVX1_535 ( .A(u2__abc_52138_new_n3980_), .Y(u2__abc_52138_new_n3981_));
INVX1 INVX1_536 ( .A(u2__abc_52138_new_n3983_), .Y(u2__abc_52138_new_n3984_));
INVX1 INVX1_537 ( .A(u2__abc_52138_new_n3535_), .Y(u2__abc_52138_new_n3992_));
INVX1 INVX1_538 ( .A(u2__abc_52138_new_n3996_), .Y(u2__abc_52138_new_n3997_));
INVX1 INVX1_539 ( .A(u2_o_246_), .Y(u2__abc_52138_new_n4003_));
INVX1 INVX1_54 ( .A(sqrto_128_), .Y(_abc_65734_new_n986_));
INVX1 INVX1_540 ( .A(u2_remHi_246_), .Y(u2__abc_52138_new_n4005_));
INVX1 INVX1_541 ( .A(u2_o_247_), .Y(u2__abc_52138_new_n4008_));
INVX1 INVX1_542 ( .A(u2_remHi_247_), .Y(u2__abc_52138_new_n4010_));
INVX1 INVX1_543 ( .A(u2_o_248_), .Y(u2__abc_52138_new_n4014_));
INVX1 INVX1_544 ( .A(u2_remHi_248_), .Y(u2__abc_52138_new_n4016_));
INVX1 INVX1_545 ( .A(u2_o_249_), .Y(u2__abc_52138_new_n4019_));
INVX1 INVX1_546 ( .A(u2_remHi_249_), .Y(u2__abc_52138_new_n4021_));
INVX1 INVX1_547 ( .A(u2_o_252_), .Y(u2__abc_52138_new_n4026_));
INVX1 INVX1_548 ( .A(u2_remHi_252_), .Y(u2__abc_52138_new_n4028_));
INVX1 INVX1_549 ( .A(u2_remHi_253_), .Y(u2__abc_52138_new_n4031_));
INVX1 INVX1_55 ( .A(sqrto_129_), .Y(_abc_65734_new_n989_));
INVX1 INVX1_550 ( .A(u2_o_253_), .Y(u2__abc_52138_new_n4033_));
INVX1 INVX1_551 ( .A(u2_o_251_), .Y(u2__abc_52138_new_n4037_));
INVX1 INVX1_552 ( .A(u2_remHi_251_), .Y(u2__abc_52138_new_n4039_));
INVX1 INVX1_553 ( .A(u2_o_250_), .Y(u2__abc_52138_new_n4042_));
INVX1 INVX1_554 ( .A(u2_remHi_250_), .Y(u2__abc_52138_new_n4044_));
INVX1 INVX1_555 ( .A(u2_o_238_), .Y(u2__abc_52138_new_n4050_));
INVX1 INVX1_556 ( .A(u2_remHi_238_), .Y(u2__abc_52138_new_n4052_));
INVX1 INVX1_557 ( .A(u2_o_239_), .Y(u2__abc_52138_new_n4055_));
INVX1 INVX1_558 ( .A(u2_remHi_239_), .Y(u2__abc_52138_new_n4057_));
INVX1 INVX1_559 ( .A(u2_o_240_), .Y(u2__abc_52138_new_n4061_));
INVX1 INVX1_56 ( .A(sqrto_130_), .Y(_abc_65734_new_n992_));
INVX1 INVX1_560 ( .A(u2_remHi_240_), .Y(u2__abc_52138_new_n4063_));
INVX1 INVX1_561 ( .A(u2_o_241_), .Y(u2__abc_52138_new_n4066_));
INVX1 INVX1_562 ( .A(u2_remHi_241_), .Y(u2__abc_52138_new_n4068_));
INVX1 INVX1_563 ( .A(u2__abc_52138_new_n4071_), .Y(u2__abc_52138_new_n4072_));
INVX1 INVX1_564 ( .A(u2_o_244_), .Y(u2__abc_52138_new_n4074_));
INVX1 INVX1_565 ( .A(u2_remHi_244_), .Y(u2__abc_52138_new_n4076_));
INVX1 INVX1_566 ( .A(u2_o_245_), .Y(u2__abc_52138_new_n4079_));
INVX1 INVX1_567 ( .A(u2_remHi_245_), .Y(u2__abc_52138_new_n4081_));
INVX1 INVX1_568 ( .A(u2_remHi_243_), .Y(u2__abc_52138_new_n4085_));
INVX1 INVX1_569 ( .A(u2_o_243_), .Y(u2__abc_52138_new_n4087_));
INVX1 INVX1_57 ( .A(sqrto_131_), .Y(_abc_65734_new_n995_));
INVX1 INVX1_570 ( .A(u2_o_242_), .Y(u2__abc_52138_new_n4090_));
INVX1 INVX1_571 ( .A(u2_remHi_242_), .Y(u2__abc_52138_new_n4092_));
INVX1 INVX1_572 ( .A(u2_o_236_), .Y(u2__abc_52138_new_n4099_));
INVX1 INVX1_573 ( .A(u2_remHi_236_), .Y(u2__abc_52138_new_n4101_));
INVX1 INVX1_574 ( .A(u2_o_237_), .Y(u2__abc_52138_new_n4104_));
INVX1 INVX1_575 ( .A(u2_remHi_237_), .Y(u2__abc_52138_new_n4106_));
INVX1 INVX1_576 ( .A(u2_o_235_), .Y(u2__abc_52138_new_n4110_));
INVX1 INVX1_577 ( .A(u2_remHi_235_), .Y(u2__abc_52138_new_n4112_));
INVX1 INVX1_578 ( .A(u2_o_234_), .Y(u2__abc_52138_new_n4115_));
INVX1 INVX1_579 ( .A(u2_remHi_234_), .Y(u2__abc_52138_new_n4117_));
INVX1 INVX1_58 ( .A(sqrto_132_), .Y(_abc_65734_new_n998_));
INVX1 INVX1_580 ( .A(u2__abc_52138_new_n4121_), .Y(u2__abc_52138_new_n4122_));
INVX1 INVX1_581 ( .A(u2_o_232_), .Y(u2__abc_52138_new_n4123_));
INVX1 INVX1_582 ( .A(u2_remHi_232_), .Y(u2__abc_52138_new_n4125_));
INVX1 INVX1_583 ( .A(u2_o_233_), .Y(u2__abc_52138_new_n4128_));
INVX1 INVX1_584 ( .A(u2_remHi_233_), .Y(u2__abc_52138_new_n4130_));
INVX1 INVX1_585 ( .A(u2_remHi_231_), .Y(u2__abc_52138_new_n4134_));
INVX1 INVX1_586 ( .A(u2__abc_52138_new_n4135_), .Y(u2__abc_52138_new_n4136_));
INVX1 INVX1_587 ( .A(u2_remHi_230_), .Y(u2__abc_52138_new_n4138_));
INVX1 INVX1_588 ( .A(u2_o_230_), .Y(u2__abc_52138_new_n4140_));
INVX1 INVX1_589 ( .A(sqrto_224_), .Y(u2__abc_52138_new_n4146_));
INVX1 INVX1_59 ( .A(sqrto_133_), .Y(_abc_65734_new_n1001_));
INVX1 INVX1_590 ( .A(u2_remHi_224_), .Y(u2__abc_52138_new_n4148_));
INVX1 INVX1_591 ( .A(sqrto_225_), .Y(u2__abc_52138_new_n4151_));
INVX1 INVX1_592 ( .A(u2_remHi_225_), .Y(u2__abc_52138_new_n4153_));
INVX1 INVX1_593 ( .A(sqrto_223_), .Y(u2__abc_52138_new_n4157_));
INVX1 INVX1_594 ( .A(u2_remHi_223_), .Y(u2__abc_52138_new_n4159_));
INVX1 INVX1_595 ( .A(sqrto_222_), .Y(u2__abc_52138_new_n4162_));
INVX1 INVX1_596 ( .A(u2_remHi_222_), .Y(u2__abc_52138_new_n4164_));
INVX1 INVX1_597 ( .A(u2_o_228_), .Y(u2__abc_52138_new_n4169_));
INVX1 INVX1_598 ( .A(u2_remHi_228_), .Y(u2__abc_52138_new_n4171_));
INVX1 INVX1_599 ( .A(u2_o_229_), .Y(u2__abc_52138_new_n4174_));
INVX1 INVX1_6 ( .A(sqrto_80_), .Y(_abc_65734_new_n842_));
INVX1 INVX1_60 ( .A(sqrto_134_), .Y(_abc_65734_new_n1004_));
INVX1 INVX1_600 ( .A(u2_remHi_229_), .Y(u2__abc_52138_new_n4176_));
INVX1 INVX1_601 ( .A(u2_remHi_227_), .Y(u2__abc_52138_new_n4180_));
INVX1 INVX1_602 ( .A(u2_o_227_), .Y(u2__abc_52138_new_n4182_));
INVX1 INVX1_603 ( .A(u2_remHi_226_), .Y(u2__abc_52138_new_n4185_));
INVX1 INVX1_604 ( .A(u2_o_226_), .Y(u2__abc_52138_new_n4187_));
INVX1 INVX1_605 ( .A(sqrto_216_), .Y(u2__abc_52138_new_n4194_));
INVX1 INVX1_606 ( .A(u2_remHi_216_), .Y(u2__abc_52138_new_n4196_));
INVX1 INVX1_607 ( .A(sqrto_217_), .Y(u2__abc_52138_new_n4199_));
INVX1 INVX1_608 ( .A(u2_remHi_217_), .Y(u2__abc_52138_new_n4201_));
INVX1 INVX1_609 ( .A(sqrto_214_), .Y(u2__abc_52138_new_n4205_));
INVX1 INVX1_61 ( .A(sqrto_135_), .Y(_abc_65734_new_n1007_));
INVX1 INVX1_610 ( .A(u2_remHi_214_), .Y(u2__abc_52138_new_n4207_));
INVX1 INVX1_611 ( .A(sqrto_215_), .Y(u2__abc_52138_new_n4210_));
INVX1 INVX1_612 ( .A(u2_remHi_215_), .Y(u2__abc_52138_new_n4212_));
INVX1 INVX1_613 ( .A(sqrto_220_), .Y(u2__abc_52138_new_n4217_));
INVX1 INVX1_614 ( .A(u2_remHi_220_), .Y(u2__abc_52138_new_n4219_));
INVX1 INVX1_615 ( .A(sqrto_221_), .Y(u2__abc_52138_new_n4222_));
INVX1 INVX1_616 ( .A(u2_remHi_221_), .Y(u2__abc_52138_new_n4224_));
INVX1 INVX1_617 ( .A(u2_remHi_219_), .Y(u2__abc_52138_new_n4228_));
INVX1 INVX1_618 ( .A(sqrto_219_), .Y(u2__abc_52138_new_n4230_));
INVX1 INVX1_619 ( .A(sqrto_218_), .Y(u2__abc_52138_new_n4233_));
INVX1 INVX1_62 ( .A(sqrto_136_), .Y(_abc_65734_new_n1010_));
INVX1 INVX1_620 ( .A(u2_remHi_218_), .Y(u2__abc_52138_new_n4235_));
INVX1 INVX1_621 ( .A(sqrto_208_), .Y(u2__abc_52138_new_n4241_));
INVX1 INVX1_622 ( .A(u2_remHi_208_), .Y(u2__abc_52138_new_n4243_));
INVX1 INVX1_623 ( .A(sqrto_209_), .Y(u2__abc_52138_new_n4246_));
INVX1 INVX1_624 ( .A(u2_remHi_209_), .Y(u2__abc_52138_new_n4248_));
INVX1 INVX1_625 ( .A(sqrto_206_), .Y(u2__abc_52138_new_n4252_));
INVX1 INVX1_626 ( .A(u2_remHi_206_), .Y(u2__abc_52138_new_n4254_));
INVX1 INVX1_627 ( .A(sqrto_207_), .Y(u2__abc_52138_new_n4257_));
INVX1 INVX1_628 ( .A(u2_remHi_207_), .Y(u2__abc_52138_new_n4259_));
INVX1 INVX1_629 ( .A(u2_remHi_212_), .Y(u2__abc_52138_new_n4264_));
INVX1 INVX1_63 ( .A(sqrto_137_), .Y(_abc_65734_new_n1013_));
INVX1 INVX1_630 ( .A(sqrto_212_), .Y(u2__abc_52138_new_n4266_));
INVX1 INVX1_631 ( .A(u2_remHi_213_), .Y(u2__abc_52138_new_n4269_));
INVX1 INVX1_632 ( .A(sqrto_213_), .Y(u2__abc_52138_new_n4271_));
INVX1 INVX1_633 ( .A(u2_remHi_211_), .Y(u2__abc_52138_new_n4275_));
INVX1 INVX1_634 ( .A(sqrto_211_), .Y(u2__abc_52138_new_n4277_));
INVX1 INVX1_635 ( .A(u2_remHi_210_), .Y(u2__abc_52138_new_n4280_));
INVX1 INVX1_636 ( .A(sqrto_210_), .Y(u2__abc_52138_new_n4282_));
INVX1 INVX1_637 ( .A(sqrto_200_), .Y(u2__abc_52138_new_n4289_));
INVX1 INVX1_638 ( .A(u2_remHi_200_), .Y(u2__abc_52138_new_n4291_));
INVX1 INVX1_639 ( .A(sqrto_201_), .Y(u2__abc_52138_new_n4294_));
INVX1 INVX1_64 ( .A(sqrto_138_), .Y(_abc_65734_new_n1016_));
INVX1 INVX1_640 ( .A(u2_remHi_201_), .Y(u2__abc_52138_new_n4296_));
INVX1 INVX1_641 ( .A(sqrto_199_), .Y(u2__abc_52138_new_n4300_));
INVX1 INVX1_642 ( .A(u2_remHi_199_), .Y(u2__abc_52138_new_n4302_));
INVX1 INVX1_643 ( .A(sqrto_198_), .Y(u2__abc_52138_new_n4305_));
INVX1 INVX1_644 ( .A(u2_remHi_198_), .Y(u2__abc_52138_new_n4307_));
INVX1 INVX1_645 ( .A(sqrto_204_), .Y(u2__abc_52138_new_n4312_));
INVX1 INVX1_646 ( .A(u2_remHi_204_), .Y(u2__abc_52138_new_n4314_));
INVX1 INVX1_647 ( .A(sqrto_205_), .Y(u2__abc_52138_new_n4317_));
INVX1 INVX1_648 ( .A(u2_remHi_205_), .Y(u2__abc_52138_new_n4319_));
INVX1 INVX1_649 ( .A(u2_remHi_203_), .Y(u2__abc_52138_new_n4323_));
INVX1 INVX1_65 ( .A(sqrto_139_), .Y(_abc_65734_new_n1019_));
INVX1 INVX1_650 ( .A(sqrto_203_), .Y(u2__abc_52138_new_n4325_));
INVX1 INVX1_651 ( .A(sqrto_196_), .Y(u2__abc_52138_new_n4331_));
INVX1 INVX1_652 ( .A(u2_remHi_196_), .Y(u2__abc_52138_new_n4333_));
INVX1 INVX1_653 ( .A(sqrto_197_), .Y(u2__abc_52138_new_n4336_));
INVX1 INVX1_654 ( .A(u2_remHi_197_), .Y(u2__abc_52138_new_n4338_));
INVX1 INVX1_655 ( .A(sqrto_195_), .Y(u2__abc_52138_new_n4342_));
INVX1 INVX1_656 ( .A(u2_remHi_195_), .Y(u2__abc_52138_new_n4344_));
INVX1 INVX1_657 ( .A(sqrto_194_), .Y(u2__abc_52138_new_n4347_));
INVX1 INVX1_658 ( .A(u2_remHi_194_), .Y(u2__abc_52138_new_n4349_));
INVX1 INVX1_659 ( .A(u2_remHi_192_), .Y(u2__abc_52138_new_n4354_));
INVX1 INVX1_66 ( .A(sqrto_140_), .Y(_abc_65734_new_n1022_));
INVX1 INVX1_660 ( .A(sqrto_192_), .Y(u2__abc_52138_new_n4356_));
INVX1 INVX1_661 ( .A(sqrto_193_), .Y(u2__abc_52138_new_n4358_));
INVX1 INVX1_662 ( .A(u2_remHi_193_), .Y(u2__abc_52138_new_n4360_));
INVX1 INVX1_663 ( .A(u2_remHi_190_), .Y(u2__abc_52138_new_n4364_));
INVX1 INVX1_664 ( .A(sqrto_190_), .Y(u2__abc_52138_new_n4366_));
INVX1 INVX1_665 ( .A(u2_remHi_191_), .Y(u2__abc_52138_new_n4369_));
INVX1 INVX1_666 ( .A(u2__abc_52138_new_n4370_), .Y(u2__abc_52138_new_n4371_));
INVX1 INVX1_667 ( .A(sqrto_191_), .Y(u2__abc_52138_new_n4372_));
INVX1 INVX1_668 ( .A(u2__abc_52138_new_n4373_), .Y(u2__abc_52138_new_n4374_));
INVX1 INVX1_669 ( .A(sqrto_182_), .Y(u2__abc_52138_new_n4382_));
INVX1 INVX1_67 ( .A(sqrto_141_), .Y(_abc_65734_new_n1025_));
INVX1 INVX1_670 ( .A(u2_remHi_182_), .Y(u2__abc_52138_new_n4384_));
INVX1 INVX1_671 ( .A(sqrto_183_), .Y(u2__abc_52138_new_n4387_));
INVX1 INVX1_672 ( .A(u2_remHi_183_), .Y(u2__abc_52138_new_n4389_));
INVX1 INVX1_673 ( .A(sqrto_184_), .Y(u2__abc_52138_new_n4393_));
INVX1 INVX1_674 ( .A(u2_remHi_184_), .Y(u2__abc_52138_new_n4395_));
INVX1 INVX1_675 ( .A(sqrto_185_), .Y(u2__abc_52138_new_n4398_));
INVX1 INVX1_676 ( .A(u2_remHi_185_), .Y(u2__abc_52138_new_n4400_));
INVX1 INVX1_677 ( .A(sqrto_188_), .Y(u2__abc_52138_new_n4405_));
INVX1 INVX1_678 ( .A(u2_remHi_188_), .Y(u2__abc_52138_new_n4407_));
INVX1 INVX1_679 ( .A(sqrto_189_), .Y(u2__abc_52138_new_n4410_));
INVX1 INVX1_68 ( .A(sqrto_142_), .Y(_abc_65734_new_n1028_));
INVX1 INVX1_680 ( .A(u2_remHi_189_), .Y(u2__abc_52138_new_n4412_));
INVX1 INVX1_681 ( .A(sqrto_187_), .Y(u2__abc_52138_new_n4416_));
INVX1 INVX1_682 ( .A(u2_remHi_187_), .Y(u2__abc_52138_new_n4418_));
INVX1 INVX1_683 ( .A(sqrto_186_), .Y(u2__abc_52138_new_n4421_));
INVX1 INVX1_684 ( .A(u2_remHi_186_), .Y(u2__abc_52138_new_n4423_));
INVX1 INVX1_685 ( .A(sqrto_180_), .Y(u2__abc_52138_new_n4429_));
INVX1 INVX1_686 ( .A(u2_remHi_180_), .Y(u2__abc_52138_new_n4431_));
INVX1 INVX1_687 ( .A(sqrto_181_), .Y(u2__abc_52138_new_n4434_));
INVX1 INVX1_688 ( .A(u2_remHi_181_), .Y(u2__abc_52138_new_n4436_));
INVX1 INVX1_689 ( .A(sqrto_179_), .Y(u2__abc_52138_new_n4440_));
INVX1 INVX1_69 ( .A(sqrto_143_), .Y(_abc_65734_new_n1031_));
INVX1 INVX1_690 ( .A(u2_remHi_179_), .Y(u2__abc_52138_new_n4442_));
INVX1 INVX1_691 ( .A(sqrto_178_), .Y(u2__abc_52138_new_n4445_));
INVX1 INVX1_692 ( .A(u2_remHi_178_), .Y(u2__abc_52138_new_n4447_));
INVX1 INVX1_693 ( .A(sqrto_176_), .Y(u2__abc_52138_new_n4452_));
INVX1 INVX1_694 ( .A(u2_remHi_176_), .Y(u2__abc_52138_new_n4454_));
INVX1 INVX1_695 ( .A(sqrto_177_), .Y(u2__abc_52138_new_n4457_));
INVX1 INVX1_696 ( .A(u2_remHi_177_), .Y(u2__abc_52138_new_n4459_));
INVX1 INVX1_697 ( .A(sqrto_174_), .Y(u2__abc_52138_new_n4463_));
INVX1 INVX1_698 ( .A(u2_remHi_174_), .Y(u2__abc_52138_new_n4465_));
INVX1 INVX1_699 ( .A(u2__abc_52138_new_n4467_), .Y(u2__abc_52138_new_n4468_));
INVX1 INVX1_7 ( .A(sqrto_81_), .Y(_abc_65734_new_n845_));
INVX1 INVX1_70 ( .A(sqrto_144_), .Y(_abc_65734_new_n1034_));
INVX1 INVX1_700 ( .A(sqrto_175_), .Y(u2__abc_52138_new_n4469_));
INVX1 INVX1_701 ( .A(u2_remHi_175_), .Y(u2__abc_52138_new_n4471_));
INVX1 INVX1_702 ( .A(u2__abc_52138_new_n4473_), .Y(u2__abc_52138_new_n4474_));
INVX1 INVX1_703 ( .A(sqrto_172_), .Y(u2__abc_52138_new_n4478_));
INVX1 INVX1_704 ( .A(u2_remHi_172_), .Y(u2__abc_52138_new_n4480_));
INVX1 INVX1_705 ( .A(sqrto_173_), .Y(u2__abc_52138_new_n4483_));
INVX1 INVX1_706 ( .A(u2_remHi_173_), .Y(u2__abc_52138_new_n4485_));
INVX1 INVX1_707 ( .A(sqrto_171_), .Y(u2__abc_52138_new_n4489_));
INVX1 INVX1_708 ( .A(u2_remHi_171_), .Y(u2__abc_52138_new_n4491_));
INVX1 INVX1_709 ( .A(sqrto_170_), .Y(u2__abc_52138_new_n4494_));
INVX1 INVX1_71 ( .A(sqrto_145_), .Y(_abc_65734_new_n1037_));
INVX1 INVX1_710 ( .A(u2_remHi_170_), .Y(u2__abc_52138_new_n4496_));
INVX1 INVX1_711 ( .A(sqrto_168_), .Y(u2__abc_52138_new_n4501_));
INVX1 INVX1_712 ( .A(u2_remHi_168_), .Y(u2__abc_52138_new_n4503_));
INVX1 INVX1_713 ( .A(sqrto_169_), .Y(u2__abc_52138_new_n4506_));
INVX1 INVX1_714 ( .A(u2_remHi_169_), .Y(u2__abc_52138_new_n4508_));
INVX1 INVX1_715 ( .A(sqrto_167_), .Y(u2__abc_52138_new_n4512_));
INVX1 INVX1_716 ( .A(u2_remHi_167_), .Y(u2__abc_52138_new_n4514_));
INVX1 INVX1_717 ( .A(u2_remHi_166_), .Y(u2__abc_52138_new_n4517_));
INVX1 INVX1_718 ( .A(sqrto_166_), .Y(u2__abc_52138_new_n4519_));
INVX1 INVX1_719 ( .A(sqrto_160_), .Y(u2__abc_52138_new_n4525_));
INVX1 INVX1_72 ( .A(sqrto_146_), .Y(_abc_65734_new_n1040_));
INVX1 INVX1_720 ( .A(u2_remHi_160_), .Y(u2__abc_52138_new_n4527_));
INVX1 INVX1_721 ( .A(sqrto_161_), .Y(u2__abc_52138_new_n4530_));
INVX1 INVX1_722 ( .A(u2_remHi_161_), .Y(u2__abc_52138_new_n4532_));
INVX1 INVX1_723 ( .A(sqrto_159_), .Y(u2__abc_52138_new_n4536_));
INVX1 INVX1_724 ( .A(u2__abc_52138_new_n4538_), .Y(u2__abc_52138_new_n4539_));
INVX1 INVX1_725 ( .A(u2_remHi_158_), .Y(u2__abc_52138_new_n4541_));
INVX1 INVX1_726 ( .A(sqrto_158_), .Y(u2__abc_52138_new_n4543_));
INVX1 INVX1_727 ( .A(sqrto_164_), .Y(u2__abc_52138_new_n4548_));
INVX1 INVX1_728 ( .A(u2_remHi_164_), .Y(u2__abc_52138_new_n4550_));
INVX1 INVX1_729 ( .A(sqrto_165_), .Y(u2__abc_52138_new_n4553_));
INVX1 INVX1_73 ( .A(sqrto_147_), .Y(_abc_65734_new_n1043_));
INVX1 INVX1_730 ( .A(u2_remHi_165_), .Y(u2__abc_52138_new_n4555_));
INVX1 INVX1_731 ( .A(sqrto_163_), .Y(u2__abc_52138_new_n4559_));
INVX1 INVX1_732 ( .A(u2_remHi_163_), .Y(u2__abc_52138_new_n4561_));
INVX1 INVX1_733 ( .A(sqrto_162_), .Y(u2__abc_52138_new_n4564_));
INVX1 INVX1_734 ( .A(u2_remHi_162_), .Y(u2__abc_52138_new_n4566_));
INVX1 INVX1_735 ( .A(sqrto_152_), .Y(u2__abc_52138_new_n4573_));
INVX1 INVX1_736 ( .A(u2_remHi_152_), .Y(u2__abc_52138_new_n4575_));
INVX1 INVX1_737 ( .A(sqrto_153_), .Y(u2__abc_52138_new_n4578_));
INVX1 INVX1_738 ( .A(u2_remHi_153_), .Y(u2__abc_52138_new_n4580_));
INVX1 INVX1_739 ( .A(sqrto_151_), .Y(u2__abc_52138_new_n4584_));
INVX1 INVX1_74 ( .A(sqrto_148_), .Y(_abc_65734_new_n1046_));
INVX1 INVX1_740 ( .A(u2_remHi_151_), .Y(u2__abc_52138_new_n4586_));
INVX1 INVX1_741 ( .A(sqrto_150_), .Y(u2__abc_52138_new_n4589_));
INVX1 INVX1_742 ( .A(u2_remHi_150_), .Y(u2__abc_52138_new_n4591_));
INVX1 INVX1_743 ( .A(sqrto_156_), .Y(u2__abc_52138_new_n4596_));
INVX1 INVX1_744 ( .A(u2_remHi_156_), .Y(u2__abc_52138_new_n4598_));
INVX1 INVX1_745 ( .A(sqrto_157_), .Y(u2__abc_52138_new_n4601_));
INVX1 INVX1_746 ( .A(u2_remHi_157_), .Y(u2__abc_52138_new_n4603_));
INVX1 INVX1_747 ( .A(u2_remHi_155_), .Y(u2__abc_52138_new_n4607_));
INVX1 INVX1_748 ( .A(sqrto_155_), .Y(u2__abc_52138_new_n4609_));
INVX1 INVX1_749 ( .A(u2_remHi_154_), .Y(u2__abc_52138_new_n4612_));
INVX1 INVX1_75 ( .A(sqrto_149_), .Y(_abc_65734_new_n1049_));
INVX1 INVX1_750 ( .A(sqrto_154_), .Y(u2__abc_52138_new_n4614_));
INVX1 INVX1_751 ( .A(sqrto_148_), .Y(u2__abc_52138_new_n4619_));
INVX1 INVX1_752 ( .A(u2_remHi_148_), .Y(u2__abc_52138_new_n4621_));
INVX1 INVX1_753 ( .A(sqrto_149_), .Y(u2__abc_52138_new_n4624_));
INVX1 INVX1_754 ( .A(u2_remHi_149_), .Y(u2__abc_52138_new_n4626_));
INVX1 INVX1_755 ( .A(sqrto_147_), .Y(u2__abc_52138_new_n4630_));
INVX1 INVX1_756 ( .A(u2_remHi_147_), .Y(u2__abc_52138_new_n4632_));
INVX1 INVX1_757 ( .A(sqrto_146_), .Y(u2__abc_52138_new_n4635_));
INVX1 INVX1_758 ( .A(u2_remHi_146_), .Y(u2__abc_52138_new_n4637_));
INVX1 INVX1_759 ( .A(sqrto_144_), .Y(u2__abc_52138_new_n4642_));
INVX1 INVX1_76 ( .A(sqrto_150_), .Y(_abc_65734_new_n1052_));
INVX1 INVX1_760 ( .A(u2_remHi_144_), .Y(u2__abc_52138_new_n4644_));
INVX1 INVX1_761 ( .A(sqrto_145_), .Y(u2__abc_52138_new_n4647_));
INVX1 INVX1_762 ( .A(u2_remHi_145_), .Y(u2__abc_52138_new_n4649_));
INVX1 INVX1_763 ( .A(u2_remHi_143_), .Y(u2__abc_52138_new_n4652_));
INVX1 INVX1_764 ( .A(u2__abc_52138_new_n4653_), .Y(u2__abc_52138_new_n4654_));
INVX1 INVX1_765 ( .A(sqrto_143_), .Y(u2__abc_52138_new_n4655_));
INVX1 INVX1_766 ( .A(u2__abc_52138_new_n4656_), .Y(u2__abc_52138_new_n4657_));
INVX1 INVX1_767 ( .A(u2_remHi_142_), .Y(u2__abc_52138_new_n4658_));
INVX1 INVX1_768 ( .A(sqrto_142_), .Y(u2__abc_52138_new_n4660_));
INVX1 INVX1_769 ( .A(sqrto_136_), .Y(u2__abc_52138_new_n4666_));
INVX1 INVX1_77 ( .A(sqrto_151_), .Y(_abc_65734_new_n1055_));
INVX1 INVX1_770 ( .A(u2_remHi_136_), .Y(u2__abc_52138_new_n4668_));
INVX1 INVX1_771 ( .A(sqrto_137_), .Y(u2__abc_52138_new_n4671_));
INVX1 INVX1_772 ( .A(u2_remHi_137_), .Y(u2__abc_52138_new_n4673_));
INVX1 INVX1_773 ( .A(sqrto_134_), .Y(u2__abc_52138_new_n4677_));
INVX1 INVX1_774 ( .A(u2_remHi_134_), .Y(u2__abc_52138_new_n4679_));
INVX1 INVX1_775 ( .A(sqrto_135_), .Y(u2__abc_52138_new_n4682_));
INVX1 INVX1_776 ( .A(u2_remHi_135_), .Y(u2__abc_52138_new_n4684_));
INVX1 INVX1_777 ( .A(sqrto_140_), .Y(u2__abc_52138_new_n4689_));
INVX1 INVX1_778 ( .A(u2_remHi_140_), .Y(u2__abc_52138_new_n4691_));
INVX1 INVX1_779 ( .A(sqrto_141_), .Y(u2__abc_52138_new_n4694_));
INVX1 INVX1_78 ( .A(sqrto_152_), .Y(_abc_65734_new_n1058_));
INVX1 INVX1_780 ( .A(u2_remHi_141_), .Y(u2__abc_52138_new_n4696_));
INVX1 INVX1_781 ( .A(sqrto_139_), .Y(u2__abc_52138_new_n4700_));
INVX1 INVX1_782 ( .A(u2_remHi_139_), .Y(u2__abc_52138_new_n4702_));
INVX1 INVX1_783 ( .A(sqrto_138_), .Y(u2__abc_52138_new_n4705_));
INVX1 INVX1_784 ( .A(u2_remHi_138_), .Y(u2__abc_52138_new_n4707_));
INVX1 INVX1_785 ( .A(sqrto_126_), .Y(u2__abc_52138_new_n4713_));
INVX1 INVX1_786 ( .A(u2_remHi_126_), .Y(u2__abc_52138_new_n4715_));
INVX1 INVX1_787 ( .A(u2__abc_52138_new_n4717_), .Y(u2__abc_52138_new_n4718_));
INVX1 INVX1_788 ( .A(sqrto_127_), .Y(u2__abc_52138_new_n4719_));
INVX1 INVX1_789 ( .A(u2_remHi_127_), .Y(u2__abc_52138_new_n4721_));
INVX1 INVX1_79 ( .A(sqrto_153_), .Y(_abc_65734_new_n1061_));
INVX1 INVX1_790 ( .A(u2__abc_52138_new_n4723_), .Y(u2__abc_52138_new_n4724_));
INVX1 INVX1_791 ( .A(sqrto_129_), .Y(u2__abc_52138_new_n4727_));
INVX1 INVX1_792 ( .A(u2_remHi_129_), .Y(u2__abc_52138_new_n4729_));
INVX1 INVX1_793 ( .A(sqrto_132_), .Y(u2__abc_52138_new_n4733_));
INVX1 INVX1_794 ( .A(u2_remHi_132_), .Y(u2__abc_52138_new_n4735_));
INVX1 INVX1_795 ( .A(sqrto_133_), .Y(u2__abc_52138_new_n4738_));
INVX1 INVX1_796 ( .A(u2_remHi_133_), .Y(u2__abc_52138_new_n4740_));
INVX1 INVX1_797 ( .A(sqrto_131_), .Y(u2__abc_52138_new_n4744_));
INVX1 INVX1_798 ( .A(u2_remHi_131_), .Y(u2__abc_52138_new_n4746_));
INVX1 INVX1_799 ( .A(u2__abc_52138_new_n4477_), .Y(u2__abc_52138_new_n4754_));
INVX1 INVX1_8 ( .A(sqrto_82_), .Y(_abc_65734_new_n848_));
INVX1 INVX1_80 ( .A(sqrto_154_), .Y(_abc_65734_new_n1064_));
INVX1 INVX1_800 ( .A(u2__abc_52138_new_n4500_), .Y(u2__abc_52138_new_n4755_));
INVX1 INVX1_801 ( .A(u2__abc_52138_new_n4716_), .Y(u2__abc_52138_new_n4767_));
INVX1 INVX1_802 ( .A(u2__abc_52138_new_n4722_), .Y(u2__abc_52138_new_n4768_));
INVX1 INVX1_803 ( .A(sqrto_128_), .Y(u2__abc_52138_new_n4770_));
INVX1 INVX1_804 ( .A(u2__abc_52138_new_n4730_), .Y(u2__abc_52138_new_n4772_));
INVX1 INVX1_805 ( .A(u2_remHi_130_), .Y(u2__abc_52138_new_n4776_));
INVX1 INVX1_806 ( .A(u2__abc_52138_new_n4778_), .Y(u2__abc_52138_new_n4779_));
INVX1 INVX1_807 ( .A(u2__abc_52138_new_n4781_), .Y(u2__abc_52138_new_n4782_));
INVX1 INVX1_808 ( .A(u2__abc_52138_new_n4680_), .Y(u2__abc_52138_new_n4786_));
INVX1 INVX1_809 ( .A(u2__abc_52138_new_n4685_), .Y(u2__abc_52138_new_n4787_));
INVX1 INVX1_81 ( .A(sqrto_155_), .Y(_abc_65734_new_n1067_));
INVX1 INVX1_810 ( .A(u2__abc_52138_new_n4790_), .Y(u2__abc_52138_new_n4791_));
INVX1 INVX1_811 ( .A(u2__abc_52138_new_n4701_), .Y(u2__abc_52138_new_n4793_));
INVX1 INVX1_812 ( .A(u2__abc_52138_new_n4796_), .Y(u2__abc_52138_new_n4797_));
INVX1 INVX1_813 ( .A(u2__abc_52138_new_n4808_), .Y(u2__abc_52138_new_n4809_));
INVX1 INVX1_814 ( .A(u2__abc_52138_new_n4617_), .Y(u2__abc_52138_new_n4815_));
INVX1 INVX1_815 ( .A(u2__abc_52138_new_n4585_), .Y(u2__abc_52138_new_n4816_));
INVX1 INVX1_816 ( .A(u2__abc_52138_new_n4819_), .Y(u2__abc_52138_new_n4820_));
INVX1 INVX1_817 ( .A(u2__abc_52138_new_n4825_), .Y(u2__abc_52138_new_n4826_));
INVX1 INVX1_818 ( .A(u2__abc_52138_new_n4834_), .Y(u2__abc_52138_new_n4835_));
INVX1 INVX1_819 ( .A(u2__abc_52138_new_n4839_), .Y(u2__abc_52138_new_n4840_));
INVX1 INVX1_82 ( .A(sqrto_156_), .Y(_abc_65734_new_n1070_));
INVX1 INVX1_820 ( .A(u2__abc_52138_new_n4841_), .Y(u2__abc_52138_new_n4842_));
INVX1 INVX1_821 ( .A(u2__abc_52138_new_n4848_), .Y(u2__abc_52138_new_n4849_));
INVX1 INVX1_822 ( .A(u2__abc_52138_new_n4481_), .Y(u2__abc_52138_new_n4853_));
INVX1 INVX1_823 ( .A(u2__abc_52138_new_n4470_), .Y(u2__abc_52138_new_n4858_));
INVX1 INVX1_824 ( .A(u2__abc_52138_new_n4435_), .Y(u2__abc_52138_new_n4862_));
INVX1 INVX1_825 ( .A(u2__abc_52138_new_n4411_), .Y(u2__abc_52138_new_n4872_));
INVX1 INVX1_826 ( .A(u2__abc_52138_new_n4875_), .Y(u2__abc_52138_new_n4876_));
INVX1 INVX1_827 ( .A(u2__abc_52138_new_n4890_), .Y(u2__abc_52138_new_n4891_));
INVX1 INVX1_828 ( .A(u2__abc_52138_new_n4893_), .Y(u2__abc_52138_new_n4894_));
INVX1 INVX1_829 ( .A(u2__abc_52138_new_n4329_), .Y(u2__abc_52138_new_n4897_));
INVX1 INVX1_83 ( .A(sqrto_157_), .Y(_abc_65734_new_n1073_));
INVX1 INVX1_830 ( .A(u2__abc_52138_new_n4301_), .Y(u2__abc_52138_new_n4898_));
INVX1 INVX1_831 ( .A(u2__abc_52138_new_n4901_), .Y(u2__abc_52138_new_n4902_));
INVX1 INVX1_832 ( .A(u2__abc_52138_new_n4326_), .Y(u2__abc_52138_new_n4904_));
INVX1 INVX1_833 ( .A(u2_remHi_202_), .Y(u2__abc_52138_new_n4905_));
INVX1 INVX1_834 ( .A(u2__abc_52138_new_n4318_), .Y(u2__abc_52138_new_n4909_));
INVX1 INVX1_835 ( .A(u2__abc_52138_new_n4255_), .Y(u2__abc_52138_new_n4914_));
INVX1 INVX1_836 ( .A(u2__abc_52138_new_n4260_), .Y(u2__abc_52138_new_n4915_));
INVX1 INVX1_837 ( .A(u2__abc_52138_new_n4244_), .Y(u2__abc_52138_new_n4917_));
INVX1 INVX1_838 ( .A(u2__abc_52138_new_n4249_), .Y(u2__abc_52138_new_n4918_));
INVX1 INVX1_839 ( .A(u2__abc_52138_new_n4276_), .Y(u2__abc_52138_new_n4921_));
INVX1 INVX1_84 ( .A(sqrto_158_), .Y(_abc_65734_new_n1076_));
INVX1 INVX1_840 ( .A(u2__abc_52138_new_n4272_), .Y(u2__abc_52138_new_n4923_));
INVX1 INVX1_841 ( .A(u2__abc_52138_new_n4931_), .Y(u2__abc_52138_new_n4932_));
INVX1 INVX1_842 ( .A(u2__abc_52138_new_n4223_), .Y(u2__abc_52138_new_n4935_));
INVX1 INVX1_843 ( .A(u2__abc_52138_new_n4231_), .Y(u2__abc_52138_new_n4937_));
INVX1 INVX1_844 ( .A(u2__abc_52138_new_n4939_), .Y(u2__abc_52138_new_n4940_));
INVX1 INVX1_845 ( .A(u2__abc_52138_new_n4190_), .Y(u2__abc_52138_new_n4944_));
INVX1 INVX1_846 ( .A(u2__abc_52138_new_n4158_), .Y(u2__abc_52138_new_n4945_));
INVX1 INVX1_847 ( .A(u2__abc_52138_new_n4948_), .Y(u2__abc_52138_new_n4949_));
INVX1 INVX1_848 ( .A(u2__abc_52138_new_n4175_), .Y(u2__abc_52138_new_n4954_));
INVX1 INVX1_849 ( .A(u2__abc_52138_new_n4955_), .Y(u2__abc_52138_new_n4956_));
INVX1 INVX1_85 ( .A(sqrto_159_), .Y(_abc_65734_new_n1079_));
INVX1 INVX1_850 ( .A(u2_o_231_), .Y(u2__abc_52138_new_n4960_));
INVX1 INVX1_851 ( .A(u2__abc_52138_new_n4968_), .Y(u2__abc_52138_new_n4969_));
INVX1 INVX1_852 ( .A(u2__abc_52138_new_n4974_), .Y(u2__abc_52138_new_n4975_));
INVX1 INVX1_853 ( .A(u2__abc_52138_new_n4979_), .Y(u2__abc_52138_new_n4980_));
INVX1 INVX1_854 ( .A(u2__abc_52138_new_n4080_), .Y(u2__abc_52138_new_n4987_));
INVX1 INVX1_855 ( .A(u2__abc_52138_new_n4088_), .Y(u2__abc_52138_new_n4989_));
INVX1 INVX1_856 ( .A(u2_remHi_380_), .Y(u2__abc_52138_new_n4999_));
INVX1 INVX1_857 ( .A(u2_o_380_), .Y(u2__abc_52138_new_n5001_));
INVX1 INVX1_858 ( .A(u2_o_381_), .Y(u2__abc_52138_new_n5004_));
INVX1 INVX1_859 ( .A(u2_remHi_381_), .Y(u2__abc_52138_new_n5006_));
INVX1 INVX1_86 ( .A(sqrto_160_), .Y(_abc_65734_new_n1082_));
INVX1 INVX1_860 ( .A(u2_remHi_379_), .Y(u2__abc_52138_new_n5011_));
INVX1 INVX1_861 ( .A(u2_o_379_), .Y(u2__abc_52138_new_n5013_));
INVX1 INVX1_862 ( .A(u2_o_374_), .Y(u2__abc_52138_new_n5018_));
INVX1 INVX1_863 ( .A(u2_remHi_374_), .Y(u2__abc_52138_new_n5020_));
INVX1 INVX1_864 ( .A(u2_remHi_375_), .Y(u2__abc_52138_new_n5023_));
INVX1 INVX1_865 ( .A(u2_o_375_), .Y(u2__abc_52138_new_n5025_));
INVX1 INVX1_866 ( .A(u2__abc_52138_new_n5027_), .Y(u2__abc_52138_new_n5028_));
INVX1 INVX1_867 ( .A(u2_remHi_376_), .Y(u2__abc_52138_new_n5030_));
INVX1 INVX1_868 ( .A(u2_o_376_), .Y(u2__abc_52138_new_n5032_));
INVX1 INVX1_869 ( .A(u2_remHi_377_), .Y(u2__abc_52138_new_n5035_));
INVX1 INVX1_87 ( .A(sqrto_161_), .Y(_abc_65734_new_n1085_));
INVX1 INVX1_870 ( .A(u2__abc_52138_new_n5036_), .Y(u2__abc_52138_new_n5037_));
INVX1 INVX1_871 ( .A(u2_o_377_), .Y(u2__abc_52138_new_n5038_));
INVX1 INVX1_872 ( .A(u2__abc_52138_new_n5039_), .Y(u2__abc_52138_new_n5040_));
INVX1 INVX1_873 ( .A(u2_remHi_368_), .Y(u2__abc_52138_new_n5045_));
INVX1 INVX1_874 ( .A(u2_o_368_), .Y(u2__abc_52138_new_n5047_));
INVX1 INVX1_875 ( .A(u2_remHi_366_), .Y(u2__abc_52138_new_n5052_));
INVX1 INVX1_876 ( .A(u2__abc_52138_new_n5053_), .Y(u2__abc_52138_new_n5054_));
INVX1 INVX1_877 ( .A(u2_o_367_), .Y(u2__abc_52138_new_n5057_));
INVX1 INVX1_878 ( .A(u2_remHi_367_), .Y(u2__abc_52138_new_n5059_));
INVX1 INVX1_879 ( .A(u2__abc_52138_new_n5061_), .Y(u2__abc_52138_new_n5062_));
INVX1 INVX1_88 ( .A(sqrto_162_), .Y(_abc_65734_new_n1088_));
INVX1 INVX1_880 ( .A(u2_remHi_372_), .Y(u2__abc_52138_new_n5065_));
INVX1 INVX1_881 ( .A(u2_o_372_), .Y(u2__abc_52138_new_n5067_));
INVX1 INVX1_882 ( .A(u2_remHi_373_), .Y(u2__abc_52138_new_n5070_));
INVX1 INVX1_883 ( .A(u2_o_373_), .Y(u2__abc_52138_new_n5072_));
INVX1 INVX1_884 ( .A(u2_o_371_), .Y(u2__abc_52138_new_n5076_));
INVX1 INVX1_885 ( .A(u2_remHi_371_), .Y(u2__abc_52138_new_n5078_));
INVX1 INVX1_886 ( .A(u2__abc_52138_new_n5080_), .Y(u2__abc_52138_new_n5081_));
INVX1 INVX1_887 ( .A(u2_o_370_), .Y(u2__abc_52138_new_n5082_));
INVX1 INVX1_888 ( .A(u2_remHi_370_), .Y(u2__abc_52138_new_n5084_));
INVX1 INVX1_889 ( .A(u2_o_358_), .Y(u2__abc_52138_new_n5091_));
INVX1 INVX1_89 ( .A(sqrto_163_), .Y(_abc_65734_new_n1091_));
INVX1 INVX1_890 ( .A(u2_remHi_358_), .Y(u2__abc_52138_new_n5093_));
INVX1 INVX1_891 ( .A(u2_remHi_359_), .Y(u2__abc_52138_new_n5096_));
INVX1 INVX1_892 ( .A(u2_o_359_), .Y(u2__abc_52138_new_n5098_));
INVX1 INVX1_893 ( .A(u2_remHi_360_), .Y(u2__abc_52138_new_n5102_));
INVX1 INVX1_894 ( .A(u2_o_360_), .Y(u2__abc_52138_new_n5104_));
INVX1 INVX1_895 ( .A(u2_o_361_), .Y(u2__abc_52138_new_n5107_));
INVX1 INVX1_896 ( .A(u2_remHi_361_), .Y(u2__abc_52138_new_n5109_));
INVX1 INVX1_897 ( .A(u2_remHi_364_), .Y(u2__abc_52138_new_n5114_));
INVX1 INVX1_898 ( .A(u2_o_364_), .Y(u2__abc_52138_new_n5116_));
INVX1 INVX1_899 ( .A(u2_remHi_365_), .Y(u2__abc_52138_new_n5119_));
INVX1 INVX1_9 ( .A(sqrto_83_), .Y(_abc_65734_new_n851_));
INVX1 INVX1_90 ( .A(sqrto_164_), .Y(_abc_65734_new_n1094_));
INVX1 INVX1_900 ( .A(u2_o_365_), .Y(u2__abc_52138_new_n5121_));
INVX1 INVX1_901 ( .A(u2_remHi_363_), .Y(u2__abc_52138_new_n5126_));
INVX1 INVX1_902 ( .A(u2_o_363_), .Y(u2__abc_52138_new_n5128_));
INVX1 INVX1_903 ( .A(u2_remHi_352_), .Y(u2__abc_52138_new_n5134_));
INVX1 INVX1_904 ( .A(u2_o_352_), .Y(u2__abc_52138_new_n5136_));
INVX1 INVX1_905 ( .A(u2_remHi_353_), .Y(u2__abc_52138_new_n5139_));
INVX1 INVX1_906 ( .A(u2_o_353_), .Y(u2__abc_52138_new_n5141_));
INVX1 INVX1_907 ( .A(u2_remHi_350_), .Y(u2__abc_52138_new_n5145_));
INVX1 INVX1_908 ( .A(u2_o_350_), .Y(u2__abc_52138_new_n5147_));
INVX1 INVX1_909 ( .A(u2_remHi_351_), .Y(u2__abc_52138_new_n5150_));
INVX1 INVX1_91 ( .A(sqrto_165_), .Y(_abc_65734_new_n1097_));
INVX1 INVX1_910 ( .A(u2_o_351_), .Y(u2__abc_52138_new_n5152_));
INVX1 INVX1_911 ( .A(u2_remHi_356_), .Y(u2__abc_52138_new_n5157_));
INVX1 INVX1_912 ( .A(u2_o_356_), .Y(u2__abc_52138_new_n5159_));
INVX1 INVX1_913 ( .A(u2_remHi_357_), .Y(u2__abc_52138_new_n5162_));
INVX1 INVX1_914 ( .A(u2_o_357_), .Y(u2__abc_52138_new_n5164_));
INVX1 INVX1_915 ( .A(u2_remHi_354_), .Y(u2__abc_52138_new_n5168_));
INVX1 INVX1_916 ( .A(u2_o_354_), .Y(u2__abc_52138_new_n5170_));
INVX1 INVX1_917 ( .A(u2_remHi_355_), .Y(u2__abc_52138_new_n5173_));
INVX1 INVX1_918 ( .A(u2_o_355_), .Y(u2__abc_52138_new_n5175_));
INVX1 INVX1_919 ( .A(u2_o_344_), .Y(u2__abc_52138_new_n5183_));
INVX1 INVX1_92 ( .A(sqrto_166_), .Y(_abc_65734_new_n1100_));
INVX1 INVX1_920 ( .A(u2_remHi_344_), .Y(u2__abc_52138_new_n5185_));
INVX1 INVX1_921 ( .A(u2_remHi_345_), .Y(u2__abc_52138_new_n5188_));
INVX1 INVX1_922 ( .A(u2_o_345_), .Y(u2__abc_52138_new_n5190_));
INVX1 INVX1_923 ( .A(u2__abc_52138_new_n5193_), .Y(u2__abc_52138_new_n5194_));
INVX1 INVX1_924 ( .A(u2_remHi_342_), .Y(u2__abc_52138_new_n5195_));
INVX1 INVX1_925 ( .A(u2_o_342_), .Y(u2__abc_52138_new_n5197_));
INVX1 INVX1_926 ( .A(u2_remHi_343_), .Y(u2__abc_52138_new_n5200_));
INVX1 INVX1_927 ( .A(u2_o_343_), .Y(u2__abc_52138_new_n5202_));
INVX1 INVX1_928 ( .A(u2_o_348_), .Y(u2__abc_52138_new_n5206_));
INVX1 INVX1_929 ( .A(u2_remHi_348_), .Y(u2__abc_52138_new_n5208_));
INVX1 INVX1_93 ( .A(sqrto_167_), .Y(_abc_65734_new_n1103_));
INVX1 INVX1_930 ( .A(u2_remHi_349_), .Y(u2__abc_52138_new_n5210_));
INVX1 INVX1_931 ( .A(u2_o_349_), .Y(u2__abc_52138_new_n5212_));
INVX1 INVX1_932 ( .A(u2_remHi_346_), .Y(u2__abc_52138_new_n5216_));
INVX1 INVX1_933 ( .A(u2_o_346_), .Y(u2__abc_52138_new_n5218_));
INVX1 INVX1_934 ( .A(u2_remHi_347_), .Y(u2__abc_52138_new_n5221_));
INVX1 INVX1_935 ( .A(u2_o_347_), .Y(u2__abc_52138_new_n5223_));
INVX1 INVX1_936 ( .A(u2_remHi_336_), .Y(u2__abc_52138_new_n5229_));
INVX1 INVX1_937 ( .A(u2_o_336_), .Y(u2__abc_52138_new_n5231_));
INVX1 INVX1_938 ( .A(u2_remHi_337_), .Y(u2__abc_52138_new_n5234_));
INVX1 INVX1_939 ( .A(u2_o_337_), .Y(u2__abc_52138_new_n5236_));
INVX1 INVX1_94 ( .A(sqrto_168_), .Y(_abc_65734_new_n1106_));
INVX1 INVX1_940 ( .A(u2__abc_52138_new_n5239_), .Y(u2__abc_52138_new_n5240_));
INVX1 INVX1_941 ( .A(u2_o_335_), .Y(u2__abc_52138_new_n5242_));
INVX1 INVX1_942 ( .A(u2_remHi_335_), .Y(u2__abc_52138_new_n5244_));
INVX1 INVX1_943 ( .A(u2__abc_52138_new_n5246_), .Y(u2__abc_52138_new_n5247_));
INVX1 INVX1_944 ( .A(u2_o_340_), .Y(u2__abc_52138_new_n5249_));
INVX1 INVX1_945 ( .A(u2_remHi_340_), .Y(u2__abc_52138_new_n5251_));
INVX1 INVX1_946 ( .A(u2_remHi_341_), .Y(u2__abc_52138_new_n5254_));
INVX1 INVX1_947 ( .A(u2_o_341_), .Y(u2__abc_52138_new_n5256_));
INVX1 INVX1_948 ( .A(u2__abc_52138_new_n5259_), .Y(u2__abc_52138_new_n5260_));
INVX1 INVX1_949 ( .A(u2_remHi_338_), .Y(u2__abc_52138_new_n5261_));
INVX1 INVX1_95 ( .A(sqrto_169_), .Y(_abc_65734_new_n1109_));
INVX1 INVX1_950 ( .A(u2__abc_52138_new_n5262_), .Y(u2__abc_52138_new_n5263_));
INVX1 INVX1_951 ( .A(u2_remHi_339_), .Y(u2__abc_52138_new_n5266_));
INVX1 INVX1_952 ( .A(u2_o_339_), .Y(u2__abc_52138_new_n5268_));
INVX1 INVX1_953 ( .A(u2_o_326_), .Y(u2__abc_52138_new_n5274_));
INVX1 INVX1_954 ( .A(u2_remHi_326_), .Y(u2__abc_52138_new_n5276_));
INVX1 INVX1_955 ( .A(u2_remHi_327_), .Y(u2__abc_52138_new_n5279_));
INVX1 INVX1_956 ( .A(u2_o_327_), .Y(u2__abc_52138_new_n5281_));
INVX1 INVX1_957 ( .A(u2_remHi_328_), .Y(u2__abc_52138_new_n5285_));
INVX1 INVX1_958 ( .A(u2_o_328_), .Y(u2__abc_52138_new_n5287_));
INVX1 INVX1_959 ( .A(u2_remHi_329_), .Y(u2__abc_52138_new_n5290_));
INVX1 INVX1_96 ( .A(sqrto_170_), .Y(_abc_65734_new_n1112_));
INVX1 INVX1_960 ( .A(u2_o_329_), .Y(u2__abc_52138_new_n5292_));
INVX1 INVX1_961 ( .A(u2_remHi_332_), .Y(u2__abc_52138_new_n5297_));
INVX1 INVX1_962 ( .A(u2_o_332_), .Y(u2__abc_52138_new_n5299_));
INVX1 INVX1_963 ( .A(u2_remHi_333_), .Y(u2__abc_52138_new_n5302_));
INVX1 INVX1_964 ( .A(u2_o_333_), .Y(u2__abc_52138_new_n5304_));
INVX1 INVX1_965 ( .A(u2_remHi_330_), .Y(u2__abc_52138_new_n5308_));
INVX1 INVX1_966 ( .A(u2_o_330_), .Y(u2__abc_52138_new_n5310_));
INVX1 INVX1_967 ( .A(u2_remHi_331_), .Y(u2__abc_52138_new_n5313_));
INVX1 INVX1_968 ( .A(u2_o_331_), .Y(u2__abc_52138_new_n5315_));
INVX1 INVX1_969 ( .A(u2_o_324_), .Y(u2__abc_52138_new_n5321_));
INVX1 INVX1_97 ( .A(sqrto_171_), .Y(_abc_65734_new_n1115_));
INVX1 INVX1_970 ( .A(u2_remHi_324_), .Y(u2__abc_52138_new_n5323_));
INVX1 INVX1_971 ( .A(u2_o_325_), .Y(u2__abc_52138_new_n5326_));
INVX1 INVX1_972 ( .A(u2_remHi_325_), .Y(u2__abc_52138_new_n5328_));
INVX1 INVX1_973 ( .A(u2_o_323_), .Y(u2__abc_52138_new_n5333_));
INVX1 INVX1_974 ( .A(u2_remHi_323_), .Y(u2__abc_52138_new_n5335_));
INVX1 INVX1_975 ( .A(u2__abc_52138_new_n5339_), .Y(u2__abc_52138_new_n5340_));
INVX1 INVX1_976 ( .A(u2_o_318_), .Y(u2__abc_52138_new_n5341_));
INVX1 INVX1_977 ( .A(u2_remHi_318_), .Y(u2__abc_52138_new_n5343_));
INVX1 INVX1_978 ( .A(u2_remHi_319_), .Y(u2__abc_52138_new_n5346_));
INVX1 INVX1_979 ( .A(u2_o_319_), .Y(u2__abc_52138_new_n5348_));
INVX1 INVX1_98 ( .A(sqrto_172_), .Y(_abc_65734_new_n1118_));
INVX1 INVX1_980 ( .A(u2_remHi_320_), .Y(u2__abc_52138_new_n5352_));
INVX1 INVX1_981 ( .A(u2_o_320_), .Y(u2__abc_52138_new_n5354_));
INVX1 INVX1_982 ( .A(u2_remHi_321_), .Y(u2__abc_52138_new_n5357_));
INVX1 INVX1_983 ( .A(u2_o_321_), .Y(u2__abc_52138_new_n5359_));
INVX1 INVX1_984 ( .A(u2_remHi_312_), .Y(u2__abc_52138_new_n5368_));
INVX1 INVX1_985 ( .A(u2_o_312_), .Y(u2__abc_52138_new_n5370_));
INVX1 INVX1_986 ( .A(u2_remHi_313_), .Y(u2__abc_52138_new_n5373_));
INVX1 INVX1_987 ( .A(u2_o_313_), .Y(u2__abc_52138_new_n5375_));
INVX1 INVX1_988 ( .A(u2_remHi_311_), .Y(u2__abc_52138_new_n5380_));
INVX1 INVX1_989 ( .A(u2_o_311_), .Y(u2__abc_52138_new_n5382_));
INVX1 INVX1_99 ( .A(sqrto_173_), .Y(_abc_65734_new_n1121_));
INVX1 INVX1_990 ( .A(u2_remHi_316_), .Y(u2__abc_52138_new_n5387_));
INVX1 INVX1_991 ( .A(u2_o_316_), .Y(u2__abc_52138_new_n5389_));
INVX1 INVX1_992 ( .A(u2_remHi_317_), .Y(u2__abc_52138_new_n5392_));
INVX1 INVX1_993 ( .A(u2_o_317_), .Y(u2__abc_52138_new_n5394_));
INVX1 INVX1_994 ( .A(u2_remHi_315_), .Y(u2__abc_52138_new_n5399_));
INVX1 INVX1_995 ( .A(u2_o_315_), .Y(u2__abc_52138_new_n5401_));
INVX1 INVX1_996 ( .A(u2_o_302_), .Y(u2__abc_52138_new_n5407_));
INVX1 INVX1_997 ( .A(u2_remHi_302_), .Y(u2__abc_52138_new_n5409_));
INVX1 INVX1_998 ( .A(u2_o_303_), .Y(u2__abc_52138_new_n5412_));
INVX1 INVX1_999 ( .A(u2_remHi_303_), .Y(u2__abc_52138_new_n5414_));
NAND2X1 NAND2X1_1 ( .A(aNan), .B(\a[0] ), .Y(_abc_65734_new_n831_));
NAND2X1 NAND2X1_10 ( .A(aNan), .B(\a[9] ), .Y(_abc_65734_new_n858_));
NAND2X1 NAND2X1_100 ( .A(aNan), .B(\a[99] ), .Y(_abc_65734_new_n1128_));
NAND2X1 NAND2X1_1000 ( .A(u2_remHi_371_), .B(u2__abc_52138_new_n5076_), .Y(u2__abc_52138_new_n5077_));
NAND2X1 NAND2X1_1001 ( .A(u2_o_371_), .B(u2__abc_52138_new_n5078_), .Y(u2__abc_52138_new_n5079_));
NAND2X1 NAND2X1_1002 ( .A(u2__abc_52138_new_n5077_), .B(u2__abc_52138_new_n5079_), .Y(u2__abc_52138_new_n5080_));
NAND2X1 NAND2X1_1003 ( .A(u2_remHi_370_), .B(u2__abc_52138_new_n5082_), .Y(u2__abc_52138_new_n5083_));
NAND2X1 NAND2X1_1004 ( .A(u2_o_370_), .B(u2__abc_52138_new_n5084_), .Y(u2__abc_52138_new_n5085_));
NAND2X1 NAND2X1_1005 ( .A(u2__abc_52138_new_n5086_), .B(u2__abc_52138_new_n5081_), .Y(u2__abc_52138_new_n5087_));
NAND2X1 NAND2X1_1006 ( .A(u2__abc_52138_new_n5088_), .B(u2__abc_52138_new_n5064_), .Y(u2__abc_52138_new_n5089_));
NAND2X1 NAND2X1_1007 ( .A(u2_o_359_), .B(u2__abc_52138_new_n5096_), .Y(u2__abc_52138_new_n5097_));
NAND2X1 NAND2X1_1008 ( .A(u2_remHi_359_), .B(u2__abc_52138_new_n5098_), .Y(u2__abc_52138_new_n5099_));
NAND2X1 NAND2X1_1009 ( .A(u2__abc_52138_new_n5100_), .B(u2__abc_52138_new_n5095_), .Y(u2__abc_52138_new_n5101_));
NAND2X1 NAND2X1_101 ( .A(aNan), .B(\a[100] ), .Y(_abc_65734_new_n1131_));
NAND2X1 NAND2X1_1010 ( .A(u2_remHi_361_), .B(u2__abc_52138_new_n5107_), .Y(u2__abc_52138_new_n5108_));
NAND2X1 NAND2X1_1011 ( .A(u2_o_361_), .B(u2__abc_52138_new_n5109_), .Y(u2__abc_52138_new_n5110_));
NAND2X1 NAND2X1_1012 ( .A(u2__abc_52138_new_n5111_), .B(u2__abc_52138_new_n5106_), .Y(u2__abc_52138_new_n5112_));
NAND2X1 NAND2X1_1013 ( .A(u2__abc_52138_new_n5118_), .B(u2__abc_52138_new_n5123_), .Y(u2__abc_52138_new_n5124_));
NAND2X1 NAND2X1_1014 ( .A(u2__abc_52138_new_n5125_), .B(u2__abc_52138_new_n5130_), .Y(u2__abc_52138_new_n5131_));
NAND2X1 NAND2X1_1015 ( .A(u2__abc_52138_new_n5138_), .B(u2__abc_52138_new_n5143_), .Y(u2__abc_52138_new_n5144_));
NAND2X1 NAND2X1_1016 ( .A(u2__abc_52138_new_n5149_), .B(u2__abc_52138_new_n5154_), .Y(u2__abc_52138_new_n5155_));
NAND2X1 NAND2X1_1017 ( .A(u2__abc_52138_new_n5161_), .B(u2__abc_52138_new_n5166_), .Y(u2__abc_52138_new_n5167_));
NAND2X1 NAND2X1_1018 ( .A(u2__abc_52138_new_n5172_), .B(u2__abc_52138_new_n5177_), .Y(u2__abc_52138_new_n5178_));
NAND2X1 NAND2X1_1019 ( .A(u2__abc_52138_new_n5156_), .B(u2__abc_52138_new_n5179_), .Y(u2__abc_52138_new_n5180_));
NAND2X1 NAND2X1_102 ( .A(aNan), .B(\a[101] ), .Y(_abc_65734_new_n1134_));
NAND2X1 NAND2X1_1020 ( .A(u2_remHi_344_), .B(u2__abc_52138_new_n5183_), .Y(u2__abc_52138_new_n5184_));
NAND2X1 NAND2X1_1021 ( .A(u2_o_344_), .B(u2__abc_52138_new_n5185_), .Y(u2__abc_52138_new_n5186_));
NAND2X1 NAND2X1_1022 ( .A(u2__abc_52138_new_n5187_), .B(u2__abc_52138_new_n5192_), .Y(u2__abc_52138_new_n5193_));
NAND2X1 NAND2X1_1023 ( .A(u2_remHi_348_), .B(u2__abc_52138_new_n5206_), .Y(u2__abc_52138_new_n5207_));
NAND2X1 NAND2X1_1024 ( .A(u2_o_348_), .B(u2__abc_52138_new_n5208_), .Y(u2__abc_52138_new_n5209_));
NAND2X1 NAND2X1_1025 ( .A(u2__abc_52138_new_n5220_), .B(u2__abc_52138_new_n5225_), .Y(u2__abc_52138_new_n5226_));
NAND2X1 NAND2X1_1026 ( .A(u2__abc_52138_new_n5233_), .B(u2__abc_52138_new_n5238_), .Y(u2__abc_52138_new_n5239_));
NAND2X1 NAND2X1_1027 ( .A(u2_remHi_335_), .B(u2__abc_52138_new_n5242_), .Y(u2__abc_52138_new_n5243_));
NAND2X1 NAND2X1_1028 ( .A(u2_o_335_), .B(u2__abc_52138_new_n5244_), .Y(u2__abc_52138_new_n5245_));
NAND2X1 NAND2X1_1029 ( .A(u2__abc_52138_new_n5243_), .B(u2__abc_52138_new_n5245_), .Y(u2__abc_52138_new_n5246_));
NAND2X1 NAND2X1_103 ( .A(aNan), .B(\a[102] ), .Y(_abc_65734_new_n1137_));
NAND2X1 NAND2X1_1030 ( .A(u2_remHi_340_), .B(u2__abc_52138_new_n5249_), .Y(u2__abc_52138_new_n5250_));
NAND2X1 NAND2X1_1031 ( .A(u2_o_340_), .B(u2__abc_52138_new_n5251_), .Y(u2__abc_52138_new_n5252_));
NAND2X1 NAND2X1_1032 ( .A(u2__abc_52138_new_n5253_), .B(u2__abc_52138_new_n5258_), .Y(u2__abc_52138_new_n5259_));
NAND2X1 NAND2X1_1033 ( .A(u2_o_338_), .B(u2__abc_52138_new_n5261_), .Y(u2__abc_52138_new_n5264_));
NAND2X1 NAND2X1_1034 ( .A(u2__abc_52138_new_n5228_), .B(u2__abc_52138_new_n5272_), .Y(u2__abc_52138_new_n5273_));
NAND2X1 NAND2X1_1035 ( .A(u2_o_327_), .B(u2__abc_52138_new_n5279_), .Y(u2__abc_52138_new_n5280_));
NAND2X1 NAND2X1_1036 ( .A(u2_remHi_327_), .B(u2__abc_52138_new_n5281_), .Y(u2__abc_52138_new_n5282_));
NAND2X1 NAND2X1_1037 ( .A(u2__abc_52138_new_n5283_), .B(u2__abc_52138_new_n5278_), .Y(u2__abc_52138_new_n5284_));
NAND2X1 NAND2X1_1038 ( .A(u2__abc_52138_new_n5289_), .B(u2__abc_52138_new_n5294_), .Y(u2__abc_52138_new_n5295_));
NAND2X1 NAND2X1_1039 ( .A(u2__abc_52138_new_n5301_), .B(u2__abc_52138_new_n5306_), .Y(u2__abc_52138_new_n5307_));
NAND2X1 NAND2X1_104 ( .A(aNan), .B(\a[103] ), .Y(_abc_65734_new_n1140_));
NAND2X1 NAND2X1_1040 ( .A(u2__abc_52138_new_n5312_), .B(u2__abc_52138_new_n5317_), .Y(u2__abc_52138_new_n5318_));
NAND2X1 NAND2X1_1041 ( .A(u2__abc_52138_new_n5325_), .B(u2__abc_52138_new_n5330_), .Y(u2__abc_52138_new_n5331_));
NAND2X1 NAND2X1_1042 ( .A(u2_remHi_323_), .B(u2__abc_52138_new_n5333_), .Y(u2__abc_52138_new_n5334_));
NAND2X1 NAND2X1_1043 ( .A(u2_o_323_), .B(u2__abc_52138_new_n5335_), .Y(u2__abc_52138_new_n5336_));
NAND2X1 NAND2X1_1044 ( .A(u2__abc_52138_new_n5332_), .B(u2__abc_52138_new_n5337_), .Y(u2__abc_52138_new_n5338_));
NAND2X1 NAND2X1_1045 ( .A(u2_o_319_), .B(u2__abc_52138_new_n5346_), .Y(u2__abc_52138_new_n5347_));
NAND2X1 NAND2X1_1046 ( .A(u2_remHi_319_), .B(u2__abc_52138_new_n5348_), .Y(u2__abc_52138_new_n5349_));
NAND2X1 NAND2X1_1047 ( .A(u2__abc_52138_new_n5350_), .B(u2__abc_52138_new_n5345_), .Y(u2__abc_52138_new_n5351_));
NAND2X1 NAND2X1_1048 ( .A(u2__abc_52138_new_n5356_), .B(u2__abc_52138_new_n5361_), .Y(u2__abc_52138_new_n5362_));
NAND2X1 NAND2X1_1049 ( .A(u2__abc_52138_new_n5320_), .B(u2__abc_52138_new_n5364_), .Y(u2__abc_52138_new_n5365_));
NAND2X1 NAND2X1_105 ( .A(aNan), .B(\a[104] ), .Y(_abc_65734_new_n1143_));
NAND2X1 NAND2X1_1050 ( .A(u2__abc_52138_new_n5366_), .B(u2__abc_52138_new_n5182_), .Y(u2__abc_52138_new_n5367_));
NAND2X1 NAND2X1_1051 ( .A(u2__abc_52138_new_n5372_), .B(u2__abc_52138_new_n5377_), .Y(u2__abc_52138_new_n5378_));
NAND2X1 NAND2X1_1052 ( .A(u2__abc_52138_new_n5379_), .B(u2__abc_52138_new_n5384_), .Y(u2__abc_52138_new_n5385_));
NAND2X1 NAND2X1_1053 ( .A(u2__abc_52138_new_n5391_), .B(u2__abc_52138_new_n5396_), .Y(u2__abc_52138_new_n5397_));
NAND2X1 NAND2X1_1054 ( .A(u2__abc_52138_new_n5398_), .B(u2__abc_52138_new_n5403_), .Y(u2__abc_52138_new_n5404_));
NAND2X1 NAND2X1_1055 ( .A(u2__abc_52138_new_n5386_), .B(u2__abc_52138_new_n5405_), .Y(u2__abc_52138_new_n5406_));
NAND2X1 NAND2X1_1056 ( .A(u2__abc_52138_new_n5411_), .B(u2__abc_52138_new_n5416_), .Y(u2__abc_52138_new_n5417_));
NAND2X1 NAND2X1_1057 ( .A(u2__abc_52138_new_n5422_), .B(u2__abc_52138_new_n5427_), .Y(u2__abc_52138_new_n5428_));
NAND2X1 NAND2X1_1058 ( .A(u2__abc_52138_new_n5434_), .B(u2__abc_52138_new_n5439_), .Y(u2__abc_52138_new_n5440_));
NAND2X1 NAND2X1_1059 ( .A(u2__abc_52138_new_n5445_), .B(u2__abc_52138_new_n5450_), .Y(u2__abc_52138_new_n5451_));
NAND2X1 NAND2X1_106 ( .A(aNan), .B(\a[105] ), .Y(_abc_65734_new_n1146_));
NAND2X1 NAND2X1_1060 ( .A(u2__abc_52138_new_n5429_), .B(u2__abc_52138_new_n5452_), .Y(u2__abc_52138_new_n5453_));
NAND2X1 NAND2X1_1061 ( .A(u2_o_295_), .B(u2__abc_52138_new_n5460_), .Y(u2__abc_52138_new_n5461_));
NAND2X1 NAND2X1_1062 ( .A(u2_remHi_295_), .B(u2__abc_52138_new_n5462_), .Y(u2__abc_52138_new_n5463_));
NAND2X1 NAND2X1_1063 ( .A(u2__abc_52138_new_n5464_), .B(u2__abc_52138_new_n5459_), .Y(u2__abc_52138_new_n5465_));
NAND2X1 NAND2X1_1064 ( .A(u2__abc_52138_new_n5470_), .B(u2__abc_52138_new_n5475_), .Y(u2__abc_52138_new_n5476_));
NAND2X1 NAND2X1_1065 ( .A(u2__abc_52138_new_n5482_), .B(u2__abc_52138_new_n5487_), .Y(u2__abc_52138_new_n5488_));
NAND2X1 NAND2X1_1066 ( .A(u2__abc_52138_new_n5493_), .B(u2__abc_52138_new_n5498_), .Y(u2__abc_52138_new_n5499_));
NAND2X1 NAND2X1_1067 ( .A(u2__abc_52138_new_n5477_), .B(u2__abc_52138_new_n5500_), .Y(u2__abc_52138_new_n5501_));
NAND2X1 NAND2X1_1068 ( .A(u2__abc_52138_new_n5506_), .B(u2__abc_52138_new_n5511_), .Y(u2__abc_52138_new_n5512_));
NAND2X1 NAND2X1_1069 ( .A(u2__abc_52138_new_n5517_), .B(u2__abc_52138_new_n5522_), .Y(u2__abc_52138_new_n5523_));
NAND2X1 NAND2X1_107 ( .A(aNan), .B(\a[106] ), .Y(_abc_65734_new_n1149_));
NAND2X1 NAND2X1_1070 ( .A(u2__abc_52138_new_n5529_), .B(u2__abc_52138_new_n5534_), .Y(u2__abc_52138_new_n5535_));
NAND2X1 NAND2X1_1071 ( .A(u2__abc_52138_new_n5536_), .B(u2__abc_52138_new_n5541_), .Y(u2__abc_52138_new_n5542_));
NAND2X1 NAND2X1_1072 ( .A(u2__abc_52138_new_n5543_), .B(u2__abc_52138_new_n5524_), .Y(u2__abc_52138_new_n5544_));
NAND2X1 NAND2X1_1073 ( .A(u2__abc_52138_new_n5454_), .B(u2__abc_52138_new_n5545_), .Y(u2__abc_52138_new_n5546_));
NAND2X1 NAND2X1_1074 ( .A(u2__abc_52138_new_n5552_), .B(u2__abc_52138_new_n5557_), .Y(u2__abc_52138_new_n5558_));
NAND2X1 NAND2X1_1075 ( .A(u2__abc_52138_new_n5563_), .B(u2__abc_52138_new_n5568_), .Y(u2__abc_52138_new_n5569_));
NAND2X1 NAND2X1_1076 ( .A(u2__abc_52138_new_n5575_), .B(u2__abc_52138_new_n5580_), .Y(u2__abc_52138_new_n5581_));
NAND2X1 NAND2X1_1077 ( .A(u2__abc_52138_new_n5586_), .B(u2__abc_52138_new_n5591_), .Y(u2__abc_52138_new_n5592_));
NAND2X1 NAND2X1_1078 ( .A(u2__abc_52138_new_n5570_), .B(u2__abc_52138_new_n5593_), .Y(u2__abc_52138_new_n5594_));
NAND2X1 NAND2X1_1079 ( .A(u2__abc_52138_new_n5599_), .B(u2__abc_52138_new_n5604_), .Y(u2__abc_52138_new_n5605_));
NAND2X1 NAND2X1_108 ( .A(aNan), .B(\a[107] ), .Y(_abc_65734_new_n1152_));
NAND2X1 NAND2X1_1080 ( .A(u2__abc_52138_new_n5610_), .B(u2__abc_52138_new_n5615_), .Y(u2__abc_52138_new_n5616_));
NAND2X1 NAND2X1_1081 ( .A(u2__abc_52138_new_n5622_), .B(u2__abc_52138_new_n5627_), .Y(u2__abc_52138_new_n5628_));
NAND2X1 NAND2X1_1082 ( .A(u2__abc_52138_new_n5629_), .B(u2__abc_52138_new_n5634_), .Y(u2__abc_52138_new_n5635_));
NAND2X1 NAND2X1_1083 ( .A(u2__abc_52138_new_n5636_), .B(u2__abc_52138_new_n5617_), .Y(u2__abc_52138_new_n5637_));
NAND2X1 NAND2X1_1084 ( .A(u2__abc_52138_new_n5644_), .B(u2__abc_52138_new_n5649_), .Y(u2__abc_52138_new_n5650_));
NAND2X1 NAND2X1_1085 ( .A(u2__abc_52138_new_n5655_), .B(u2__abc_52138_new_n5660_), .Y(u2__abc_52138_new_n5661_));
NAND2X1 NAND2X1_1086 ( .A(u2__abc_52138_new_n5667_), .B(u2__abc_52138_new_n5672_), .Y(u2__abc_52138_new_n5673_));
NAND2X1 NAND2X1_1087 ( .A(u2__abc_52138_new_n5678_), .B(u2__abc_52138_new_n5683_), .Y(u2__abc_52138_new_n5684_));
NAND2X1 NAND2X1_1088 ( .A(u2__abc_52138_new_n5662_), .B(u2__abc_52138_new_n5685_), .Y(u2__abc_52138_new_n5686_));
NAND2X1 NAND2X1_1089 ( .A(u2_o_255_), .B(u2__abc_52138_new_n5688_), .Y(u2__abc_52138_new_n5689_));
NAND2X1 NAND2X1_109 ( .A(aNan), .B(\a[108] ), .Y(_abc_65734_new_n1155_));
NAND2X1 NAND2X1_1090 ( .A(u2_remHi_255_), .B(u2__abc_52138_new_n5692_), .Y(u2__abc_52138_new_n5693_));
NAND2X1 NAND2X1_1091 ( .A(u2__abc_52138_new_n5701_), .B(u2__abc_52138_new_n5706_), .Y(u2__abc_52138_new_n5707_));
NAND2X1 NAND2X1_1092 ( .A(u2__abc_52138_new_n5713_), .B(u2__abc_52138_new_n5718_), .Y(u2__abc_52138_new_n5719_));
NAND2X1 NAND2X1_1093 ( .A(u2__abc_52138_new_n5724_), .B(u2__abc_52138_new_n5729_), .Y(u2__abc_52138_new_n5730_));
NAND2X1 NAND2X1_1094 ( .A(u2__abc_52138_new_n5731_), .B(u2__abc_52138_new_n5708_), .Y(u2__abc_52138_new_n5732_));
NAND2X1 NAND2X1_1095 ( .A(u2__abc_52138_new_n5547_), .B(u2__abc_52138_new_n5734_), .Y(u2__abc_52138_new_n5735_));
NAND2X1 NAND2X1_1096 ( .A(u2__abc_52138_new_n5662_), .B(u2__abc_52138_new_n5749_), .Y(u2__abc_52138_new_n5750_));
NAND2X1 NAND2X1_1097 ( .A(u2_o_275_), .B(u2__abc_52138_new_n5630_), .Y(u2__abc_52138_new_n5762_));
NAND2X1 NAND2X1_1098 ( .A(u2__abc_52138_new_n5593_), .B(u2__abc_52138_new_n5772_), .Y(u2__abc_52138_new_n5773_));
NAND2X1 NAND2X1_1099 ( .A(u2__abc_52138_new_n5780_), .B(u2__abc_52138_new_n5755_), .Y(u2__abc_52138_new_n5781_));
NAND2X1 NAND2X1_11 ( .A(aNan), .B(\a[10] ), .Y(_abc_65734_new_n861_));
NAND2X1 NAND2X1_110 ( .A(aNan), .B(\a[109] ), .Y(_abc_65734_new_n1158_));
NAND2X1 NAND2X1_1100 ( .A(u2__abc_52138_new_n5500_), .B(u2__abc_52138_new_n5799_), .Y(u2__abc_52138_new_n5800_));
NAND2X1 NAND2X1_1101 ( .A(u2__abc_52138_new_n5492_), .B(u2__abc_52138_new_n5498_), .Y(u2__abc_52138_new_n5802_));
NAND2X1 NAND2X1_1102 ( .A(u2__abc_52138_new_n5801_), .B(u2__abc_52138_new_n5803_), .Y(u2__abc_52138_new_n5804_));
NAND2X1 NAND2X1_1103 ( .A(u2__abc_52138_new_n5405_), .B(u2__abc_52138_new_n5816_), .Y(u2__abc_52138_new_n5817_));
NAND2X1 NAND2X1_1104 ( .A(u2_o_314_), .B(u2__abc_52138_new_n5818_), .Y(u2__abc_52138_new_n5819_));
NAND2X1 NAND2X1_1105 ( .A(u2__abc_52138_new_n5833_), .B(u2__abc_52138_new_n5807_), .Y(u2__abc_52138_new_n5834_));
NAND2X1 NAND2X1_1106 ( .A(u2__abc_52138_new_n5339_), .B(u2__abc_52138_new_n5840_), .Y(u2__abc_52138_new_n5841_));
NAND2X1 NAND2X1_1107 ( .A(u2__abc_52138_new_n5319_), .B(u2__abc_52138_new_n5852_), .Y(u2__abc_52138_new_n5853_));
NAND2X1 NAND2X1_1108 ( .A(u2__abc_52138_new_n5198_), .B(u2__abc_52138_new_n5204_), .Y(u2__abc_52138_new_n5860_));
NAND2X1 NAND2X1_1109 ( .A(u2__abc_52138_new_n5219_), .B(u2__abc_52138_new_n5225_), .Y(u2__abc_52138_new_n5866_));
NAND2X1 NAND2X1_111 ( .A(aNan), .B(\a[110] ), .Y(_abc_65734_new_n1161_));
NAND2X1 NAND2X1_1110 ( .A(u2_o_334_), .B(u2__abc_52138_new_n5874_), .Y(u2__abc_52138_new_n5875_));
NAND2X1 NAND2X1_1111 ( .A(u2_o_369_), .B(u2__abc_52138_new_n5886_), .Y(u2__abc_52138_new_n5887_));
NAND2X1 NAND2X1_1112 ( .A(u2__abc_52138_new_n5896_), .B(u2__abc_52138_new_n5895_), .Y(u2__abc_52138_new_n5897_));
NAND2X1 NAND2X1_1113 ( .A(u2__abc_52138_new_n5907_), .B(u2__abc_52138_new_n5902_), .Y(u2__abc_52138_new_n5908_));
NAND2X1 NAND2X1_1114 ( .A(u2__abc_52138_new_n5948_), .B(u2__abc_52138_new_n5953_), .Y(u2__abc_52138_new_n5954_));
NAND2X1 NAND2X1_1115 ( .A(u2__abc_52138_new_n5959_), .B(u2__abc_52138_new_n5964_), .Y(u2__abc_52138_new_n5965_));
NAND2X1 NAND2X1_1116 ( .A(u2__abc_52138_new_n5972_), .B(u2__abc_52138_new_n5971_), .Y(u2__abc_52138_new_n5973_));
NAND2X1 NAND2X1_1117 ( .A(u2__abc_52138_new_n5978_), .B(u2__abc_52138_new_n5983_), .Y(u2__abc_52138_new_n5984_));
NAND2X1 NAND2X1_1118 ( .A(u2__abc_52138_new_n5985_), .B(u2__abc_52138_new_n5966_), .Y(u2__abc_52138_new_n5986_));
NAND2X1 NAND2X1_1119 ( .A(u2__abc_52138_new_n5991_), .B(u2__abc_52138_new_n5996_), .Y(u2__abc_52138_new_n5997_));
NAND2X1 NAND2X1_112 ( .A(aNan), .B(\a[111] ), .Y(_abc_65734_new_n1164_));
NAND2X1 NAND2X1_1120 ( .A(u2__abc_52138_new_n6002_), .B(u2__abc_52138_new_n6007_), .Y(u2__abc_52138_new_n6008_));
NAND2X1 NAND2X1_1121 ( .A(u2__abc_52138_new_n6014_), .B(u2__abc_52138_new_n6019_), .Y(u2__abc_52138_new_n6020_));
NAND2X1 NAND2X1_1122 ( .A(u2__abc_52138_new_n6025_), .B(u2__abc_52138_new_n6030_), .Y(u2__abc_52138_new_n6031_));
NAND2X1 NAND2X1_1123 ( .A(u2__abc_52138_new_n6009_), .B(u2__abc_52138_new_n6032_), .Y(u2__abc_52138_new_n6033_));
NAND2X1 NAND2X1_1124 ( .A(u2_remHi_424_), .B(u2__abc_52138_new_n6036_), .Y(u2__abc_52138_new_n6037_));
NAND2X1 NAND2X1_1125 ( .A(u2_o_424_), .B(u2__abc_52138_new_n6038_), .Y(u2__abc_52138_new_n6039_));
NAND2X1 NAND2X1_1126 ( .A(u2__abc_52138_new_n6037_), .B(u2__abc_52138_new_n6039_), .Y(u2__abc_52138_new_n6040_));
NAND2X1 NAND2X1_1127 ( .A(u2_o_425_), .B(u2__abc_52138_new_n6041_), .Y(u2__abc_52138_new_n6042_));
NAND2X1 NAND2X1_1128 ( .A(u2_remHi_425_), .B(u2__abc_52138_new_n6043_), .Y(u2__abc_52138_new_n6044_));
NAND2X1 NAND2X1_1129 ( .A(u2__abc_52138_new_n6042_), .B(u2__abc_52138_new_n6044_), .Y(u2__abc_52138_new_n6045_));
NAND2X1 NAND2X1_113 ( .A(\a[112] ), .B(\a[1] ), .Y(_abc_65734_new_n1171_));
NAND2X1 NAND2X1_1130 ( .A(u2_remHi_428_), .B(u2__abc_52138_new_n6058_), .Y(u2__abc_52138_new_n6059_));
NAND2X1 NAND2X1_1131 ( .A(u2_o_428_), .B(u2__abc_52138_new_n6060_), .Y(u2__abc_52138_new_n6061_));
NAND2X1 NAND2X1_1132 ( .A(u2__abc_52138_new_n6059_), .B(u2__abc_52138_new_n6061_), .Y(u2__abc_52138_new_n6062_));
NAND2X1 NAND2X1_1133 ( .A(u2_remHi_429_), .B(u2__abc_52138_new_n6063_), .Y(u2__abc_52138_new_n6064_));
NAND2X1 NAND2X1_1134 ( .A(u2_o_429_), .B(u2__abc_52138_new_n6065_), .Y(u2__abc_52138_new_n6066_));
NAND2X1 NAND2X1_1135 ( .A(u2__abc_52138_new_n6064_), .B(u2__abc_52138_new_n6066_), .Y(u2__abc_52138_new_n6067_));
NAND2X1 NAND2X1_1136 ( .A(u2__abc_52138_new_n6074_), .B(u2__abc_52138_new_n6079_), .Y(u2__abc_52138_new_n6080_));
NAND2X1 NAND2X1_1137 ( .A(u2_remHi_420_), .B(u2__abc_52138_new_n6084_), .Y(u2__abc_52138_new_n6085_));
NAND2X1 NAND2X1_1138 ( .A(u2_o_420_), .B(u2__abc_52138_new_n6086_), .Y(u2__abc_52138_new_n6087_));
NAND2X1 NAND2X1_1139 ( .A(u2__abc_52138_new_n6085_), .B(u2__abc_52138_new_n6087_), .Y(u2__abc_52138_new_n6088_));
NAND2X1 NAND2X1_114 ( .A(\a[1] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1174_));
NAND2X1 NAND2X1_1140 ( .A(u2_remHi_421_), .B(u2__abc_52138_new_n6089_), .Y(u2__abc_52138_new_n6090_));
NAND2X1 NAND2X1_1141 ( .A(u2_o_421_), .B(u2__abc_52138_new_n6091_), .Y(u2__abc_52138_new_n6092_));
NAND2X1 NAND2X1_1142 ( .A(u2__abc_52138_new_n6090_), .B(u2__abc_52138_new_n6092_), .Y(u2__abc_52138_new_n6093_));
NAND2X1 NAND2X1_1143 ( .A(u2__abc_52138_new_n6100_), .B(u2__abc_52138_new_n6105_), .Y(u2__abc_52138_new_n6106_));
NAND2X1 NAND2X1_1144 ( .A(u2_remHi_416_), .B(u2__abc_52138_new_n6108_), .Y(u2__abc_52138_new_n6109_));
NAND2X1 NAND2X1_1145 ( .A(u2_o_416_), .B(u2__abc_52138_new_n6110_), .Y(u2__abc_52138_new_n6111_));
NAND2X1 NAND2X1_1146 ( .A(u2__abc_52138_new_n6109_), .B(u2__abc_52138_new_n6111_), .Y(u2__abc_52138_new_n6112_));
NAND2X1 NAND2X1_1147 ( .A(u2_o_417_), .B(u2__abc_52138_new_n6113_), .Y(u2__abc_52138_new_n6114_));
NAND2X1 NAND2X1_1148 ( .A(u2_remHi_417_), .B(u2__abc_52138_new_n6115_), .Y(u2__abc_52138_new_n6116_));
NAND2X1 NAND2X1_1149 ( .A(u2__abc_52138_new_n6114_), .B(u2__abc_52138_new_n6116_), .Y(u2__abc_52138_new_n6117_));
NAND2X1 NAND2X1_115 ( .A(\a[112] ), .B(\a[3] ), .Y(_abc_65734_new_n1176_));
NAND2X1 NAND2X1_1150 ( .A(u2__abc_52138_new_n6124_), .B(u2__abc_52138_new_n6129_), .Y(u2__abc_52138_new_n6130_));
NAND2X1 NAND2X1_1151 ( .A(u2__abc_52138_new_n6107_), .B(u2__abc_52138_new_n6131_), .Y(u2__abc_52138_new_n6132_));
NAND2X1 NAND2X1_1152 ( .A(u2__abc_52138_new_n6133_), .B(u2__abc_52138_new_n6083_), .Y(u2__abc_52138_new_n6134_));
NAND2X1 NAND2X1_1153 ( .A(u2__abc_52138_new_n6140_), .B(u2__abc_52138_new_n6145_), .Y(u2__abc_52138_new_n6146_));
NAND2X1 NAND2X1_1154 ( .A(u2__abc_52138_new_n6151_), .B(u2__abc_52138_new_n6156_), .Y(u2__abc_52138_new_n6157_));
NAND2X1 NAND2X1_1155 ( .A(u2__abc_52138_new_n6164_), .B(u2__abc_52138_new_n6169_), .Y(u2__abc_52138_new_n6170_));
NAND2X1 NAND2X1_1156 ( .A(u2__abc_52138_new_n6175_), .B(u2__abc_52138_new_n6180_), .Y(u2__abc_52138_new_n6181_));
NAND2X1 NAND2X1_1157 ( .A(u2__abc_52138_new_n6189_), .B(u2__abc_52138_new_n6194_), .Y(u2__abc_52138_new_n6195_));
NAND2X1 NAND2X1_1158 ( .A(u2__abc_52138_new_n6200_), .B(u2__abc_52138_new_n6205_), .Y(u2__abc_52138_new_n6206_));
NAND2X1 NAND2X1_1159 ( .A(u2__abc_52138_new_n6212_), .B(u2__abc_52138_new_n6217_), .Y(u2__abc_52138_new_n6218_));
NAND2X1 NAND2X1_116 ( .A(\a[3] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1179_));
NAND2X1 NAND2X1_1160 ( .A(u2__abc_52138_new_n6223_), .B(u2__abc_52138_new_n6228_), .Y(u2__abc_52138_new_n6229_));
NAND2X1 NAND2X1_1161 ( .A(u2__abc_52138_new_n6207_), .B(u2__abc_52138_new_n6230_), .Y(u2__abc_52138_new_n6231_));
NAND2X1 NAND2X1_1162 ( .A(u2__abc_52138_new_n6236_), .B(u2__abc_52138_new_n6241_), .Y(u2__abc_52138_new_n6242_));
NAND2X1 NAND2X1_1163 ( .A(u2__abc_52138_new_n6247_), .B(u2__abc_52138_new_n6252_), .Y(u2__abc_52138_new_n6253_));
NAND2X1 NAND2X1_1164 ( .A(u2__abc_52138_new_n6259_), .B(u2__abc_52138_new_n6264_), .Y(u2__abc_52138_new_n6265_));
NAND2X1 NAND2X1_1165 ( .A(u2__abc_52138_new_n6270_), .B(u2__abc_52138_new_n6275_), .Y(u2__abc_52138_new_n6276_));
NAND2X1 NAND2X1_1166 ( .A(u2__abc_52138_new_n6254_), .B(u2__abc_52138_new_n6277_), .Y(u2__abc_52138_new_n6278_));
NAND2X1 NAND2X1_1167 ( .A(u2_remHi_393_), .B(u2__abc_52138_new_n6285_), .Y(u2__abc_52138_new_n6288_));
NAND2X1 NAND2X1_1168 ( .A(u2__abc_52138_new_n6288_), .B(u2__abc_52138_new_n6287_), .Y(u2__abc_52138_new_n6289_));
NAND2X1 NAND2X1_1169 ( .A(u2__abc_52138_new_n6284_), .B(u2__abc_52138_new_n6290_), .Y(u2__abc_52138_new_n6291_));
NAND2X1 NAND2X1_117 ( .A(\a[112] ), .B(\a[5] ), .Y(_abc_65734_new_n1181_));
NAND2X1 NAND2X1_1170 ( .A(u2_o_390_), .B(u2__abc_52138_new_n6292_), .Y(u2__abc_52138_new_n6294_));
NAND2X1 NAND2X1_1171 ( .A(u2_o_391_), .B(u2__abc_52138_new_n6297_), .Y(u2__abc_52138_new_n6298_));
NAND2X1 NAND2X1_1172 ( .A(u2__abc_52138_new_n6301_), .B(u2__abc_52138_new_n6296_), .Y(u2__abc_52138_new_n6302_));
NAND2X1 NAND2X1_1173 ( .A(u2__abc_52138_new_n6308_), .B(u2__abc_52138_new_n6313_), .Y(u2__abc_52138_new_n6314_));
NAND2X1 NAND2X1_1174 ( .A(u2_o_394_), .B(u2__abc_52138_new_n6320_), .Y(u2__abc_52138_new_n6323_));
NAND2X1 NAND2X1_1175 ( .A(u2__abc_52138_new_n6319_), .B(u2__abc_52138_new_n6324_), .Y(u2__abc_52138_new_n6325_));
NAND2X1 NAND2X1_1176 ( .A(u2__abc_52138_new_n6326_), .B(u2__abc_52138_new_n6303_), .Y(u2__abc_52138_new_n6327_));
NAND2X1 NAND2X1_1177 ( .A(u2__abc_52138_new_n6279_), .B(u2__abc_52138_new_n6328_), .Y(u2__abc_52138_new_n6329_));
NAND2X1 NAND2X1_1178 ( .A(u2__abc_52138_new_n6135_), .B(u2__abc_52138_new_n6331_), .Y(u2__abc_52138_new_n6332_));
NAND2X1 NAND2X1_1179 ( .A(u2__abc_52138_new_n6347_), .B(u2__abc_52138_new_n6345_), .Y(u2__abc_52138_new_n6348_));
NAND2X1 NAND2X1_118 ( .A(\a[5] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1184_));
NAND2X1 NAND2X1_1180 ( .A(u2__abc_52138_new_n6230_), .B(u2__abc_52138_new_n6362_), .Y(u2__abc_52138_new_n6363_));
NAND2X1 NAND2X1_1181 ( .A(u2__abc_52138_new_n6371_), .B(u2__abc_52138_new_n6363_), .Y(u2__abc_52138_new_n6372_));
NAND2X1 NAND2X1_1182 ( .A(u2__abc_52138_new_n6410_), .B(u2__abc_52138_new_n6405_), .Y(u2__abc_52138_new_n6411_));
NAND2X1 NAND2X1_1183 ( .A(u2__abc_52138_new_n6438_), .B(u2__abc_52138_new_n6412_), .Y(u2__abc_52138_new_n6439_));
NAND2X1 NAND2X1_1184 ( .A(u2__abc_52138_new_n3015_), .B(u2__abc_52138_new_n6441_), .Y(u2__abc_52138_new_n6442_));
NAND2X1 NAND2X1_1185 ( .A(u2_remHiShift_0_), .B(u2__abc_52138_new_n6455_), .Y(u2__abc_52138_new_n6456_));
NAND2X1 NAND2X1_1186 ( .A(u2_remHi_4_), .B(u2__abc_52138_new_n6458_), .Y(u2__abc_52138_new_n6459_));
NAND2X1 NAND2X1_1187 ( .A(u2__abc_52138_new_n6459_), .B(u2__abc_52138_new_n3087_), .Y(u2__abc_52138_new_n6460_));
NAND2X1 NAND2X1_1188 ( .A(u2__abc_52138_new_n3055_), .B(u2__abc_52138_new_n3057_), .Y(u2__abc_52138_new_n6461_));
NAND2X1 NAND2X1_1189 ( .A(u2__abc_52138_new_n3080_), .B(u2__abc_52138_new_n3082_), .Y(u2__abc_52138_new_n6463_));
NAND2X1 NAND2X1_119 ( .A(\a[112] ), .B(\a[7] ), .Y(_abc_65734_new_n1186_));
NAND2X1 NAND2X1_1190 ( .A(u2__abc_52138_new_n3061_), .B(u2__abc_52138_new_n3063_), .Y(u2__abc_52138_new_n6464_));
NAND2X1 NAND2X1_1191 ( .A(u2__abc_52138_new_n6462_), .B(u2__abc_52138_new_n6465_), .Y(u2__abc_52138_new_n6466_));
NAND2X1 NAND2X1_1192 ( .A(u2__abc_52138_new_n4341_), .B(u2__abc_52138_new_n4352_), .Y(u2__abc_52138_new_n6467_));
NAND2X1 NAND2X1_1193 ( .A(u2__abc_52138_new_n6034_), .B(u2__abc_52138_new_n6473_), .Y(u2__abc_52138_new_n6474_));
NAND2X1 NAND2X1_1194 ( .A(u2__abc_52138_new_n4758_), .B(u2__abc_52138_new_n5090_), .Y(u2__abc_52138_new_n6475_));
NAND2X1 NAND2X1_1195 ( .A(u2__abc_52138_new_n6184_), .B(u2__abc_52138_new_n6083_), .Y(u2__abc_52138_new_n6480_));
NAND2X1 NAND2X1_1196 ( .A(u2__abc_52138_new_n3526_), .B(u2__abc_52138_new_n3515_), .Y(u2__abc_52138_new_n6487_));
NAND2X1 NAND2X1_1197 ( .A(u2__abc_52138_new_n6511_), .B(u2__abc_52138_new_n6456_), .Y(u2__abc_52138_new_n6512_));
NAND2X1 NAND2X1_1198 ( .A(u2_remHiShift_1_), .B(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n6513_));
NAND2X1 NAND2X1_1199 ( .A(u2__abc_52138_new_n3066_), .B(u2__abc_52138_new_n6520_), .Y(u2__abc_52138_new_n6521_));
NAND2X1 NAND2X1_12 ( .A(aNan), .B(\a[11] ), .Y(_abc_65734_new_n864_));
NAND2X1 NAND2X1_120 ( .A(\a[7] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1189_));
NAND2X1 NAND2X1_1200 ( .A(u2__abc_52138_new_n3067_), .B(u2__abc_52138_new_n6529_), .Y(u2__abc_52138_new_n6531_));
NAND2X1 NAND2X1_1201 ( .A(u2__abc_52138_new_n6497_), .B(u2__abc_52138_new_n6479_), .Y(u2__abc_52138_new_n6540_));
NAND2X1 NAND2X1_1202 ( .A(u2__abc_52138_new_n6599_), .B(u2__abc_52138_new_n6604_), .Y(u2__abc_52138_new_n6605_));
NAND2X1 NAND2X1_1203 ( .A(u2__abc_52138_new_n3036_), .B(u2__abc_52138_new_n3038_), .Y(u2__abc_52138_new_n6614_));
NAND2X1 NAND2X1_1204 ( .A(u2_remHi_8_), .B(u2__abc_52138_new_n3096_), .Y(u2__abc_52138_new_n6615_));
NAND2X1 NAND2X1_1205 ( .A(u2__abc_52138_new_n3031_), .B(u2__abc_52138_new_n6626_), .Y(u2__abc_52138_new_n6628_));
NAND2X1 NAND2X1_1206 ( .A(u2__abc_52138_new_n3018_), .B(u2__abc_52138_new_n3020_), .Y(u2__abc_52138_new_n6653_));
NAND2X1 NAND2X1_1207 ( .A(u2_remHi_12_), .B(u2__abc_52138_new_n6654_), .Y(u2__abc_52138_new_n6655_));
NAND2X1 NAND2X1_1208 ( .A(u2__abc_52138_new_n6665_), .B(u2__abc_52138_new_n3033_), .Y(u2__abc_52138_new_n6666_));
NAND2X1 NAND2X1_1209 ( .A(u2__abc_52138_new_n6655_), .B(u2__abc_52138_new_n3102_), .Y(u2__abc_52138_new_n6667_));
NAND2X1 NAND2X1_121 ( .A(\a[112] ), .B(\a[9] ), .Y(_abc_65734_new_n1191_));
NAND2X1 NAND2X1_1210 ( .A(u2__abc_52138_new_n3190_), .B(u2__abc_52138_new_n3192_), .Y(u2__abc_52138_new_n6711_));
NAND2X1 NAND2X1_1211 ( .A(u2__abc_52138_new_n6711_), .B(u2__abc_52138_new_n6716_), .Y(u2__abc_52138_new_n6717_));
NAND2X1 NAND2X1_1212 ( .A(u2_remHi_20_), .B(u2__abc_52138_new_n6733_), .Y(u2__abc_52138_new_n6734_));
NAND2X1 NAND2X1_1213 ( .A(u2__abc_52138_new_n6734_), .B(u2__abc_52138_new_n3212_), .Y(u2__abc_52138_new_n6735_));
NAND2X1 NAND2X1_1214 ( .A(u2__abc_52138_new_n6735_), .B(u2__abc_52138_new_n6738_), .Y(u2__abc_52138_new_n6739_));
NAND2X1 NAND2X1_1215 ( .A(u2__abc_52138_new_n3184_), .B(u2__abc_52138_new_n3186_), .Y(u2__abc_52138_new_n6747_));
NAND2X1 NAND2X1_1216 ( .A(u2__abc_52138_new_n3194_), .B(u2__abc_52138_new_n6715_), .Y(u2__abc_52138_new_n6757_));
NAND2X1 NAND2X1_1217 ( .A(u2__abc_52138_new_n6737_), .B(u2__abc_52138_new_n6758_), .Y(u2__abc_52138_new_n6759_));
NAND2X1 NAND2X1_1218 ( .A(u2__abc_52138_new_n3132_), .B(u2__abc_52138_new_n6763_), .Y(u2__abc_52138_new_n6764_));
NAND2X1 NAND2X1_1219 ( .A(u2__abc_52138_new_n6782_), .B(u2__abc_52138_new_n6783_), .Y(u2__abc_52138_new_n6784_));
NAND2X1 NAND2X1_122 ( .A(\a[9] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1194_));
NAND2X1 NAND2X1_1220 ( .A(u2__abc_52138_new_n3219_), .B(u2__abc_52138_new_n6784_), .Y(u2__abc_52138_new_n6786_));
NAND2X1 NAND2X1_1221 ( .A(u2__abc_52138_new_n3155_), .B(u2__abc_52138_new_n6806_), .Y(u2__abc_52138_new_n6807_));
NAND2X1 NAND2X1_1222 ( .A(u2__abc_52138_new_n3432_), .B(u2__abc_52138_new_n6863_), .Y(u2__abc_52138_new_n6865_));
NAND2X1 NAND2X1_1223 ( .A(u2_remHi_32_), .B(u2__abc_52138_new_n3437_), .Y(u2__abc_52138_new_n6882_));
NAND2X1 NAND2X1_1224 ( .A(u2__abc_52138_new_n3417_), .B(u2__abc_52138_new_n6885_), .Y(u2__abc_52138_new_n6887_));
NAND2X1 NAND2X1_1225 ( .A(u2__abc_52138_new_n3413_), .B(u2__abc_52138_new_n3415_), .Y(u2__abc_52138_new_n6895_));
NAND2X1 NAND2X1_1226 ( .A(u2__abc_52138_new_n3419_), .B(u2__abc_52138_new_n6844_), .Y(u2__abc_52138_new_n6928_));
NAND2X1 NAND2X1_1227 ( .A(u2__abc_52138_new_n6927_), .B(u2__abc_52138_new_n6928_), .Y(u2__abc_52138_new_n6929_));
NAND2X1 NAND2X1_1228 ( .A(u2__abc_52138_new_n6923_), .B(u2__abc_52138_new_n6929_), .Y(u2__abc_52138_new_n6931_));
NAND2X1 NAND2X1_1229 ( .A(u2__abc_52138_new_n3378_), .B(u2__abc_52138_new_n6971_), .Y(u2__abc_52138_new_n6972_));
NAND2X1 NAND2X1_123 ( .A(\a[112] ), .B(\a[11] ), .Y(_abc_65734_new_n1196_));
NAND2X1 NAND2X1_1230 ( .A(u2_remHi_48_), .B(u2__abc_52138_new_n3289_), .Y(u2__abc_52138_new_n7034_));
NAND2X1 NAND2X1_1231 ( .A(u2__abc_52138_new_n7034_), .B(u2__abc_52138_new_n3472_), .Y(u2__abc_52138_new_n7035_));
NAND2X1 NAND2X1_1232 ( .A(u2_remHi_49_), .B(u2__abc_52138_new_n3294_), .Y(u2__abc_52138_new_n7052_));
NAND2X1 NAND2X1_1233 ( .A(u2__abc_52138_new_n3331_), .B(u2__abc_52138_new_n7056_), .Y(u2__abc_52138_new_n7057_));
NAND2X1 NAND2X1_1234 ( .A(u2__abc_52138_new_n3321_), .B(u2__abc_52138_new_n3332_), .Y(u2__abc_52138_new_n7093_));
NAND2X1 NAND2X1_1235 ( .A(u2__abc_52138_new_n3255_), .B(u2__abc_52138_new_n7100_), .Y(u2__abc_52138_new_n7101_));
NAND2X1 NAND2X1_1236 ( .A(u2__abc_52138_new_n7135_), .B(u2__abc_52138_new_n7139_), .Y(u2__abc_52138_new_n7140_));
NAND2X1 NAND2X1_1237 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7144_), .Y(u2__abc_52138_new_n7145_));
NAND2X1 NAND2X1_1238 ( .A(u2__abc_52138_new_n7146_), .B(u2__abc_52138_new_n7145_), .Y(u2__abc_52138_new_n7147_));
NAND2X1 NAND2X1_1239 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7154_), .Y(u2__abc_52138_new_n7155_));
NAND2X1 NAND2X1_124 ( .A(\a[11] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1199_));
NAND2X1 NAND2X1_1240 ( .A(u2__abc_52138_new_n7156_), .B(u2__abc_52138_new_n7155_), .Y(u2__abc_52138_new_n7157_));
NAND2X1 NAND2X1_1241 ( .A(u2__abc_52138_new_n3836_), .B(u2__abc_52138_new_n7186_), .Y(u2__abc_52138_new_n7187_));
NAND2X1 NAND2X1_1242 ( .A(u2__abc_52138_new_n3863_), .B(u2__abc_52138_new_n3865_), .Y(u2__abc_52138_new_n7222_));
NAND2X1 NAND2X1_1243 ( .A(u2__abc_52138_new_n3861_), .B(u2__abc_52138_new_n7235_), .Y(u2__abc_52138_new_n7243_));
NAND2X1 NAND2X1_1244 ( .A(u2__abc_52138_new_n3857_), .B(u2__abc_52138_new_n3859_), .Y(u2__abc_52138_new_n7252_));
NAND2X1 NAND2X1_1245 ( .A(u2__abc_52138_new_n3855_), .B(u2__abc_52138_new_n7244_), .Y(u2__abc_52138_new_n7253_));
NAND2X1 NAND2X1_1246 ( .A(u2_remHi_68_), .B(u2__abc_52138_new_n7264_), .Y(u2__abc_52138_new_n7265_));
NAND2X1 NAND2X1_1247 ( .A(u2__abc_52138_new_n3790_), .B(u2__abc_52138_new_n7270_), .Y(u2__abc_52138_new_n7273_));
NAND2X1 NAND2X1_1248 ( .A(u2__abc_52138_new_n3803_), .B(u2__abc_52138_new_n3805_), .Y(u2__abc_52138_new_n7298_));
NAND2X1 NAND2X1_1249 ( .A(u2__abc_52138_new_n3801_), .B(u2__abc_52138_new_n7290_), .Y(u2__abc_52138_new_n7299_));
NAND2X1 NAND2X1_125 ( .A(\a[112] ), .B(\a[13] ), .Y(_abc_65734_new_n1201_));
NAND2X1 NAND2X1_1250 ( .A(u2__abc_52138_new_n3798_), .B(u2__abc_52138_new_n3800_), .Y(u2__abc_52138_new_n7308_));
NAND2X1 NAND2X1_1251 ( .A(u2__abc_52138_new_n3828_), .B(u2__abc_52138_new_n7314_), .Y(u2__abc_52138_new_n7315_));
NAND2X1 NAND2X1_1252 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7319_), .Y(u2__abc_52138_new_n7320_));
NAND2X1 NAND2X1_1253 ( .A(u2__abc_52138_new_n7321_), .B(u2__abc_52138_new_n7320_), .Y(u2__abc_52138_new_n7322_));
NAND2X1 NAND2X1_1254 ( .A(sqrto_77_), .B(u2__abc_52138_new_n3813_), .Y(u2__abc_52138_new_n7352_));
NAND2X1 NAND2X1_1255 ( .A(u2__abc_52138_new_n3903_), .B(u2__abc_52138_new_n7352_), .Y(u2__abc_52138_new_n7353_));
NAND2X1 NAND2X1_1256 ( .A(u2__abc_52138_new_n3753_), .B(u2__abc_52138_new_n7382_), .Y(u2__abc_52138_new_n7390_));
NAND2X1 NAND2X1_1257 ( .A(u2__abc_52138_new_n3750_), .B(u2__abc_52138_new_n3752_), .Y(u2__abc_52138_new_n7401_));
NAND2X1 NAND2X1_1258 ( .A(u2__abc_52138_new_n3755_), .B(u2__abc_52138_new_n3757_), .Y(u2__abc_52138_new_n7402_));
NAND2X1 NAND2X1_1259 ( .A(u2__abc_52138_new_n7399_), .B(u2__abc_52138_new_n7406_), .Y(u2__abc_52138_new_n7407_));
NAND2X1 NAND2X1_126 ( .A(\a[13] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1204_));
NAND2X1 NAND2X1_1260 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7411_), .Y(u2__abc_52138_new_n7412_));
NAND2X1 NAND2X1_1261 ( .A(u2__abc_52138_new_n7413_), .B(u2__abc_52138_new_n7412_), .Y(u2__abc_52138_new_n7414_));
NAND2X1 NAND2X1_1262 ( .A(u2__abc_52138_new_n3765_), .B(u2__abc_52138_new_n7426_), .Y(u2__abc_52138_new_n7428_));
NAND2X1 NAND2X1_1263 ( .A(u2__abc_52138_new_n3771_), .B(u2__abc_52138_new_n3782_), .Y(u2__abc_52138_new_n7447_));
NAND2X1 NAND2X1_1264 ( .A(u2__abc_52138_new_n3734_), .B(u2__abc_52138_new_n7451_), .Y(u2__abc_52138_new_n7452_));
NAND2X1 NAND2X1_1265 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7456_), .Y(u2__abc_52138_new_n7457_));
NAND2X1 NAND2X1_1266 ( .A(u2__abc_52138_new_n7458_), .B(u2__abc_52138_new_n7457_), .Y(u2__abc_52138_new_n7459_));
NAND2X1 NAND2X1_1267 ( .A(u2__abc_52138_new_n3726_), .B(u2__abc_52138_new_n3729_), .Y(u2__abc_52138_new_n7462_));
NAND2X1 NAND2X1_1268 ( .A(u2__abc_52138_new_n7472_), .B(u2__abc_52138_new_n7473_), .Y(u2__abc_52138_new_n7474_));
NAND2X1 NAND2X1_1269 ( .A(u2__abc_52138_new_n3703_), .B(u2__abc_52138_new_n3705_), .Y(u2__abc_52138_new_n7503_));
NAND2X1 NAND2X1_127 ( .A(\a[112] ), .B(\a[15] ), .Y(_abc_65734_new_n1206_));
NAND2X1 NAND2X1_1270 ( .A(u2__abc_52138_new_n3785_), .B(u2__abc_52138_new_n7362_), .Y(u2__abc_52138_new_n7531_));
NAND2X1 NAND2X1_1271 ( .A(u2__abc_52138_new_n3662_), .B(u2__abc_52138_new_n7541_), .Y(u2__abc_52138_new_n7542_));
NAND2X1 NAND2X1_1272 ( .A(u2_remHi_97_), .B(u2__abc_52138_new_n3649_), .Y(u2__abc_52138_new_n7569_));
NAND2X1 NAND2X1_1273 ( .A(u2__abc_52138_new_n7569_), .B(u2__abc_52138_new_n3943_), .Y(u2__abc_52138_new_n7570_));
NAND2X1 NAND2X1_1274 ( .A(u2_remHi_96_), .B(u2__abc_52138_new_n3644_), .Y(u2__abc_52138_new_n7580_));
NAND2X1 NAND2X1_1275 ( .A(u2__abc_52138_new_n7584_), .B(u2__abc_52138_new_n7585_), .Y(u2__abc_52138_new_n7586_));
NAND2X1 NAND2X1_1276 ( .A(u2__abc_52138_new_n7579_), .B(u2__abc_52138_new_n7586_), .Y(u2__abc_52138_new_n7587_));
NAND2X1 NAND2X1_1277 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7591_), .Y(u2__abc_52138_new_n7592_));
NAND2X1 NAND2X1_1278 ( .A(u2__abc_52138_new_n7593_), .B(u2__abc_52138_new_n7592_), .Y(u2__abc_52138_new_n7594_));
NAND2X1 NAND2X1_1279 ( .A(u2__abc_52138_new_n3669_), .B(u2__abc_52138_new_n7606_), .Y(u2__abc_52138_new_n7608_));
NAND2X1 NAND2X1_128 ( .A(\a[15] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1209_));
NAND2X1 NAND2X1_1280 ( .A(u2__abc_52138_new_n3675_), .B(u2__abc_52138_new_n3686_), .Y(u2__abc_52138_new_n7625_));
NAND2X1 NAND2X1_1281 ( .A(u2__abc_52138_new_n3616_), .B(u2__abc_52138_new_n7631_), .Y(u2__abc_52138_new_n7632_));
NAND2X1 NAND2X1_1282 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7636_), .Y(u2__abc_52138_new_n7637_));
NAND2X1 NAND2X1_1283 ( .A(u2__abc_52138_new_n7638_), .B(u2__abc_52138_new_n7637_), .Y(u2__abc_52138_new_n7639_));
NAND2X1 NAND2X1_1284 ( .A(u2__abc_52138_new_n3609_), .B(u2__abc_52138_new_n3611_), .Y(u2__abc_52138_new_n7642_));
NAND2X1 NAND2X1_1285 ( .A(u2__abc_52138_new_n3601_), .B(u2__abc_52138_new_n7652_), .Y(u2__abc_52138_new_n7654_));
NAND2X1 NAND2X1_1286 ( .A(u2__abc_52138_new_n7719_), .B(u2__abc_52138_new_n7720_), .Y(u2__abc_52138_new_n7721_));
NAND2X1 NAND2X1_1287 ( .A(u2__abc_52138_new_n3565_), .B(u2__abc_52138_new_n7739_), .Y(u2__abc_52138_new_n7741_));
NAND2X1 NAND2X1_1288 ( .A(u2__abc_52138_new_n3592_), .B(u2__abc_52138_new_n7761_), .Y(u2__abc_52138_new_n7763_));
NAND2X1 NAND2X1_1289 ( .A(u2__abc_52138_new_n7771_), .B(u2__abc_52138_new_n7772_), .Y(u2__abc_52138_new_n7781_));
NAND2X1 NAND2X1_129 ( .A(\a[112] ), .B(\a[17] ), .Y(_abc_65734_new_n1211_));
NAND2X1 NAND2X1_1290 ( .A(u2__abc_52138_new_n3577_), .B(u2__abc_52138_new_n7782_), .Y(u2__abc_52138_new_n7783_));
NAND2X1 NAND2X1_1291 ( .A(u2__abc_52138_new_n3579_), .B(u2__abc_52138_new_n3581_), .Y(u2__abc_52138_new_n7792_));
NAND2X1 NAND2X1_1292 ( .A(u2__abc_52138_new_n3594_), .B(u2__abc_52138_new_n7760_), .Y(u2__abc_52138_new_n7801_));
NAND2X1 NAND2X1_1293 ( .A(u2__abc_52138_new_n7804_), .B(u2__abc_52138_new_n7803_), .Y(u2__abc_52138_new_n7805_));
NAND2X1 NAND2X1_1294 ( .A(u2__abc_52138_new_n7830_), .B(u2__abc_52138_new_n7831_), .Y(u2__abc_52138_new_n7832_));
NAND2X1 NAND2X1_1295 ( .A(u2__abc_52138_new_n7828_), .B(u2__abc_52138_new_n7832_), .Y(u2__abc_52138_new_n7840_));
NAND2X1 NAND2X1_1296 ( .A(u2__abc_52138_new_n3546_), .B(u2__abc_52138_new_n7851_), .Y(u2__abc_52138_new_n7852_));
NAND2X1 NAND2X1_1297 ( .A(u2__abc_52138_new_n3539_), .B(u2__abc_52138_new_n3541_), .Y(u2__abc_52138_new_n7862_));
NAND2X1 NAND2X1_1298 ( .A(u2__abc_52138_new_n6483_), .B(u2__abc_52138_new_n6489_), .Y(u2__abc_52138_new_n7893_));
NAND2X1 NAND2X1_1299 ( .A(u2__abc_52138_new_n7891_), .B(u2__abc_52138_new_n7898_), .Y(u2__abc_52138_new_n7899_));
NAND2X1 NAND2X1_13 ( .A(aNan), .B(\a[12] ), .Y(_abc_65734_new_n867_));
NAND2X1 NAND2X1_130 ( .A(\a[17] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1214_));
NAND2X1 NAND2X1_1300 ( .A(u2__abc_52138_new_n4717_), .B(u2__abc_52138_new_n7901_), .Y(u2__abc_52138_new_n7902_));
NAND2X1 NAND2X1_1301 ( .A(u2__abc_52138_new_n4728_), .B(u2__abc_52138_new_n4730_), .Y(u2__abc_52138_new_n7928_));
NAND2X1 NAND2X1_1302 ( .A(u2__abc_52138_new_n4726_), .B(u2__abc_52138_new_n7920_), .Y(u2__abc_52138_new_n7929_));
NAND2X1 NAND2X1_1303 ( .A(u2_remHi_128_), .B(u2__abc_52138_new_n4770_), .Y(u2__abc_52138_new_n7940_));
NAND2X1 NAND2X1_1304 ( .A(u2__abc_52138_new_n4749_), .B(u2__abc_52138_new_n7943_), .Y(u2__abc_52138_new_n7944_));
NAND2X1 NAND2X1_1305 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7948_), .Y(u2__abc_52138_new_n7949_));
NAND2X1 NAND2X1_1306 ( .A(u2__abc_52138_new_n7950_), .B(u2__abc_52138_new_n7949_), .Y(u2__abc_52138_new_n7951_));
NAND2X1 NAND2X1_1307 ( .A(u2__abc_52138_new_n4737_), .B(u2__abc_52138_new_n7963_), .Y(u2__abc_52138_new_n7965_));
NAND2X1 NAND2X1_1308 ( .A(u2__abc_52138_new_n7981_), .B(u2__abc_52138_new_n7988_), .Y(u2__abc_52138_new_n7989_));
NAND2X1 NAND2X1_1309 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n7993_), .Y(u2__abc_52138_new_n7994_));
NAND2X1 NAND2X1_131 ( .A(\a[112] ), .B(\a[19] ), .Y(_abc_65734_new_n1216_));
NAND2X1 NAND2X1_1310 ( .A(u2__abc_52138_new_n7995_), .B(u2__abc_52138_new_n7994_), .Y(u2__abc_52138_new_n7996_));
NAND2X1 NAND2X1_1311 ( .A(u2__abc_52138_new_n4709_), .B(u2__abc_52138_new_n8034_), .Y(u2__abc_52138_new_n8036_));
NAND2X1 NAND2X1_1312 ( .A(u2__abc_52138_new_n4676_), .B(u2__abc_52138_new_n4687_), .Y(u2__abc_52138_new_n8069_));
NAND2X1 NAND2X1_1313 ( .A(u2__abc_52138_new_n4699_), .B(u2__abc_52138_new_n4710_), .Y(u2__abc_52138_new_n8070_));
NAND2X1 NAND2X1_1314 ( .A(u2__abc_52138_new_n4711_), .B(u2__abc_52138_new_n8033_), .Y(u2__abc_52138_new_n8073_));
NAND2X1 NAND2X1_1315 ( .A(u2__abc_52138_new_n8076_), .B(u2__abc_52138_new_n8073_), .Y(u2__abc_52138_new_n8077_));
NAND2X1 NAND2X1_1316 ( .A(u2__abc_52138_new_n8078_), .B(u2__abc_52138_new_n8080_), .Y(u2__abc_52138_new_n8081_));
NAND2X1 NAND2X1_1317 ( .A(u2__abc_52138_new_n4662_), .B(u2__abc_52138_new_n8081_), .Y(u2__abc_52138_new_n8082_));
NAND2X1 NAND2X1_1318 ( .A(u2__abc_52138_new_n2978_), .B(u2__abc_52138_new_n8086_), .Y(u2__abc_52138_new_n8087_));
NAND2X1 NAND2X1_1319 ( .A(u2__abc_52138_new_n8088_), .B(u2__abc_52138_new_n8087_), .Y(u2__abc_52138_new_n8089_));
NAND2X1 NAND2X1_132 ( .A(\a[19] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1219_));
NAND2X1 NAND2X1_1320 ( .A(u2__abc_52138_new_n4643_), .B(u2__abc_52138_new_n4645_), .Y(u2__abc_52138_new_n8101_));
NAND2X1 NAND2X1_1321 ( .A(u2__abc_52138_new_n8101_), .B(u2__abc_52138_new_n8102_), .Y(u2__abc_52138_new_n8104_));
NAND2X1 NAND2X1_1322 ( .A(u2__abc_52138_new_n4648_), .B(u2__abc_52138_new_n4650_), .Y(u2__abc_52138_new_n8112_));
NAND2X1 NAND2X1_1323 ( .A(u2__abc_52138_new_n4639_), .B(u2__abc_52138_new_n8122_), .Y(u2__abc_52138_new_n8124_));
NAND2X1 NAND2X1_1324 ( .A(u2__abc_52138_new_n8132_), .B(u2__abc_52138_new_n8133_), .Y(u2__abc_52138_new_n8143_));
NAND2X1 NAND2X1_1325 ( .A(u2__abc_52138_new_n8142_), .B(u2__abc_52138_new_n8144_), .Y(u2__abc_52138_new_n8145_));
NAND2X1 NAND2X1_1326 ( .A(u2__abc_52138_new_n8164_), .B(u2__abc_52138_new_n8169_), .Y(u2__abc_52138_new_n8170_));
NAND2X1 NAND2X1_1327 ( .A(u2__abc_52138_new_n4593_), .B(u2__abc_52138_new_n8173_), .Y(u2__abc_52138_new_n8174_));
NAND2X1 NAND2X1_1328 ( .A(u2__abc_52138_new_n4616_), .B(u2__abc_52138_new_n8210_), .Y(u2__abc_52138_new_n8211_));
NAND2X1 NAND2X1_1329 ( .A(u2__abc_52138_new_n8254_), .B(u2__abc_52138_new_n8255_), .Y(u2__abc_52138_new_n8256_));
NAND2X1 NAND2X1_133 ( .A(\a[112] ), .B(\a[21] ), .Y(_abc_65734_new_n1221_));
NAND2X1 NAND2X1_1330 ( .A(u2__abc_52138_new_n8260_), .B(u2__abc_52138_new_n8259_), .Y(u2__abc_52138_new_n8261_));
NAND2X1 NAND2X1_1331 ( .A(u2__abc_52138_new_n4568_), .B(u2__abc_52138_new_n8302_), .Y(u2__abc_52138_new_n8305_));
NAND2X1 NAND2X1_1332 ( .A(u2__abc_52138_new_n4505_), .B(u2__abc_52138_new_n8364_), .Y(u2__abc_52138_new_n8366_));
NAND2X1 NAND2X1_1333 ( .A(u2__abc_52138_new_n8448_), .B(u2__abc_52138_new_n8453_), .Y(u2__abc_52138_new_n8454_));
NAND2X1 NAND2X1_1334 ( .A(u2__abc_52138_new_n8513_), .B(u2__abc_52138_new_n8514_), .Y(u2__abc_52138_new_n8515_));
NAND2X1 NAND2X1_1335 ( .A(u2__abc_52138_new_n4392_), .B(u2__abc_52138_new_n8515_), .Y(u2__abc_52138_new_n8534_));
NAND2X1 NAND2X1_1336 ( .A(u2__abc_52138_new_n8533_), .B(u2__abc_52138_new_n8534_), .Y(u2__abc_52138_new_n8535_));
NAND2X1 NAND2X1_1337 ( .A(u2__abc_52138_new_n4425_), .B(u2__abc_52138_new_n8555_), .Y(u2__abc_52138_new_n8557_));
NAND2X1 NAND2X1_1338 ( .A(u2__abc_52138_new_n4572_), .B(u2__abc_52138_new_n4752_), .Y(u2__abc_52138_new_n8590_));
NAND2X1 NAND2X1_1339 ( .A(u2__abc_52138_new_n8607_), .B(u2__abc_52138_new_n8606_), .Y(u2__abc_52138_new_n8608_));
NAND2X1 NAND2X1_134 ( .A(\a[21] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1224_));
NAND2X1 NAND2X1_1340 ( .A(u2__abc_52138_new_n4880_), .B(u2__abc_52138_new_n8624_), .Y(u2__abc_52138_new_n8625_));
NAND2X1 NAND2X1_1341 ( .A(u2__abc_52138_new_n4351_), .B(u2__abc_52138_new_n8644_), .Y(u2__abc_52138_new_n8646_));
NAND2X1 NAND2X1_1342 ( .A(u2__abc_52138_new_n8654_), .B(u2__abc_52138_new_n8655_), .Y(u2__abc_52138_new_n8666_));
NAND2X1 NAND2X1_1343 ( .A(u2__abc_52138_new_n8665_), .B(u2__abc_52138_new_n8667_), .Y(u2__abc_52138_new_n8668_));
NAND2X1 NAND2X1_1344 ( .A(u2__abc_52138_new_n4353_), .B(u2__abc_52138_new_n8643_), .Y(u2__abc_52138_new_n8686_));
NAND2X1 NAND2X1_1345 ( .A(u2__abc_52138_new_n4341_), .B(u2__abc_52138_new_n8687_), .Y(u2__abc_52138_new_n8688_));
NAND2X1 NAND2X1_1346 ( .A(u2__abc_52138_new_n4309_), .B(u2__abc_52138_new_n8693_), .Y(u2__abc_52138_new_n8694_));
NAND2X1 NAND2X1_1347 ( .A(u2__abc_52138_new_n4328_), .B(u2__abc_52138_new_n8730_), .Y(u2__abc_52138_new_n8731_));
NAND2X1 NAND2X1_1348 ( .A(u2__abc_52138_new_n8768_), .B(u2__abc_52138_new_n8690_), .Y(u2__abc_52138_new_n8769_));
NAND2X1 NAND2X1_1349 ( .A(u2__abc_52138_new_n8814_), .B(u2__abc_52138_new_n8815_), .Y(u2__abc_52138_new_n8816_));
NAND2X1 NAND2X1_135 ( .A(\a[112] ), .B(\a[23] ), .Y(_abc_65734_new_n1226_));
NAND2X1 NAND2X1_1350 ( .A(u2__abc_52138_new_n4284_), .B(u2__abc_52138_new_n8816_), .Y(u2__abc_52138_new_n8817_));
NAND2X1 NAND2X1_1351 ( .A(u2__abc_52138_new_n4279_), .B(u2__abc_52138_new_n8826_), .Y(u2__abc_52138_new_n8834_));
NAND2X1 NAND2X1_1352 ( .A(u2__abc_52138_new_n4288_), .B(u2__abc_52138_new_n8774_), .Y(u2__abc_52138_new_n8936_));
NAND2X1 NAND2X1_1353 ( .A(u2__abc_52138_new_n4189_), .B(u2__abc_52138_new_n8982_), .Y(u2__abc_52138_new_n8983_));
NAND2X1 NAND2X1_1354 ( .A(u2__abc_52138_new_n4142_), .B(u2__abc_52138_new_n9024_), .Y(u2__abc_52138_new_n9025_));
NAND2X1 NAND2X1_1355 ( .A(u2__abc_52138_new_n4137_), .B(u2__abc_52138_new_n4136_), .Y(u2__abc_52138_new_n9034_));
NAND2X1 NAND2X1_1356 ( .A(u2__abc_52138_new_n4127_), .B(u2__abc_52138_new_n9043_), .Y(u2__abc_52138_new_n9045_));
NAND2X1 NAND2X1_1357 ( .A(u2__abc_52138_new_n4119_), .B(u2__abc_52138_new_n9062_), .Y(u2__abc_52138_new_n9064_));
NAND2X1 NAND2X1_1358 ( .A(u2__abc_52138_new_n9105_), .B(u2__abc_52138_new_n9106_), .Y(u2__abc_52138_new_n9107_));
NAND2X1 NAND2X1_1359 ( .A(u2__abc_52138_new_n4089_), .B(u2__abc_52138_new_n9155_), .Y(u2__abc_52138_new_n9164_));
NAND2X1 NAND2X1_136 ( .A(\a[23] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1229_));
NAND2X1 NAND2X1_1360 ( .A(u2__abc_52138_new_n9207_), .B(u2__abc_52138_new_n9208_), .Y(u2__abc_52138_new_n9209_));
NAND2X1 NAND2X1_1361 ( .A(u2__abc_52138_new_n9205_), .B(u2__abc_52138_new_n9209_), .Y(u2__abc_52138_new_n9217_));
NAND2X1 NAND2X1_1362 ( .A(u2__abc_52138_new_n9226_), .B(u2__abc_52138_new_n9229_), .Y(u2__abc_52138_new_n9230_));
NAND2X1 NAND2X1_1363 ( .A(u2__abc_52138_new_n5724_), .B(u2__abc_52138_new_n9321_), .Y(u2__abc_52138_new_n9322_));
NAND2X1 NAND2X1_1364 ( .A(u2__abc_52138_new_n5667_), .B(u2__abc_52138_new_n9383_), .Y(u2__abc_52138_new_n9391_));
NAND2X1 NAND2X1_1365 ( .A(u2__abc_52138_new_n5629_), .B(u2__abc_52138_new_n9490_), .Y(u2__abc_52138_new_n9491_));
NAND2X1 NAND2X1_1366 ( .A(u2__abc_52138_new_n5563_), .B(u2__abc_52138_new_n9532_), .Y(u2__abc_52138_new_n9533_));
NAND2X1 NAND2X1_1367 ( .A(u2__abc_52138_new_n5586_), .B(u2__abc_52138_new_n9574_), .Y(u2__abc_52138_new_n9575_));
NAND2X1 NAND2X1_1368 ( .A(u2_remHi_284_), .B(u2__abc_52138_new_n5573_), .Y(u2__abc_52138_new_n9604_));
NAND2X1 NAND2X1_1369 ( .A(u2__abc_52138_new_n5536_), .B(u2__abc_52138_new_n9666_), .Y(u2__abc_52138_new_n9667_));
NAND2X1 NAND2X1_137 ( .A(\a[112] ), .B(\a[25] ), .Y(_abc_65734_new_n1231_));
NAND2X1 NAND2X1_1370 ( .A(u2__abc_52138_new_n5470_), .B(u2__abc_52138_new_n9728_), .Y(u2__abc_52138_new_n9736_));
NAND2X1 NAND2X1_1371 ( .A(u2__abc_52138_new_n5493_), .B(u2__abc_52138_new_n9748_), .Y(u2__abc_52138_new_n9749_));
NAND2X1 NAND2X1_1372 ( .A(u2_remHi_300_), .B(u2__abc_52138_new_n5480_), .Y(u2__abc_52138_new_n9778_));
NAND2X1 NAND2X1_1373 ( .A(u2__abc_52138_new_n5500_), .B(u2__abc_52138_new_n9746_), .Y(u2__abc_52138_new_n9788_));
NAND2X1 NAND2X1_1374 ( .A(u2__abc_52138_new_n9792_), .B(u2__abc_52138_new_n9793_), .Y(u2__abc_52138_new_n9794_));
NAND2X1 NAND2X1_1375 ( .A(u2__abc_52138_new_n5422_), .B(u2__abc_52138_new_n9813_), .Y(u2__abc_52138_new_n9821_));
NAND2X1 NAND2X1_1376 ( .A(u2__abc_52138_new_n5450_), .B(u2__abc_52138_new_n9834_), .Y(u2__abc_52138_new_n9835_));
NAND2X1 NAND2X1_1377 ( .A(u2__abc_52138_new_n5379_), .B(u2__abc_52138_new_n9876_), .Y(u2__abc_52138_new_n9877_));
NAND2X1 NAND2X1_1378 ( .A(u2__abc_52138_new_n5386_), .B(u2__abc_52138_new_n9876_), .Y(u2__abc_52138_new_n9918_));
NAND2X1 NAND2X1_1379 ( .A(u2__abc_52138_new_n9917_), .B(u2__abc_52138_new_n9918_), .Y(u2__abc_52138_new_n9919_));
NAND2X1 NAND2X1_138 ( .A(\a[25] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1234_));
NAND2X1 NAND2X1_1380 ( .A(u2__abc_52138_new_n5398_), .B(u2__abc_52138_new_n9919_), .Y(u2__abc_52138_new_n9920_));
NAND2X1 NAND2X1_1381 ( .A(u2__abc_52138_new_n5405_), .B(u2__abc_52138_new_n9916_), .Y(u2__abc_52138_new_n9958_));
NAND2X1 NAND2X1_1382 ( .A(u2__abc_52138_new_n5347_), .B(u2__abc_52138_new_n5349_), .Y(u2__abc_52138_new_n9985_));
NAND2X1 NAND2X1_1383 ( .A(u2__abc_52138_new_n5356_), .B(u2__abc_52138_new_n9988_), .Y(u2__abc_52138_new_n9997_));
NAND2X1 NAND2X1_1384 ( .A(u2__abc_52138_new_n5332_), .B(u2__abc_52138_new_n10009_), .Y(u2__abc_52138_new_n10010_));
NAND2X1 NAND2X1_1385 ( .A(u2__abc_52138_new_n10050_), .B(u2__abc_52138_new_n10051_), .Y(u2__abc_52138_new_n10052_));
NAND2X1 NAND2X1_1386 ( .A(u2__abc_52138_new_n5289_), .B(u2__abc_52138_new_n10072_), .Y(u2__abc_52138_new_n10080_));
NAND2X1 NAND2X1_1387 ( .A(u2__abc_52138_new_n5312_), .B(u2__abc_52138_new_n10092_), .Y(u2__abc_52138_new_n10093_));
NAND2X1 NAND2X1_1388 ( .A(u2_remHi_332_), .B(u2__abc_52138_new_n5299_), .Y(u2__abc_52138_new_n10122_));
NAND2X1 NAND2X1_1389 ( .A(u2__abc_52138_new_n5241_), .B(u2__abc_52138_new_n10137_), .Y(u2__abc_52138_new_n10138_));
NAND2X1 NAND2X1_139 ( .A(\a[112] ), .B(\a[27] ), .Y(_abc_65734_new_n1236_));
NAND2X1 NAND2X1_1390 ( .A(u2__abc_52138_new_n5265_), .B(u2__abc_52138_new_n10180_), .Y(u2__abc_52138_new_n10181_));
NAND2X1 NAND2X1_1391 ( .A(u2__abc_52138_new_n5199_), .B(u2__abc_52138_new_n10223_), .Y(u2__abc_52138_new_n10224_));
NAND2X1 NAND2X1_1392 ( .A(u2__abc_52138_new_n5220_), .B(u2__abc_52138_new_n10267_), .Y(u2__abc_52138_new_n10268_));
NAND2X1 NAND2X1_1393 ( .A(u2__abc_52138_new_n5207_), .B(u2__abc_52138_new_n5209_), .Y(u2__abc_52138_new_n10285_));
NAND2X1 NAND2X1_1394 ( .A(u2__abc_52138_new_n10285_), .B(u2__abc_52138_new_n10287_), .Y(u2__abc_52138_new_n10289_));
NAND2X1 NAND2X1_1395 ( .A(u2__abc_52138_new_n10311_), .B(u2__abc_52138_new_n10312_), .Y(u2__abc_52138_new_n10313_));
NAND2X1 NAND2X1_1396 ( .A(u2__abc_52138_new_n5149_), .B(u2__abc_52138_new_n10313_), .Y(u2__abc_52138_new_n10314_));
NAND2X1 NAND2X1_1397 ( .A(u2__abc_52138_new_n5172_), .B(u2__abc_52138_new_n10355_), .Y(u2__abc_52138_new_n10356_));
NAND2X1 NAND2X1_1398 ( .A(u2__abc_52138_new_n5094_), .B(u2__abc_52138_new_n5100_), .Y(u2__abc_52138_new_n10418_));
NAND2X1 NAND2X1_1399 ( .A(u2__abc_52138_new_n5106_), .B(u2__abc_52138_new_n10421_), .Y(u2__abc_52138_new_n10430_));
NAND2X1 NAND2X1_14 ( .A(aNan), .B(\a[13] ), .Y(_abc_65734_new_n870_));
NAND2X1 NAND2X1_140 ( .A(\a[27] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1239_));
NAND2X1 NAND2X1_1400 ( .A(u2__abc_52138_new_n5125_), .B(u2__abc_52138_new_n10443_), .Y(u2__abc_52138_new_n10444_));
NAND2X1 NAND2X1_1401 ( .A(u2__abc_52138_new_n10526_), .B(u2__abc_52138_new_n10527_), .Y(u2__abc_52138_new_n10528_));
NAND2X1 NAND2X1_1402 ( .A(u2__abc_52138_new_n5086_), .B(u2__abc_52138_new_n10528_), .Y(u2__abc_52138_new_n10536_));
NAND2X1 NAND2X1_1403 ( .A(u2__abc_52138_new_n5069_), .B(u2__abc_52138_new_n10546_), .Y(u2__abc_52138_new_n10554_));
NAND2X1 NAND2X1_1404 ( .A(u2__abc_52138_new_n5022_), .B(u2__abc_52138_new_n10568_), .Y(u2__abc_52138_new_n10576_));
NAND2X1 NAND2X1_1405 ( .A(u2__abc_52138_new_n5010_), .B(u2__abc_52138_new_n10608_), .Y(u2__abc_52138_new_n10609_));
NAND2X1 NAND2X1_1406 ( .A(u2__abc_52138_new_n10648_), .B(u2__abc_52138_new_n9965_), .Y(u2__abc_52138_new_n10649_));
NAND2X1 NAND2X1_1407 ( .A(u2__abc_52138_new_n6156_), .B(u2__abc_52138_new_n10704_), .Y(u2__abc_52138_new_n10705_));
NAND2X1 NAND2X1_1408 ( .A(u2__abc_52138_new_n10749_), .B(u2__abc_52138_new_n10750_), .Y(u2__abc_52138_new_n10751_));
NAND2X1 NAND2X1_1409 ( .A(u2__abc_52138_new_n6296_), .B(u2__abc_52138_new_n10751_), .Y(u2__abc_52138_new_n10759_));
NAND2X1 NAND2X1_141 ( .A(\a[112] ), .B(\a[29] ), .Y(_abc_65734_new_n1241_));
NAND2X1 NAND2X1_1410 ( .A(u2__abc_52138_new_n6301_), .B(u2__abc_52138_new_n10762_), .Y(u2__abc_52138_new_n10763_));
NAND2X1 NAND2X1_1411 ( .A(u2__abc_52138_new_n6284_), .B(u2__abc_52138_new_n10770_), .Y(u2__abc_52138_new_n10778_));
NAND2X1 NAND2X1_1412 ( .A(u2__abc_52138_new_n6324_), .B(u2__abc_52138_new_n10793_), .Y(u2__abc_52138_new_n10794_));
NAND2X1 NAND2X1_1413 ( .A(u2_remHi_396_), .B(u2__abc_52138_new_n6306_), .Y(u2__abc_52138_new_n10821_));
NAND2X1 NAND2X1_1414 ( .A(u2__abc_52138_new_n6247_), .B(u2__abc_52138_new_n10855_), .Y(u2__abc_52138_new_n10863_));
NAND2X1 NAND2X1_1415 ( .A(u2__abc_52138_new_n6275_), .B(u2__abc_52138_new_n10877_), .Y(u2__abc_52138_new_n10878_));
NAND2X1 NAND2X1_1416 ( .A(u2__abc_52138_new_n6205_), .B(u2__abc_52138_new_n10921_), .Y(u2__abc_52138_new_n10922_));
NAND2X1 NAND2X1_1417 ( .A(u2__abc_52138_new_n6228_), .B(u2__abc_52138_new_n10964_), .Y(u2__abc_52138_new_n10965_));
NAND2X1 NAND2X1_1418 ( .A(u2__abc_52138_new_n6279_), .B(u2__abc_52138_new_n10833_), .Y(u2__abc_52138_new_n11008_));
NAND2X1 NAND2X1_1419 ( .A(u2__abc_52138_new_n11010_), .B(u2__abc_52138_new_n11002_), .Y(u2__abc_52138_new_n11011_));
NAND2X1 NAND2X1_142 ( .A(\a[29] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1244_));
NAND2X1 NAND2X1_1420 ( .A(u2__abc_52138_new_n6129_), .B(u2__abc_52138_new_n11011_), .Y(u2__abc_52138_new_n11012_));
NAND2X1 NAND2X1_1421 ( .A(u2__abc_52138_new_n6112_), .B(u2__abc_52138_new_n11031_), .Y(u2__abc_52138_new_n11033_));
NAND2X1 NAND2X1_1422 ( .A(u2__abc_52138_new_n6105_), .B(u2__abc_52138_new_n11055_), .Y(u2__abc_52138_new_n11056_));
NAND2X1 NAND2X1_1423 ( .A(u2__abc_52138_new_n6088_), .B(u2__abc_52138_new_n11075_), .Y(u2__abc_52138_new_n11077_));
NAND2X1 NAND2X1_1424 ( .A(u2__abc_52138_new_n6040_), .B(u2__abc_52138_new_n11118_), .Y(u2__abc_52138_new_n11120_));
NAND2X1 NAND2X1_1425 ( .A(u2__abc_52138_new_n6079_), .B(u2__abc_52138_new_n11140_), .Y(u2__abc_52138_new_n11141_));
NAND2X1 NAND2X1_1426 ( .A(u2__abc_52138_new_n6062_), .B(u2__abc_52138_new_n11160_), .Y(u2__abc_52138_new_n11162_));
NAND2X1 NAND2X1_1427 ( .A(u2__abc_52138_new_n6025_), .B(u2__abc_52138_new_n11205_), .Y(u2__abc_52138_new_n11206_));
NAND2X1 NAND2X1_1428 ( .A(u2__abc_52138_new_n6002_), .B(u2__abc_52138_new_n11235_), .Y(u2__abc_52138_new_n11236_));
NAND2X1 NAND2X1_1429 ( .A(u2__abc_52138_new_n5971_), .B(u2__abc_52138_new_n11269_), .Y(u2__abc_52138_new_n11277_));
NAND2X1 NAND2X1_143 ( .A(\a[112] ), .B(\a[31] ), .Y(_abc_65734_new_n1246_));
NAND2X1 NAND2X1_1430 ( .A(u2__abc_52138_new_n5985_), .B(u2__abc_52138_new_n11269_), .Y(u2__abc_52138_new_n11312_));
NAND2X1 NAND2X1_1431 ( .A(u2__abc_52138_new_n11311_), .B(u2__abc_52138_new_n11312_), .Y(u2__abc_52138_new_n11313_));
NAND2X1 NAND2X1_1432 ( .A(u2__abc_52138_new_n5964_), .B(u2__abc_52138_new_n11313_), .Y(u2__abc_52138_new_n11314_));
NAND2X1 NAND2X1_1433 ( .A(u2_cnt_2_), .B(u2__abc_52138_new_n11382_), .Y(u2__abc_52138_new_n11388_));
NAND2X1 NAND2X1_1434 ( .A(u2_cnt_3_), .B(u2__abc_52138_new_n11391_), .Y(u2__abc_52138_new_n11392_));
NAND2X1 NAND2X1_1435 ( .A(u2_cnt_5_), .B(u2__abc_52138_new_n11398_), .Y(u2__abc_52138_new_n11401_));
NAND2X1 NAND2X1_1436 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11514_));
NAND2X1 NAND2X1_1437 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11526_));
NAND2X1 NAND2X1_1438 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11565_));
NAND2X1 NAND2X1_1439 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11625_));
NAND2X1 NAND2X1_144 ( .A(\a[31] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1249_));
NAND2X1 NAND2X1_1440 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11655_));
NAND2X1 NAND2X1_1441 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11730_));
NAND2X1 NAND2X1_1442 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11784_));
NAND2X1 NAND2X1_1443 ( .A(1'h0), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11832_));
NAND2X1 NAND2X1_1444 ( .A(fracta1_19_), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n11932_));
NAND2X1 NAND2X1_1445 ( .A(fracta1_51_), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n12032_));
NAND2X1 NAND2X1_1446 ( .A(fracta1_60_), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n12062_));
NAND2X1 NAND2X1_1447 ( .A(fracta1_83_), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n12135_));
NAND2X1 NAND2X1_1448 ( .A(fracta1_84_), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n12141_));
NAND2X1 NAND2X1_1449 ( .A(u2__abc_52138_new_n3023_), .B(u2__abc_52138_new_n3025_), .Y(u2__abc_52138_new_n12833_));
NAND2X1 NAND2X1_145 ( .A(\a[112] ), .B(\a[33] ), .Y(_abc_65734_new_n1251_));
NAND2X1 NAND2X1_1450 ( .A(u2__abc_52138_new_n7052_), .B(u2__abc_52138_new_n3473_), .Y(u2__abc_52138_new_n12872_));
NAND2X1 NAND2X1_1451 ( .A(u2__abc_52138_new_n6484_), .B(u2__abc_52138_new_n12887_), .Y(u2__abc_52138_new_n12888_));
NAND2X1 NAND2X1_1452 ( .A(u2__abc_52138_new_n7265_), .B(u2__abc_52138_new_n3889_), .Y(u2__abc_52138_new_n12894_));
NAND2X1 NAND2X1_1453 ( .A(u2__abc_52138_new_n3882_), .B(u2__abc_52138_new_n3884_), .Y(u2__abc_52138_new_n12896_));
NAND2X1 NAND2X1_1454 ( .A(u2__abc_52138_new_n3928_), .B(u2__abc_52138_new_n12916_), .Y(u2__abc_52138_new_n12917_));
NAND2X1 NAND2X1_1455 ( .A(u2__abc_52138_new_n7580_), .B(u2__abc_52138_new_n3942_), .Y(u2__abc_52138_new_n12926_));
NAND2X1 NAND2X1_1456 ( .A(u2__abc_52138_new_n12941_), .B(u2__abc_52138_new_n7803_), .Y(u2__abc_52138_new_n12942_));
NAND2X1 NAND2X1_1457 ( .A(u2__abc_52138_new_n4629_), .B(u2__abc_52138_new_n4640_), .Y(u2__abc_52138_new_n12967_));
NAND2X1 NAND2X1_1458 ( .A(u2__abc_52138_new_n4558_), .B(u2__abc_52138_new_n4569_), .Y(u2__abc_52138_new_n12981_));
NAND2X1 NAND2X1_1459 ( .A(u2__abc_52138_new_n4979_), .B(u2__abc_52138_new_n13025_), .Y(u2__abc_52138_new_n13026_));
NAND2X1 NAND2X1_146 ( .A(\a[33] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1254_));
NAND2X1 NAND2X1_1460 ( .A(u2__abc_52138_new_n5182_), .B(u2__abc_52138_new_n5885_), .Y(u2__abc_52138_new_n13035_));
NAND2X1 NAND2X1_1461 ( .A(u2__abc_52138_new_n13047_), .B(u2__abc_52138_new_n13046_), .Y(u2__abc_52138_new_n13048_));
NAND2X1 NAND2X1_1462 ( .A(u2__abc_52138_new_n13054_), .B(u2__abc_52138_new_n13053_), .Y(u2__abc_52138_new_n13055_));
NAND2X1 NAND2X1_1463 ( .A(u2__abc_52138_new_n13062_), .B(u2__abc_52138_new_n13061_), .Y(u2__abc_52138_new_n13063_));
NAND2X1 NAND2X1_1464 ( .A(u2__abc_52138_new_n13070_), .B(u2__abc_52138_new_n13069_), .Y(u2__abc_52138_new_n13071_));
NAND2X1 NAND2X1_1465 ( .A(u2__abc_52138_new_n13078_), .B(u2__abc_52138_new_n13077_), .Y(u2__abc_52138_new_n13079_));
NAND2X1 NAND2X1_1466 ( .A(u2__abc_52138_new_n13085_), .B(u2__abc_52138_new_n13084_), .Y(u2__abc_52138_new_n13086_));
NAND2X1 NAND2X1_1467 ( .A(u2__abc_52138_new_n13093_), .B(u2__abc_52138_new_n13092_), .Y(u2__abc_52138_new_n13094_));
NAND2X1 NAND2X1_1468 ( .A(u2__abc_52138_new_n13101_), .B(u2__abc_52138_new_n13100_), .Y(u2__abc_52138_new_n13102_));
NAND2X1 NAND2X1_1469 ( .A(u2__abc_52138_new_n13109_), .B(u2__abc_52138_new_n13108_), .Y(u2__abc_52138_new_n13110_));
NAND2X1 NAND2X1_147 ( .A(\a[112] ), .B(\a[35] ), .Y(_abc_65734_new_n1256_));
NAND2X1 NAND2X1_1470 ( .A(u2__abc_52138_new_n13116_), .B(u2__abc_52138_new_n13115_), .Y(u2__abc_52138_new_n13117_));
NAND2X1 NAND2X1_1471 ( .A(u2__abc_52138_new_n13124_), .B(u2__abc_52138_new_n13123_), .Y(u2__abc_52138_new_n13125_));
NAND2X1 NAND2X1_1472 ( .A(u2__abc_52138_new_n13132_), .B(u2__abc_52138_new_n13131_), .Y(u2__abc_52138_new_n13133_));
NAND2X1 NAND2X1_1473 ( .A(u2__abc_52138_new_n13140_), .B(u2__abc_52138_new_n13139_), .Y(u2__abc_52138_new_n13141_));
NAND2X1 NAND2X1_1474 ( .A(u2__abc_52138_new_n13147_), .B(u2__abc_52138_new_n13146_), .Y(u2__abc_52138_new_n13148_));
NAND2X1 NAND2X1_1475 ( .A(u2__abc_52138_new_n13155_), .B(u2__abc_52138_new_n13154_), .Y(u2__abc_52138_new_n13156_));
NAND2X1 NAND2X1_1476 ( .A(u2__abc_52138_new_n13163_), .B(u2__abc_52138_new_n13162_), .Y(u2__abc_52138_new_n13164_));
NAND2X1 NAND2X1_1477 ( .A(u2__abc_52138_new_n13171_), .B(u2__abc_52138_new_n13170_), .Y(u2__abc_52138_new_n13172_));
NAND2X1 NAND2X1_1478 ( .A(u2__abc_52138_new_n13178_), .B(u2__abc_52138_new_n13177_), .Y(u2__abc_52138_new_n13179_));
NAND2X1 NAND2X1_1479 ( .A(u2__abc_52138_new_n13186_), .B(u2__abc_52138_new_n13185_), .Y(u2__abc_52138_new_n13187_));
NAND2X1 NAND2X1_148 ( .A(\a[35] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1259_));
NAND2X1 NAND2X1_1480 ( .A(u2__abc_52138_new_n13194_), .B(u2__abc_52138_new_n13193_), .Y(u2__abc_52138_new_n13195_));
NAND2X1 NAND2X1_1481 ( .A(u2__abc_52138_new_n13202_), .B(u2__abc_52138_new_n13201_), .Y(u2__abc_52138_new_n13203_));
NAND2X1 NAND2X1_1482 ( .A(u2__abc_52138_new_n13209_), .B(u2__abc_52138_new_n13208_), .Y(u2__abc_52138_new_n13210_));
NAND2X1 NAND2X1_1483 ( .A(u2__abc_52138_new_n13217_), .B(u2__abc_52138_new_n13216_), .Y(u2__abc_52138_new_n13218_));
NAND2X1 NAND2X1_1484 ( .A(u2__abc_52138_new_n13225_), .B(u2__abc_52138_new_n13224_), .Y(u2__abc_52138_new_n13226_));
NAND2X1 NAND2X1_1485 ( .A(u2__abc_52138_new_n13233_), .B(u2__abc_52138_new_n13232_), .Y(u2__abc_52138_new_n13234_));
NAND2X1 NAND2X1_1486 ( .A(u2__abc_52138_new_n13240_), .B(u2__abc_52138_new_n13239_), .Y(u2__abc_52138_new_n13241_));
NAND2X1 NAND2X1_1487 ( .A(u2__abc_52138_new_n13248_), .B(u2__abc_52138_new_n13247_), .Y(u2__abc_52138_new_n13249_));
NAND2X1 NAND2X1_1488 ( .A(u2__abc_52138_new_n13256_), .B(u2__abc_52138_new_n13255_), .Y(u2__abc_52138_new_n13257_));
NAND2X1 NAND2X1_1489 ( .A(u2__abc_52138_new_n13264_), .B(u2__abc_52138_new_n13263_), .Y(u2__abc_52138_new_n13265_));
NAND2X1 NAND2X1_149 ( .A(\a[112] ), .B(\a[37] ), .Y(_abc_65734_new_n1261_));
NAND2X1 NAND2X1_1490 ( .A(u2__abc_52138_new_n13271_), .B(u2__abc_52138_new_n13270_), .Y(u2__abc_52138_new_n13272_));
NAND2X1 NAND2X1_1491 ( .A(u2__abc_52138_new_n13279_), .B(u2__abc_52138_new_n13278_), .Y(u2__abc_52138_new_n13280_));
NAND2X1 NAND2X1_1492 ( .A(u2__abc_52138_new_n13287_), .B(u2__abc_52138_new_n13286_), .Y(u2__abc_52138_new_n13288_));
NAND2X1 NAND2X1_1493 ( .A(u2__abc_52138_new_n13295_), .B(u2__abc_52138_new_n13294_), .Y(u2__abc_52138_new_n13296_));
NAND2X1 NAND2X1_1494 ( .A(u2__abc_52138_new_n13302_), .B(u2__abc_52138_new_n13301_), .Y(u2__abc_52138_new_n13303_));
NAND2X1 NAND2X1_1495 ( .A(u2__abc_52138_new_n13311_), .B(u2__abc_52138_new_n13309_), .Y(u2__abc_52138_new_n13312_));
NAND2X1 NAND2X1_1496 ( .A(u2__abc_52138_new_n13319_), .B(u2__abc_52138_new_n13318_), .Y(u2__abc_52138_new_n13320_));
NAND2X1 NAND2X1_1497 ( .A(u2__abc_52138_new_n13327_), .B(u2__abc_52138_new_n13326_), .Y(u2__abc_52138_new_n13328_));
NAND2X1 NAND2X1_1498 ( .A(u2__abc_52138_new_n13334_), .B(u2__abc_52138_new_n13333_), .Y(u2__abc_52138_new_n13335_));
NAND2X1 NAND2X1_1499 ( .A(u2__abc_52138_new_n13342_), .B(u2__abc_52138_new_n13341_), .Y(u2__abc_52138_new_n13343_));
NAND2X1 NAND2X1_15 ( .A(aNan), .B(\a[14] ), .Y(_abc_65734_new_n873_));
NAND2X1 NAND2X1_150 ( .A(\a[37] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1264_));
NAND2X1 NAND2X1_1500 ( .A(u2__abc_52138_new_n13350_), .B(u2__abc_52138_new_n13349_), .Y(u2__abc_52138_new_n13351_));
NAND2X1 NAND2X1_1501 ( .A(u2__abc_52138_new_n13358_), .B(u2__abc_52138_new_n13357_), .Y(u2__abc_52138_new_n13359_));
NAND2X1 NAND2X1_1502 ( .A(u2__abc_52138_new_n13365_), .B(u2__abc_52138_new_n13364_), .Y(u2__abc_52138_new_n13366_));
NAND2X1 NAND2X1_1503 ( .A(u2__abc_52138_new_n13373_), .B(u2__abc_52138_new_n13372_), .Y(u2__abc_52138_new_n13374_));
NAND2X1 NAND2X1_1504 ( .A(u2__abc_52138_new_n13381_), .B(u2__abc_52138_new_n13380_), .Y(u2__abc_52138_new_n13382_));
NAND2X1 NAND2X1_1505 ( .A(u2__abc_52138_new_n13389_), .B(u2__abc_52138_new_n13388_), .Y(u2__abc_52138_new_n13390_));
NAND2X1 NAND2X1_1506 ( .A(u2__abc_52138_new_n13396_), .B(u2__abc_52138_new_n13395_), .Y(u2__abc_52138_new_n13397_));
NAND2X1 NAND2X1_1507 ( .A(u2__abc_52138_new_n13404_), .B(u2__abc_52138_new_n13403_), .Y(u2__abc_52138_new_n13405_));
NAND2X1 NAND2X1_1508 ( .A(u2__abc_52138_new_n13412_), .B(u2__abc_52138_new_n13411_), .Y(u2__abc_52138_new_n13413_));
NAND2X1 NAND2X1_1509 ( .A(u2__abc_52138_new_n13420_), .B(u2__abc_52138_new_n13419_), .Y(u2__abc_52138_new_n13421_));
NAND2X1 NAND2X1_151 ( .A(\a[112] ), .B(\a[39] ), .Y(_abc_65734_new_n1266_));
NAND2X1 NAND2X1_1510 ( .A(u2__abc_52138_new_n13427_), .B(u2__abc_52138_new_n13426_), .Y(u2__abc_52138_new_n13428_));
NAND2X1 NAND2X1_1511 ( .A(u2__abc_52138_new_n13435_), .B(u2__abc_52138_new_n13434_), .Y(u2__abc_52138_new_n13436_));
NAND2X1 NAND2X1_1512 ( .A(u2__abc_52138_new_n13443_), .B(u2__abc_52138_new_n13442_), .Y(u2__abc_52138_new_n13444_));
NAND2X1 NAND2X1_1513 ( .A(u2__abc_52138_new_n13451_), .B(u2__abc_52138_new_n13450_), .Y(u2__abc_52138_new_n13452_));
NAND2X1 NAND2X1_1514 ( .A(u2__abc_52138_new_n13458_), .B(u2__abc_52138_new_n13457_), .Y(u2__abc_52138_new_n13459_));
NAND2X1 NAND2X1_1515 ( .A(u2__abc_52138_new_n13466_), .B(u2__abc_52138_new_n13465_), .Y(u2__abc_52138_new_n13467_));
NAND2X1 NAND2X1_1516 ( .A(u2__abc_52138_new_n13474_), .B(u2__abc_52138_new_n13473_), .Y(u2__abc_52138_new_n13475_));
NAND2X1 NAND2X1_1517 ( .A(u2__abc_52138_new_n13482_), .B(u2__abc_52138_new_n13481_), .Y(u2__abc_52138_new_n13483_));
NAND2X1 NAND2X1_1518 ( .A(u2__abc_52138_new_n13489_), .B(u2__abc_52138_new_n13488_), .Y(u2__abc_52138_new_n13490_));
NAND2X1 NAND2X1_1519 ( .A(u2__abc_52138_new_n13497_), .B(u2__abc_52138_new_n13496_), .Y(u2__abc_52138_new_n13498_));
NAND2X1 NAND2X1_152 ( .A(\a[39] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1269_));
NAND2X1 NAND2X1_1520 ( .A(u2__abc_52138_new_n13505_), .B(u2__abc_52138_new_n13504_), .Y(u2__abc_52138_new_n13506_));
NAND2X1 NAND2X1_1521 ( .A(u2__abc_52138_new_n13513_), .B(u2__abc_52138_new_n13512_), .Y(u2__abc_52138_new_n13514_));
NAND2X1 NAND2X1_1522 ( .A(u2__abc_52138_new_n13520_), .B(u2__abc_52138_new_n13519_), .Y(u2__abc_52138_new_n13521_));
NAND2X1 NAND2X1_1523 ( .A(u2__abc_52138_new_n13528_), .B(u2__abc_52138_new_n13527_), .Y(u2__abc_52138_new_n13529_));
NAND2X1 NAND2X1_1524 ( .A(u2__abc_52138_new_n13536_), .B(u2__abc_52138_new_n13535_), .Y(u2__abc_52138_new_n13537_));
NAND2X1 NAND2X1_1525 ( .A(u2__abc_52138_new_n13544_), .B(u2__abc_52138_new_n13543_), .Y(u2__abc_52138_new_n13545_));
NAND2X1 NAND2X1_1526 ( .A(u2__abc_52138_new_n13551_), .B(u2__abc_52138_new_n13550_), .Y(u2__abc_52138_new_n13552_));
NAND2X1 NAND2X1_1527 ( .A(u2__abc_52138_new_n13559_), .B(u2__abc_52138_new_n13558_), .Y(u2__abc_52138_new_n13560_));
NAND2X1 NAND2X1_1528 ( .A(u2__abc_52138_new_n13567_), .B(u2__abc_52138_new_n13566_), .Y(u2__abc_52138_new_n13568_));
NAND2X1 NAND2X1_1529 ( .A(u2__abc_52138_new_n13575_), .B(u2__abc_52138_new_n13574_), .Y(u2__abc_52138_new_n13576_));
NAND2X1 NAND2X1_153 ( .A(\a[112] ), .B(\a[41] ), .Y(_abc_65734_new_n1271_));
NAND2X1 NAND2X1_1530 ( .A(u2__abc_52138_new_n13582_), .B(u2__abc_52138_new_n13581_), .Y(u2__abc_52138_new_n13583_));
NAND2X1 NAND2X1_1531 ( .A(u2__abc_52138_new_n13590_), .B(u2__abc_52138_new_n13589_), .Y(u2__abc_52138_new_n13591_));
NAND2X1 NAND2X1_1532 ( .A(u2__abc_52138_new_n13598_), .B(u2__abc_52138_new_n13597_), .Y(u2__abc_52138_new_n13599_));
NAND2X1 NAND2X1_1533 ( .A(u2__abc_52138_new_n13606_), .B(u2__abc_52138_new_n13605_), .Y(u2__abc_52138_new_n13607_));
NAND2X1 NAND2X1_1534 ( .A(u2__abc_52138_new_n13613_), .B(u2__abc_52138_new_n13612_), .Y(u2__abc_52138_new_n13614_));
NAND2X1 NAND2X1_1535 ( .A(u2__abc_52138_new_n13621_), .B(u2__abc_52138_new_n13620_), .Y(u2__abc_52138_new_n13622_));
NAND2X1 NAND2X1_1536 ( .A(u2__abc_52138_new_n13629_), .B(u2__abc_52138_new_n13628_), .Y(u2__abc_52138_new_n13630_));
NAND2X1 NAND2X1_1537 ( .A(u2__abc_52138_new_n13637_), .B(u2__abc_52138_new_n13636_), .Y(u2__abc_52138_new_n13638_));
NAND2X1 NAND2X1_1538 ( .A(u2__abc_52138_new_n13644_), .B(u2__abc_52138_new_n13643_), .Y(u2__abc_52138_new_n13645_));
NAND2X1 NAND2X1_1539 ( .A(u2__abc_52138_new_n13652_), .B(u2__abc_52138_new_n13651_), .Y(u2__abc_52138_new_n13653_));
NAND2X1 NAND2X1_154 ( .A(\a[41] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1274_));
NAND2X1 NAND2X1_1540 ( .A(u2__abc_52138_new_n13660_), .B(u2__abc_52138_new_n13659_), .Y(u2__abc_52138_new_n13661_));
NAND2X1 NAND2X1_1541 ( .A(u2__abc_52138_new_n13668_), .B(u2__abc_52138_new_n13667_), .Y(u2__abc_52138_new_n13669_));
NAND2X1 NAND2X1_1542 ( .A(u2__abc_52138_new_n13675_), .B(u2__abc_52138_new_n13674_), .Y(u2__abc_52138_new_n13676_));
NAND2X1 NAND2X1_1543 ( .A(u2__abc_52138_new_n13683_), .B(u2__abc_52138_new_n13682_), .Y(u2__abc_52138_new_n13684_));
NAND2X1 NAND2X1_1544 ( .A(u2__abc_52138_new_n13691_), .B(u2__abc_52138_new_n13690_), .Y(u2__abc_52138_new_n13692_));
NAND2X1 NAND2X1_1545 ( .A(u2__abc_52138_new_n13699_), .B(u2__abc_52138_new_n13698_), .Y(u2__abc_52138_new_n13700_));
NAND2X1 NAND2X1_1546 ( .A(u2__abc_52138_new_n13706_), .B(u2__abc_52138_new_n13705_), .Y(u2__abc_52138_new_n13707_));
NAND2X1 NAND2X1_1547 ( .A(u2__abc_52138_new_n13714_), .B(u2__abc_52138_new_n13713_), .Y(u2__abc_52138_new_n13715_));
NAND2X1 NAND2X1_1548 ( .A(u2__abc_52138_new_n13722_), .B(u2__abc_52138_new_n13721_), .Y(u2__abc_52138_new_n13723_));
NAND2X1 NAND2X1_1549 ( .A(u2__abc_52138_new_n13730_), .B(u2__abc_52138_new_n13729_), .Y(u2__abc_52138_new_n13731_));
NAND2X1 NAND2X1_155 ( .A(\a[112] ), .B(\a[43] ), .Y(_abc_65734_new_n1276_));
NAND2X1 NAND2X1_1550 ( .A(u2__abc_52138_new_n13737_), .B(u2__abc_52138_new_n13736_), .Y(u2__abc_52138_new_n13738_));
NAND2X1 NAND2X1_1551 ( .A(u2__abc_52138_new_n13745_), .B(u2__abc_52138_new_n13744_), .Y(u2__abc_52138_new_n13746_));
NAND2X1 NAND2X1_1552 ( .A(u2__abc_52138_new_n13753_), .B(u2__abc_52138_new_n13752_), .Y(u2__abc_52138_new_n13754_));
NAND2X1 NAND2X1_1553 ( .A(u2__abc_52138_new_n13761_), .B(u2__abc_52138_new_n13760_), .Y(u2__abc_52138_new_n13762_));
NAND2X1 NAND2X1_1554 ( .A(u2__abc_52138_new_n13768_), .B(u2__abc_52138_new_n13767_), .Y(u2__abc_52138_new_n13769_));
NAND2X1 NAND2X1_1555 ( .A(u2__abc_52138_new_n13776_), .B(u2__abc_52138_new_n13775_), .Y(u2__abc_52138_new_n13777_));
NAND2X1 NAND2X1_1556 ( .A(u2__abc_52138_new_n13784_), .B(u2__abc_52138_new_n13783_), .Y(u2__abc_52138_new_n13785_));
NAND2X1 NAND2X1_1557 ( .A(u2__abc_52138_new_n13792_), .B(u2__abc_52138_new_n13791_), .Y(u2__abc_52138_new_n13793_));
NAND2X1 NAND2X1_1558 ( .A(u2__abc_52138_new_n13799_), .B(u2__abc_52138_new_n13798_), .Y(u2__abc_52138_new_n13800_));
NAND2X1 NAND2X1_1559 ( .A(u2__abc_52138_new_n13807_), .B(u2__abc_52138_new_n13806_), .Y(u2__abc_52138_new_n13808_));
NAND2X1 NAND2X1_156 ( .A(\a[43] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1279_));
NAND2X1 NAND2X1_1560 ( .A(u2__abc_52138_new_n13815_), .B(u2__abc_52138_new_n13814_), .Y(u2__abc_52138_new_n13816_));
NAND2X1 NAND2X1_1561 ( .A(u2__abc_52138_new_n13823_), .B(u2__abc_52138_new_n13822_), .Y(u2__abc_52138_new_n13824_));
NAND2X1 NAND2X1_1562 ( .A(u2__abc_52138_new_n13830_), .B(u2__abc_52138_new_n13829_), .Y(u2__abc_52138_new_n13831_));
NAND2X1 NAND2X1_1563 ( .A(u2__abc_52138_new_n13838_), .B(u2__abc_52138_new_n13837_), .Y(u2__abc_52138_new_n13839_));
NAND2X1 NAND2X1_1564 ( .A(u2__abc_52138_new_n13846_), .B(u2__abc_52138_new_n13845_), .Y(u2__abc_52138_new_n13847_));
NAND2X1 NAND2X1_1565 ( .A(u2__abc_52138_new_n13854_), .B(u2__abc_52138_new_n13853_), .Y(u2__abc_52138_new_n13855_));
NAND2X1 NAND2X1_1566 ( .A(u2__abc_52138_new_n13861_), .B(u2__abc_52138_new_n13860_), .Y(u2__abc_52138_new_n13862_));
NAND2X1 NAND2X1_1567 ( .A(u2__abc_52138_new_n13869_), .B(u2__abc_52138_new_n13868_), .Y(u2__abc_52138_new_n13870_));
NAND2X1 NAND2X1_1568 ( .A(u2__abc_52138_new_n13877_), .B(u2__abc_52138_new_n13876_), .Y(u2__abc_52138_new_n13878_));
NAND2X1 NAND2X1_1569 ( .A(u2__abc_52138_new_n13885_), .B(u2__abc_52138_new_n13884_), .Y(u2__abc_52138_new_n13886_));
NAND2X1 NAND2X1_157 ( .A(\a[112] ), .B(\a[45] ), .Y(_abc_65734_new_n1281_));
NAND2X1 NAND2X1_1570 ( .A(u2__abc_52138_new_n13892_), .B(u2__abc_52138_new_n13891_), .Y(u2__abc_52138_new_n13893_));
NAND2X1 NAND2X1_1571 ( .A(u2__abc_52138_new_n13900_), .B(u2__abc_52138_new_n13899_), .Y(u2__abc_52138_new_n13901_));
NAND2X1 NAND2X1_1572 ( .A(u2__abc_52138_new_n13908_), .B(u2__abc_52138_new_n13907_), .Y(u2__abc_52138_new_n13909_));
NAND2X1 NAND2X1_1573 ( .A(u2__abc_52138_new_n13916_), .B(u2__abc_52138_new_n13915_), .Y(u2__abc_52138_new_n13917_));
NAND2X1 NAND2X1_1574 ( .A(u2__abc_52138_new_n13923_), .B(u2__abc_52138_new_n13922_), .Y(u2__abc_52138_new_n13924_));
NAND2X1 NAND2X1_1575 ( .A(u2__abc_52138_new_n13931_), .B(u2__abc_52138_new_n13930_), .Y(u2__abc_52138_new_n13932_));
NAND2X1 NAND2X1_1576 ( .A(u2__abc_52138_new_n13939_), .B(u2__abc_52138_new_n13938_), .Y(u2__abc_52138_new_n13940_));
NAND2X1 NAND2X1_1577 ( .A(u2__abc_52138_new_n13947_), .B(u2__abc_52138_new_n13946_), .Y(u2__abc_52138_new_n13948_));
NAND2X1 NAND2X1_1578 ( .A(u2__abc_52138_new_n13954_), .B(u2__abc_52138_new_n13953_), .Y(u2__abc_52138_new_n13955_));
NAND2X1 NAND2X1_1579 ( .A(u2__abc_52138_new_n13963_), .B(u2__abc_52138_new_n13961_), .Y(u2__abc_52138_new_n13964_));
NAND2X1 NAND2X1_158 ( .A(\a[45] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1284_));
NAND2X1 NAND2X1_1580 ( .A(u2__abc_52138_new_n13971_), .B(u2__abc_52138_new_n13970_), .Y(u2__abc_52138_new_n13972_));
NAND2X1 NAND2X1_1581 ( .A(u2__abc_52138_new_n13979_), .B(u2__abc_52138_new_n13978_), .Y(u2__abc_52138_new_n13980_));
NAND2X1 NAND2X1_1582 ( .A(u2__abc_52138_new_n13986_), .B(u2__abc_52138_new_n13985_), .Y(u2__abc_52138_new_n13987_));
NAND2X1 NAND2X1_1583 ( .A(u2__abc_52138_new_n13994_), .B(u2__abc_52138_new_n13993_), .Y(u2__abc_52138_new_n13995_));
NAND2X1 NAND2X1_1584 ( .A(u2__abc_52138_new_n14002_), .B(u2__abc_52138_new_n14001_), .Y(u2__abc_52138_new_n14003_));
NAND2X1 NAND2X1_1585 ( .A(u2__abc_52138_new_n14010_), .B(u2__abc_52138_new_n14009_), .Y(u2__abc_52138_new_n14011_));
NAND2X1 NAND2X1_1586 ( .A(u2__abc_52138_new_n14017_), .B(u2__abc_52138_new_n14016_), .Y(u2__abc_52138_new_n14018_));
NAND2X1 NAND2X1_1587 ( .A(u2__abc_52138_new_n14025_), .B(u2__abc_52138_new_n14024_), .Y(u2__abc_52138_new_n14026_));
NAND2X1 NAND2X1_1588 ( .A(u2__abc_52138_new_n14033_), .B(u2__abc_52138_new_n14032_), .Y(u2__abc_52138_new_n14034_));
NAND2X1 NAND2X1_1589 ( .A(u2__abc_52138_new_n14041_), .B(u2__abc_52138_new_n14040_), .Y(u2__abc_52138_new_n14042_));
NAND2X1 NAND2X1_159 ( .A(\a[112] ), .B(\a[47] ), .Y(_abc_65734_new_n1286_));
NAND2X1 NAND2X1_1590 ( .A(u2__abc_52138_new_n14048_), .B(u2__abc_52138_new_n14047_), .Y(u2__abc_52138_new_n14049_));
NAND2X1 NAND2X1_1591 ( .A(u2__abc_52138_new_n14057_), .B(u2__abc_52138_new_n14055_), .Y(u2__abc_52138_new_n14058_));
NAND2X1 NAND2X1_1592 ( .A(u2__abc_52138_new_n14065_), .B(u2__abc_52138_new_n14064_), .Y(u2__abc_52138_new_n14066_));
NAND2X1 NAND2X1_1593 ( .A(u2__abc_52138_new_n14073_), .B(u2__abc_52138_new_n14072_), .Y(u2__abc_52138_new_n14074_));
NAND2X1 NAND2X1_1594 ( .A(u2__abc_52138_new_n14080_), .B(u2__abc_52138_new_n14079_), .Y(u2__abc_52138_new_n14081_));
NAND2X1 NAND2X1_1595 ( .A(u2__abc_52138_new_n14088_), .B(u2__abc_52138_new_n14087_), .Y(u2__abc_52138_new_n14089_));
NAND2X1 NAND2X1_1596 ( .A(u2__abc_52138_new_n14096_), .B(u2__abc_52138_new_n14095_), .Y(u2__abc_52138_new_n14097_));
NAND2X1 NAND2X1_1597 ( .A(u2__abc_52138_new_n14104_), .B(u2__abc_52138_new_n14103_), .Y(u2__abc_52138_new_n14105_));
NAND2X1 NAND2X1_1598 ( .A(u2__abc_52138_new_n14111_), .B(u2__abc_52138_new_n14110_), .Y(u2__abc_52138_new_n14112_));
NAND2X1 NAND2X1_1599 ( .A(u2__abc_52138_new_n14119_), .B(u2__abc_52138_new_n14118_), .Y(u2__abc_52138_new_n14120_));
NAND2X1 NAND2X1_16 ( .A(aNan), .B(\a[15] ), .Y(_abc_65734_new_n876_));
NAND2X1 NAND2X1_160 ( .A(\a[47] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1289_));
NAND2X1 NAND2X1_1600 ( .A(u2__abc_52138_new_n14127_), .B(u2__abc_52138_new_n14126_), .Y(u2__abc_52138_new_n14128_));
NAND2X1 NAND2X1_1601 ( .A(u2__abc_52138_new_n14135_), .B(u2__abc_52138_new_n14134_), .Y(u2__abc_52138_new_n14136_));
NAND2X1 NAND2X1_1602 ( .A(u2__abc_52138_new_n14142_), .B(u2__abc_52138_new_n14141_), .Y(u2__abc_52138_new_n14143_));
NAND2X1 NAND2X1_1603 ( .A(u2__abc_52138_new_n14150_), .B(u2__abc_52138_new_n14149_), .Y(u2__abc_52138_new_n14151_));
NAND2X1 NAND2X1_1604 ( .A(u2__abc_52138_new_n14158_), .B(u2__abc_52138_new_n14157_), .Y(u2__abc_52138_new_n14159_));
NAND2X1 NAND2X1_1605 ( .A(u2__abc_52138_new_n14166_), .B(u2__abc_52138_new_n14165_), .Y(u2__abc_52138_new_n14167_));
NAND2X1 NAND2X1_1606 ( .A(u2__abc_52138_new_n14173_), .B(u2__abc_52138_new_n14172_), .Y(u2__abc_52138_new_n14174_));
NAND2X1 NAND2X1_1607 ( .A(u2__abc_52138_new_n14181_), .B(u2__abc_52138_new_n14180_), .Y(u2__abc_52138_new_n14182_));
NAND2X1 NAND2X1_1608 ( .A(u2__abc_52138_new_n14189_), .B(u2__abc_52138_new_n14188_), .Y(u2__abc_52138_new_n14190_));
NAND2X1 NAND2X1_1609 ( .A(u2__abc_52138_new_n14197_), .B(u2__abc_52138_new_n14196_), .Y(u2__abc_52138_new_n14198_));
NAND2X1 NAND2X1_161 ( .A(\a[112] ), .B(\a[49] ), .Y(_abc_65734_new_n1291_));
NAND2X1 NAND2X1_1610 ( .A(u2__abc_52138_new_n14204_), .B(u2__abc_52138_new_n14203_), .Y(u2__abc_52138_new_n14205_));
NAND2X1 NAND2X1_1611 ( .A(u2__abc_52138_new_n14212_), .B(u2__abc_52138_new_n14211_), .Y(u2__abc_52138_new_n14213_));
NAND2X1 NAND2X1_1612 ( .A(u2__abc_52138_new_n14220_), .B(u2__abc_52138_new_n14219_), .Y(u2__abc_52138_new_n14221_));
NAND2X1 NAND2X1_1613 ( .A(u2__abc_52138_new_n14228_), .B(u2__abc_52138_new_n14227_), .Y(u2__abc_52138_new_n14229_));
NAND2X1 NAND2X1_1614 ( .A(u2__abc_52138_new_n14235_), .B(u2__abc_52138_new_n14234_), .Y(u2__abc_52138_new_n14236_));
NAND2X1 NAND2X1_1615 ( .A(u2__abc_52138_new_n14243_), .B(u2__abc_52138_new_n14242_), .Y(u2__abc_52138_new_n14244_));
NAND2X1 NAND2X1_1616 ( .A(u2__abc_52138_new_n14251_), .B(u2__abc_52138_new_n14250_), .Y(u2__abc_52138_new_n14252_));
NAND2X1 NAND2X1_1617 ( .A(u2__abc_52138_new_n14259_), .B(u2__abc_52138_new_n14258_), .Y(u2__abc_52138_new_n14260_));
NAND2X1 NAND2X1_1618 ( .A(u2__abc_52138_new_n14266_), .B(u2__abc_52138_new_n14265_), .Y(u2__abc_52138_new_n14267_));
NAND2X1 NAND2X1_1619 ( .A(u2__abc_52138_new_n14274_), .B(u2__abc_52138_new_n14273_), .Y(u2__abc_52138_new_n14275_));
NAND2X1 NAND2X1_162 ( .A(\a[49] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1294_));
NAND2X1 NAND2X1_1620 ( .A(u2__abc_52138_new_n14282_), .B(u2__abc_52138_new_n14281_), .Y(u2__abc_52138_new_n14283_));
NAND2X1 NAND2X1_1621 ( .A(u2__abc_52138_new_n14290_), .B(u2__abc_52138_new_n14289_), .Y(u2__abc_52138_new_n14291_));
NAND2X1 NAND2X1_1622 ( .A(u2__abc_52138_new_n14297_), .B(u2__abc_52138_new_n14296_), .Y(u2__abc_52138_new_n14298_));
NAND2X1 NAND2X1_1623 ( .A(u2__abc_52138_new_n14305_), .B(u2__abc_52138_new_n14304_), .Y(u2__abc_52138_new_n14306_));
NAND2X1 NAND2X1_1624 ( .A(u2__abc_52138_new_n14313_), .B(u2__abc_52138_new_n14312_), .Y(u2__abc_52138_new_n14314_));
NAND2X1 NAND2X1_1625 ( .A(u2__abc_52138_new_n14321_), .B(u2__abc_52138_new_n14320_), .Y(u2__abc_52138_new_n14322_));
NAND2X1 NAND2X1_1626 ( .A(u2__abc_52138_new_n14328_), .B(u2__abc_52138_new_n14327_), .Y(u2__abc_52138_new_n14329_));
NAND2X1 NAND2X1_1627 ( .A(u2__abc_52138_new_n14336_), .B(u2__abc_52138_new_n14335_), .Y(u2__abc_52138_new_n14337_));
NAND2X1 NAND2X1_1628 ( .A(u2__abc_52138_new_n14344_), .B(u2__abc_52138_new_n14343_), .Y(u2__abc_52138_new_n14345_));
NAND2X1 NAND2X1_1629 ( .A(u2__abc_52138_new_n14352_), .B(u2__abc_52138_new_n14351_), .Y(u2__abc_52138_new_n14353_));
NAND2X1 NAND2X1_163 ( .A(\a[112] ), .B(\a[51] ), .Y(_abc_65734_new_n1296_));
NAND2X1 NAND2X1_1630 ( .A(u2__abc_52138_new_n14359_), .B(u2__abc_52138_new_n14358_), .Y(u2__abc_52138_new_n14360_));
NAND2X1 NAND2X1_1631 ( .A(u2__abc_52138_new_n14367_), .B(u2__abc_52138_new_n14366_), .Y(u2__abc_52138_new_n14368_));
NAND2X1 NAND2X1_1632 ( .A(u2__abc_52138_new_n14375_), .B(u2__abc_52138_new_n14374_), .Y(u2__abc_52138_new_n14376_));
NAND2X1 NAND2X1_1633 ( .A(u2__abc_52138_new_n14383_), .B(u2__abc_52138_new_n14382_), .Y(u2__abc_52138_new_n14384_));
NAND2X1 NAND2X1_1634 ( .A(u2__abc_52138_new_n14390_), .B(u2__abc_52138_new_n14389_), .Y(u2__abc_52138_new_n14391_));
NAND2X1 NAND2X1_1635 ( .A(u2__abc_52138_new_n14398_), .B(u2__abc_52138_new_n14397_), .Y(u2__abc_52138_new_n14399_));
NAND2X1 NAND2X1_1636 ( .A(u2__abc_52138_new_n14406_), .B(u2__abc_52138_new_n14405_), .Y(u2__abc_52138_new_n14407_));
NAND2X1 NAND2X1_1637 ( .A(u2__abc_52138_new_n14414_), .B(u2__abc_52138_new_n14413_), .Y(u2__abc_52138_new_n14415_));
NAND2X1 NAND2X1_1638 ( .A(u2__abc_52138_new_n14421_), .B(u2__abc_52138_new_n14420_), .Y(u2__abc_52138_new_n14422_));
NAND2X1 NAND2X1_1639 ( .A(u2__abc_52138_new_n14429_), .B(u2__abc_52138_new_n14428_), .Y(u2__abc_52138_new_n14430_));
NAND2X1 NAND2X1_164 ( .A(\a[51] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1299_));
NAND2X1 NAND2X1_1640 ( .A(u2__abc_52138_new_n14437_), .B(u2__abc_52138_new_n14436_), .Y(u2__abc_52138_new_n14438_));
NAND2X1 NAND2X1_1641 ( .A(u2__abc_52138_new_n14445_), .B(u2__abc_52138_new_n14444_), .Y(u2__abc_52138_new_n14446_));
NAND2X1 NAND2X1_1642 ( .A(u2__abc_52138_new_n14452_), .B(u2__abc_52138_new_n14451_), .Y(u2__abc_52138_new_n14453_));
NAND2X1 NAND2X1_1643 ( .A(u2__abc_52138_new_n14460_), .B(u2__abc_52138_new_n14459_), .Y(u2__abc_52138_new_n14461_));
NAND2X1 NAND2X1_1644 ( .A(u2__abc_52138_new_n14468_), .B(u2__abc_52138_new_n14467_), .Y(u2__abc_52138_new_n14469_));
NAND2X1 NAND2X1_1645 ( .A(u2__abc_52138_new_n14476_), .B(u2__abc_52138_new_n14475_), .Y(u2__abc_52138_new_n14477_));
NAND2X1 NAND2X1_1646 ( .A(u2__abc_52138_new_n14483_), .B(u2__abc_52138_new_n14482_), .Y(u2__abc_52138_new_n14484_));
NAND2X1 NAND2X1_1647 ( .A(u2__abc_52138_new_n14491_), .B(u2__abc_52138_new_n14490_), .Y(u2__abc_52138_new_n14492_));
NAND2X1 NAND2X1_1648 ( .A(u2__abc_52138_new_n14499_), .B(u2__abc_52138_new_n14498_), .Y(u2__abc_52138_new_n14500_));
NAND2X1 NAND2X1_1649 ( .A(u2__abc_52138_new_n14507_), .B(u2__abc_52138_new_n14506_), .Y(u2__abc_52138_new_n14508_));
NAND2X1 NAND2X1_165 ( .A(\a[112] ), .B(\a[53] ), .Y(_abc_65734_new_n1301_));
NAND2X1 NAND2X1_1650 ( .A(u2__abc_52138_new_n14514_), .B(u2__abc_52138_new_n14513_), .Y(u2__abc_52138_new_n14515_));
NAND2X1 NAND2X1_1651 ( .A(u2__abc_52138_new_n14522_), .B(u2__abc_52138_new_n14521_), .Y(u2__abc_52138_new_n14523_));
NAND2X1 NAND2X1_1652 ( .A(u2__abc_52138_new_n14530_), .B(u2__abc_52138_new_n14529_), .Y(u2__abc_52138_new_n14531_));
NAND2X1 NAND2X1_1653 ( .A(u2__abc_52138_new_n14538_), .B(u2__abc_52138_new_n14537_), .Y(u2__abc_52138_new_n14539_));
NAND2X1 NAND2X1_1654 ( .A(u2__abc_52138_new_n14545_), .B(u2__abc_52138_new_n14544_), .Y(u2__abc_52138_new_n14546_));
NAND2X1 NAND2X1_1655 ( .A(u2__abc_52138_new_n14553_), .B(u2__abc_52138_new_n14552_), .Y(u2__abc_52138_new_n14554_));
NAND2X1 NAND2X1_1656 ( .A(u2__abc_52138_new_n14561_), .B(u2__abc_52138_new_n14560_), .Y(u2__abc_52138_new_n14562_));
NAND2X1 NAND2X1_1657 ( .A(u2__abc_52138_new_n14569_), .B(u2__abc_52138_new_n14568_), .Y(u2__abc_52138_new_n14570_));
NAND2X1 NAND2X1_1658 ( .A(u2__abc_52138_new_n14576_), .B(u2__abc_52138_new_n14575_), .Y(u2__abc_52138_new_n14577_));
NAND2X1 NAND2X1_1659 ( .A(u2__abc_52138_new_n14584_), .B(u2__abc_52138_new_n14583_), .Y(u2__abc_52138_new_n14585_));
NAND2X1 NAND2X1_166 ( .A(\a[53] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1304_));
NAND2X1 NAND2X1_1660 ( .A(u2__abc_52138_new_n14592_), .B(u2__abc_52138_new_n14591_), .Y(u2__abc_52138_new_n14593_));
NAND2X1 NAND2X1_1661 ( .A(u2__abc_52138_new_n14600_), .B(u2__abc_52138_new_n14599_), .Y(u2__abc_52138_new_n14601_));
NAND2X1 NAND2X1_1662 ( .A(u2__abc_52138_new_n14607_), .B(u2__abc_52138_new_n14606_), .Y(u2__abc_52138_new_n14608_));
NAND2X1 NAND2X1_1663 ( .A(u2__abc_52138_new_n14616_), .B(u2__abc_52138_new_n14614_), .Y(u2__abc_52138_new_n14617_));
NAND2X1 NAND2X1_1664 ( .A(u2__abc_52138_new_n14624_), .B(u2__abc_52138_new_n14623_), .Y(u2__abc_52138_new_n14625_));
NAND2X1 NAND2X1_1665 ( .A(u2__abc_52138_new_n14632_), .B(u2__abc_52138_new_n14631_), .Y(u2__abc_52138_new_n14633_));
NAND2X1 NAND2X1_1666 ( .A(u2__abc_52138_new_n14639_), .B(u2__abc_52138_new_n14638_), .Y(u2__abc_52138_new_n14640_));
NAND2X1 NAND2X1_1667 ( .A(u2__abc_52138_new_n14647_), .B(u2__abc_52138_new_n14646_), .Y(u2__abc_52138_new_n14648_));
NAND2X1 NAND2X1_1668 ( .A(u2__abc_52138_new_n14655_), .B(u2__abc_52138_new_n14654_), .Y(u2__abc_52138_new_n14656_));
NAND2X1 NAND2X1_1669 ( .A(u2__abc_52138_new_n14663_), .B(u2__abc_52138_new_n14662_), .Y(u2__abc_52138_new_n14664_));
NAND2X1 NAND2X1_167 ( .A(\a[112] ), .B(\a[55] ), .Y(_abc_65734_new_n1306_));
NAND2X1 NAND2X1_1670 ( .A(u2__abc_52138_new_n14670_), .B(u2__abc_52138_new_n14669_), .Y(u2__abc_52138_new_n14671_));
NAND2X1 NAND2X1_1671 ( .A(u2__abc_52138_new_n14678_), .B(u2__abc_52138_new_n14677_), .Y(u2__abc_52138_new_n14679_));
NAND2X1 NAND2X1_1672 ( .A(u2__abc_52138_new_n14686_), .B(u2__abc_52138_new_n14685_), .Y(u2__abc_52138_new_n14687_));
NAND2X1 NAND2X1_1673 ( .A(u2__abc_52138_new_n14694_), .B(u2__abc_52138_new_n14693_), .Y(u2__abc_52138_new_n14695_));
NAND2X1 NAND2X1_1674 ( .A(u2__abc_52138_new_n14701_), .B(u2__abc_52138_new_n14700_), .Y(u2__abc_52138_new_n14702_));
NAND2X1 NAND2X1_1675 ( .A(u2__abc_52138_new_n14709_), .B(u2__abc_52138_new_n14708_), .Y(u2__abc_52138_new_n14710_));
NAND2X1 NAND2X1_1676 ( .A(u2__abc_52138_new_n14717_), .B(u2__abc_52138_new_n14716_), .Y(u2__abc_52138_new_n14718_));
NAND2X1 NAND2X1_1677 ( .A(u2__abc_52138_new_n14725_), .B(u2__abc_52138_new_n14724_), .Y(u2__abc_52138_new_n14726_));
NAND2X1 NAND2X1_1678 ( .A(u2__abc_52138_new_n14732_), .B(u2__abc_52138_new_n14731_), .Y(u2__abc_52138_new_n14733_));
NAND2X1 NAND2X1_1679 ( .A(u2__abc_52138_new_n14740_), .B(u2__abc_52138_new_n14739_), .Y(u2__abc_52138_new_n14741_));
NAND2X1 NAND2X1_168 ( .A(\a[55] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1309_));
NAND2X1 NAND2X1_1680 ( .A(u2__abc_52138_new_n14748_), .B(u2__abc_52138_new_n14747_), .Y(u2__abc_52138_new_n14749_));
NAND2X1 NAND2X1_1681 ( .A(u2__abc_52138_new_n14756_), .B(u2__abc_52138_new_n14755_), .Y(u2__abc_52138_new_n14757_));
NAND2X1 NAND2X1_1682 ( .A(u2__abc_52138_new_n14763_), .B(u2__abc_52138_new_n14762_), .Y(u2__abc_52138_new_n14764_));
NAND2X1 NAND2X1_1683 ( .A(u2__abc_52138_new_n14771_), .B(u2__abc_52138_new_n14770_), .Y(u2__abc_52138_new_n14772_));
NAND2X1 NAND2X1_1684 ( .A(u2__abc_52138_new_n14779_), .B(u2__abc_52138_new_n14778_), .Y(u2__abc_52138_new_n14780_));
NAND2X1 NAND2X1_1685 ( .A(u2__abc_52138_new_n14787_), .B(u2__abc_52138_new_n14786_), .Y(u2__abc_52138_new_n14788_));
NAND2X1 NAND2X1_1686 ( .A(u2__abc_52138_new_n14794_), .B(u2__abc_52138_new_n14793_), .Y(u2__abc_52138_new_n14795_));
NAND2X1 NAND2X1_1687 ( .A(u2__abc_52138_new_n14802_), .B(u2__abc_52138_new_n14801_), .Y(u2__abc_52138_new_n14803_));
NAND2X1 NAND2X1_1688 ( .A(u2__abc_52138_new_n14810_), .B(u2__abc_52138_new_n14809_), .Y(u2__abc_52138_new_n14811_));
NAND2X1 NAND2X1_1689 ( .A(u2__abc_52138_new_n14818_), .B(u2__abc_52138_new_n14817_), .Y(u2__abc_52138_new_n14819_));
NAND2X1 NAND2X1_169 ( .A(\a[112] ), .B(\a[57] ), .Y(_abc_65734_new_n1311_));
NAND2X1 NAND2X1_1690 ( .A(u2__abc_52138_new_n14825_), .B(u2__abc_52138_new_n14824_), .Y(u2__abc_52138_new_n14826_));
NAND2X1 NAND2X1_1691 ( .A(u2__abc_52138_new_n14833_), .B(u2__abc_52138_new_n14832_), .Y(u2__abc_52138_new_n14834_));
NAND2X1 NAND2X1_1692 ( .A(u2__abc_52138_new_n14841_), .B(u2__abc_52138_new_n14840_), .Y(u2__abc_52138_new_n14842_));
NAND2X1 NAND2X1_1693 ( .A(u2__abc_52138_new_n14849_), .B(u2__abc_52138_new_n14848_), .Y(u2__abc_52138_new_n14850_));
NAND2X1 NAND2X1_1694 ( .A(u2__abc_52138_new_n14856_), .B(u2__abc_52138_new_n14855_), .Y(u2__abc_52138_new_n14857_));
NAND2X1 NAND2X1_1695 ( .A(u2__abc_52138_new_n14864_), .B(u2__abc_52138_new_n14863_), .Y(u2__abc_52138_new_n14865_));
NAND2X1 NAND2X1_1696 ( .A(u2__abc_52138_new_n14872_), .B(u2__abc_52138_new_n14871_), .Y(u2__abc_52138_new_n14873_));
NAND2X1 NAND2X1_1697 ( .A(u2__abc_52138_new_n14880_), .B(u2__abc_52138_new_n14879_), .Y(u2__abc_52138_new_n14881_));
NAND2X1 NAND2X1_1698 ( .A(u2__abc_52138_new_n14887_), .B(u2__abc_52138_new_n14886_), .Y(u2__abc_52138_new_n14888_));
NAND2X1 NAND2X1_1699 ( .A(u2__abc_52138_new_n14895_), .B(u2__abc_52138_new_n14894_), .Y(u2__abc_52138_new_n14896_));
NAND2X1 NAND2X1_17 ( .A(aNan), .B(\a[16] ), .Y(_abc_65734_new_n879_));
NAND2X1 NAND2X1_170 ( .A(\a[57] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1314_));
NAND2X1 NAND2X1_1700 ( .A(u2__abc_52138_new_n14903_), .B(u2__abc_52138_new_n14902_), .Y(u2__abc_52138_new_n14904_));
NAND2X1 NAND2X1_1701 ( .A(u2__abc_52138_new_n14911_), .B(u2__abc_52138_new_n14910_), .Y(u2__abc_52138_new_n14912_));
NAND2X1 NAND2X1_1702 ( .A(u2__abc_52138_new_n14918_), .B(u2__abc_52138_new_n14917_), .Y(u2__abc_52138_new_n14919_));
NAND2X1 NAND2X1_1703 ( .A(u2__abc_52138_new_n14926_), .B(u2__abc_52138_new_n14925_), .Y(u2__abc_52138_new_n14927_));
NAND2X1 NAND2X1_1704 ( .A(u2__abc_52138_new_n14934_), .B(u2__abc_52138_new_n14933_), .Y(u2__abc_52138_new_n14935_));
NAND2X1 NAND2X1_1705 ( .A(u2__abc_52138_new_n14942_), .B(u2__abc_52138_new_n14941_), .Y(u2__abc_52138_new_n14943_));
NAND2X1 NAND2X1_1706 ( .A(u2__abc_52138_new_n14949_), .B(u2__abc_52138_new_n14948_), .Y(u2__abc_52138_new_n14950_));
NAND2X1 NAND2X1_1707 ( .A(u2__abc_52138_new_n14957_), .B(u2__abc_52138_new_n14956_), .Y(u2__abc_52138_new_n14958_));
NAND2X1 NAND2X1_1708 ( .A(u2__abc_52138_new_n14965_), .B(u2__abc_52138_new_n14964_), .Y(u2__abc_52138_new_n14966_));
NAND2X1 NAND2X1_1709 ( .A(u2__abc_52138_new_n14973_), .B(u2__abc_52138_new_n14972_), .Y(u2__abc_52138_new_n14974_));
NAND2X1 NAND2X1_171 ( .A(\a[112] ), .B(\a[59] ), .Y(_abc_65734_new_n1316_));
NAND2X1 NAND2X1_1710 ( .A(u2__abc_52138_new_n14980_), .B(u2__abc_52138_new_n14979_), .Y(u2__abc_52138_new_n14981_));
NAND2X1 NAND2X1_1711 ( .A(u2__abc_52138_new_n14988_), .B(u2__abc_52138_new_n14987_), .Y(u2__abc_52138_new_n14989_));
NAND2X1 NAND2X1_1712 ( .A(u2__abc_52138_new_n14996_), .B(u2__abc_52138_new_n14995_), .Y(u2__abc_52138_new_n14997_));
NAND2X1 NAND2X1_1713 ( .A(u2__abc_52138_new_n15004_), .B(u2__abc_52138_new_n15003_), .Y(u2__abc_52138_new_n15005_));
NAND2X1 NAND2X1_1714 ( .A(u2__abc_52138_new_n15011_), .B(u2__abc_52138_new_n15010_), .Y(u2__abc_52138_new_n15012_));
NAND2X1 NAND2X1_1715 ( .A(u2__abc_52138_new_n15019_), .B(u2__abc_52138_new_n15018_), .Y(u2__abc_52138_new_n15020_));
NAND2X1 NAND2X1_1716 ( .A(u2__abc_52138_new_n15027_), .B(u2__abc_52138_new_n15026_), .Y(u2__abc_52138_new_n15028_));
NAND2X1 NAND2X1_1717 ( .A(u2__abc_52138_new_n15035_), .B(u2__abc_52138_new_n15034_), .Y(u2__abc_52138_new_n15036_));
NAND2X1 NAND2X1_1718 ( .A(u2__abc_52138_new_n15042_), .B(u2__abc_52138_new_n15041_), .Y(u2__abc_52138_new_n15043_));
NAND2X1 NAND2X1_1719 ( .A(u2__abc_52138_new_n15050_), .B(u2__abc_52138_new_n15049_), .Y(u2__abc_52138_new_n15051_));
NAND2X1 NAND2X1_172 ( .A(\a[59] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1319_));
NAND2X1 NAND2X1_1720 ( .A(u2__abc_52138_new_n15058_), .B(u2__abc_52138_new_n15057_), .Y(u2__abc_52138_new_n15059_));
NAND2X1 NAND2X1_1721 ( .A(u2__abc_52138_new_n15066_), .B(u2__abc_52138_new_n15065_), .Y(u2__abc_52138_new_n15067_));
NAND2X1 NAND2X1_1722 ( .A(u2__abc_52138_new_n15073_), .B(u2__abc_52138_new_n15072_), .Y(u2__abc_52138_new_n15074_));
NAND2X1 NAND2X1_1723 ( .A(u2__abc_52138_new_n15081_), .B(u2__abc_52138_new_n15080_), .Y(u2__abc_52138_new_n15082_));
NAND2X1 NAND2X1_1724 ( .A(u2__abc_52138_new_n15089_), .B(u2__abc_52138_new_n15088_), .Y(u2__abc_52138_new_n15090_));
NAND2X1 NAND2X1_1725 ( .A(u2__abc_52138_new_n15097_), .B(u2__abc_52138_new_n15096_), .Y(u2__abc_52138_new_n15098_));
NAND2X1 NAND2X1_1726 ( .A(u2__abc_52138_new_n15104_), .B(u2__abc_52138_new_n15103_), .Y(u2__abc_52138_new_n15105_));
NAND2X1 NAND2X1_1727 ( .A(u2__abc_52138_new_n15112_), .B(u2__abc_52138_new_n15111_), .Y(u2__abc_52138_new_n15113_));
NAND2X1 NAND2X1_1728 ( .A(u2__abc_52138_new_n15120_), .B(u2__abc_52138_new_n15119_), .Y(u2__abc_52138_new_n15121_));
NAND2X1 NAND2X1_1729 ( .A(u2__abc_52138_new_n15128_), .B(u2__abc_52138_new_n15127_), .Y(u2__abc_52138_new_n15129_));
NAND2X1 NAND2X1_173 ( .A(\a[112] ), .B(\a[61] ), .Y(_abc_65734_new_n1321_));
NAND2X1 NAND2X1_1730 ( .A(u2__abc_52138_new_n15135_), .B(u2__abc_52138_new_n15134_), .Y(u2__abc_52138_new_n15136_));
NAND2X1 NAND2X1_1731 ( .A(u2__abc_52138_new_n15143_), .B(u2__abc_52138_new_n15142_), .Y(u2__abc_52138_new_n15144_));
NAND2X1 NAND2X1_1732 ( .A(u2__abc_52138_new_n15151_), .B(u2__abc_52138_new_n15150_), .Y(u2__abc_52138_new_n15152_));
NAND2X1 NAND2X1_1733 ( .A(u2__abc_52138_new_n15159_), .B(u2__abc_52138_new_n15158_), .Y(u2__abc_52138_new_n15160_));
NAND2X1 NAND2X1_1734 ( .A(u2__abc_52138_new_n15166_), .B(u2__abc_52138_new_n15165_), .Y(u2__abc_52138_new_n15167_));
NAND2X1 NAND2X1_1735 ( .A(u2__abc_52138_new_n15174_), .B(u2__abc_52138_new_n15173_), .Y(u2__abc_52138_new_n15175_));
NAND2X1 NAND2X1_1736 ( .A(u2__abc_52138_new_n15182_), .B(u2__abc_52138_new_n15181_), .Y(u2__abc_52138_new_n15183_));
NAND2X1 NAND2X1_1737 ( .A(u2__abc_52138_new_n15190_), .B(u2__abc_52138_new_n15189_), .Y(u2__abc_52138_new_n15191_));
NAND2X1 NAND2X1_1738 ( .A(u2__abc_52138_new_n15197_), .B(u2__abc_52138_new_n15196_), .Y(u2__abc_52138_new_n15198_));
NAND2X1 NAND2X1_1739 ( .A(u2__abc_52138_new_n15205_), .B(u2__abc_52138_new_n15204_), .Y(u2__abc_52138_new_n15206_));
NAND2X1 NAND2X1_174 ( .A(\a[61] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1324_));
NAND2X1 NAND2X1_1740 ( .A(u2__abc_52138_new_n15213_), .B(u2__abc_52138_new_n15212_), .Y(u2__abc_52138_new_n15214_));
NAND2X1 NAND2X1_1741 ( .A(u2__abc_52138_new_n15221_), .B(u2__abc_52138_new_n15220_), .Y(u2__abc_52138_new_n15222_));
NAND2X1 NAND2X1_1742 ( .A(u2__abc_52138_new_n15228_), .B(u2__abc_52138_new_n15227_), .Y(u2__abc_52138_new_n15229_));
NAND2X1 NAND2X1_1743 ( .A(u2__abc_52138_new_n15236_), .B(u2__abc_52138_new_n15235_), .Y(u2__abc_52138_new_n15237_));
NAND2X1 NAND2X1_1744 ( .A(u2__abc_52138_new_n15244_), .B(u2__abc_52138_new_n15243_), .Y(u2__abc_52138_new_n15245_));
NAND2X1 NAND2X1_1745 ( .A(u2__abc_52138_new_n15252_), .B(u2__abc_52138_new_n15251_), .Y(u2__abc_52138_new_n15253_));
NAND2X1 NAND2X1_1746 ( .A(u2__abc_52138_new_n15259_), .B(u2__abc_52138_new_n15258_), .Y(u2__abc_52138_new_n15260_));
NAND2X1 NAND2X1_1747 ( .A(u2__abc_52138_new_n15267_), .B(u2__abc_52138_new_n15266_), .Y(u2__abc_52138_new_n15268_));
NAND2X1 NAND2X1_1748 ( .A(u2__abc_52138_new_n15275_), .B(u2__abc_52138_new_n15274_), .Y(u2__abc_52138_new_n15276_));
NAND2X1 NAND2X1_1749 ( .A(u2__abc_52138_new_n15283_), .B(u2__abc_52138_new_n15282_), .Y(u2__abc_52138_new_n15284_));
NAND2X1 NAND2X1_175 ( .A(\a[112] ), .B(\a[63] ), .Y(_abc_65734_new_n1326_));
NAND2X1 NAND2X1_1750 ( .A(u2__abc_52138_new_n15290_), .B(u2__abc_52138_new_n15289_), .Y(u2__abc_52138_new_n15291_));
NAND2X1 NAND2X1_1751 ( .A(u2__abc_52138_new_n15298_), .B(u2__abc_52138_new_n15297_), .Y(u2__abc_52138_new_n15299_));
NAND2X1 NAND2X1_1752 ( .A(u2__abc_52138_new_n15306_), .B(u2__abc_52138_new_n15305_), .Y(u2__abc_52138_new_n15307_));
NAND2X1 NAND2X1_1753 ( .A(u2__abc_52138_new_n15314_), .B(u2__abc_52138_new_n15313_), .Y(u2__abc_52138_new_n15315_));
NAND2X1 NAND2X1_1754 ( .A(u2__abc_52138_new_n15321_), .B(u2__abc_52138_new_n15320_), .Y(u2__abc_52138_new_n15322_));
NAND2X1 NAND2X1_1755 ( .A(u2__abc_52138_new_n15329_), .B(u2__abc_52138_new_n15328_), .Y(u2__abc_52138_new_n15330_));
NAND2X1 NAND2X1_1756 ( .A(u2__abc_52138_new_n15337_), .B(u2__abc_52138_new_n15336_), .Y(u2__abc_52138_new_n15338_));
NAND2X1 NAND2X1_1757 ( .A(u2__abc_52138_new_n15345_), .B(u2__abc_52138_new_n15344_), .Y(u2__abc_52138_new_n15346_));
NAND2X1 NAND2X1_1758 ( .A(u2__abc_52138_new_n15352_), .B(u2__abc_52138_new_n15351_), .Y(u2__abc_52138_new_n15353_));
NAND2X1 NAND2X1_1759 ( .A(u2__abc_52138_new_n15360_), .B(u2__abc_52138_new_n15359_), .Y(u2__abc_52138_new_n15361_));
NAND2X1 NAND2X1_176 ( .A(\a[63] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1329_));
NAND2X1 NAND2X1_1760 ( .A(u2__abc_52138_new_n15368_), .B(u2__abc_52138_new_n15367_), .Y(u2__abc_52138_new_n15369_));
NAND2X1 NAND2X1_1761 ( .A(u2__abc_52138_new_n15376_), .B(u2__abc_52138_new_n15375_), .Y(u2__abc_52138_new_n15377_));
NAND2X1 NAND2X1_1762 ( .A(u2__abc_52138_new_n15383_), .B(u2__abc_52138_new_n15382_), .Y(u2__abc_52138_new_n15384_));
NAND2X1 NAND2X1_1763 ( .A(u2__abc_52138_new_n15391_), .B(u2__abc_52138_new_n15390_), .Y(u2__abc_52138_new_n15392_));
NAND2X1 NAND2X1_1764 ( .A(u2__abc_52138_new_n15399_), .B(u2__abc_52138_new_n15398_), .Y(u2__abc_52138_new_n15400_));
NAND2X1 NAND2X1_1765 ( .A(u2__abc_52138_new_n15407_), .B(u2__abc_52138_new_n15406_), .Y(u2__abc_52138_new_n15408_));
NAND2X1 NAND2X1_1766 ( .A(u2__abc_52138_new_n15414_), .B(u2__abc_52138_new_n15413_), .Y(u2__abc_52138_new_n15415_));
NAND2X1 NAND2X1_1767 ( .A(u2__abc_52138_new_n15422_), .B(u2__abc_52138_new_n15421_), .Y(u2__abc_52138_new_n15423_));
NAND2X1 NAND2X1_1768 ( .A(u2__abc_52138_new_n15430_), .B(u2__abc_52138_new_n15429_), .Y(u2__abc_52138_new_n15431_));
NAND2X1 NAND2X1_1769 ( .A(u2__abc_52138_new_n15438_), .B(u2__abc_52138_new_n15437_), .Y(u2__abc_52138_new_n15439_));
NAND2X1 NAND2X1_177 ( .A(\a[112] ), .B(\a[65] ), .Y(_abc_65734_new_n1331_));
NAND2X1 NAND2X1_1770 ( .A(u2__abc_52138_new_n15445_), .B(u2__abc_52138_new_n15444_), .Y(u2__abc_52138_new_n15446_));
NAND2X1 NAND2X1_1771 ( .A(u2__abc_52138_new_n15453_), .B(u2__abc_52138_new_n15452_), .Y(u2__abc_52138_new_n15454_));
NAND2X1 NAND2X1_1772 ( .A(u2__abc_52138_new_n15461_), .B(u2__abc_52138_new_n15460_), .Y(u2__abc_52138_new_n15462_));
NAND2X1 NAND2X1_1773 ( .A(u2__abc_52138_new_n15469_), .B(u2__abc_52138_new_n15468_), .Y(u2__abc_52138_new_n15470_));
NAND2X1 NAND2X1_1774 ( .A(u2__abc_52138_new_n15476_), .B(u2__abc_52138_new_n15475_), .Y(u2__abc_52138_new_n15477_));
NAND2X1 NAND2X1_1775 ( .A(u2__abc_52138_new_n15485_), .B(u2__abc_52138_new_n15483_), .Y(u2__abc_52138_new_n15486_));
NAND2X1 NAND2X1_1776 ( .A(u2__abc_52138_new_n15493_), .B(u2__abc_52138_new_n15492_), .Y(u2__abc_52138_new_n15494_));
NAND2X1 NAND2X1_1777 ( .A(u2__abc_52138_new_n15501_), .B(u2__abc_52138_new_n15500_), .Y(u2__abc_52138_new_n15502_));
NAND2X1 NAND2X1_1778 ( .A(u2__abc_52138_new_n15508_), .B(u2__abc_52138_new_n15507_), .Y(u2__abc_52138_new_n15509_));
NAND2X1 NAND2X1_1779 ( .A(u2__abc_52138_new_n15516_), .B(u2__abc_52138_new_n15515_), .Y(u2__abc_52138_new_n15517_));
NAND2X1 NAND2X1_178 ( .A(\a[65] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1334_));
NAND2X1 NAND2X1_1780 ( .A(u2__abc_52138_new_n15524_), .B(u2__abc_52138_new_n15523_), .Y(u2__abc_52138_new_n15525_));
NAND2X1 NAND2X1_1781 ( .A(u2__abc_52138_new_n15532_), .B(u2__abc_52138_new_n15531_), .Y(u2__abc_52138_new_n15533_));
NAND2X1 NAND2X1_1782 ( .A(u2__abc_52138_new_n15539_), .B(u2__abc_52138_new_n15538_), .Y(u2__abc_52138_new_n15540_));
NAND2X1 NAND2X1_1783 ( .A(u2__abc_52138_new_n15547_), .B(u2__abc_52138_new_n15546_), .Y(u2__abc_52138_new_n15548_));
NAND2X1 NAND2X1_1784 ( .A(u2__abc_52138_new_n15555_), .B(u2__abc_52138_new_n15554_), .Y(u2__abc_52138_new_n15556_));
NAND2X1 NAND2X1_1785 ( .A(u2__abc_52138_new_n15563_), .B(u2__abc_52138_new_n15562_), .Y(u2__abc_52138_new_n15564_));
NAND2X1 NAND2X1_1786 ( .A(u2__abc_52138_new_n15570_), .B(u2__abc_52138_new_n15569_), .Y(u2__abc_52138_new_n15571_));
NAND2X1 NAND2X1_1787 ( .A(u2__abc_52138_new_n15578_), .B(u2__abc_52138_new_n15577_), .Y(u2__abc_52138_new_n15579_));
NAND2X1 NAND2X1_1788 ( .A(u2__abc_52138_new_n15586_), .B(u2__abc_52138_new_n15585_), .Y(u2__abc_52138_new_n15587_));
NAND2X1 NAND2X1_1789 ( .A(u2__abc_52138_new_n15594_), .B(u2__abc_52138_new_n15593_), .Y(u2__abc_52138_new_n15595_));
NAND2X1 NAND2X1_179 ( .A(\a[112] ), .B(\a[67] ), .Y(_abc_65734_new_n1336_));
NAND2X1 NAND2X1_1790 ( .A(u2__abc_52138_new_n15601_), .B(u2__abc_52138_new_n15600_), .Y(u2__abc_52138_new_n15602_));
NAND2X1 NAND2X1_1791 ( .A(u2__abc_52138_new_n15609_), .B(u2__abc_52138_new_n15608_), .Y(u2__abc_52138_new_n15610_));
NAND2X1 NAND2X1_1792 ( .A(u2__abc_52138_new_n15617_), .B(u2__abc_52138_new_n15616_), .Y(u2__abc_52138_new_n15618_));
NAND2X1 NAND2X1_1793 ( .A(u2__abc_52138_new_n15625_), .B(u2__abc_52138_new_n15624_), .Y(u2__abc_52138_new_n15626_));
NAND2X1 NAND2X1_1794 ( .A(u2__abc_52138_new_n15632_), .B(u2__abc_52138_new_n15631_), .Y(u2__abc_52138_new_n15633_));
NAND2X1 NAND2X1_1795 ( .A(u2__abc_52138_new_n15641_), .B(u2__abc_52138_new_n15639_), .Y(u2__abc_52138_new_n15642_));
NAND2X1 NAND2X1_1796 ( .A(u2__abc_52138_new_n15649_), .B(u2__abc_52138_new_n15648_), .Y(u2__abc_52138_new_n15650_));
NAND2X1 NAND2X1_1797 ( .A(u2__abc_52138_new_n15657_), .B(u2__abc_52138_new_n15656_), .Y(u2__abc_52138_new_n15658_));
NAND2X1 NAND2X1_1798 ( .A(u2__abc_52138_new_n15664_), .B(u2__abc_52138_new_n15663_), .Y(u2__abc_52138_new_n15665_));
NAND2X1 NAND2X1_1799 ( .A(u2__abc_52138_new_n15673_), .B(u2__abc_52138_new_n15671_), .Y(u2__abc_52138_new_n15674_));
NAND2X1 NAND2X1_18 ( .A(aNan), .B(\a[17] ), .Y(_abc_65734_new_n882_));
NAND2X1 NAND2X1_180 ( .A(\a[67] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1339_));
NAND2X1 NAND2X1_1800 ( .A(u2__abc_52138_new_n15681_), .B(u2__abc_52138_new_n15680_), .Y(u2__abc_52138_new_n15682_));
NAND2X1 NAND2X1_1801 ( .A(u2__abc_52138_new_n15689_), .B(u2__abc_52138_new_n15688_), .Y(u2__abc_52138_new_n15690_));
NAND2X1 NAND2X1_1802 ( .A(u2__abc_52138_new_n15696_), .B(u2__abc_52138_new_n15695_), .Y(u2__abc_52138_new_n15697_));
NAND2X1 NAND2X1_1803 ( .A(u2__abc_52138_new_n15704_), .B(u2__abc_52138_new_n15703_), .Y(u2__abc_52138_new_n15705_));
NAND2X1 NAND2X1_1804 ( .A(u2__abc_52138_new_n15712_), .B(u2__abc_52138_new_n15711_), .Y(u2__abc_52138_new_n15713_));
NAND2X1 NAND2X1_1805 ( .A(u2__abc_52138_new_n15720_), .B(u2__abc_52138_new_n15719_), .Y(u2__abc_52138_new_n15721_));
NAND2X1 NAND2X1_1806 ( .A(u2__abc_52138_new_n15727_), .B(u2__abc_52138_new_n15726_), .Y(u2__abc_52138_new_n15728_));
NAND2X1 NAND2X1_1807 ( .A(u2__abc_52138_new_n15735_), .B(u2__abc_52138_new_n15734_), .Y(u2__abc_52138_new_n15736_));
NAND2X1 NAND2X1_1808 ( .A(u2__abc_52138_new_n15743_), .B(u2__abc_52138_new_n15742_), .Y(u2__abc_52138_new_n15744_));
NAND2X1 NAND2X1_1809 ( .A(u2__abc_52138_new_n15751_), .B(u2__abc_52138_new_n15750_), .Y(u2__abc_52138_new_n15752_));
NAND2X1 NAND2X1_181 ( .A(\a[112] ), .B(\a[69] ), .Y(_abc_65734_new_n1341_));
NAND2X1 NAND2X1_1810 ( .A(u2__abc_52138_new_n15758_), .B(u2__abc_52138_new_n15757_), .Y(u2__abc_52138_new_n15759_));
NAND2X1 NAND2X1_1811 ( .A(u2__abc_52138_new_n15766_), .B(u2__abc_52138_new_n15765_), .Y(u2__abc_52138_new_n15767_));
NAND2X1 NAND2X1_1812 ( .A(u2__abc_52138_new_n15774_), .B(u2__abc_52138_new_n15773_), .Y(u2__abc_52138_new_n15775_));
NAND2X1 NAND2X1_1813 ( .A(u2__abc_52138_new_n15782_), .B(u2__abc_52138_new_n15781_), .Y(u2__abc_52138_new_n15783_));
NAND2X1 NAND2X1_1814 ( .A(u2__abc_52138_new_n15789_), .B(u2__abc_52138_new_n15788_), .Y(u2__abc_52138_new_n15790_));
NAND2X1 NAND2X1_1815 ( .A(u2__abc_52138_new_n15797_), .B(u2__abc_52138_new_n15796_), .Y(u2__abc_52138_new_n15798_));
NAND2X1 NAND2X1_1816 ( .A(u2__abc_52138_new_n15805_), .B(u2__abc_52138_new_n15804_), .Y(u2__abc_52138_new_n15806_));
NAND2X1 NAND2X1_1817 ( .A(u2__abc_52138_new_n15813_), .B(u2__abc_52138_new_n15812_), .Y(u2__abc_52138_new_n15814_));
NAND2X1 NAND2X1_1818 ( .A(u2__abc_52138_new_n15820_), .B(u2__abc_52138_new_n15819_), .Y(u2__abc_52138_new_n15821_));
NAND2X1 NAND2X1_1819 ( .A(u2__abc_52138_new_n15828_), .B(u2__abc_52138_new_n15827_), .Y(u2__abc_52138_new_n15829_));
NAND2X1 NAND2X1_182 ( .A(\a[69] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1344_));
NAND2X1 NAND2X1_1820 ( .A(u2__abc_52138_new_n15836_), .B(u2__abc_52138_new_n15835_), .Y(u2__abc_52138_new_n15837_));
NAND2X1 NAND2X1_1821 ( .A(u2__abc_52138_new_n15844_), .B(u2__abc_52138_new_n15843_), .Y(u2__abc_52138_new_n15845_));
NAND2X1 NAND2X1_1822 ( .A(u2__abc_52138_new_n15851_), .B(u2__abc_52138_new_n15850_), .Y(u2__abc_52138_new_n15852_));
NAND2X1 NAND2X1_1823 ( .A(u2__abc_52138_new_n15859_), .B(u2__abc_52138_new_n15858_), .Y(u2__abc_52138_new_n15860_));
NAND2X1 NAND2X1_1824 ( .A(u2__abc_52138_new_n15867_), .B(u2__abc_52138_new_n15866_), .Y(u2__abc_52138_new_n15868_));
NAND2X1 NAND2X1_1825 ( .A(u2__abc_52138_new_n15875_), .B(u2__abc_52138_new_n15874_), .Y(u2__abc_52138_new_n15876_));
NAND2X1 NAND2X1_1826 ( .A(u2__abc_52138_new_n15882_), .B(u2__abc_52138_new_n15881_), .Y(u2__abc_52138_new_n15883_));
NAND2X1 NAND2X1_1827 ( .A(u2__abc_52138_new_n15890_), .B(u2__abc_52138_new_n15889_), .Y(u2__abc_52138_new_n15891_));
NAND2X1 NAND2X1_1828 ( .A(u2__abc_52138_new_n15898_), .B(u2__abc_52138_new_n15897_), .Y(u2__abc_52138_new_n15899_));
NAND2X1 NAND2X1_1829 ( .A(u2__abc_52138_new_n15906_), .B(u2__abc_52138_new_n15905_), .Y(u2__abc_52138_new_n15907_));
NAND2X1 NAND2X1_183 ( .A(\a[112] ), .B(\a[71] ), .Y(_abc_65734_new_n1346_));
NAND2X1 NAND2X1_1830 ( .A(u2__abc_52138_new_n15914_), .B(u2__abc_52138_new_n15912_), .Y(u2__abc_52138_new_n15915_));
NAND2X1 NAND2X1_1831 ( .A(u2__abc_52138_new_n15922_), .B(u2__abc_52138_new_n15921_), .Y(u2__abc_52138_new_n15923_));
NAND2X1 NAND2X1_1832 ( .A(u2__abc_52138_new_n15930_), .B(u2__abc_52138_new_n15929_), .Y(u2__abc_52138_new_n15931_));
NAND2X1 NAND2X1_1833 ( .A(u2__abc_52138_new_n15938_), .B(u2__abc_52138_new_n15937_), .Y(u2__abc_52138_new_n15939_));
NAND2X1 NAND2X1_1834 ( .A(u2__abc_52138_new_n15945_), .B(u2__abc_52138_new_n15944_), .Y(u2__abc_52138_new_n15946_));
NAND2X1 NAND2X1_1835 ( .A(u2__abc_52138_new_n15953_), .B(u2__abc_52138_new_n15952_), .Y(u2__abc_52138_new_n15954_));
NAND2X1 NAND2X1_1836 ( .A(u2__abc_52138_new_n15961_), .B(u2__abc_52138_new_n15960_), .Y(u2__abc_52138_new_n15962_));
NAND2X1 NAND2X1_1837 ( .A(u2__abc_52138_new_n15969_), .B(u2__abc_52138_new_n15968_), .Y(u2__abc_52138_new_n15970_));
NAND2X1 NAND2X1_1838 ( .A(u2__abc_52138_new_n15976_), .B(u2__abc_52138_new_n15975_), .Y(u2__abc_52138_new_n15977_));
NAND2X1 NAND2X1_1839 ( .A(u2__abc_52138_new_n15984_), .B(u2__abc_52138_new_n15983_), .Y(u2__abc_52138_new_n15985_));
NAND2X1 NAND2X1_184 ( .A(\a[71] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1349_));
NAND2X1 NAND2X1_1840 ( .A(u2__abc_52138_new_n15992_), .B(u2__abc_52138_new_n15991_), .Y(u2__abc_52138_new_n15993_));
NAND2X1 NAND2X1_1841 ( .A(u2__abc_52138_new_n16000_), .B(u2__abc_52138_new_n15999_), .Y(u2__abc_52138_new_n16001_));
NAND2X1 NAND2X1_1842 ( .A(u2__abc_52138_new_n16007_), .B(u2__abc_52138_new_n16006_), .Y(u2__abc_52138_new_n16008_));
NAND2X1 NAND2X1_1843 ( .A(u2__abc_52138_new_n16015_), .B(u2__abc_52138_new_n16014_), .Y(u2__abc_52138_new_n16016_));
NAND2X1 NAND2X1_1844 ( .A(u2__abc_52138_new_n16023_), .B(u2__abc_52138_new_n16022_), .Y(u2__abc_52138_new_n16024_));
NAND2X1 NAND2X1_1845 ( .A(u2__abc_52138_new_n16031_), .B(u2__abc_52138_new_n16030_), .Y(u2__abc_52138_new_n16032_));
NAND2X1 NAND2X1_1846 ( .A(u2__abc_52138_new_n16038_), .B(u2__abc_52138_new_n16037_), .Y(u2__abc_52138_new_n16039_));
NAND2X1 NAND2X1_1847 ( .A(u2__abc_52138_new_n16046_), .B(u2__abc_52138_new_n16045_), .Y(u2__abc_52138_new_n16047_));
NAND2X1 NAND2X1_1848 ( .A(u2__abc_52138_new_n16054_), .B(u2__abc_52138_new_n16053_), .Y(u2__abc_52138_new_n16055_));
NAND2X1 NAND2X1_1849 ( .A(u2__abc_52138_new_n16062_), .B(u2__abc_52138_new_n16061_), .Y(u2__abc_52138_new_n16063_));
NAND2X1 NAND2X1_185 ( .A(\a[112] ), .B(\a[73] ), .Y(_abc_65734_new_n1351_));
NAND2X1 NAND2X1_1850 ( .A(u2__abc_52138_new_n16069_), .B(u2__abc_52138_new_n16068_), .Y(u2__abc_52138_new_n16070_));
NAND2X1 NAND2X1_1851 ( .A(u2__abc_52138_new_n16078_), .B(u2__abc_52138_new_n16076_), .Y(u2__abc_52138_new_n16079_));
NAND2X1 NAND2X1_1852 ( .A(u2__abc_52138_new_n16087_), .B(u2__abc_52138_new_n16085_), .Y(u2__abc_52138_new_n16088_));
NAND2X1 NAND2X1_1853 ( .A(u2__abc_52138_new_n16095_), .B(u2__abc_52138_new_n16094_), .Y(u2__abc_52138_new_n16096_));
NAND2X1 NAND2X1_1854 ( .A(u2__abc_52138_new_n16102_), .B(u2__abc_52138_new_n16101_), .Y(u2__abc_52138_new_n16103_));
NAND2X1 NAND2X1_1855 ( .A(u2__abc_52138_new_n16111_), .B(u2__abc_52138_new_n16109_), .Y(u2__abc_52138_new_n16112_));
NAND2X1 NAND2X1_1856 ( .A(u2__abc_52138_new_n16119_), .B(u2__abc_52138_new_n16118_), .Y(u2__abc_52138_new_n16120_));
NAND2X1 NAND2X1_1857 ( .A(u2__abc_52138_new_n16127_), .B(u2__abc_52138_new_n16126_), .Y(u2__abc_52138_new_n16128_));
NAND2X1 NAND2X1_1858 ( .A(u2__abc_52138_new_n16134_), .B(u2__abc_52138_new_n16133_), .Y(u2__abc_52138_new_n16135_));
NAND2X1 NAND2X1_1859 ( .A(u2__abc_52138_new_n16142_), .B(u2__abc_52138_new_n16141_), .Y(u2__abc_52138_new_n16143_));
NAND2X1 NAND2X1_186 ( .A(\a[73] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1354_));
NAND2X1 NAND2X1_1860 ( .A(u2__abc_52138_new_n16150_), .B(u2__abc_52138_new_n16149_), .Y(u2__abc_52138_new_n16151_));
NAND2X1 NAND2X1_1861 ( .A(u2__abc_52138_new_n16158_), .B(u2__abc_52138_new_n16157_), .Y(u2__abc_52138_new_n16159_));
NAND2X1 NAND2X1_1862 ( .A(u2__abc_52138_new_n16165_), .B(u2__abc_52138_new_n16164_), .Y(u2__abc_52138_new_n16166_));
NAND2X1 NAND2X1_1863 ( .A(u2__abc_52138_new_n16173_), .B(u2__abc_52138_new_n16172_), .Y(u2__abc_52138_new_n16174_));
NAND2X1 NAND2X1_1864 ( .A(u2__abc_52138_new_n16181_), .B(u2__abc_52138_new_n16180_), .Y(u2__abc_52138_new_n16182_));
NAND2X1 NAND2X1_1865 ( .A(u2__abc_52138_new_n16189_), .B(u2__abc_52138_new_n16188_), .Y(u2__abc_52138_new_n16190_));
NAND2X1 NAND2X1_1866 ( .A(u2__abc_52138_new_n16196_), .B(u2__abc_52138_new_n16195_), .Y(u2__abc_52138_new_n16197_));
NAND2X1 NAND2X1_1867 ( .A(u2__abc_52138_new_n16204_), .B(u2__abc_52138_new_n16203_), .Y(u2__abc_52138_new_n16205_));
NAND2X1 NAND2X1_1868 ( .A(u2__abc_52138_new_n16212_), .B(u2__abc_52138_new_n16211_), .Y(u2__abc_52138_new_n16213_));
NAND2X1 NAND2X1_1869 ( .A(u2__abc_52138_new_n16220_), .B(u2__abc_52138_new_n16219_), .Y(u2__abc_52138_new_n16221_));
NAND2X1 NAND2X1_187 ( .A(\a[112] ), .B(\a[75] ), .Y(_abc_65734_new_n1356_));
NAND2X1 NAND2X1_1870 ( .A(u2__abc_52138_new_n16227_), .B(u2__abc_52138_new_n16226_), .Y(u2__abc_52138_new_n16228_));
NAND2X1 NAND2X1_1871 ( .A(u2__abc_52138_new_n16235_), .B(u2__abc_52138_new_n16234_), .Y(u2__abc_52138_new_n16236_));
NAND2X1 NAND2X1_1872 ( .A(u2__abc_52138_new_n16243_), .B(u2__abc_52138_new_n16242_), .Y(u2__abc_52138_new_n16244_));
NAND2X1 NAND2X1_1873 ( .A(u2__abc_52138_new_n16251_), .B(u2__abc_52138_new_n16250_), .Y(u2__abc_52138_new_n16252_));
NAND2X1 NAND2X1_1874 ( .A(u2__abc_52138_new_n16258_), .B(u2__abc_52138_new_n16257_), .Y(u2__abc_52138_new_n16259_));
NAND2X1 NAND2X1_1875 ( .A(u2__abc_52138_new_n16266_), .B(u2__abc_52138_new_n16265_), .Y(u2__abc_52138_new_n16267_));
NAND2X1 NAND2X1_1876 ( .A(u2__abc_52138_new_n16274_), .B(u2__abc_52138_new_n16273_), .Y(u2__abc_52138_new_n16275_));
NAND2X1 NAND2X1_1877 ( .A(u2__abc_52138_new_n16282_), .B(u2__abc_52138_new_n16281_), .Y(u2__abc_52138_new_n16283_));
NAND2X1 NAND2X1_1878 ( .A(u2__abc_52138_new_n16289_), .B(u2__abc_52138_new_n16288_), .Y(u2__abc_52138_new_n16290_));
NAND2X1 NAND2X1_1879 ( .A(u2__abc_52138_new_n16297_), .B(u2__abc_52138_new_n16296_), .Y(u2__abc_52138_new_n16298_));
NAND2X1 NAND2X1_188 ( .A(\a[75] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1359_));
NAND2X1 NAND2X1_1880 ( .A(u2__abc_52138_new_n16305_), .B(u2__abc_52138_new_n16304_), .Y(u2__abc_52138_new_n16306_));
NAND2X1 NAND2X1_1881 ( .A(u2__abc_52138_new_n16313_), .B(u2__abc_52138_new_n16312_), .Y(u2__abc_52138_new_n16314_));
NAND2X1 NAND2X1_1882 ( .A(u2__abc_52138_new_n16320_), .B(u2__abc_52138_new_n16319_), .Y(u2__abc_52138_new_n16321_));
NAND2X1 NAND2X1_1883 ( .A(u2__abc_52138_new_n16328_), .B(u2__abc_52138_new_n16327_), .Y(u2__abc_52138_new_n16329_));
NAND2X1 NAND2X1_1884 ( .A(u2__abc_52138_new_n16336_), .B(u2__abc_52138_new_n16335_), .Y(u2__abc_52138_new_n16337_));
NAND2X1 NAND2X1_1885 ( .A(u2__abc_52138_new_n16344_), .B(u2__abc_52138_new_n16343_), .Y(u2__abc_52138_new_n16345_));
NAND2X1 NAND2X1_1886 ( .A(u2__abc_52138_new_n16351_), .B(u2__abc_52138_new_n16350_), .Y(u2__abc_52138_new_n16352_));
NAND2X1 NAND2X1_1887 ( .A(u2__abc_52138_new_n16359_), .B(u2__abc_52138_new_n16358_), .Y(u2__abc_52138_new_n16360_));
NAND2X1 NAND2X1_1888 ( .A(u2__abc_52138_new_n16367_), .B(u2__abc_52138_new_n16366_), .Y(u2__abc_52138_new_n16368_));
NAND2X1 NAND2X1_1889 ( .A(u2__abc_52138_new_n16375_), .B(u2__abc_52138_new_n16374_), .Y(u2__abc_52138_new_n16376_));
NAND2X1 NAND2X1_189 ( .A(\a[112] ), .B(\a[77] ), .Y(_abc_65734_new_n1361_));
NAND2X1 NAND2X1_1890 ( .A(u2__abc_52138_new_n16382_), .B(u2__abc_52138_new_n16381_), .Y(u2__abc_52138_new_n16383_));
NAND2X1 NAND2X1_1891 ( .A(u2__abc_52138_new_n16390_), .B(u2__abc_52138_new_n16389_), .Y(u2__abc_52138_new_n16391_));
NAND2X1 NAND2X1_1892 ( .A(u2__abc_52138_new_n16398_), .B(u2__abc_52138_new_n16397_), .Y(u2__abc_52138_new_n16399_));
NAND2X1 NAND2X1_1893 ( .A(u2__abc_52138_new_n16406_), .B(u2__abc_52138_new_n16405_), .Y(u2__abc_52138_new_n16407_));
NAND2X1 NAND2X1_1894 ( .A(u2__abc_52138_new_n16413_), .B(u2__abc_52138_new_n16412_), .Y(u2__abc_52138_new_n16414_));
NAND2X1 NAND2X1_1895 ( .A(u2__abc_52138_new_n16421_), .B(u2__abc_52138_new_n16420_), .Y(u2__abc_52138_new_n16422_));
NAND2X1 NAND2X1_1896 ( .A(u2__abc_52138_new_n16429_), .B(u2__abc_52138_new_n16428_), .Y(u2__abc_52138_new_n16430_));
NAND2X1 NAND2X1_1897 ( .A(u2__abc_52138_new_n16437_), .B(u2__abc_52138_new_n16436_), .Y(u2__abc_52138_new_n16438_));
NAND2X1 NAND2X1_1898 ( .A(u2__abc_52138_new_n16444_), .B(u2__abc_52138_new_n16443_), .Y(u2__abc_52138_new_n16445_));
NAND2X1 NAND2X1_1899 ( .A(u2__abc_52138_new_n16452_), .B(u2__abc_52138_new_n16451_), .Y(u2__abc_52138_new_n16453_));
NAND2X1 NAND2X1_19 ( .A(aNan), .B(\a[18] ), .Y(_abc_65734_new_n885_));
NAND2X1 NAND2X1_190 ( .A(\a[77] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1364_));
NAND2X1 NAND2X1_1900 ( .A(u2__abc_52138_new_n16460_), .B(u2__abc_52138_new_n16459_), .Y(u2__abc_52138_new_n16461_));
NAND2X1 NAND2X1_1901 ( .A(u2__abc_52138_new_n16468_), .B(u2__abc_52138_new_n16467_), .Y(u2__abc_52138_new_n16469_));
NAND2X1 NAND2X1_1902 ( .A(u2__abc_52138_new_n16475_), .B(u2__abc_52138_new_n16474_), .Y(u2__abc_52138_new_n16476_));
NAND2X1 NAND2X1_1903 ( .A(u2__abc_52138_new_n16483_), .B(u2__abc_52138_new_n16482_), .Y(u2__abc_52138_new_n16484_));
NAND2X1 NAND2X1_1904 ( .A(u2__abc_52138_new_n16491_), .B(u2__abc_52138_new_n16490_), .Y(u2__abc_52138_new_n16492_));
NAND2X1 NAND2X1_1905 ( .A(u2__abc_52138_new_n16499_), .B(u2__abc_52138_new_n16498_), .Y(u2__abc_52138_new_n16500_));
NAND2X1 NAND2X1_1906 ( .A(u2__abc_52138_new_n16506_), .B(u2__abc_52138_new_n16505_), .Y(u2__abc_52138_new_n16507_));
NAND2X1 NAND2X1_1907 ( .A(u2__abc_52138_new_n16514_), .B(u2__abc_52138_new_n16513_), .Y(u2__abc_52138_new_n16515_));
NAND2X1 NAND2X1_1908 ( .A(u2__abc_52138_new_n16522_), .B(u2__abc_52138_new_n16521_), .Y(u2__abc_52138_new_n16523_));
NAND2X1 NAND2X1_1909 ( .A(u2__abc_52138_new_n16530_), .B(u2__abc_52138_new_n16529_), .Y(u2__abc_52138_new_n16531_));
NAND2X1 NAND2X1_191 ( .A(\a[112] ), .B(\a[79] ), .Y(_abc_65734_new_n1366_));
NAND2X1 NAND2X1_1910 ( .A(u2__abc_52138_new_n16537_), .B(u2__abc_52138_new_n16536_), .Y(u2__abc_52138_new_n16538_));
NAND2X1 NAND2X1_192 ( .A(\a[79] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1369_));
NAND2X1 NAND2X1_193 ( .A(\a[112] ), .B(\a[81] ), .Y(_abc_65734_new_n1371_));
NAND2X1 NAND2X1_194 ( .A(\a[81] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1374_));
NAND2X1 NAND2X1_195 ( .A(\a[112] ), .B(\a[83] ), .Y(_abc_65734_new_n1376_));
NAND2X1 NAND2X1_196 ( .A(\a[83] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1379_));
NAND2X1 NAND2X1_197 ( .A(\a[112] ), .B(\a[85] ), .Y(_abc_65734_new_n1381_));
NAND2X1 NAND2X1_198 ( .A(\a[85] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1384_));
NAND2X1 NAND2X1_199 ( .A(\a[112] ), .B(\a[87] ), .Y(_abc_65734_new_n1386_));
NAND2X1 NAND2X1_2 ( .A(aNan), .B(\a[1] ), .Y(_abc_65734_new_n834_));
NAND2X1 NAND2X1_20 ( .A(aNan), .B(\a[19] ), .Y(_abc_65734_new_n888_));
NAND2X1 NAND2X1_200 ( .A(\a[87] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1389_));
NAND2X1 NAND2X1_201 ( .A(\a[112] ), .B(\a[89] ), .Y(_abc_65734_new_n1391_));
NAND2X1 NAND2X1_202 ( .A(\a[89] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1394_));
NAND2X1 NAND2X1_203 ( .A(\a[112] ), .B(\a[91] ), .Y(_abc_65734_new_n1396_));
NAND2X1 NAND2X1_204 ( .A(\a[91] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1399_));
NAND2X1 NAND2X1_205 ( .A(\a[112] ), .B(\a[93] ), .Y(_abc_65734_new_n1401_));
NAND2X1 NAND2X1_206 ( .A(\a[93] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1404_));
NAND2X1 NAND2X1_207 ( .A(\a[112] ), .B(\a[95] ), .Y(_abc_65734_new_n1406_));
NAND2X1 NAND2X1_208 ( .A(\a[95] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1409_));
NAND2X1 NAND2X1_209 ( .A(\a[112] ), .B(\a[97] ), .Y(_abc_65734_new_n1411_));
NAND2X1 NAND2X1_21 ( .A(aNan), .B(\a[20] ), .Y(_abc_65734_new_n891_));
NAND2X1 NAND2X1_210 ( .A(\a[97] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1414_));
NAND2X1 NAND2X1_211 ( .A(\a[112] ), .B(\a[99] ), .Y(_abc_65734_new_n1416_));
NAND2X1 NAND2X1_212 ( .A(\a[99] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1419_));
NAND2X1 NAND2X1_213 ( .A(\a[112] ), .B(\a[101] ), .Y(_abc_65734_new_n1421_));
NAND2X1 NAND2X1_214 ( .A(\a[101] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1424_));
NAND2X1 NAND2X1_215 ( .A(\a[112] ), .B(\a[103] ), .Y(_abc_65734_new_n1426_));
NAND2X1 NAND2X1_216 ( .A(\a[103] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1429_));
NAND2X1 NAND2X1_217 ( .A(\a[112] ), .B(\a[105] ), .Y(_abc_65734_new_n1431_));
NAND2X1 NAND2X1_218 ( .A(\a[105] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1434_));
NAND2X1 NAND2X1_219 ( .A(\a[112] ), .B(\a[107] ), .Y(_abc_65734_new_n1436_));
NAND2X1 NAND2X1_22 ( .A(aNan), .B(\a[21] ), .Y(_abc_65734_new_n894_));
NAND2X1 NAND2X1_220 ( .A(\a[107] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1439_));
NAND2X1 NAND2X1_221 ( .A(\a[112] ), .B(\a[109] ), .Y(_abc_65734_new_n1441_));
NAND2X1 NAND2X1_222 ( .A(\a[109] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1444_));
NAND2X1 NAND2X1_223 ( .A(\a[112] ), .B(\a[111] ), .Y(_abc_65734_new_n1446_));
NAND2X1 NAND2X1_224 ( .A(\a[111] ), .B(_abc_65734_new_n1168_), .Y(_abc_65734_new_n1449_));
NAND2X1 NAND2X1_225 ( .A(\a[112] ), .B(\a[113] ), .Y(_abc_65734_new_n1461_));
NAND2X1 NAND2X1_226 ( .A(\a[114] ), .B(\a[115] ), .Y(_abc_65734_new_n1462_));
NAND2X1 NAND2X1_227 ( .A(_abc_65734_new_n1452_), .B(_abc_65734_new_n1470_), .Y(_abc_65734_new_n1471_));
NAND2X1 NAND2X1_228 ( .A(\a[117] ), .B(_abc_65734_new_n1486_), .Y(_abc_65734_new_n1487_));
NAND2X1 NAND2X1_229 ( .A(_abc_65734_new_n1485_), .B(_abc_65734_new_n1487_), .Y(_abc_65734_new_n1488_));
NAND2X1 NAND2X1_23 ( .A(aNan), .B(\a[22] ), .Y(_abc_65734_new_n897_));
NAND2X1 NAND2X1_230 ( .A(_abc_65734_new_n1492_), .B(_abc_65734_new_n1494_), .Y(_abc_65734_new_n1496_));
NAND2X1 NAND2X1_231 ( .A(_abc_65734_new_n1502_), .B(_abc_65734_new_n1501_), .Y(_abc_65734_new_n1503_));
NAND2X1 NAND2X1_232 ( .A(_abc_65734_new_n1513_), .B(_abc_65734_new_n1512_), .Y(_abc_65734_new_n1514_));
NAND2X1 NAND2X1_233 ( .A(_abc_65734_new_n1517_), .B(_abc_65734_new_n1516_), .Y(_abc_65734_new_n1518_));
NAND2X1 NAND2X1_234 ( .A(_abc_65734_new_n1525_), .B(_abc_65734_new_n1526_), .Y(_abc_65734_new_n1527_));
NAND2X1 NAND2X1_235 ( .A(\a[120] ), .B(\a[121] ), .Y(_abc_65734_new_n1534_));
NAND2X1 NAND2X1_236 ( .A(_abc_65734_new_n1536_), .B(_abc_65734_new_n1537_), .Y(_abc_65734_new_n1538_));
NAND2X1 NAND2X1_237 ( .A(_abc_65734_new_n1549_), .B(_abc_65734_new_n1547_), .Y(_abc_65734_new_n1550_));
NAND2X1 NAND2X1_238 ( .A(aNan), .B(\a[122] ), .Y(_abc_65734_new_n1552_));
NAND2X1 NAND2X1_239 ( .A(aNan), .B(\a[123] ), .Y(_abc_65734_new_n1554_));
NAND2X1 NAND2X1_24 ( .A(aNan), .B(\a[23] ), .Y(_abc_65734_new_n900_));
NAND2X1 NAND2X1_240 ( .A(_abc_65734_new_n1564_), .B(_abc_65734_new_n1566_), .Y(_abc_65734_new_n1567_));
NAND2X1 NAND2X1_241 ( .A(aNan), .B(\a[124] ), .Y(_abc_65734_new_n1569_));
NAND2X1 NAND2X1_242 ( .A(aNan), .B(\a[125] ), .Y(_abc_65734_new_n1578_));
NAND2X1 NAND2X1_243 ( .A(_abc_65734_new_n1578_), .B(_abc_65734_new_n1577_), .Y(\o[239] ));
NAND2X1 NAND2X1_244 ( .A(\a[126] ), .B(_abc_65734_new_n1583_), .Y(_abc_65734_new_n1584_));
NAND2X1 NAND2X1_245 ( .A(u1__abc_51895_new_n137_), .B(u1__abc_51895_new_n138_), .Y(u1__abc_51895_new_n139_));
NAND2X1 NAND2X1_246 ( .A(u1__abc_51895_new_n140_), .B(u1__abc_51895_new_n141_), .Y(u1__abc_51895_new_n142_));
NAND2X1 NAND2X1_247 ( .A(u1__abc_51895_new_n144_), .B(u1__abc_51895_new_n145_), .Y(u1__abc_51895_new_n146_));
NAND2X1 NAND2X1_248 ( .A(u1__abc_51895_new_n147_), .B(u1__abc_51895_new_n148_), .Y(u1__abc_51895_new_n149_));
NAND2X1 NAND2X1_249 ( .A(u1__abc_51895_new_n150_), .B(u1__abc_51895_new_n143_), .Y(fracta_112_));
NAND2X1 NAND2X1_25 ( .A(aNan), .B(\a[24] ), .Y(_abc_65734_new_n903_));
NAND2X1 NAND2X1_250 ( .A(\a[121] ), .B(\a[122] ), .Y(u1__abc_51895_new_n153_));
NAND2X1 NAND2X1_251 ( .A(\a[119] ), .B(\a[120] ), .Y(u1__abc_51895_new_n154_));
NAND2X1 NAND2X1_252 ( .A(\a[125] ), .B(\a[126] ), .Y(u1__abc_51895_new_n156_));
NAND2X1 NAND2X1_253 ( .A(\a[123] ), .B(\a[124] ), .Y(u1__abc_51895_new_n157_));
NAND2X1 NAND2X1_254 ( .A(u1__abc_51895_new_n155_), .B(u1__abc_51895_new_n158_), .Y(u1__abc_51895_new_n159_));
NAND2X1 NAND2X1_255 ( .A(\a[117] ), .B(\a[118] ), .Y(u1__abc_51895_new_n161_));
NAND2X1 NAND2X1_256 ( .A(\a[115] ), .B(\a[116] ), .Y(u1__abc_51895_new_n162_));
NAND2X1 NAND2X1_257 ( .A(u1__abc_51895_new_n166_), .B(u1__abc_51895_new_n167_), .Y(u1__abc_51895_new_n168_));
NAND2X1 NAND2X1_258 ( .A(u1__abc_51895_new_n169_), .B(u1__abc_51895_new_n170_), .Y(u1__abc_51895_new_n171_));
NAND2X1 NAND2X1_259 ( .A(u1__abc_51895_new_n173_), .B(u1__abc_51895_new_n174_), .Y(u1__abc_51895_new_n175_));
NAND2X1 NAND2X1_26 ( .A(aNan), .B(\a[25] ), .Y(_abc_65734_new_n906_));
NAND2X1 NAND2X1_260 ( .A(u1__abc_51895_new_n176_), .B(u1__abc_51895_new_n177_), .Y(u1__abc_51895_new_n178_));
NAND2X1 NAND2X1_261 ( .A(u1__abc_51895_new_n172_), .B(u1__abc_51895_new_n179_), .Y(u1__abc_51895_new_n180_));
NAND2X1 NAND2X1_262 ( .A(u1__abc_51895_new_n282_), .B(u1__abc_51895_new_n283_), .Y(u1__abc_51895_new_n284_));
NAND2X1 NAND2X1_263 ( .A(u1__abc_51895_new_n285_), .B(u1__abc_51895_new_n286_), .Y(u1__abc_51895_new_n287_));
NAND2X1 NAND2X1_264 ( .A(u1__abc_51895_new_n289_), .B(u1__abc_51895_new_n290_), .Y(u1__abc_51895_new_n291_));
NAND2X1 NAND2X1_265 ( .A(u1__abc_51895_new_n292_), .B(u1__abc_51895_new_n293_), .Y(u1__abc_51895_new_n294_));
NAND2X1 NAND2X1_266 ( .A(u1__abc_51895_new_n288_), .B(u1__abc_51895_new_n295_), .Y(u1__abc_51895_new_n296_));
NAND2X1 NAND2X1_267 ( .A(u1__abc_51895_new_n298_), .B(u1__abc_51895_new_n299_), .Y(u1__abc_51895_new_n300_));
NAND2X1 NAND2X1_268 ( .A(u1__abc_51895_new_n301_), .B(u1__abc_51895_new_n302_), .Y(u1__abc_51895_new_n303_));
NAND2X1 NAND2X1_269 ( .A(u1__abc_51895_new_n305_), .B(u1__abc_51895_new_n306_), .Y(u1__abc_51895_new_n307_));
NAND2X1 NAND2X1_27 ( .A(aNan), .B(\a[26] ), .Y(_abc_65734_new_n909_));
NAND2X1 NAND2X1_270 ( .A(u1__abc_51895_new_n308_), .B(u1__abc_51895_new_n309_), .Y(u1__abc_51895_new_n310_));
NAND2X1 NAND2X1_271 ( .A(u1__abc_51895_new_n304_), .B(u1__abc_51895_new_n311_), .Y(u1__abc_51895_new_n312_));
NAND2X1 NAND2X1_272 ( .A(u1__abc_51895_new_n313_), .B(u1__abc_51895_new_n314_), .Y(u1__abc_51895_new_n315_));
NAND2X1 NAND2X1_273 ( .A(u1__abc_51895_new_n316_), .B(u1__abc_51895_new_n317_), .Y(u1__abc_51895_new_n318_));
NAND2X1 NAND2X1_274 ( .A(u1__abc_51895_new_n320_), .B(u1__abc_51895_new_n321_), .Y(u1__abc_51895_new_n322_));
NAND2X1 NAND2X1_275 ( .A(u1__abc_51895_new_n323_), .B(u1__abc_51895_new_n324_), .Y(u1__abc_51895_new_n325_));
NAND2X1 NAND2X1_276 ( .A(u1__abc_51895_new_n319_), .B(u1__abc_51895_new_n326_), .Y(u1__abc_51895_new_n327_));
NAND2X1 NAND2X1_277 ( .A(u1__abc_51895_new_n330_), .B(u1__abc_51895_new_n331_), .Y(u1__abc_51895_new_n332_));
NAND2X1 NAND2X1_278 ( .A(u1__abc_51895_new_n333_), .B(u1__abc_51895_new_n334_), .Y(u1__abc_51895_new_n335_));
NAND2X1 NAND2X1_279 ( .A(u1__abc_51895_new_n337_), .B(u1__abc_51895_new_n338_), .Y(u1__abc_51895_new_n339_));
NAND2X1 NAND2X1_28 ( .A(aNan), .B(\a[27] ), .Y(_abc_65734_new_n912_));
NAND2X1 NAND2X1_280 ( .A(u1__abc_51895_new_n340_), .B(u1__abc_51895_new_n341_), .Y(u1__abc_51895_new_n342_));
NAND2X1 NAND2X1_281 ( .A(u1__abc_51895_new_n336_), .B(u1__abc_51895_new_n343_), .Y(u1__abc_51895_new_n344_));
NAND2X1 NAND2X1_282 ( .A(u1__abc_51895_new_n345_), .B(u1__abc_51895_new_n346_), .Y(u1__abc_51895_new_n347_));
NAND2X1 NAND2X1_283 ( .A(u1__abc_51895_new_n348_), .B(u1__abc_51895_new_n349_), .Y(u1__abc_51895_new_n350_));
NAND2X1 NAND2X1_284 ( .A(u1__abc_51895_new_n352_), .B(u1__abc_51895_new_n353_), .Y(u1__abc_51895_new_n354_));
NAND2X1 NAND2X1_285 ( .A(u1__abc_51895_new_n355_), .B(u1__abc_51895_new_n356_), .Y(u1__abc_51895_new_n357_));
NAND2X1 NAND2X1_286 ( .A(u1__abc_51895_new_n351_), .B(u1__abc_51895_new_n358_), .Y(u1__abc_51895_new_n359_));
NAND2X1 NAND2X1_287 ( .A(u1__abc_51895_new_n360_), .B(u1__abc_51895_new_n361_), .Y(u1__abc_51895_new_n362_));
NAND2X1 NAND2X1_288 ( .A(u1__abc_51895_new_n363_), .B(u1__abc_51895_new_n364_), .Y(u1__abc_51895_new_n365_));
NAND2X1 NAND2X1_289 ( .A(u1__abc_51895_new_n367_), .B(u1__abc_51895_new_n368_), .Y(u1__abc_51895_new_n369_));
NAND2X1 NAND2X1_29 ( .A(aNan), .B(\a[28] ), .Y(_abc_65734_new_n915_));
NAND2X1 NAND2X1_290 ( .A(u1__abc_51895_new_n370_), .B(u1__abc_51895_new_n371_), .Y(u1__abc_51895_new_n372_));
NAND2X1 NAND2X1_291 ( .A(u1__abc_51895_new_n366_), .B(u1__abc_51895_new_n373_), .Y(u1__abc_51895_new_n374_));
NAND2X1 NAND2X1_292 ( .A(ce), .B(u2__abc_52138_new_n2964_), .Y(u2__abc_52138_new_n2965_));
NAND2X1 NAND2X1_293 ( .A(u2_cnt_7_), .B(u2__abc_52138_new_n2967_), .Y(u2__abc_52138_new_n2968_));
NAND2X1 NAND2X1_294 ( .A(u2__abc_52138_new_n2971_), .B(u2__abc_52138_new_n2977_), .Y(u2__abc_52138_new_n2978_));
NAND2X1 NAND2X1_295 ( .A(done), .B(u2__abc_52138_new_n2982_), .Y(u2__abc_52138_new_n2987_));
NAND2X1 NAND2X1_296 ( .A(u2__abc_52138_new_n2988_), .B(u2__abc_52138_new_n2989_), .Y(u2__abc_52138_new_n2990_));
NAND2X1 NAND2X1_297 ( .A(u2_state_2_), .B(u2__abc_52138_new_n2991_), .Y(u2__abc_52138_new_n2992_));
NAND2X1 NAND2X1_298 ( .A(u2__abc_52138_new_n3013_), .B(u2__abc_52138_new_n3002_), .Y(u2__abc_52138_new_n3014_));
NAND2X1 NAND2X1_299 ( .A(sqrto_13_), .B(u2__abc_52138_new_n3017_), .Y(u2__abc_52138_new_n3018_));
NAND2X1 NAND2X1_3 ( .A(aNan), .B(\a[2] ), .Y(_abc_65734_new_n837_));
NAND2X1 NAND2X1_30 ( .A(aNan), .B(\a[29] ), .Y(_abc_65734_new_n918_));
NAND2X1 NAND2X1_300 ( .A(u2_remHi_13_), .B(u2__abc_52138_new_n3019_), .Y(u2__abc_52138_new_n3020_));
NAND2X1 NAND2X1_301 ( .A(u2_remHi_11_), .B(u2__abc_52138_new_n3022_), .Y(u2__abc_52138_new_n3023_));
NAND2X1 NAND2X1_302 ( .A(sqrto_11_), .B(u2__abc_52138_new_n3024_), .Y(u2__abc_52138_new_n3025_));
NAND2X1 NAND2X1_303 ( .A(u2_remHi_10_), .B(u2__abc_52138_new_n3027_), .Y(u2__abc_52138_new_n3028_));
NAND2X1 NAND2X1_304 ( .A(sqrto_10_), .B(u2__abc_52138_new_n3029_), .Y(u2__abc_52138_new_n3030_));
NAND2X1 NAND2X1_305 ( .A(u2__abc_52138_new_n3026_), .B(u2__abc_52138_new_n3031_), .Y(u2__abc_52138_new_n3032_));
NAND2X1 NAND2X1_306 ( .A(u2_remHi_9_), .B(u2__abc_52138_new_n3035_), .Y(u2__abc_52138_new_n3036_));
NAND2X1 NAND2X1_307 ( .A(sqrto_9_), .B(u2__abc_52138_new_n3037_), .Y(u2__abc_52138_new_n3038_));
NAND2X1 NAND2X1_308 ( .A(u2_remHi_7_), .B(u2__abc_52138_new_n3040_), .Y(u2__abc_52138_new_n3041_));
NAND2X1 NAND2X1_309 ( .A(sqrto_7_), .B(u2__abc_52138_new_n3042_), .Y(u2__abc_52138_new_n3043_));
NAND2X1 NAND2X1_31 ( .A(aNan), .B(\a[30] ), .Y(_abc_65734_new_n921_));
NAND2X1 NAND2X1_310 ( .A(u2_remHi_6_), .B(u2__abc_52138_new_n3045_), .Y(u2__abc_52138_new_n3046_));
NAND2X1 NAND2X1_311 ( .A(sqrto_6_), .B(u2__abc_52138_new_n3047_), .Y(u2__abc_52138_new_n3048_));
NAND2X1 NAND2X1_312 ( .A(u2__abc_52138_new_n3044_), .B(u2__abc_52138_new_n3049_), .Y(u2__abc_52138_new_n3050_));
NAND2X1 NAND2X1_313 ( .A(u2__abc_52138_new_n3033_), .B(u2__abc_52138_new_n3051_), .Y(u2__abc_52138_new_n3052_));
NAND2X1 NAND2X1_314 ( .A(sqrto_5_), .B(u2__abc_52138_new_n3054_), .Y(u2__abc_52138_new_n3055_));
NAND2X1 NAND2X1_315 ( .A(u2_remHi_5_), .B(u2__abc_52138_new_n3056_), .Y(u2__abc_52138_new_n3057_));
NAND2X1 NAND2X1_316 ( .A(u2_remHi_2_), .B(u2__abc_52138_new_n3060_), .Y(u2__abc_52138_new_n3061_));
NAND2X1 NAND2X1_317 ( .A(sqrto_2_), .B(u2__abc_52138_new_n3062_), .Y(u2__abc_52138_new_n3063_));
NAND2X1 NAND2X1_318 ( .A(u2__abc_52138_new_n3066_), .B(u2__abc_52138_new_n3067_), .Y(u2__abc_52138_new_n3068_));
NAND2X1 NAND2X1_319 ( .A(u2_remHiShift_1_), .B(u2__abc_52138_new_n3069_), .Y(u2__abc_52138_new_n3070_));
NAND2X1 NAND2X1_32 ( .A(aNan), .B(\a[31] ), .Y(_abc_65734_new_n924_));
NAND2X1 NAND2X1_320 ( .A(u2_remHi_1_), .B(u2__abc_52138_new_n3074_), .Y(u2__abc_52138_new_n3076_));
NAND2X1 NAND2X1_321 ( .A(u2_remHi_3_), .B(u2__abc_52138_new_n3079_), .Y(u2__abc_52138_new_n3080_));
NAND2X1 NAND2X1_322 ( .A(sqrto_3_), .B(u2__abc_52138_new_n3081_), .Y(u2__abc_52138_new_n3082_));
NAND2X1 NAND2X1_323 ( .A(sqrto_4_), .B(u2__abc_52138_new_n3086_), .Y(u2__abc_52138_new_n3087_));
NAND2X1 NAND2X1_324 ( .A(sqrto_12_), .B(u2__abc_52138_new_n3101_), .Y(u2__abc_52138_new_n3102_));
NAND2X1 NAND2X1_325 ( .A(u2_remHi_24_), .B(u2__abc_52138_new_n3112_), .Y(u2__abc_52138_new_n3113_));
NAND2X1 NAND2X1_326 ( .A(sqrto_24_), .B(u2__abc_52138_new_n3114_), .Y(u2__abc_52138_new_n3115_));
NAND2X1 NAND2X1_327 ( .A(u2__abc_52138_new_n3113_), .B(u2__abc_52138_new_n3115_), .Y(u2__abc_52138_new_n3116_));
NAND2X1 NAND2X1_328 ( .A(u2_remHi_25_), .B(u2__abc_52138_new_n3117_), .Y(u2__abc_52138_new_n3118_));
NAND2X1 NAND2X1_329 ( .A(sqrto_25_), .B(u2__abc_52138_new_n3119_), .Y(u2__abc_52138_new_n3120_));
NAND2X1 NAND2X1_33 ( .A(aNan), .B(\a[32] ), .Y(_abc_65734_new_n927_));
NAND2X1 NAND2X1_330 ( .A(u2__abc_52138_new_n3118_), .B(u2__abc_52138_new_n3120_), .Y(u2__abc_52138_new_n3121_));
NAND2X1 NAND2X1_331 ( .A(u2_remHi_23_), .B(u2__abc_52138_new_n3123_), .Y(u2__abc_52138_new_n3124_));
NAND2X1 NAND2X1_332 ( .A(sqrto_23_), .B(u2__abc_52138_new_n3125_), .Y(u2__abc_52138_new_n3126_));
NAND2X1 NAND2X1_333 ( .A(u2__abc_52138_new_n3124_), .B(u2__abc_52138_new_n3126_), .Y(u2__abc_52138_new_n3127_));
NAND2X1 NAND2X1_334 ( .A(u2_remHi_22_), .B(u2__abc_52138_new_n3128_), .Y(u2__abc_52138_new_n3129_));
NAND2X1 NAND2X1_335 ( .A(sqrto_22_), .B(u2__abc_52138_new_n3130_), .Y(u2__abc_52138_new_n3131_));
NAND2X1 NAND2X1_336 ( .A(u2__abc_52138_new_n3129_), .B(u2__abc_52138_new_n3131_), .Y(u2__abc_52138_new_n3132_));
NAND2X1 NAND2X1_337 ( .A(u2__abc_52138_new_n3122_), .B(u2__abc_52138_new_n3133_), .Y(u2__abc_52138_new_n3134_));
NAND2X1 NAND2X1_338 ( .A(u2_remHi_28_), .B(u2__abc_52138_new_n3135_), .Y(u2__abc_52138_new_n3136_));
NAND2X1 NAND2X1_339 ( .A(sqrto_28_), .B(u2__abc_52138_new_n3137_), .Y(u2__abc_52138_new_n3138_));
NAND2X1 NAND2X1_34 ( .A(aNan), .B(\a[33] ), .Y(_abc_65734_new_n930_));
NAND2X1 NAND2X1_340 ( .A(u2__abc_52138_new_n3136_), .B(u2__abc_52138_new_n3138_), .Y(u2__abc_52138_new_n3139_));
NAND2X1 NAND2X1_341 ( .A(sqrto_29_), .B(u2__abc_52138_new_n3140_), .Y(u2__abc_52138_new_n3141_));
NAND2X1 NAND2X1_342 ( .A(u2_remHi_29_), .B(u2__abc_52138_new_n3142_), .Y(u2__abc_52138_new_n3143_));
NAND2X1 NAND2X1_343 ( .A(u2__abc_52138_new_n3141_), .B(u2__abc_52138_new_n3143_), .Y(u2__abc_52138_new_n3144_));
NAND2X1 NAND2X1_344 ( .A(u2_remHi_27_), .B(u2__abc_52138_new_n3146_), .Y(u2__abc_52138_new_n3147_));
NAND2X1 NAND2X1_345 ( .A(sqrto_27_), .B(u2__abc_52138_new_n3148_), .Y(u2__abc_52138_new_n3149_));
NAND2X1 NAND2X1_346 ( .A(u2__abc_52138_new_n3147_), .B(u2__abc_52138_new_n3149_), .Y(u2__abc_52138_new_n3150_));
NAND2X1 NAND2X1_347 ( .A(u2_remHi_26_), .B(u2__abc_52138_new_n3151_), .Y(u2__abc_52138_new_n3152_));
NAND2X1 NAND2X1_348 ( .A(sqrto_26_), .B(u2__abc_52138_new_n3153_), .Y(u2__abc_52138_new_n3154_));
NAND2X1 NAND2X1_349 ( .A(u2__abc_52138_new_n3152_), .B(u2__abc_52138_new_n3154_), .Y(u2__abc_52138_new_n3155_));
NAND2X1 NAND2X1_35 ( .A(aNan), .B(\a[34] ), .Y(_abc_65734_new_n933_));
NAND2X1 NAND2X1_350 ( .A(u2__abc_52138_new_n3145_), .B(u2__abc_52138_new_n3156_), .Y(u2__abc_52138_new_n3157_));
NAND2X1 NAND2X1_351 ( .A(u2_remHi_16_), .B(u2__abc_52138_new_n3159_), .Y(u2__abc_52138_new_n3160_));
NAND2X1 NAND2X1_352 ( .A(sqrto_16_), .B(u2__abc_52138_new_n3161_), .Y(u2__abc_52138_new_n3162_));
NAND2X1 NAND2X1_353 ( .A(u2__abc_52138_new_n3160_), .B(u2__abc_52138_new_n3162_), .Y(u2__abc_52138_new_n3163_));
NAND2X1 NAND2X1_354 ( .A(u2_remHi_17_), .B(u2__abc_52138_new_n3164_), .Y(u2__abc_52138_new_n3165_));
NAND2X1 NAND2X1_355 ( .A(sqrto_17_), .B(u2__abc_52138_new_n3166_), .Y(u2__abc_52138_new_n3167_));
NAND2X1 NAND2X1_356 ( .A(u2__abc_52138_new_n3165_), .B(u2__abc_52138_new_n3167_), .Y(u2__abc_52138_new_n3168_));
NAND2X1 NAND2X1_357 ( .A(u2_remHi_14_), .B(u2__abc_52138_new_n3170_), .Y(u2__abc_52138_new_n3171_));
NAND2X1 NAND2X1_358 ( .A(sqrto_14_), .B(u2__abc_52138_new_n3172_), .Y(u2__abc_52138_new_n3173_));
NAND2X1 NAND2X1_359 ( .A(u2__abc_52138_new_n3171_), .B(u2__abc_52138_new_n3173_), .Y(u2__abc_52138_new_n3174_));
NAND2X1 NAND2X1_36 ( .A(aNan), .B(\a[35] ), .Y(_abc_65734_new_n936_));
NAND2X1 NAND2X1_360 ( .A(u2_remHi_15_), .B(u2__abc_52138_new_n3175_), .Y(u2__abc_52138_new_n3176_));
NAND2X1 NAND2X1_361 ( .A(sqrto_15_), .B(u2__abc_52138_new_n3177_), .Y(u2__abc_52138_new_n3178_));
NAND2X1 NAND2X1_362 ( .A(u2__abc_52138_new_n3176_), .B(u2__abc_52138_new_n3178_), .Y(u2__abc_52138_new_n3179_));
NAND2X1 NAND2X1_363 ( .A(u2_remHi_21_), .B(u2__abc_52138_new_n3183_), .Y(u2__abc_52138_new_n3184_));
NAND2X1 NAND2X1_364 ( .A(sqrto_21_), .B(u2__abc_52138_new_n3185_), .Y(u2__abc_52138_new_n3186_));
NAND2X1 NAND2X1_365 ( .A(u2_remHi_18_), .B(u2__abc_52138_new_n3189_), .Y(u2__abc_52138_new_n3190_));
NAND2X1 NAND2X1_366 ( .A(sqrto_18_), .B(u2__abc_52138_new_n3191_), .Y(u2__abc_52138_new_n3192_));
NAND2X1 NAND2X1_367 ( .A(u2__abc_52138_new_n3194_), .B(u2__abc_52138_new_n3181_), .Y(u2__abc_52138_new_n3195_));
NAND2X1 NAND2X1_368 ( .A(u2_remHi_19_), .B(u2__abc_52138_new_n3206_), .Y(u2__abc_52138_new_n3207_));
NAND2X1 NAND2X1_369 ( .A(sqrto_20_), .B(u2__abc_52138_new_n3211_), .Y(u2__abc_52138_new_n3212_));
NAND2X1 NAND2X1_37 ( .A(aNan), .B(\a[36] ), .Y(_abc_65734_new_n939_));
NAND2X1 NAND2X1_370 ( .A(u2__abc_52138_new_n3219_), .B(u2__abc_52138_new_n3220_), .Y(u2__abc_52138_new_n3221_));
NAND2X1 NAND2X1_371 ( .A(u2_remHi_56_), .B(u2__abc_52138_new_n3240_), .Y(u2__abc_52138_new_n3241_));
NAND2X1 NAND2X1_372 ( .A(sqrto_56_), .B(u2__abc_52138_new_n3242_), .Y(u2__abc_52138_new_n3243_));
NAND2X1 NAND2X1_373 ( .A(u2__abc_52138_new_n3241_), .B(u2__abc_52138_new_n3243_), .Y(u2__abc_52138_new_n3244_));
NAND2X1 NAND2X1_374 ( .A(u2_remHi_57_), .B(u2__abc_52138_new_n3245_), .Y(u2__abc_52138_new_n3246_));
NAND2X1 NAND2X1_375 ( .A(sqrto_57_), .B(u2__abc_52138_new_n3247_), .Y(u2__abc_52138_new_n3248_));
NAND2X1 NAND2X1_376 ( .A(u2__abc_52138_new_n3246_), .B(u2__abc_52138_new_n3248_), .Y(u2__abc_52138_new_n3249_));
NAND2X1 NAND2X1_377 ( .A(u2_remHi_54_), .B(u2__abc_52138_new_n3251_), .Y(u2__abc_52138_new_n3252_));
NAND2X1 NAND2X1_378 ( .A(sqrto_54_), .B(u2__abc_52138_new_n3253_), .Y(u2__abc_52138_new_n3254_));
NAND2X1 NAND2X1_379 ( .A(u2__abc_52138_new_n3252_), .B(u2__abc_52138_new_n3254_), .Y(u2__abc_52138_new_n3255_));
NAND2X1 NAND2X1_38 ( .A(aNan), .B(\a[37] ), .Y(_abc_65734_new_n942_));
NAND2X1 NAND2X1_380 ( .A(u2_remHi_55_), .B(u2__abc_52138_new_n3256_), .Y(u2__abc_52138_new_n3257_));
NAND2X1 NAND2X1_381 ( .A(sqrto_55_), .B(u2__abc_52138_new_n3258_), .Y(u2__abc_52138_new_n3259_));
NAND2X1 NAND2X1_382 ( .A(u2__abc_52138_new_n3257_), .B(u2__abc_52138_new_n3259_), .Y(u2__abc_52138_new_n3260_));
NAND2X1 NAND2X1_383 ( .A(u2__abc_52138_new_n3250_), .B(u2__abc_52138_new_n3261_), .Y(u2__abc_52138_new_n3262_));
NAND2X1 NAND2X1_384 ( .A(u2_remHi_60_), .B(u2__abc_52138_new_n3263_), .Y(u2__abc_52138_new_n3264_));
NAND2X1 NAND2X1_385 ( .A(sqrto_60_), .B(u2__abc_52138_new_n3265_), .Y(u2__abc_52138_new_n3266_));
NAND2X1 NAND2X1_386 ( .A(u2__abc_52138_new_n3264_), .B(u2__abc_52138_new_n3266_), .Y(u2__abc_52138_new_n3267_));
NAND2X1 NAND2X1_387 ( .A(sqrto_61_), .B(u2__abc_52138_new_n3268_), .Y(u2__abc_52138_new_n3269_));
NAND2X1 NAND2X1_388 ( .A(u2_remHi_61_), .B(u2__abc_52138_new_n3270_), .Y(u2__abc_52138_new_n3271_));
NAND2X1 NAND2X1_389 ( .A(u2__abc_52138_new_n3269_), .B(u2__abc_52138_new_n3271_), .Y(u2__abc_52138_new_n3272_));
NAND2X1 NAND2X1_39 ( .A(aNan), .B(\a[38] ), .Y(_abc_65734_new_n945_));
NAND2X1 NAND2X1_390 ( .A(u2_remHi_59_), .B(u2__abc_52138_new_n3274_), .Y(u2__abc_52138_new_n3275_));
NAND2X1 NAND2X1_391 ( .A(sqrto_59_), .B(u2__abc_52138_new_n3276_), .Y(u2__abc_52138_new_n3277_));
NAND2X1 NAND2X1_392 ( .A(u2__abc_52138_new_n3275_), .B(u2__abc_52138_new_n3277_), .Y(u2__abc_52138_new_n3278_));
NAND2X1 NAND2X1_393 ( .A(u2_remHi_58_), .B(u2__abc_52138_new_n3279_), .Y(u2__abc_52138_new_n3280_));
NAND2X1 NAND2X1_394 ( .A(sqrto_58_), .B(u2__abc_52138_new_n3281_), .Y(u2__abc_52138_new_n3282_));
NAND2X1 NAND2X1_395 ( .A(u2__abc_52138_new_n3280_), .B(u2__abc_52138_new_n3282_), .Y(u2__abc_52138_new_n3283_));
NAND2X1 NAND2X1_396 ( .A(u2__abc_52138_new_n3273_), .B(u2__abc_52138_new_n3284_), .Y(u2__abc_52138_new_n3285_));
NAND2X1 NAND2X1_397 ( .A(u2__abc_52138_new_n3291_), .B(u2__abc_52138_new_n3296_), .Y(u2__abc_52138_new_n3297_));
NAND2X1 NAND2X1_398 ( .A(u2_remHi_46_), .B(u2__abc_52138_new_n3303_), .Y(u2__abc_52138_new_n3304_));
NAND2X1 NAND2X1_399 ( .A(sqrto_46_), .B(u2__abc_52138_new_n3305_), .Y(u2__abc_52138_new_n3306_));
NAND2X1 NAND2X1_4 ( .A(aNan), .B(\a[3] ), .Y(_abc_65734_new_n840_));
NAND2X1 NAND2X1_40 ( .A(aNan), .B(\a[39] ), .Y(_abc_65734_new_n948_));
NAND2X1 NAND2X1_400 ( .A(u2__abc_52138_new_n3304_), .B(u2__abc_52138_new_n3306_), .Y(u2__abc_52138_new_n3307_));
NAND2X1 NAND2X1_401 ( .A(u2__abc_52138_new_n3302_), .B(u2__abc_52138_new_n3308_), .Y(u2__abc_52138_new_n3309_));
NAND2X1 NAND2X1_402 ( .A(u2_remHi_52_), .B(u2__abc_52138_new_n3311_), .Y(u2__abc_52138_new_n3312_));
NAND2X1 NAND2X1_403 ( .A(sqrto_52_), .B(u2__abc_52138_new_n3313_), .Y(u2__abc_52138_new_n3314_));
NAND2X1 NAND2X1_404 ( .A(u2__abc_52138_new_n3312_), .B(u2__abc_52138_new_n3314_), .Y(u2__abc_52138_new_n3315_));
NAND2X1 NAND2X1_405 ( .A(u2_remHi_53_), .B(u2__abc_52138_new_n3316_), .Y(u2__abc_52138_new_n3317_));
NAND2X1 NAND2X1_406 ( .A(sqrto_53_), .B(u2__abc_52138_new_n3318_), .Y(u2__abc_52138_new_n3319_));
NAND2X1 NAND2X1_407 ( .A(u2__abc_52138_new_n3317_), .B(u2__abc_52138_new_n3319_), .Y(u2__abc_52138_new_n3320_));
NAND2X1 NAND2X1_408 ( .A(u2_remHi_51_), .B(u2__abc_52138_new_n3322_), .Y(u2__abc_52138_new_n3323_));
NAND2X1 NAND2X1_409 ( .A(sqrto_51_), .B(u2__abc_52138_new_n3324_), .Y(u2__abc_52138_new_n3325_));
NAND2X1 NAND2X1_41 ( .A(aNan), .B(\a[40] ), .Y(_abc_65734_new_n951_));
NAND2X1 NAND2X1_410 ( .A(u2__abc_52138_new_n3323_), .B(u2__abc_52138_new_n3325_), .Y(u2__abc_52138_new_n3326_));
NAND2X1 NAND2X1_411 ( .A(u2_remHi_50_), .B(u2__abc_52138_new_n3327_), .Y(u2__abc_52138_new_n3328_));
NAND2X1 NAND2X1_412 ( .A(sqrto_50_), .B(u2__abc_52138_new_n3329_), .Y(u2__abc_52138_new_n3330_));
NAND2X1 NAND2X1_413 ( .A(u2__abc_52138_new_n3328_), .B(u2__abc_52138_new_n3330_), .Y(u2__abc_52138_new_n3331_));
NAND2X1 NAND2X1_414 ( .A(u2_remHi_40_), .B(u2__abc_52138_new_n3335_), .Y(u2__abc_52138_new_n3336_));
NAND2X1 NAND2X1_415 ( .A(sqrto_40_), .B(u2__abc_52138_new_n3337_), .Y(u2__abc_52138_new_n3338_));
NAND2X1 NAND2X1_416 ( .A(u2__abc_52138_new_n3336_), .B(u2__abc_52138_new_n3338_), .Y(u2__abc_52138_new_n3339_));
NAND2X1 NAND2X1_417 ( .A(u2_remHi_41_), .B(u2__abc_52138_new_n3340_), .Y(u2__abc_52138_new_n3341_));
NAND2X1 NAND2X1_418 ( .A(sqrto_41_), .B(u2__abc_52138_new_n3342_), .Y(u2__abc_52138_new_n3343_));
NAND2X1 NAND2X1_419 ( .A(u2__abc_52138_new_n3341_), .B(u2__abc_52138_new_n3343_), .Y(u2__abc_52138_new_n3344_));
NAND2X1 NAND2X1_42 ( .A(aNan), .B(\a[41] ), .Y(_abc_65734_new_n954_));
NAND2X1 NAND2X1_420 ( .A(u2_remHi_38_), .B(u2__abc_52138_new_n3346_), .Y(u2__abc_52138_new_n3347_));
NAND2X1 NAND2X1_421 ( .A(sqrto_38_), .B(u2__abc_52138_new_n3348_), .Y(u2__abc_52138_new_n3349_));
NAND2X1 NAND2X1_422 ( .A(u2__abc_52138_new_n3347_), .B(u2__abc_52138_new_n3349_), .Y(u2__abc_52138_new_n3350_));
NAND2X1 NAND2X1_423 ( .A(u2_remHi_39_), .B(u2__abc_52138_new_n3351_), .Y(u2__abc_52138_new_n3352_));
NAND2X1 NAND2X1_424 ( .A(sqrto_39_), .B(u2__abc_52138_new_n3353_), .Y(u2__abc_52138_new_n3354_));
NAND2X1 NAND2X1_425 ( .A(u2__abc_52138_new_n3352_), .B(u2__abc_52138_new_n3354_), .Y(u2__abc_52138_new_n3355_));
NAND2X1 NAND2X1_426 ( .A(u2__abc_52138_new_n3345_), .B(u2__abc_52138_new_n3356_), .Y(u2__abc_52138_new_n3357_));
NAND2X1 NAND2X1_427 ( .A(u2_remHi_44_), .B(u2__abc_52138_new_n3358_), .Y(u2__abc_52138_new_n3359_));
NAND2X1 NAND2X1_428 ( .A(sqrto_44_), .B(u2__abc_52138_new_n3360_), .Y(u2__abc_52138_new_n3361_));
NAND2X1 NAND2X1_429 ( .A(u2__abc_52138_new_n3359_), .B(u2__abc_52138_new_n3361_), .Y(u2__abc_52138_new_n3362_));
NAND2X1 NAND2X1_43 ( .A(aNan), .B(\a[42] ), .Y(_abc_65734_new_n957_));
NAND2X1 NAND2X1_430 ( .A(u2_remHi_45_), .B(u2__abc_52138_new_n3363_), .Y(u2__abc_52138_new_n3364_));
NAND2X1 NAND2X1_431 ( .A(sqrto_45_), .B(u2__abc_52138_new_n3365_), .Y(u2__abc_52138_new_n3366_));
NAND2X1 NAND2X1_432 ( .A(u2__abc_52138_new_n3364_), .B(u2__abc_52138_new_n3366_), .Y(u2__abc_52138_new_n3367_));
NAND2X1 NAND2X1_433 ( .A(u2_remHi_43_), .B(u2__abc_52138_new_n3369_), .Y(u2__abc_52138_new_n3370_));
NAND2X1 NAND2X1_434 ( .A(sqrto_43_), .B(u2__abc_52138_new_n3371_), .Y(u2__abc_52138_new_n3372_));
NAND2X1 NAND2X1_435 ( .A(u2__abc_52138_new_n3370_), .B(u2__abc_52138_new_n3372_), .Y(u2__abc_52138_new_n3373_));
NAND2X1 NAND2X1_436 ( .A(u2_remHi_42_), .B(u2__abc_52138_new_n3374_), .Y(u2__abc_52138_new_n3375_));
NAND2X1 NAND2X1_437 ( .A(sqrto_42_), .B(u2__abc_52138_new_n3376_), .Y(u2__abc_52138_new_n3377_));
NAND2X1 NAND2X1_438 ( .A(u2__abc_52138_new_n3375_), .B(u2__abc_52138_new_n3377_), .Y(u2__abc_52138_new_n3378_));
NAND2X1 NAND2X1_439 ( .A(u2__abc_52138_new_n3368_), .B(u2__abc_52138_new_n3379_), .Y(u2__abc_52138_new_n3380_));
NAND2X1 NAND2X1_44 ( .A(aNan), .B(\a[43] ), .Y(_abc_65734_new_n960_));
NAND2X1 NAND2X1_440 ( .A(u2_remHi_33_), .B(u2__abc_52138_new_n3383_), .Y(u2__abc_52138_new_n3384_));
NAND2X1 NAND2X1_441 ( .A(sqrto_33_), .B(u2__abc_52138_new_n3385_), .Y(u2__abc_52138_new_n3386_));
NAND2X1 NAND2X1_442 ( .A(u2__abc_52138_new_n3384_), .B(u2__abc_52138_new_n3386_), .Y(u2__abc_52138_new_n3387_));
NAND2X1 NAND2X1_443 ( .A(u2_remHi_30_), .B(u2__abc_52138_new_n3389_), .Y(u2__abc_52138_new_n3390_));
NAND2X1 NAND2X1_444 ( .A(sqrto_30_), .B(u2__abc_52138_new_n3391_), .Y(u2__abc_52138_new_n3392_));
NAND2X1 NAND2X1_445 ( .A(u2__abc_52138_new_n3390_), .B(u2__abc_52138_new_n3392_), .Y(u2__abc_52138_new_n3393_));
NAND2X1 NAND2X1_446 ( .A(u2_remHi_31_), .B(u2__abc_52138_new_n3394_), .Y(u2__abc_52138_new_n3395_));
NAND2X1 NAND2X1_447 ( .A(sqrto_31_), .B(u2__abc_52138_new_n3396_), .Y(u2__abc_52138_new_n3397_));
NAND2X1 NAND2X1_448 ( .A(u2__abc_52138_new_n3395_), .B(u2__abc_52138_new_n3397_), .Y(u2__abc_52138_new_n3398_));
NAND2X1 NAND2X1_449 ( .A(u2__abc_52138_new_n3388_), .B(u2__abc_52138_new_n3399_), .Y(u2__abc_52138_new_n3400_));
NAND2X1 NAND2X1_45 ( .A(aNan), .B(\a[44] ), .Y(_abc_65734_new_n963_));
NAND2X1 NAND2X1_450 ( .A(u2_remHi_36_), .B(u2__abc_52138_new_n3401_), .Y(u2__abc_52138_new_n3402_));
NAND2X1 NAND2X1_451 ( .A(sqrto_36_), .B(u2__abc_52138_new_n3403_), .Y(u2__abc_52138_new_n3404_));
NAND2X1 NAND2X1_452 ( .A(u2__abc_52138_new_n3402_), .B(u2__abc_52138_new_n3404_), .Y(u2__abc_52138_new_n3405_));
NAND2X1 NAND2X1_453 ( .A(u2_remHi_37_), .B(u2__abc_52138_new_n3406_), .Y(u2__abc_52138_new_n3407_));
NAND2X1 NAND2X1_454 ( .A(sqrto_37_), .B(u2__abc_52138_new_n3408_), .Y(u2__abc_52138_new_n3409_));
NAND2X1 NAND2X1_455 ( .A(u2__abc_52138_new_n3407_), .B(u2__abc_52138_new_n3409_), .Y(u2__abc_52138_new_n3410_));
NAND2X1 NAND2X1_456 ( .A(u2_remHi_35_), .B(u2__abc_52138_new_n3412_), .Y(u2__abc_52138_new_n3413_));
NAND2X1 NAND2X1_457 ( .A(sqrto_35_), .B(u2__abc_52138_new_n3414_), .Y(u2__abc_52138_new_n3415_));
NAND2X1 NAND2X1_458 ( .A(u2__abc_52138_new_n3381_), .B(u2__abc_52138_new_n3419_), .Y(u2__abc_52138_new_n3420_));
NAND2X1 NAND2X1_459 ( .A(u2__abc_52138_new_n3333_), .B(u2__abc_52138_new_n3310_), .Y(u2__abc_52138_new_n3423_));
NAND2X1 NAND2X1_46 ( .A(aNan), .B(\a[45] ), .Y(_abc_65734_new_n966_));
NAND2X1 NAND2X1_460 ( .A(u2__abc_52138_new_n3425_), .B(u2__abc_52138_new_n3426_), .Y(u2__abc_52138_new_n3427_));
NAND2X1 NAND2X1_461 ( .A(u2__abc_52138_new_n3417_), .B(u2__abc_52138_new_n3416_), .Y(u2__abc_52138_new_n3430_));
NAND2X1 NAND2X1_462 ( .A(sqrto_34_), .B(u2__abc_52138_new_n3443_), .Y(u2__abc_52138_new_n3444_));
NAND2X1 NAND2X1_463 ( .A(u2__abc_52138_new_n3461_), .B(u2__abc_52138_new_n3368_), .Y(u2__abc_52138_new_n3462_));
NAND2X1 NAND2X1_464 ( .A(u2__abc_52138_new_n3465_), .B(u2__abc_52138_new_n3462_), .Y(u2__abc_52138_new_n3466_));
NAND2X1 NAND2X1_465 ( .A(sqrto_48_), .B(u2__abc_52138_new_n3287_), .Y(u2__abc_52138_new_n3472_));
NAND2X1 NAND2X1_466 ( .A(sqrto_49_), .B(u2__abc_52138_new_n3292_), .Y(u2__abc_52138_new_n3473_));
NAND2X1 NAND2X1_467 ( .A(u2__abc_52138_new_n3495_), .B(u2__abc_52138_new_n3273_), .Y(u2__abc_52138_new_n3496_));
NAND2X1 NAND2X1_468 ( .A(sqrto_118_), .B(u2__abc_52138_new_n3503_), .Y(u2__abc_52138_new_n3506_));
NAND2X1 NAND2X1_469 ( .A(u2__abc_52138_new_n3506_), .B(u2__abc_52138_new_n3505_), .Y(u2__abc_52138_new_n3507_));
NAND2X1 NAND2X1_47 ( .A(aNan), .B(\a[46] ), .Y(_abc_65734_new_n969_));
NAND2X1 NAND2X1_470 ( .A(u2__abc_52138_new_n3510_), .B(u2__abc_52138_new_n3513_), .Y(u2__abc_52138_new_n3514_));
NAND2X1 NAND2X1_471 ( .A(u2_remHi_120_), .B(u2__abc_52138_new_n3516_), .Y(u2__abc_52138_new_n3517_));
NAND2X1 NAND2X1_472 ( .A(sqrto_120_), .B(u2__abc_52138_new_n3518_), .Y(u2__abc_52138_new_n3519_));
NAND2X1 NAND2X1_473 ( .A(u2__abc_52138_new_n3517_), .B(u2__abc_52138_new_n3519_), .Y(u2__abc_52138_new_n3520_));
NAND2X1 NAND2X1_474 ( .A(u2_remHi_121_), .B(u2__abc_52138_new_n3521_), .Y(u2__abc_52138_new_n3522_));
NAND2X1 NAND2X1_475 ( .A(sqrto_121_), .B(u2__abc_52138_new_n3523_), .Y(u2__abc_52138_new_n3524_));
NAND2X1 NAND2X1_476 ( .A(u2__abc_52138_new_n3522_), .B(u2__abc_52138_new_n3524_), .Y(u2__abc_52138_new_n3525_));
NAND2X1 NAND2X1_477 ( .A(u2_remHi_124_), .B(u2__abc_52138_new_n3527_), .Y(u2__abc_52138_new_n3528_));
NAND2X1 NAND2X1_478 ( .A(sqrto_124_), .B(u2__abc_52138_new_n3529_), .Y(u2__abc_52138_new_n3530_));
NAND2X1 NAND2X1_479 ( .A(u2__abc_52138_new_n3528_), .B(u2__abc_52138_new_n3530_), .Y(u2__abc_52138_new_n3531_));
NAND2X1 NAND2X1_48 ( .A(aNan), .B(\a[47] ), .Y(_abc_65734_new_n972_));
NAND2X1 NAND2X1_480 ( .A(sqrto_125_), .B(u2__abc_52138_new_n3532_), .Y(u2__abc_52138_new_n3533_));
NAND2X1 NAND2X1_481 ( .A(u2_remHi_125_), .B(u2__abc_52138_new_n3534_), .Y(u2__abc_52138_new_n3535_));
NAND2X1 NAND2X1_482 ( .A(u2__abc_52138_new_n3533_), .B(u2__abc_52138_new_n3535_), .Y(u2__abc_52138_new_n3536_));
NAND2X1 NAND2X1_483 ( .A(u2_remHi_123_), .B(u2__abc_52138_new_n3538_), .Y(u2__abc_52138_new_n3539_));
NAND2X1 NAND2X1_484 ( .A(sqrto_123_), .B(u2__abc_52138_new_n3540_), .Y(u2__abc_52138_new_n3541_));
NAND2X1 NAND2X1_485 ( .A(u2_remHi_110_), .B(u2__abc_52138_new_n3550_), .Y(u2__abc_52138_new_n3551_));
NAND2X1 NAND2X1_486 ( .A(sqrto_110_), .B(u2__abc_52138_new_n3552_), .Y(u2__abc_52138_new_n3553_));
NAND2X1 NAND2X1_487 ( .A(u2__abc_52138_new_n3551_), .B(u2__abc_52138_new_n3553_), .Y(u2__abc_52138_new_n3554_));
NAND2X1 NAND2X1_488 ( .A(u2_remHi_111_), .B(u2__abc_52138_new_n3555_), .Y(u2__abc_52138_new_n3556_));
NAND2X1 NAND2X1_489 ( .A(sqrto_111_), .B(u2__abc_52138_new_n3557_), .Y(u2__abc_52138_new_n3558_));
NAND2X1 NAND2X1_49 ( .A(aNan), .B(\a[48] ), .Y(_abc_65734_new_n975_));
NAND2X1 NAND2X1_490 ( .A(u2__abc_52138_new_n3556_), .B(u2__abc_52138_new_n3558_), .Y(u2__abc_52138_new_n3559_));
NAND2X1 NAND2X1_491 ( .A(u2_remHi_112_), .B(u2__abc_52138_new_n3561_), .Y(u2__abc_52138_new_n3562_));
NAND2X1 NAND2X1_492 ( .A(sqrto_112_), .B(u2__abc_52138_new_n3563_), .Y(u2__abc_52138_new_n3564_));
NAND2X1 NAND2X1_493 ( .A(u2__abc_52138_new_n3562_), .B(u2__abc_52138_new_n3564_), .Y(u2__abc_52138_new_n3565_));
NAND2X1 NAND2X1_494 ( .A(u2_remHi_113_), .B(u2__abc_52138_new_n3566_), .Y(u2__abc_52138_new_n3567_));
NAND2X1 NAND2X1_495 ( .A(sqrto_113_), .B(u2__abc_52138_new_n3568_), .Y(u2__abc_52138_new_n3569_));
NAND2X1 NAND2X1_496 ( .A(u2__abc_52138_new_n3567_), .B(u2__abc_52138_new_n3569_), .Y(u2__abc_52138_new_n3570_));
NAND2X1 NAND2X1_497 ( .A(u2_remHi_117_), .B(u2__abc_52138_new_n3578_), .Y(u2__abc_52138_new_n3579_));
NAND2X1 NAND2X1_498 ( .A(sqrto_117_), .B(u2__abc_52138_new_n3580_), .Y(u2__abc_52138_new_n3581_));
NAND2X1 NAND2X1_499 ( .A(u2_remHi_115_), .B(u2__abc_52138_new_n3583_), .Y(u2__abc_52138_new_n3584_));
NAND2X1 NAND2X1_5 ( .A(aNan), .B(\a[4] ), .Y(_abc_65734_new_n843_));
NAND2X1 NAND2X1_50 ( .A(aNan), .B(\a[49] ), .Y(_abc_65734_new_n978_));
NAND2X1 NAND2X1_500 ( .A(sqrto_115_), .B(u2__abc_52138_new_n3585_), .Y(u2__abc_52138_new_n3586_));
NAND2X1 NAND2X1_501 ( .A(u2__abc_52138_new_n3584_), .B(u2__abc_52138_new_n3586_), .Y(u2__abc_52138_new_n3587_));
NAND2X1 NAND2X1_502 ( .A(u2_remHi_114_), .B(u2__abc_52138_new_n3588_), .Y(u2__abc_52138_new_n3589_));
NAND2X1 NAND2X1_503 ( .A(sqrto_114_), .B(u2__abc_52138_new_n3590_), .Y(u2__abc_52138_new_n3591_));
NAND2X1 NAND2X1_504 ( .A(u2__abc_52138_new_n3589_), .B(u2__abc_52138_new_n3591_), .Y(u2__abc_52138_new_n3592_));
NAND2X1 NAND2X1_505 ( .A(u2__abc_52138_new_n3572_), .B(u2__abc_52138_new_n3594_), .Y(u2__abc_52138_new_n3595_));
NAND2X1 NAND2X1_506 ( .A(u2_remHi_104_), .B(u2__abc_52138_new_n3597_), .Y(u2__abc_52138_new_n3598_));
NAND2X1 NAND2X1_507 ( .A(sqrto_104_), .B(u2__abc_52138_new_n3599_), .Y(u2__abc_52138_new_n3600_));
NAND2X1 NAND2X1_508 ( .A(u2__abc_52138_new_n3598_), .B(u2__abc_52138_new_n3600_), .Y(u2__abc_52138_new_n3601_));
NAND2X1 NAND2X1_509 ( .A(u2_remHi_105_), .B(u2__abc_52138_new_n3602_), .Y(u2__abc_52138_new_n3603_));
NAND2X1 NAND2X1_51 ( .A(aNan), .B(\a[50] ), .Y(_abc_65734_new_n981_));
NAND2X1 NAND2X1_510 ( .A(sqrto_105_), .B(u2__abc_52138_new_n3604_), .Y(u2__abc_52138_new_n3605_));
NAND2X1 NAND2X1_511 ( .A(u2__abc_52138_new_n3603_), .B(u2__abc_52138_new_n3605_), .Y(u2__abc_52138_new_n3606_));
NAND2X1 NAND2X1_512 ( .A(u2_remHi_103_), .B(u2__abc_52138_new_n3608_), .Y(u2__abc_52138_new_n3609_));
NAND2X1 NAND2X1_513 ( .A(sqrto_103_), .B(u2__abc_52138_new_n3610_), .Y(u2__abc_52138_new_n3611_));
NAND2X1 NAND2X1_514 ( .A(u2_remHi_108_), .B(u2__abc_52138_new_n3619_), .Y(u2__abc_52138_new_n3620_));
NAND2X1 NAND2X1_515 ( .A(sqrto_108_), .B(u2__abc_52138_new_n3621_), .Y(u2__abc_52138_new_n3622_));
NAND2X1 NAND2X1_516 ( .A(u2__abc_52138_new_n3620_), .B(u2__abc_52138_new_n3622_), .Y(u2__abc_52138_new_n3623_));
NAND2X1 NAND2X1_517 ( .A(u2_remHi_109_), .B(u2__abc_52138_new_n3624_), .Y(u2__abc_52138_new_n3625_));
NAND2X1 NAND2X1_518 ( .A(sqrto_109_), .B(u2__abc_52138_new_n3626_), .Y(u2__abc_52138_new_n3627_));
NAND2X1 NAND2X1_519 ( .A(u2__abc_52138_new_n3625_), .B(u2__abc_52138_new_n3627_), .Y(u2__abc_52138_new_n3628_));
NAND2X1 NAND2X1_52 ( .A(aNan), .B(\a[51] ), .Y(_abc_65734_new_n984_));
NAND2X1 NAND2X1_520 ( .A(u2_remHi_107_), .B(u2__abc_52138_new_n3630_), .Y(u2__abc_52138_new_n3631_));
NAND2X1 NAND2X1_521 ( .A(sqrto_107_), .B(u2__abc_52138_new_n3632_), .Y(u2__abc_52138_new_n3633_));
NAND2X1 NAND2X1_522 ( .A(u2__abc_52138_new_n3618_), .B(u2__abc_52138_new_n3640_), .Y(u2__abc_52138_new_n3641_));
NAND2X1 NAND2X1_523 ( .A(u2__abc_52138_new_n3646_), .B(u2__abc_52138_new_n3651_), .Y(u2__abc_52138_new_n3652_));
NAND2X1 NAND2X1_524 ( .A(u2_remHi_95_), .B(u2__abc_52138_new_n3653_), .Y(u2__abc_52138_new_n3654_));
NAND2X1 NAND2X1_525 ( .A(sqrto_95_), .B(u2__abc_52138_new_n3655_), .Y(u2__abc_52138_new_n3656_));
NAND2X1 NAND2X1_526 ( .A(u2__abc_52138_new_n3654_), .B(u2__abc_52138_new_n3656_), .Y(u2__abc_52138_new_n3657_));
NAND2X1 NAND2X1_527 ( .A(u2_remHi_94_), .B(u2__abc_52138_new_n3658_), .Y(u2__abc_52138_new_n3659_));
NAND2X1 NAND2X1_528 ( .A(sqrto_94_), .B(u2__abc_52138_new_n3660_), .Y(u2__abc_52138_new_n3661_));
NAND2X1 NAND2X1_529 ( .A(u2__abc_52138_new_n3659_), .B(u2__abc_52138_new_n3661_), .Y(u2__abc_52138_new_n3662_));
NAND2X1 NAND2X1_53 ( .A(aNan), .B(\a[52] ), .Y(_abc_65734_new_n987_));
NAND2X1 NAND2X1_530 ( .A(u2_remHi_100_), .B(u2__abc_52138_new_n3665_), .Y(u2__abc_52138_new_n3666_));
NAND2X1 NAND2X1_531 ( .A(sqrto_100_), .B(u2__abc_52138_new_n3667_), .Y(u2__abc_52138_new_n3668_));
NAND2X1 NAND2X1_532 ( .A(u2__abc_52138_new_n3666_), .B(u2__abc_52138_new_n3668_), .Y(u2__abc_52138_new_n3669_));
NAND2X1 NAND2X1_533 ( .A(u2_remHi_101_), .B(u2__abc_52138_new_n3670_), .Y(u2__abc_52138_new_n3671_));
NAND2X1 NAND2X1_534 ( .A(sqrto_101_), .B(u2__abc_52138_new_n3672_), .Y(u2__abc_52138_new_n3673_));
NAND2X1 NAND2X1_535 ( .A(u2__abc_52138_new_n3671_), .B(u2__abc_52138_new_n3673_), .Y(u2__abc_52138_new_n3674_));
NAND2X1 NAND2X1_536 ( .A(u2_remHi_99_), .B(u2__abc_52138_new_n3676_), .Y(u2__abc_52138_new_n3677_));
NAND2X1 NAND2X1_537 ( .A(sqrto_99_), .B(u2__abc_52138_new_n3678_), .Y(u2__abc_52138_new_n3679_));
NAND2X1 NAND2X1_538 ( .A(u2__abc_52138_new_n3677_), .B(u2__abc_52138_new_n3679_), .Y(u2__abc_52138_new_n3680_));
NAND2X1 NAND2X1_539 ( .A(u2_remHi_98_), .B(u2__abc_52138_new_n3681_), .Y(u2__abc_52138_new_n3682_));
NAND2X1 NAND2X1_54 ( .A(aNan), .B(\a[53] ), .Y(_abc_65734_new_n990_));
NAND2X1 NAND2X1_540 ( .A(sqrto_98_), .B(u2__abc_52138_new_n3683_), .Y(u2__abc_52138_new_n3684_));
NAND2X1 NAND2X1_541 ( .A(u2__abc_52138_new_n3682_), .B(u2__abc_52138_new_n3684_), .Y(u2__abc_52138_new_n3685_));
NAND2X1 NAND2X1_542 ( .A(u2__abc_52138_new_n3687_), .B(u2__abc_52138_new_n3664_), .Y(u2__abc_52138_new_n3688_));
NAND2X1 NAND2X1_543 ( .A(u2__abc_52138_new_n3689_), .B(u2__abc_52138_new_n3596_), .Y(u2__abc_52138_new_n3690_));
NAND2X1 NAND2X1_544 ( .A(u2_remHi_92_), .B(u2__abc_52138_new_n3691_), .Y(u2__abc_52138_new_n3692_));
NAND2X1 NAND2X1_545 ( .A(sqrto_92_), .B(u2__abc_52138_new_n3693_), .Y(u2__abc_52138_new_n3694_));
NAND2X1 NAND2X1_546 ( .A(u2__abc_52138_new_n3692_), .B(u2__abc_52138_new_n3694_), .Y(u2__abc_52138_new_n3695_));
NAND2X1 NAND2X1_547 ( .A(u2_remHi_93_), .B(u2__abc_52138_new_n3696_), .Y(u2__abc_52138_new_n3697_));
NAND2X1 NAND2X1_548 ( .A(sqrto_93_), .B(u2__abc_52138_new_n3698_), .Y(u2__abc_52138_new_n3699_));
NAND2X1 NAND2X1_549 ( .A(u2__abc_52138_new_n3697_), .B(u2__abc_52138_new_n3699_), .Y(u2__abc_52138_new_n3700_));
NAND2X1 NAND2X1_55 ( .A(aNan), .B(\a[54] ), .Y(_abc_65734_new_n993_));
NAND2X1 NAND2X1_550 ( .A(u2_remHi_91_), .B(u2__abc_52138_new_n3702_), .Y(u2__abc_52138_new_n3703_));
NAND2X1 NAND2X1_551 ( .A(sqrto_91_), .B(u2__abc_52138_new_n3704_), .Y(u2__abc_52138_new_n3705_));
NAND2X1 NAND2X1_552 ( .A(u2_remHi_88_), .B(u2__abc_52138_new_n3713_), .Y(u2__abc_52138_new_n3714_));
NAND2X1 NAND2X1_553 ( .A(sqrto_88_), .B(u2__abc_52138_new_n3715_), .Y(u2__abc_52138_new_n3716_));
NAND2X1 NAND2X1_554 ( .A(u2__abc_52138_new_n3714_), .B(u2__abc_52138_new_n3716_), .Y(u2__abc_52138_new_n3717_));
NAND2X1 NAND2X1_555 ( .A(u2_remHi_89_), .B(u2__abc_52138_new_n3718_), .Y(u2__abc_52138_new_n3719_));
NAND2X1 NAND2X1_556 ( .A(sqrto_89_), .B(u2__abc_52138_new_n3720_), .Y(u2__abc_52138_new_n3721_));
NAND2X1 NAND2X1_557 ( .A(u2__abc_52138_new_n3719_), .B(u2__abc_52138_new_n3721_), .Y(u2__abc_52138_new_n3722_));
NAND2X1 NAND2X1_558 ( .A(u2__abc_52138_new_n3712_), .B(u2__abc_52138_new_n3736_), .Y(u2__abc_52138_new_n3737_));
NAND2X1 NAND2X1_559 ( .A(u2_remHi_78_), .B(u2__abc_52138_new_n3738_), .Y(u2__abc_52138_new_n3739_));
NAND2X1 NAND2X1_56 ( .A(aNan), .B(\a[55] ), .Y(_abc_65734_new_n996_));
NAND2X1 NAND2X1_560 ( .A(sqrto_78_), .B(u2__abc_52138_new_n3740_), .Y(u2__abc_52138_new_n3741_));
NAND2X1 NAND2X1_561 ( .A(u2__abc_52138_new_n3739_), .B(u2__abc_52138_new_n3741_), .Y(u2__abc_52138_new_n3742_));
NAND2X1 NAND2X1_562 ( .A(u2_remHi_79_), .B(u2__abc_52138_new_n3743_), .Y(u2__abc_52138_new_n3744_));
NAND2X1 NAND2X1_563 ( .A(sqrto_79_), .B(u2__abc_52138_new_n3745_), .Y(u2__abc_52138_new_n3746_));
NAND2X1 NAND2X1_564 ( .A(u2__abc_52138_new_n3744_), .B(u2__abc_52138_new_n3746_), .Y(u2__abc_52138_new_n3747_));
NAND2X1 NAND2X1_565 ( .A(u2_remHi_80_), .B(u2__abc_52138_new_n3749_), .Y(u2__abc_52138_new_n3750_));
NAND2X1 NAND2X1_566 ( .A(sqrto_80_), .B(u2__abc_52138_new_n3751_), .Y(u2__abc_52138_new_n3752_));
NAND2X1 NAND2X1_567 ( .A(u2_remHi_81_), .B(u2__abc_52138_new_n3754_), .Y(u2__abc_52138_new_n3755_));
NAND2X1 NAND2X1_568 ( .A(sqrto_81_), .B(u2__abc_52138_new_n3756_), .Y(u2__abc_52138_new_n3757_));
NAND2X1 NAND2X1_569 ( .A(u2__abc_52138_new_n3753_), .B(u2__abc_52138_new_n3758_), .Y(u2__abc_52138_new_n3759_));
NAND2X1 NAND2X1_57 ( .A(aNan), .B(\a[56] ), .Y(_abc_65734_new_n999_));
NAND2X1 NAND2X1_570 ( .A(u2_remHi_84_), .B(u2__abc_52138_new_n3761_), .Y(u2__abc_52138_new_n3762_));
NAND2X1 NAND2X1_571 ( .A(sqrto_84_), .B(u2__abc_52138_new_n3763_), .Y(u2__abc_52138_new_n3764_));
NAND2X1 NAND2X1_572 ( .A(u2__abc_52138_new_n3762_), .B(u2__abc_52138_new_n3764_), .Y(u2__abc_52138_new_n3765_));
NAND2X1 NAND2X1_573 ( .A(u2_remHi_85_), .B(u2__abc_52138_new_n3766_), .Y(u2__abc_52138_new_n3767_));
NAND2X1 NAND2X1_574 ( .A(sqrto_85_), .B(u2__abc_52138_new_n3768_), .Y(u2__abc_52138_new_n3769_));
NAND2X1 NAND2X1_575 ( .A(u2__abc_52138_new_n3767_), .B(u2__abc_52138_new_n3769_), .Y(u2__abc_52138_new_n3770_));
NAND2X1 NAND2X1_576 ( .A(u2_remHi_83_), .B(u2__abc_52138_new_n3772_), .Y(u2__abc_52138_new_n3773_));
NAND2X1 NAND2X1_577 ( .A(sqrto_83_), .B(u2__abc_52138_new_n3774_), .Y(u2__abc_52138_new_n3775_));
NAND2X1 NAND2X1_578 ( .A(u2__abc_52138_new_n3773_), .B(u2__abc_52138_new_n3775_), .Y(u2__abc_52138_new_n3776_));
NAND2X1 NAND2X1_579 ( .A(u2_remHi_82_), .B(u2__abc_52138_new_n3777_), .Y(u2__abc_52138_new_n3778_));
NAND2X1 NAND2X1_58 ( .A(aNan), .B(\a[57] ), .Y(_abc_65734_new_n1002_));
NAND2X1 NAND2X1_580 ( .A(sqrto_82_), .B(u2__abc_52138_new_n3779_), .Y(u2__abc_52138_new_n3780_));
NAND2X1 NAND2X1_581 ( .A(u2__abc_52138_new_n3778_), .B(u2__abc_52138_new_n3780_), .Y(u2__abc_52138_new_n3781_));
NAND2X1 NAND2X1_582 ( .A(u2__abc_52138_new_n3783_), .B(u2__abc_52138_new_n3760_), .Y(u2__abc_52138_new_n3784_));
NAND2X1 NAND2X1_583 ( .A(u2__abc_52138_new_n3790_), .B(u2__abc_52138_new_n3795_), .Y(u2__abc_52138_new_n3796_));
NAND2X1 NAND2X1_584 ( .A(u2_remHi_72_), .B(u2__abc_52138_new_n3797_), .Y(u2__abc_52138_new_n3798_));
NAND2X1 NAND2X1_585 ( .A(sqrto_72_), .B(u2__abc_52138_new_n3799_), .Y(u2__abc_52138_new_n3800_));
NAND2X1 NAND2X1_586 ( .A(u2_remHi_73_), .B(u2__abc_52138_new_n3802_), .Y(u2__abc_52138_new_n3803_));
NAND2X1 NAND2X1_587 ( .A(sqrto_73_), .B(u2__abc_52138_new_n3804_), .Y(u2__abc_52138_new_n3805_));
NAND2X1 NAND2X1_588 ( .A(u2__abc_52138_new_n3812_), .B(u2__abc_52138_new_n3817_), .Y(u2__abc_52138_new_n3818_));
NAND2X1 NAND2X1_589 ( .A(u2__abc_52138_new_n3823_), .B(u2__abc_52138_new_n3828_), .Y(u2__abc_52138_new_n3829_));
NAND2X1 NAND2X1_59 ( .A(aNan), .B(\a[58] ), .Y(_abc_65734_new_n1005_));
NAND2X1 NAND2X1_590 ( .A(u2__abc_52138_new_n3807_), .B(u2__abc_52138_new_n3830_), .Y(u2__abc_52138_new_n3831_));
NAND2X1 NAND2X1_591 ( .A(u2_remHi_62_), .B(u2__abc_52138_new_n3832_), .Y(u2__abc_52138_new_n3833_));
NAND2X1 NAND2X1_592 ( .A(sqrto_62_), .B(u2__abc_52138_new_n3834_), .Y(u2__abc_52138_new_n3835_));
NAND2X1 NAND2X1_593 ( .A(u2__abc_52138_new_n3833_), .B(u2__abc_52138_new_n3835_), .Y(u2__abc_52138_new_n3836_));
NAND2X1 NAND2X1_594 ( .A(u2_remHi_63_), .B(u2__abc_52138_new_n3837_), .Y(u2__abc_52138_new_n3838_));
NAND2X1 NAND2X1_595 ( .A(sqrto_63_), .B(u2__abc_52138_new_n3839_), .Y(u2__abc_52138_new_n3840_));
NAND2X1 NAND2X1_596 ( .A(u2__abc_52138_new_n3838_), .B(u2__abc_52138_new_n3840_), .Y(u2__abc_52138_new_n3841_));
NAND2X1 NAND2X1_597 ( .A(u2_remHi_64_), .B(u2__abc_52138_new_n3843_), .Y(u2__abc_52138_new_n3844_));
NAND2X1 NAND2X1_598 ( .A(sqrto_64_), .B(u2__abc_52138_new_n3845_), .Y(u2__abc_52138_new_n3846_));
NAND2X1 NAND2X1_599 ( .A(u2__abc_52138_new_n3844_), .B(u2__abc_52138_new_n3846_), .Y(u2__abc_52138_new_n3847_));
NAND2X1 NAND2X1_6 ( .A(aNan), .B(\a[5] ), .Y(_abc_65734_new_n846_));
NAND2X1 NAND2X1_60 ( .A(aNan), .B(\a[59] ), .Y(_abc_65734_new_n1008_));
NAND2X1 NAND2X1_600 ( .A(u2_remHi_65_), .B(u2__abc_52138_new_n3848_), .Y(u2__abc_52138_new_n3849_));
NAND2X1 NAND2X1_601 ( .A(sqrto_65_), .B(u2__abc_52138_new_n3850_), .Y(u2__abc_52138_new_n3851_));
NAND2X1 NAND2X1_602 ( .A(u2__abc_52138_new_n3849_), .B(u2__abc_52138_new_n3851_), .Y(u2__abc_52138_new_n3852_));
NAND2X1 NAND2X1_603 ( .A(u2_remHi_69_), .B(u2__abc_52138_new_n3856_), .Y(u2__abc_52138_new_n3857_));
NAND2X1 NAND2X1_604 ( .A(sqrto_69_), .B(u2__abc_52138_new_n3858_), .Y(u2__abc_52138_new_n3859_));
NAND2X1 NAND2X1_605 ( .A(u2_remHi_66_), .B(u2__abc_52138_new_n3862_), .Y(u2__abc_52138_new_n3863_));
NAND2X1 NAND2X1_606 ( .A(sqrto_66_), .B(u2__abc_52138_new_n3864_), .Y(u2__abc_52138_new_n3865_));
NAND2X1 NAND2X1_607 ( .A(u2__abc_52138_new_n3867_), .B(u2__abc_52138_new_n3854_), .Y(u2__abc_52138_new_n3868_));
NAND2X1 NAND2X1_608 ( .A(u2__abc_52138_new_n3869_), .B(u2__abc_52138_new_n3785_), .Y(u2__abc_52138_new_n3870_));
NAND2X1 NAND2X1_609 ( .A(u2_remHi_67_), .B(u2__abc_52138_new_n3881_), .Y(u2__abc_52138_new_n3882_));
NAND2X1 NAND2X1_61 ( .A(aNan), .B(\a[60] ), .Y(_abc_65734_new_n1011_));
NAND2X1 NAND2X1_610 ( .A(sqrto_67_), .B(u2__abc_52138_new_n3883_), .Y(u2__abc_52138_new_n3884_));
NAND2X1 NAND2X1_611 ( .A(sqrto_68_), .B(u2__abc_52138_new_n3888_), .Y(u2__abc_52138_new_n3889_));
NAND2X1 NAND2X1_612 ( .A(u2_remHi_77_), .B(u2__abc_52138_new_n3815_), .Y(u2__abc_52138_new_n3903_));
NAND2X1 NAND2X1_613 ( .A(u2__abc_52138_new_n3928_), .B(u2__abc_52138_new_n3930_), .Y(u2__abc_52138_new_n3931_));
NAND2X1 NAND2X1_614 ( .A(u2__abc_52138_new_n3934_), .B(u2__abc_52138_new_n3931_), .Y(u2__abc_52138_new_n3935_));
NAND2X1 NAND2X1_615 ( .A(sqrto_96_), .B(u2__abc_52138_new_n3642_), .Y(u2__abc_52138_new_n3942_));
NAND2X1 NAND2X1_616 ( .A(sqrto_97_), .B(u2__abc_52138_new_n3647_), .Y(u2__abc_52138_new_n3943_));
NAND2X1 NAND2X1_617 ( .A(u2__abc_52138_new_n3962_), .B(u2__abc_52138_new_n3964_), .Y(u2__abc_52138_new_n3965_));
NAND2X1 NAND2X1_618 ( .A(u2__abc_52138_new_n3987_), .B(u2__abc_52138_new_n3526_), .Y(u2__abc_52138_new_n3988_));
NAND2X1 NAND2X1_619 ( .A(u2_remHi_246_), .B(u2__abc_52138_new_n4003_), .Y(u2__abc_52138_new_n4004_));
NAND2X1 NAND2X1_62 ( .A(aNan), .B(\a[61] ), .Y(_abc_65734_new_n1014_));
NAND2X1 NAND2X1_620 ( .A(u2_o_246_), .B(u2__abc_52138_new_n4005_), .Y(u2__abc_52138_new_n4006_));
NAND2X1 NAND2X1_621 ( .A(u2__abc_52138_new_n4004_), .B(u2__abc_52138_new_n4006_), .Y(u2__abc_52138_new_n4007_));
NAND2X1 NAND2X1_622 ( .A(u2_remHi_247_), .B(u2__abc_52138_new_n4008_), .Y(u2__abc_52138_new_n4009_));
NAND2X1 NAND2X1_623 ( .A(u2_o_247_), .B(u2__abc_52138_new_n4010_), .Y(u2__abc_52138_new_n4011_));
NAND2X1 NAND2X1_624 ( .A(u2__abc_52138_new_n4009_), .B(u2__abc_52138_new_n4011_), .Y(u2__abc_52138_new_n4012_));
NAND2X1 NAND2X1_625 ( .A(u2_remHi_248_), .B(u2__abc_52138_new_n4014_), .Y(u2__abc_52138_new_n4015_));
NAND2X1 NAND2X1_626 ( .A(u2_o_248_), .B(u2__abc_52138_new_n4016_), .Y(u2__abc_52138_new_n4017_));
NAND2X1 NAND2X1_627 ( .A(u2__abc_52138_new_n4015_), .B(u2__abc_52138_new_n4017_), .Y(u2__abc_52138_new_n4018_));
NAND2X1 NAND2X1_628 ( .A(u2_remHi_249_), .B(u2__abc_52138_new_n4019_), .Y(u2__abc_52138_new_n4020_));
NAND2X1 NAND2X1_629 ( .A(u2_o_249_), .B(u2__abc_52138_new_n4021_), .Y(u2__abc_52138_new_n4022_));
NAND2X1 NAND2X1_63 ( .A(aNan), .B(\a[62] ), .Y(_abc_65734_new_n1017_));
NAND2X1 NAND2X1_630 ( .A(u2__abc_52138_new_n4020_), .B(u2__abc_52138_new_n4022_), .Y(u2__abc_52138_new_n4023_));
NAND2X1 NAND2X1_631 ( .A(u2__abc_52138_new_n4013_), .B(u2__abc_52138_new_n4024_), .Y(u2__abc_52138_new_n4025_));
NAND2X1 NAND2X1_632 ( .A(u2_remHi_252_), .B(u2__abc_52138_new_n4026_), .Y(u2__abc_52138_new_n4027_));
NAND2X1 NAND2X1_633 ( .A(u2_o_252_), .B(u2__abc_52138_new_n4028_), .Y(u2__abc_52138_new_n4029_));
NAND2X1 NAND2X1_634 ( .A(u2__abc_52138_new_n4027_), .B(u2__abc_52138_new_n4029_), .Y(u2__abc_52138_new_n4030_));
NAND2X1 NAND2X1_635 ( .A(u2_o_253_), .B(u2__abc_52138_new_n4031_), .Y(u2__abc_52138_new_n4032_));
NAND2X1 NAND2X1_636 ( .A(u2_remHi_253_), .B(u2__abc_52138_new_n4033_), .Y(u2__abc_52138_new_n4034_));
NAND2X1 NAND2X1_637 ( .A(u2__abc_52138_new_n4032_), .B(u2__abc_52138_new_n4034_), .Y(u2__abc_52138_new_n4035_));
NAND2X1 NAND2X1_638 ( .A(u2_remHi_251_), .B(u2__abc_52138_new_n4037_), .Y(u2__abc_52138_new_n4038_));
NAND2X1 NAND2X1_639 ( .A(u2_o_251_), .B(u2__abc_52138_new_n4039_), .Y(u2__abc_52138_new_n4040_));
NAND2X1 NAND2X1_64 ( .A(aNan), .B(\a[63] ), .Y(_abc_65734_new_n1020_));
NAND2X1 NAND2X1_640 ( .A(u2__abc_52138_new_n4038_), .B(u2__abc_52138_new_n4040_), .Y(u2__abc_52138_new_n4041_));
NAND2X1 NAND2X1_641 ( .A(u2_remHi_250_), .B(u2__abc_52138_new_n4042_), .Y(u2__abc_52138_new_n4043_));
NAND2X1 NAND2X1_642 ( .A(u2_o_250_), .B(u2__abc_52138_new_n4044_), .Y(u2__abc_52138_new_n4045_));
NAND2X1 NAND2X1_643 ( .A(u2__abc_52138_new_n4043_), .B(u2__abc_52138_new_n4045_), .Y(u2__abc_52138_new_n4046_));
NAND2X1 NAND2X1_644 ( .A(u2__abc_52138_new_n4036_), .B(u2__abc_52138_new_n4047_), .Y(u2__abc_52138_new_n4048_));
NAND2X1 NAND2X1_645 ( .A(u2_remHi_238_), .B(u2__abc_52138_new_n4050_), .Y(u2__abc_52138_new_n4051_));
NAND2X1 NAND2X1_646 ( .A(u2_o_238_), .B(u2__abc_52138_new_n4052_), .Y(u2__abc_52138_new_n4053_));
NAND2X1 NAND2X1_647 ( .A(u2__abc_52138_new_n4051_), .B(u2__abc_52138_new_n4053_), .Y(u2__abc_52138_new_n4054_));
NAND2X1 NAND2X1_648 ( .A(u2_remHi_239_), .B(u2__abc_52138_new_n4055_), .Y(u2__abc_52138_new_n4056_));
NAND2X1 NAND2X1_649 ( .A(u2_o_239_), .B(u2__abc_52138_new_n4057_), .Y(u2__abc_52138_new_n4058_));
NAND2X1 NAND2X1_65 ( .A(aNan), .B(\a[64] ), .Y(_abc_65734_new_n1023_));
NAND2X1 NAND2X1_650 ( .A(u2__abc_52138_new_n4056_), .B(u2__abc_52138_new_n4058_), .Y(u2__abc_52138_new_n4059_));
NAND2X1 NAND2X1_651 ( .A(u2_remHi_240_), .B(u2__abc_52138_new_n4061_), .Y(u2__abc_52138_new_n4062_));
NAND2X1 NAND2X1_652 ( .A(u2_o_240_), .B(u2__abc_52138_new_n4063_), .Y(u2__abc_52138_new_n4064_));
NAND2X1 NAND2X1_653 ( .A(u2__abc_52138_new_n4062_), .B(u2__abc_52138_new_n4064_), .Y(u2__abc_52138_new_n4065_));
NAND2X1 NAND2X1_654 ( .A(u2_remHi_241_), .B(u2__abc_52138_new_n4066_), .Y(u2__abc_52138_new_n4067_));
NAND2X1 NAND2X1_655 ( .A(u2_o_241_), .B(u2__abc_52138_new_n4068_), .Y(u2__abc_52138_new_n4069_));
NAND2X1 NAND2X1_656 ( .A(u2__abc_52138_new_n4067_), .B(u2__abc_52138_new_n4069_), .Y(u2__abc_52138_new_n4070_));
NAND2X1 NAND2X1_657 ( .A(u2_remHi_244_), .B(u2__abc_52138_new_n4074_), .Y(u2__abc_52138_new_n4075_));
NAND2X1 NAND2X1_658 ( .A(u2_o_244_), .B(u2__abc_52138_new_n4076_), .Y(u2__abc_52138_new_n4077_));
NAND2X1 NAND2X1_659 ( .A(u2__abc_52138_new_n4075_), .B(u2__abc_52138_new_n4077_), .Y(u2__abc_52138_new_n4078_));
NAND2X1 NAND2X1_66 ( .A(aNan), .B(\a[65] ), .Y(_abc_65734_new_n1026_));
NAND2X1 NAND2X1_660 ( .A(u2_remHi_245_), .B(u2__abc_52138_new_n4079_), .Y(u2__abc_52138_new_n4080_));
NAND2X1 NAND2X1_661 ( .A(u2_o_245_), .B(u2__abc_52138_new_n4081_), .Y(u2__abc_52138_new_n4082_));
NAND2X1 NAND2X1_662 ( .A(u2__abc_52138_new_n4080_), .B(u2__abc_52138_new_n4082_), .Y(u2__abc_52138_new_n4083_));
NAND2X1 NAND2X1_663 ( .A(u2_remHi_242_), .B(u2__abc_52138_new_n4090_), .Y(u2__abc_52138_new_n4091_));
NAND2X1 NAND2X1_664 ( .A(u2_o_242_), .B(u2__abc_52138_new_n4092_), .Y(u2__abc_52138_new_n4093_));
NAND2X1 NAND2X1_665 ( .A(u2__abc_52138_new_n4096_), .B(u2__abc_52138_new_n4073_), .Y(u2__abc_52138_new_n4097_));
NAND2X1 NAND2X1_666 ( .A(u2_remHi_236_), .B(u2__abc_52138_new_n4099_), .Y(u2__abc_52138_new_n4100_));
NAND2X1 NAND2X1_667 ( .A(u2_o_236_), .B(u2__abc_52138_new_n4101_), .Y(u2__abc_52138_new_n4102_));
NAND2X1 NAND2X1_668 ( .A(u2__abc_52138_new_n4100_), .B(u2__abc_52138_new_n4102_), .Y(u2__abc_52138_new_n4103_));
NAND2X1 NAND2X1_669 ( .A(u2_remHi_237_), .B(u2__abc_52138_new_n4104_), .Y(u2__abc_52138_new_n4105_));
NAND2X1 NAND2X1_67 ( .A(aNan), .B(\a[66] ), .Y(_abc_65734_new_n1029_));
NAND2X1 NAND2X1_670 ( .A(u2_o_237_), .B(u2__abc_52138_new_n4106_), .Y(u2__abc_52138_new_n4107_));
NAND2X1 NAND2X1_671 ( .A(u2__abc_52138_new_n4105_), .B(u2__abc_52138_new_n4107_), .Y(u2__abc_52138_new_n4108_));
NAND2X1 NAND2X1_672 ( .A(u2_remHi_235_), .B(u2__abc_52138_new_n4110_), .Y(u2__abc_52138_new_n4111_));
NAND2X1 NAND2X1_673 ( .A(u2_o_235_), .B(u2__abc_52138_new_n4112_), .Y(u2__abc_52138_new_n4113_));
NAND2X1 NAND2X1_674 ( .A(u2__abc_52138_new_n4111_), .B(u2__abc_52138_new_n4113_), .Y(u2__abc_52138_new_n4114_));
NAND2X1 NAND2X1_675 ( .A(u2_remHi_234_), .B(u2__abc_52138_new_n4115_), .Y(u2__abc_52138_new_n4116_));
NAND2X1 NAND2X1_676 ( .A(u2_o_234_), .B(u2__abc_52138_new_n4117_), .Y(u2__abc_52138_new_n4118_));
NAND2X1 NAND2X1_677 ( .A(u2__abc_52138_new_n4116_), .B(u2__abc_52138_new_n4118_), .Y(u2__abc_52138_new_n4119_));
NAND2X1 NAND2X1_678 ( .A(u2__abc_52138_new_n4109_), .B(u2__abc_52138_new_n4120_), .Y(u2__abc_52138_new_n4121_));
NAND2X1 NAND2X1_679 ( .A(u2_remHi_232_), .B(u2__abc_52138_new_n4123_), .Y(u2__abc_52138_new_n4124_));
NAND2X1 NAND2X1_68 ( .A(aNan), .B(\a[67] ), .Y(_abc_65734_new_n1032_));
NAND2X1 NAND2X1_680 ( .A(u2_o_232_), .B(u2__abc_52138_new_n4125_), .Y(u2__abc_52138_new_n4126_));
NAND2X1 NAND2X1_681 ( .A(u2__abc_52138_new_n4124_), .B(u2__abc_52138_new_n4126_), .Y(u2__abc_52138_new_n4127_));
NAND2X1 NAND2X1_682 ( .A(u2_remHi_233_), .B(u2__abc_52138_new_n4128_), .Y(u2__abc_52138_new_n4129_));
NAND2X1 NAND2X1_683 ( .A(u2_o_233_), .B(u2__abc_52138_new_n4130_), .Y(u2__abc_52138_new_n4131_));
NAND2X1 NAND2X1_684 ( .A(u2__abc_52138_new_n4129_), .B(u2__abc_52138_new_n4131_), .Y(u2__abc_52138_new_n4132_));
NAND2X1 NAND2X1_685 ( .A(u2_o_231_), .B(u2__abc_52138_new_n4134_), .Y(u2__abc_52138_new_n4137_));
NAND2X1 NAND2X1_686 ( .A(u2__abc_52138_new_n4144_), .B(u2__abc_52138_new_n4122_), .Y(u2__abc_52138_new_n4145_));
NAND2X1 NAND2X1_687 ( .A(u2_remHi_224_), .B(u2__abc_52138_new_n4146_), .Y(u2__abc_52138_new_n4147_));
NAND2X1 NAND2X1_688 ( .A(sqrto_224_), .B(u2__abc_52138_new_n4148_), .Y(u2__abc_52138_new_n4149_));
NAND2X1 NAND2X1_689 ( .A(u2__abc_52138_new_n4147_), .B(u2__abc_52138_new_n4149_), .Y(u2__abc_52138_new_n4150_));
NAND2X1 NAND2X1_69 ( .A(aNan), .B(\a[68] ), .Y(_abc_65734_new_n1035_));
NAND2X1 NAND2X1_690 ( .A(u2_remHi_225_), .B(u2__abc_52138_new_n4151_), .Y(u2__abc_52138_new_n4152_));
NAND2X1 NAND2X1_691 ( .A(sqrto_225_), .B(u2__abc_52138_new_n4153_), .Y(u2__abc_52138_new_n4154_));
NAND2X1 NAND2X1_692 ( .A(u2__abc_52138_new_n4152_), .B(u2__abc_52138_new_n4154_), .Y(u2__abc_52138_new_n4155_));
NAND2X1 NAND2X1_693 ( .A(u2_remHi_223_), .B(u2__abc_52138_new_n4157_), .Y(u2__abc_52138_new_n4158_));
NAND2X1 NAND2X1_694 ( .A(sqrto_223_), .B(u2__abc_52138_new_n4159_), .Y(u2__abc_52138_new_n4160_));
NAND2X1 NAND2X1_695 ( .A(u2__abc_52138_new_n4158_), .B(u2__abc_52138_new_n4160_), .Y(u2__abc_52138_new_n4161_));
NAND2X1 NAND2X1_696 ( .A(u2_remHi_222_), .B(u2__abc_52138_new_n4162_), .Y(u2__abc_52138_new_n4163_));
NAND2X1 NAND2X1_697 ( .A(sqrto_222_), .B(u2__abc_52138_new_n4164_), .Y(u2__abc_52138_new_n4165_));
NAND2X1 NAND2X1_698 ( .A(u2__abc_52138_new_n4163_), .B(u2__abc_52138_new_n4165_), .Y(u2__abc_52138_new_n4166_));
NAND2X1 NAND2X1_699 ( .A(u2__abc_52138_new_n4156_), .B(u2__abc_52138_new_n4167_), .Y(u2__abc_52138_new_n4168_));
NAND2X1 NAND2X1_7 ( .A(aNan), .B(\a[6] ), .Y(_abc_65734_new_n849_));
NAND2X1 NAND2X1_70 ( .A(aNan), .B(\a[69] ), .Y(_abc_65734_new_n1038_));
NAND2X1 NAND2X1_700 ( .A(u2_remHi_228_), .B(u2__abc_52138_new_n4169_), .Y(u2__abc_52138_new_n4170_));
NAND2X1 NAND2X1_701 ( .A(u2_o_228_), .B(u2__abc_52138_new_n4171_), .Y(u2__abc_52138_new_n4172_));
NAND2X1 NAND2X1_702 ( .A(u2__abc_52138_new_n4170_), .B(u2__abc_52138_new_n4172_), .Y(u2__abc_52138_new_n4173_));
NAND2X1 NAND2X1_703 ( .A(u2_remHi_229_), .B(u2__abc_52138_new_n4174_), .Y(u2__abc_52138_new_n4175_));
NAND2X1 NAND2X1_704 ( .A(u2_o_229_), .B(u2__abc_52138_new_n4176_), .Y(u2__abc_52138_new_n4177_));
NAND2X1 NAND2X1_705 ( .A(u2__abc_52138_new_n4175_), .B(u2__abc_52138_new_n4177_), .Y(u2__abc_52138_new_n4178_));
NAND2X1 NAND2X1_706 ( .A(u2__abc_52138_new_n4192_), .B(u2__abc_52138_new_n4098_), .Y(u2__abc_52138_new_n4193_));
NAND2X1 NAND2X1_707 ( .A(u2_remHi_216_), .B(u2__abc_52138_new_n4194_), .Y(u2__abc_52138_new_n4195_));
NAND2X1 NAND2X1_708 ( .A(sqrto_216_), .B(u2__abc_52138_new_n4196_), .Y(u2__abc_52138_new_n4197_));
NAND2X1 NAND2X1_709 ( .A(u2__abc_52138_new_n4195_), .B(u2__abc_52138_new_n4197_), .Y(u2__abc_52138_new_n4198_));
NAND2X1 NAND2X1_71 ( .A(aNan), .B(\a[70] ), .Y(_abc_65734_new_n1041_));
NAND2X1 NAND2X1_710 ( .A(u2_remHi_217_), .B(u2__abc_52138_new_n4199_), .Y(u2__abc_52138_new_n4200_));
NAND2X1 NAND2X1_711 ( .A(sqrto_217_), .B(u2__abc_52138_new_n4201_), .Y(u2__abc_52138_new_n4202_));
NAND2X1 NAND2X1_712 ( .A(u2__abc_52138_new_n4200_), .B(u2__abc_52138_new_n4202_), .Y(u2__abc_52138_new_n4203_));
NAND2X1 NAND2X1_713 ( .A(u2_remHi_214_), .B(u2__abc_52138_new_n4205_), .Y(u2__abc_52138_new_n4206_));
NAND2X1 NAND2X1_714 ( .A(sqrto_214_), .B(u2__abc_52138_new_n4207_), .Y(u2__abc_52138_new_n4208_));
NAND2X1 NAND2X1_715 ( .A(u2__abc_52138_new_n4206_), .B(u2__abc_52138_new_n4208_), .Y(u2__abc_52138_new_n4209_));
NAND2X1 NAND2X1_716 ( .A(u2_remHi_215_), .B(u2__abc_52138_new_n4210_), .Y(u2__abc_52138_new_n4211_));
NAND2X1 NAND2X1_717 ( .A(sqrto_215_), .B(u2__abc_52138_new_n4212_), .Y(u2__abc_52138_new_n4213_));
NAND2X1 NAND2X1_718 ( .A(u2__abc_52138_new_n4211_), .B(u2__abc_52138_new_n4213_), .Y(u2__abc_52138_new_n4214_));
NAND2X1 NAND2X1_719 ( .A(u2_remHi_220_), .B(u2__abc_52138_new_n4217_), .Y(u2__abc_52138_new_n4218_));
NAND2X1 NAND2X1_72 ( .A(aNan), .B(\a[71] ), .Y(_abc_65734_new_n1044_));
NAND2X1 NAND2X1_720 ( .A(sqrto_220_), .B(u2__abc_52138_new_n4219_), .Y(u2__abc_52138_new_n4220_));
NAND2X1 NAND2X1_721 ( .A(u2__abc_52138_new_n4218_), .B(u2__abc_52138_new_n4220_), .Y(u2__abc_52138_new_n4221_));
NAND2X1 NAND2X1_722 ( .A(u2_remHi_221_), .B(u2__abc_52138_new_n4222_), .Y(u2__abc_52138_new_n4223_));
NAND2X1 NAND2X1_723 ( .A(sqrto_221_), .B(u2__abc_52138_new_n4224_), .Y(u2__abc_52138_new_n4225_));
NAND2X1 NAND2X1_724 ( .A(u2__abc_52138_new_n4223_), .B(u2__abc_52138_new_n4225_), .Y(u2__abc_52138_new_n4226_));
NAND2X1 NAND2X1_725 ( .A(u2_remHi_218_), .B(u2__abc_52138_new_n4233_), .Y(u2__abc_52138_new_n4234_));
NAND2X1 NAND2X1_726 ( .A(sqrto_218_), .B(u2__abc_52138_new_n4235_), .Y(u2__abc_52138_new_n4236_));
NAND2X1 NAND2X1_727 ( .A(u2__abc_52138_new_n4237_), .B(u2__abc_52138_new_n4232_), .Y(u2__abc_52138_new_n4238_));
NAND2X1 NAND2X1_728 ( .A(u2__abc_52138_new_n4239_), .B(u2__abc_52138_new_n4216_), .Y(u2__abc_52138_new_n4240_));
NAND2X1 NAND2X1_729 ( .A(u2_remHi_208_), .B(u2__abc_52138_new_n4241_), .Y(u2__abc_52138_new_n4242_));
NAND2X1 NAND2X1_73 ( .A(aNan), .B(\a[72] ), .Y(_abc_65734_new_n1047_));
NAND2X1 NAND2X1_730 ( .A(sqrto_208_), .B(u2__abc_52138_new_n4243_), .Y(u2__abc_52138_new_n4244_));
NAND2X1 NAND2X1_731 ( .A(u2__abc_52138_new_n4242_), .B(u2__abc_52138_new_n4244_), .Y(u2__abc_52138_new_n4245_));
NAND2X1 NAND2X1_732 ( .A(u2_remHi_209_), .B(u2__abc_52138_new_n4246_), .Y(u2__abc_52138_new_n4247_));
NAND2X1 NAND2X1_733 ( .A(sqrto_209_), .B(u2__abc_52138_new_n4248_), .Y(u2__abc_52138_new_n4249_));
NAND2X1 NAND2X1_734 ( .A(u2__abc_52138_new_n4247_), .B(u2__abc_52138_new_n4249_), .Y(u2__abc_52138_new_n4250_));
NAND2X1 NAND2X1_735 ( .A(u2_remHi_206_), .B(u2__abc_52138_new_n4252_), .Y(u2__abc_52138_new_n4253_));
NAND2X1 NAND2X1_736 ( .A(sqrto_206_), .B(u2__abc_52138_new_n4254_), .Y(u2__abc_52138_new_n4255_));
NAND2X1 NAND2X1_737 ( .A(u2__abc_52138_new_n4253_), .B(u2__abc_52138_new_n4255_), .Y(u2__abc_52138_new_n4256_));
NAND2X1 NAND2X1_738 ( .A(u2_remHi_207_), .B(u2__abc_52138_new_n4257_), .Y(u2__abc_52138_new_n4258_));
NAND2X1 NAND2X1_739 ( .A(sqrto_207_), .B(u2__abc_52138_new_n4259_), .Y(u2__abc_52138_new_n4260_));
NAND2X1 NAND2X1_74 ( .A(aNan), .B(\a[73] ), .Y(_abc_65734_new_n1050_));
NAND2X1 NAND2X1_740 ( .A(u2__abc_52138_new_n4258_), .B(u2__abc_52138_new_n4260_), .Y(u2__abc_52138_new_n4261_));
NAND2X1 NAND2X1_741 ( .A(u2__abc_52138_new_n4268_), .B(u2__abc_52138_new_n4273_), .Y(u2__abc_52138_new_n4274_));
NAND2X1 NAND2X1_742 ( .A(u2__abc_52138_new_n4279_), .B(u2__abc_52138_new_n4284_), .Y(u2__abc_52138_new_n4285_));
NAND2X1 NAND2X1_743 ( .A(u2__abc_52138_new_n4286_), .B(u2__abc_52138_new_n4263_), .Y(u2__abc_52138_new_n4287_));
NAND2X1 NAND2X1_744 ( .A(u2_remHi_200_), .B(u2__abc_52138_new_n4289_), .Y(u2__abc_52138_new_n4290_));
NAND2X1 NAND2X1_745 ( .A(sqrto_200_), .B(u2__abc_52138_new_n4291_), .Y(u2__abc_52138_new_n4292_));
NAND2X1 NAND2X1_746 ( .A(u2__abc_52138_new_n4290_), .B(u2__abc_52138_new_n4292_), .Y(u2__abc_52138_new_n4293_));
NAND2X1 NAND2X1_747 ( .A(u2_remHi_201_), .B(u2__abc_52138_new_n4294_), .Y(u2__abc_52138_new_n4295_));
NAND2X1 NAND2X1_748 ( .A(sqrto_201_), .B(u2__abc_52138_new_n4296_), .Y(u2__abc_52138_new_n4297_));
NAND2X1 NAND2X1_749 ( .A(u2__abc_52138_new_n4295_), .B(u2__abc_52138_new_n4297_), .Y(u2__abc_52138_new_n4298_));
NAND2X1 NAND2X1_75 ( .A(aNan), .B(\a[74] ), .Y(_abc_65734_new_n1053_));
NAND2X1 NAND2X1_750 ( .A(u2_remHi_199_), .B(u2__abc_52138_new_n4300_), .Y(u2__abc_52138_new_n4301_));
NAND2X1 NAND2X1_751 ( .A(sqrto_199_), .B(u2__abc_52138_new_n4302_), .Y(u2__abc_52138_new_n4303_));
NAND2X1 NAND2X1_752 ( .A(u2__abc_52138_new_n4301_), .B(u2__abc_52138_new_n4303_), .Y(u2__abc_52138_new_n4304_));
NAND2X1 NAND2X1_753 ( .A(u2_remHi_198_), .B(u2__abc_52138_new_n4305_), .Y(u2__abc_52138_new_n4306_));
NAND2X1 NAND2X1_754 ( .A(sqrto_198_), .B(u2__abc_52138_new_n4307_), .Y(u2__abc_52138_new_n4308_));
NAND2X1 NAND2X1_755 ( .A(u2__abc_52138_new_n4306_), .B(u2__abc_52138_new_n4308_), .Y(u2__abc_52138_new_n4309_));
NAND2X1 NAND2X1_756 ( .A(u2__abc_52138_new_n4299_), .B(u2__abc_52138_new_n4310_), .Y(u2__abc_52138_new_n4311_));
NAND2X1 NAND2X1_757 ( .A(u2_remHi_204_), .B(u2__abc_52138_new_n4312_), .Y(u2__abc_52138_new_n4313_));
NAND2X1 NAND2X1_758 ( .A(sqrto_204_), .B(u2__abc_52138_new_n4314_), .Y(u2__abc_52138_new_n4315_));
NAND2X1 NAND2X1_759 ( .A(u2__abc_52138_new_n4313_), .B(u2__abc_52138_new_n4315_), .Y(u2__abc_52138_new_n4316_));
NAND2X1 NAND2X1_76 ( .A(aNan), .B(\a[75] ), .Y(_abc_65734_new_n1056_));
NAND2X1 NAND2X1_760 ( .A(u2_remHi_205_), .B(u2__abc_52138_new_n4317_), .Y(u2__abc_52138_new_n4318_));
NAND2X1 NAND2X1_761 ( .A(sqrto_205_), .B(u2__abc_52138_new_n4319_), .Y(u2__abc_52138_new_n4320_));
NAND2X1 NAND2X1_762 ( .A(u2__abc_52138_new_n4318_), .B(u2__abc_52138_new_n4320_), .Y(u2__abc_52138_new_n4321_));
NAND2X1 NAND2X1_763 ( .A(u2_remHi_196_), .B(u2__abc_52138_new_n4331_), .Y(u2__abc_52138_new_n4332_));
NAND2X1 NAND2X1_764 ( .A(sqrto_196_), .B(u2__abc_52138_new_n4333_), .Y(u2__abc_52138_new_n4334_));
NAND2X1 NAND2X1_765 ( .A(u2__abc_52138_new_n4332_), .B(u2__abc_52138_new_n4334_), .Y(u2__abc_52138_new_n4335_));
NAND2X1 NAND2X1_766 ( .A(u2_remHi_197_), .B(u2__abc_52138_new_n4336_), .Y(u2__abc_52138_new_n4337_));
NAND2X1 NAND2X1_767 ( .A(sqrto_197_), .B(u2__abc_52138_new_n4338_), .Y(u2__abc_52138_new_n4339_));
NAND2X1 NAND2X1_768 ( .A(u2__abc_52138_new_n4337_), .B(u2__abc_52138_new_n4339_), .Y(u2__abc_52138_new_n4340_));
NAND2X1 NAND2X1_769 ( .A(u2_remHi_195_), .B(u2__abc_52138_new_n4342_), .Y(u2__abc_52138_new_n4343_));
NAND2X1 NAND2X1_77 ( .A(aNan), .B(\a[76] ), .Y(_abc_65734_new_n1059_));
NAND2X1 NAND2X1_770 ( .A(sqrto_195_), .B(u2__abc_52138_new_n4344_), .Y(u2__abc_52138_new_n4345_));
NAND2X1 NAND2X1_771 ( .A(u2__abc_52138_new_n4343_), .B(u2__abc_52138_new_n4345_), .Y(u2__abc_52138_new_n4346_));
NAND2X1 NAND2X1_772 ( .A(u2_remHi_194_), .B(u2__abc_52138_new_n4347_), .Y(u2__abc_52138_new_n4348_));
NAND2X1 NAND2X1_773 ( .A(sqrto_194_), .B(u2__abc_52138_new_n4349_), .Y(u2__abc_52138_new_n4350_));
NAND2X1 NAND2X1_774 ( .A(u2__abc_52138_new_n4348_), .B(u2__abc_52138_new_n4350_), .Y(u2__abc_52138_new_n4351_));
NAND2X1 NAND2X1_775 ( .A(u2_remHi_193_), .B(u2__abc_52138_new_n4358_), .Y(u2__abc_52138_new_n4359_));
NAND2X1 NAND2X1_776 ( .A(sqrto_193_), .B(u2__abc_52138_new_n4360_), .Y(u2__abc_52138_new_n4361_));
NAND2X1 NAND2X1_777 ( .A(u2__abc_52138_new_n4359_), .B(u2__abc_52138_new_n4361_), .Y(u2__abc_52138_new_n4362_));
NAND2X1 NAND2X1_778 ( .A(u2__abc_52138_new_n4371_), .B(u2__abc_52138_new_n4374_), .Y(u2__abc_52138_new_n4375_));
NAND2X1 NAND2X1_779 ( .A(u2__abc_52138_new_n4353_), .B(u2__abc_52138_new_n4377_), .Y(u2__abc_52138_new_n4378_));
NAND2X1 NAND2X1_78 ( .A(aNan), .B(\a[77] ), .Y(_abc_65734_new_n1062_));
NAND2X1 NAND2X1_780 ( .A(u2__abc_52138_new_n4288_), .B(u2__abc_52138_new_n4379_), .Y(u2__abc_52138_new_n4380_));
NAND2X1 NAND2X1_781 ( .A(u2_remHi_182_), .B(u2__abc_52138_new_n4382_), .Y(u2__abc_52138_new_n4383_));
NAND2X1 NAND2X1_782 ( .A(sqrto_182_), .B(u2__abc_52138_new_n4384_), .Y(u2__abc_52138_new_n4385_));
NAND2X1 NAND2X1_783 ( .A(u2__abc_52138_new_n4383_), .B(u2__abc_52138_new_n4385_), .Y(u2__abc_52138_new_n4386_));
NAND2X1 NAND2X1_784 ( .A(u2_remHi_183_), .B(u2__abc_52138_new_n4387_), .Y(u2__abc_52138_new_n4388_));
NAND2X1 NAND2X1_785 ( .A(sqrto_183_), .B(u2__abc_52138_new_n4389_), .Y(u2__abc_52138_new_n4390_));
NAND2X1 NAND2X1_786 ( .A(u2__abc_52138_new_n4388_), .B(u2__abc_52138_new_n4390_), .Y(u2__abc_52138_new_n4391_));
NAND2X1 NAND2X1_787 ( .A(u2_remHi_184_), .B(u2__abc_52138_new_n4393_), .Y(u2__abc_52138_new_n4394_));
NAND2X1 NAND2X1_788 ( .A(sqrto_184_), .B(u2__abc_52138_new_n4395_), .Y(u2__abc_52138_new_n4396_));
NAND2X1 NAND2X1_789 ( .A(u2__abc_52138_new_n4394_), .B(u2__abc_52138_new_n4396_), .Y(u2__abc_52138_new_n4397_));
NAND2X1 NAND2X1_79 ( .A(aNan), .B(\a[78] ), .Y(_abc_65734_new_n1065_));
NAND2X1 NAND2X1_790 ( .A(u2_remHi_185_), .B(u2__abc_52138_new_n4398_), .Y(u2__abc_52138_new_n4399_));
NAND2X1 NAND2X1_791 ( .A(sqrto_185_), .B(u2__abc_52138_new_n4400_), .Y(u2__abc_52138_new_n4401_));
NAND2X1 NAND2X1_792 ( .A(u2__abc_52138_new_n4399_), .B(u2__abc_52138_new_n4401_), .Y(u2__abc_52138_new_n4402_));
NAND2X1 NAND2X1_793 ( .A(u2__abc_52138_new_n4392_), .B(u2__abc_52138_new_n4403_), .Y(u2__abc_52138_new_n4404_));
NAND2X1 NAND2X1_794 ( .A(u2_remHi_188_), .B(u2__abc_52138_new_n4405_), .Y(u2__abc_52138_new_n4406_));
NAND2X1 NAND2X1_795 ( .A(sqrto_188_), .B(u2__abc_52138_new_n4407_), .Y(u2__abc_52138_new_n4408_));
NAND2X1 NAND2X1_796 ( .A(u2__abc_52138_new_n4406_), .B(u2__abc_52138_new_n4408_), .Y(u2__abc_52138_new_n4409_));
NAND2X1 NAND2X1_797 ( .A(u2_remHi_189_), .B(u2__abc_52138_new_n4410_), .Y(u2__abc_52138_new_n4411_));
NAND2X1 NAND2X1_798 ( .A(sqrto_189_), .B(u2__abc_52138_new_n4412_), .Y(u2__abc_52138_new_n4413_));
NAND2X1 NAND2X1_799 ( .A(u2__abc_52138_new_n4411_), .B(u2__abc_52138_new_n4413_), .Y(u2__abc_52138_new_n4414_));
NAND2X1 NAND2X1_8 ( .A(aNan), .B(\a[7] ), .Y(_abc_65734_new_n852_));
NAND2X1 NAND2X1_80 ( .A(aNan), .B(\a[79] ), .Y(_abc_65734_new_n1068_));
NAND2X1 NAND2X1_800 ( .A(u2_remHi_187_), .B(u2__abc_52138_new_n4416_), .Y(u2__abc_52138_new_n4417_));
NAND2X1 NAND2X1_801 ( .A(sqrto_187_), .B(u2__abc_52138_new_n4418_), .Y(u2__abc_52138_new_n4419_));
NAND2X1 NAND2X1_802 ( .A(u2__abc_52138_new_n4417_), .B(u2__abc_52138_new_n4419_), .Y(u2__abc_52138_new_n4420_));
NAND2X1 NAND2X1_803 ( .A(u2_remHi_186_), .B(u2__abc_52138_new_n4421_), .Y(u2__abc_52138_new_n4422_));
NAND2X1 NAND2X1_804 ( .A(sqrto_186_), .B(u2__abc_52138_new_n4423_), .Y(u2__abc_52138_new_n4424_));
NAND2X1 NAND2X1_805 ( .A(u2__abc_52138_new_n4422_), .B(u2__abc_52138_new_n4424_), .Y(u2__abc_52138_new_n4425_));
NAND2X1 NAND2X1_806 ( .A(u2__abc_52138_new_n4415_), .B(u2__abc_52138_new_n4426_), .Y(u2__abc_52138_new_n4427_));
NAND2X1 NAND2X1_807 ( .A(u2_remHi_180_), .B(u2__abc_52138_new_n4429_), .Y(u2__abc_52138_new_n4430_));
NAND2X1 NAND2X1_808 ( .A(sqrto_180_), .B(u2__abc_52138_new_n4431_), .Y(u2__abc_52138_new_n4432_));
NAND2X1 NAND2X1_809 ( .A(u2__abc_52138_new_n4430_), .B(u2__abc_52138_new_n4432_), .Y(u2__abc_52138_new_n4433_));
NAND2X1 NAND2X1_81 ( .A(aNan), .B(\a[80] ), .Y(_abc_65734_new_n1071_));
NAND2X1 NAND2X1_810 ( .A(u2_remHi_181_), .B(u2__abc_52138_new_n4434_), .Y(u2__abc_52138_new_n4435_));
NAND2X1 NAND2X1_811 ( .A(sqrto_181_), .B(u2__abc_52138_new_n4436_), .Y(u2__abc_52138_new_n4437_));
NAND2X1 NAND2X1_812 ( .A(u2__abc_52138_new_n4435_), .B(u2__abc_52138_new_n4437_), .Y(u2__abc_52138_new_n4438_));
NAND2X1 NAND2X1_813 ( .A(u2_remHi_179_), .B(u2__abc_52138_new_n4440_), .Y(u2__abc_52138_new_n4441_));
NAND2X1 NAND2X1_814 ( .A(sqrto_179_), .B(u2__abc_52138_new_n4442_), .Y(u2__abc_52138_new_n4443_));
NAND2X1 NAND2X1_815 ( .A(u2__abc_52138_new_n4441_), .B(u2__abc_52138_new_n4443_), .Y(u2__abc_52138_new_n4444_));
NAND2X1 NAND2X1_816 ( .A(u2_remHi_178_), .B(u2__abc_52138_new_n4445_), .Y(u2__abc_52138_new_n4446_));
NAND2X1 NAND2X1_817 ( .A(sqrto_178_), .B(u2__abc_52138_new_n4447_), .Y(u2__abc_52138_new_n4448_));
NAND2X1 NAND2X1_818 ( .A(u2__abc_52138_new_n4446_), .B(u2__abc_52138_new_n4448_), .Y(u2__abc_52138_new_n4449_));
NAND2X1 NAND2X1_819 ( .A(u2__abc_52138_new_n4439_), .B(u2__abc_52138_new_n4450_), .Y(u2__abc_52138_new_n4451_));
NAND2X1 NAND2X1_82 ( .A(aNan), .B(\a[81] ), .Y(_abc_65734_new_n1074_));
NAND2X1 NAND2X1_820 ( .A(u2_remHi_176_), .B(u2__abc_52138_new_n4452_), .Y(u2__abc_52138_new_n4453_));
NAND2X1 NAND2X1_821 ( .A(sqrto_176_), .B(u2__abc_52138_new_n4454_), .Y(u2__abc_52138_new_n4455_));
NAND2X1 NAND2X1_822 ( .A(u2__abc_52138_new_n4453_), .B(u2__abc_52138_new_n4455_), .Y(u2__abc_52138_new_n4456_));
NAND2X1 NAND2X1_823 ( .A(u2_remHi_177_), .B(u2__abc_52138_new_n4457_), .Y(u2__abc_52138_new_n4458_));
NAND2X1 NAND2X1_824 ( .A(sqrto_177_), .B(u2__abc_52138_new_n4459_), .Y(u2__abc_52138_new_n4460_));
NAND2X1 NAND2X1_825 ( .A(u2__abc_52138_new_n4458_), .B(u2__abc_52138_new_n4460_), .Y(u2__abc_52138_new_n4461_));
NAND2X1 NAND2X1_826 ( .A(u2_remHi_174_), .B(u2__abc_52138_new_n4463_), .Y(u2__abc_52138_new_n4464_));
NAND2X1 NAND2X1_827 ( .A(sqrto_174_), .B(u2__abc_52138_new_n4465_), .Y(u2__abc_52138_new_n4466_));
NAND2X1 NAND2X1_828 ( .A(u2__abc_52138_new_n4464_), .B(u2__abc_52138_new_n4466_), .Y(u2__abc_52138_new_n4467_));
NAND2X1 NAND2X1_829 ( .A(u2_remHi_175_), .B(u2__abc_52138_new_n4469_), .Y(u2__abc_52138_new_n4470_));
NAND2X1 NAND2X1_83 ( .A(aNan), .B(\a[82] ), .Y(_abc_65734_new_n1077_));
NAND2X1 NAND2X1_830 ( .A(sqrto_175_), .B(u2__abc_52138_new_n4471_), .Y(u2__abc_52138_new_n4472_));
NAND2X1 NAND2X1_831 ( .A(u2__abc_52138_new_n4470_), .B(u2__abc_52138_new_n4472_), .Y(u2__abc_52138_new_n4473_));
NAND2X1 NAND2X1_832 ( .A(u2__abc_52138_new_n4428_), .B(u2__abc_52138_new_n4476_), .Y(u2__abc_52138_new_n4477_));
NAND2X1 NAND2X1_833 ( .A(u2_remHi_172_), .B(u2__abc_52138_new_n4478_), .Y(u2__abc_52138_new_n4479_));
NAND2X1 NAND2X1_834 ( .A(sqrto_172_), .B(u2__abc_52138_new_n4480_), .Y(u2__abc_52138_new_n4481_));
NAND2X1 NAND2X1_835 ( .A(u2__abc_52138_new_n4479_), .B(u2__abc_52138_new_n4481_), .Y(u2__abc_52138_new_n4482_));
NAND2X1 NAND2X1_836 ( .A(u2_remHi_173_), .B(u2__abc_52138_new_n4483_), .Y(u2__abc_52138_new_n4484_));
NAND2X1 NAND2X1_837 ( .A(sqrto_173_), .B(u2__abc_52138_new_n4485_), .Y(u2__abc_52138_new_n4486_));
NAND2X1 NAND2X1_838 ( .A(u2__abc_52138_new_n4484_), .B(u2__abc_52138_new_n4486_), .Y(u2__abc_52138_new_n4487_));
NAND2X1 NAND2X1_839 ( .A(u2_remHi_171_), .B(u2__abc_52138_new_n4489_), .Y(u2__abc_52138_new_n4490_));
NAND2X1 NAND2X1_84 ( .A(aNan), .B(\a[83] ), .Y(_abc_65734_new_n1080_));
NAND2X1 NAND2X1_840 ( .A(sqrto_171_), .B(u2__abc_52138_new_n4491_), .Y(u2__abc_52138_new_n4492_));
NAND2X1 NAND2X1_841 ( .A(u2__abc_52138_new_n4490_), .B(u2__abc_52138_new_n4492_), .Y(u2__abc_52138_new_n4493_));
NAND2X1 NAND2X1_842 ( .A(u2_remHi_170_), .B(u2__abc_52138_new_n4494_), .Y(u2__abc_52138_new_n4495_));
NAND2X1 NAND2X1_843 ( .A(sqrto_170_), .B(u2__abc_52138_new_n4496_), .Y(u2__abc_52138_new_n4497_));
NAND2X1 NAND2X1_844 ( .A(u2__abc_52138_new_n4495_), .B(u2__abc_52138_new_n4497_), .Y(u2__abc_52138_new_n4498_));
NAND2X1 NAND2X1_845 ( .A(u2__abc_52138_new_n4488_), .B(u2__abc_52138_new_n4499_), .Y(u2__abc_52138_new_n4500_));
NAND2X1 NAND2X1_846 ( .A(u2_remHi_168_), .B(u2__abc_52138_new_n4501_), .Y(u2__abc_52138_new_n4502_));
NAND2X1 NAND2X1_847 ( .A(sqrto_168_), .B(u2__abc_52138_new_n4503_), .Y(u2__abc_52138_new_n4504_));
NAND2X1 NAND2X1_848 ( .A(u2__abc_52138_new_n4502_), .B(u2__abc_52138_new_n4504_), .Y(u2__abc_52138_new_n4505_));
NAND2X1 NAND2X1_849 ( .A(u2_remHi_169_), .B(u2__abc_52138_new_n4506_), .Y(u2__abc_52138_new_n4507_));
NAND2X1 NAND2X1_85 ( .A(aNan), .B(\a[84] ), .Y(_abc_65734_new_n1083_));
NAND2X1 NAND2X1_850 ( .A(sqrto_169_), .B(u2__abc_52138_new_n4508_), .Y(u2__abc_52138_new_n4509_));
NAND2X1 NAND2X1_851 ( .A(u2__abc_52138_new_n4507_), .B(u2__abc_52138_new_n4509_), .Y(u2__abc_52138_new_n4510_));
NAND2X1 NAND2X1_852 ( .A(u2_remHi_167_), .B(u2__abc_52138_new_n4512_), .Y(u2__abc_52138_new_n4513_));
NAND2X1 NAND2X1_853 ( .A(sqrto_167_), .B(u2__abc_52138_new_n4514_), .Y(u2__abc_52138_new_n4515_));
NAND2X1 NAND2X1_854 ( .A(u2__abc_52138_new_n4513_), .B(u2__abc_52138_new_n4515_), .Y(u2__abc_52138_new_n4516_));
NAND2X1 NAND2X1_855 ( .A(u2__abc_52138_new_n4511_), .B(u2__abc_52138_new_n4522_), .Y(u2__abc_52138_new_n4523_));
NAND2X1 NAND2X1_856 ( .A(u2_remHi_160_), .B(u2__abc_52138_new_n4525_), .Y(u2__abc_52138_new_n4526_));
NAND2X1 NAND2X1_857 ( .A(sqrto_160_), .B(u2__abc_52138_new_n4527_), .Y(u2__abc_52138_new_n4528_));
NAND2X1 NAND2X1_858 ( .A(u2__abc_52138_new_n4526_), .B(u2__abc_52138_new_n4528_), .Y(u2__abc_52138_new_n4529_));
NAND2X1 NAND2X1_859 ( .A(u2_remHi_161_), .B(u2__abc_52138_new_n4530_), .Y(u2__abc_52138_new_n4531_));
NAND2X1 NAND2X1_86 ( .A(aNan), .B(\a[85] ), .Y(_abc_65734_new_n1086_));
NAND2X1 NAND2X1_860 ( .A(sqrto_161_), .B(u2__abc_52138_new_n4532_), .Y(u2__abc_52138_new_n4533_));
NAND2X1 NAND2X1_861 ( .A(u2__abc_52138_new_n4531_), .B(u2__abc_52138_new_n4533_), .Y(u2__abc_52138_new_n4534_));
NAND2X1 NAND2X1_862 ( .A(u2_remHi_159_), .B(u2__abc_52138_new_n4536_), .Y(u2__abc_52138_new_n4537_));
NAND2X1 NAND2X1_863 ( .A(u2__abc_52138_new_n4537_), .B(u2__abc_52138_new_n4539_), .Y(u2__abc_52138_new_n4540_));
NAND2X1 NAND2X1_864 ( .A(u2_remHi_164_), .B(u2__abc_52138_new_n4548_), .Y(u2__abc_52138_new_n4549_));
NAND2X1 NAND2X1_865 ( .A(sqrto_164_), .B(u2__abc_52138_new_n4550_), .Y(u2__abc_52138_new_n4551_));
NAND2X1 NAND2X1_866 ( .A(u2__abc_52138_new_n4549_), .B(u2__abc_52138_new_n4551_), .Y(u2__abc_52138_new_n4552_));
NAND2X1 NAND2X1_867 ( .A(u2_remHi_165_), .B(u2__abc_52138_new_n4553_), .Y(u2__abc_52138_new_n4554_));
NAND2X1 NAND2X1_868 ( .A(sqrto_165_), .B(u2__abc_52138_new_n4555_), .Y(u2__abc_52138_new_n4556_));
NAND2X1 NAND2X1_869 ( .A(u2__abc_52138_new_n4554_), .B(u2__abc_52138_new_n4556_), .Y(u2__abc_52138_new_n4557_));
NAND2X1 NAND2X1_87 ( .A(aNan), .B(\a[86] ), .Y(_abc_65734_new_n1089_));
NAND2X1 NAND2X1_870 ( .A(u2_remHi_163_), .B(u2__abc_52138_new_n4559_), .Y(u2__abc_52138_new_n4560_));
NAND2X1 NAND2X1_871 ( .A(sqrto_163_), .B(u2__abc_52138_new_n4561_), .Y(u2__abc_52138_new_n4562_));
NAND2X1 NAND2X1_872 ( .A(u2__abc_52138_new_n4560_), .B(u2__abc_52138_new_n4562_), .Y(u2__abc_52138_new_n4563_));
NAND2X1 NAND2X1_873 ( .A(u2_remHi_162_), .B(u2__abc_52138_new_n4564_), .Y(u2__abc_52138_new_n4565_));
NAND2X1 NAND2X1_874 ( .A(sqrto_162_), .B(u2__abc_52138_new_n4566_), .Y(u2__abc_52138_new_n4567_));
NAND2X1 NAND2X1_875 ( .A(u2__abc_52138_new_n4565_), .B(u2__abc_52138_new_n4567_), .Y(u2__abc_52138_new_n4568_));
NAND2X1 NAND2X1_876 ( .A(u2_remHi_152_), .B(u2__abc_52138_new_n4573_), .Y(u2__abc_52138_new_n4574_));
NAND2X1 NAND2X1_877 ( .A(sqrto_152_), .B(u2__abc_52138_new_n4575_), .Y(u2__abc_52138_new_n4576_));
NAND2X1 NAND2X1_878 ( .A(u2__abc_52138_new_n4574_), .B(u2__abc_52138_new_n4576_), .Y(u2__abc_52138_new_n4577_));
NAND2X1 NAND2X1_879 ( .A(u2_remHi_153_), .B(u2__abc_52138_new_n4578_), .Y(u2__abc_52138_new_n4579_));
NAND2X1 NAND2X1_88 ( .A(aNan), .B(\a[87] ), .Y(_abc_65734_new_n1092_));
NAND2X1 NAND2X1_880 ( .A(sqrto_153_), .B(u2__abc_52138_new_n4580_), .Y(u2__abc_52138_new_n4581_));
NAND2X1 NAND2X1_881 ( .A(u2__abc_52138_new_n4579_), .B(u2__abc_52138_new_n4581_), .Y(u2__abc_52138_new_n4582_));
NAND2X1 NAND2X1_882 ( .A(u2_remHi_151_), .B(u2__abc_52138_new_n4584_), .Y(u2__abc_52138_new_n4585_));
NAND2X1 NAND2X1_883 ( .A(sqrto_151_), .B(u2__abc_52138_new_n4586_), .Y(u2__abc_52138_new_n4587_));
NAND2X1 NAND2X1_884 ( .A(u2__abc_52138_new_n4585_), .B(u2__abc_52138_new_n4587_), .Y(u2__abc_52138_new_n4588_));
NAND2X1 NAND2X1_885 ( .A(u2_remHi_150_), .B(u2__abc_52138_new_n4589_), .Y(u2__abc_52138_new_n4590_));
NAND2X1 NAND2X1_886 ( .A(sqrto_150_), .B(u2__abc_52138_new_n4591_), .Y(u2__abc_52138_new_n4592_));
NAND2X1 NAND2X1_887 ( .A(u2__abc_52138_new_n4590_), .B(u2__abc_52138_new_n4592_), .Y(u2__abc_52138_new_n4593_));
NAND2X1 NAND2X1_888 ( .A(u2__abc_52138_new_n4583_), .B(u2__abc_52138_new_n4594_), .Y(u2__abc_52138_new_n4595_));
NAND2X1 NAND2X1_889 ( .A(u2_remHi_156_), .B(u2__abc_52138_new_n4596_), .Y(u2__abc_52138_new_n4597_));
NAND2X1 NAND2X1_89 ( .A(aNan), .B(\a[88] ), .Y(_abc_65734_new_n1095_));
NAND2X1 NAND2X1_890 ( .A(sqrto_156_), .B(u2__abc_52138_new_n4598_), .Y(u2__abc_52138_new_n4599_));
NAND2X1 NAND2X1_891 ( .A(u2__abc_52138_new_n4597_), .B(u2__abc_52138_new_n4599_), .Y(u2__abc_52138_new_n4600_));
NAND2X1 NAND2X1_892 ( .A(u2_remHi_157_), .B(u2__abc_52138_new_n4601_), .Y(u2__abc_52138_new_n4602_));
NAND2X1 NAND2X1_893 ( .A(sqrto_157_), .B(u2__abc_52138_new_n4603_), .Y(u2__abc_52138_new_n4604_));
NAND2X1 NAND2X1_894 ( .A(u2__abc_52138_new_n4602_), .B(u2__abc_52138_new_n4604_), .Y(u2__abc_52138_new_n4605_));
NAND2X1 NAND2X1_895 ( .A(u2_remHi_148_), .B(u2__abc_52138_new_n4619_), .Y(u2__abc_52138_new_n4620_));
NAND2X1 NAND2X1_896 ( .A(sqrto_148_), .B(u2__abc_52138_new_n4621_), .Y(u2__abc_52138_new_n4622_));
NAND2X1 NAND2X1_897 ( .A(u2__abc_52138_new_n4620_), .B(u2__abc_52138_new_n4622_), .Y(u2__abc_52138_new_n4623_));
NAND2X1 NAND2X1_898 ( .A(u2_remHi_149_), .B(u2__abc_52138_new_n4624_), .Y(u2__abc_52138_new_n4625_));
NAND2X1 NAND2X1_899 ( .A(sqrto_149_), .B(u2__abc_52138_new_n4626_), .Y(u2__abc_52138_new_n4627_));
NAND2X1 NAND2X1_9 ( .A(aNan), .B(\a[8] ), .Y(_abc_65734_new_n855_));
NAND2X1 NAND2X1_90 ( .A(aNan), .B(\a[89] ), .Y(_abc_65734_new_n1098_));
NAND2X1 NAND2X1_900 ( .A(u2__abc_52138_new_n4625_), .B(u2__abc_52138_new_n4627_), .Y(u2__abc_52138_new_n4628_));
NAND2X1 NAND2X1_901 ( .A(u2_remHi_147_), .B(u2__abc_52138_new_n4630_), .Y(u2__abc_52138_new_n4631_));
NAND2X1 NAND2X1_902 ( .A(sqrto_147_), .B(u2__abc_52138_new_n4632_), .Y(u2__abc_52138_new_n4633_));
NAND2X1 NAND2X1_903 ( .A(u2__abc_52138_new_n4631_), .B(u2__abc_52138_new_n4633_), .Y(u2__abc_52138_new_n4634_));
NAND2X1 NAND2X1_904 ( .A(u2_remHi_146_), .B(u2__abc_52138_new_n4635_), .Y(u2__abc_52138_new_n4636_));
NAND2X1 NAND2X1_905 ( .A(sqrto_146_), .B(u2__abc_52138_new_n4637_), .Y(u2__abc_52138_new_n4638_));
NAND2X1 NAND2X1_906 ( .A(u2__abc_52138_new_n4636_), .B(u2__abc_52138_new_n4638_), .Y(u2__abc_52138_new_n4639_));
NAND2X1 NAND2X1_907 ( .A(u2_remHi_144_), .B(u2__abc_52138_new_n4642_), .Y(u2__abc_52138_new_n4643_));
NAND2X1 NAND2X1_908 ( .A(sqrto_144_), .B(u2__abc_52138_new_n4644_), .Y(u2__abc_52138_new_n4645_));
NAND2X1 NAND2X1_909 ( .A(u2_remHi_145_), .B(u2__abc_52138_new_n4647_), .Y(u2__abc_52138_new_n4648_));
NAND2X1 NAND2X1_91 ( .A(aNan), .B(\a[90] ), .Y(_abc_65734_new_n1101_));
NAND2X1 NAND2X1_910 ( .A(sqrto_145_), .B(u2__abc_52138_new_n4649_), .Y(u2__abc_52138_new_n4650_));
NAND2X1 NAND2X1_911 ( .A(u2_remHi_136_), .B(u2__abc_52138_new_n4666_), .Y(u2__abc_52138_new_n4667_));
NAND2X1 NAND2X1_912 ( .A(sqrto_136_), .B(u2__abc_52138_new_n4668_), .Y(u2__abc_52138_new_n4669_));
NAND2X1 NAND2X1_913 ( .A(u2__abc_52138_new_n4667_), .B(u2__abc_52138_new_n4669_), .Y(u2__abc_52138_new_n4670_));
NAND2X1 NAND2X1_914 ( .A(u2_remHi_137_), .B(u2__abc_52138_new_n4671_), .Y(u2__abc_52138_new_n4672_));
NAND2X1 NAND2X1_915 ( .A(sqrto_137_), .B(u2__abc_52138_new_n4673_), .Y(u2__abc_52138_new_n4674_));
NAND2X1 NAND2X1_916 ( .A(u2__abc_52138_new_n4672_), .B(u2__abc_52138_new_n4674_), .Y(u2__abc_52138_new_n4675_));
NAND2X1 NAND2X1_917 ( .A(u2_remHi_134_), .B(u2__abc_52138_new_n4677_), .Y(u2__abc_52138_new_n4678_));
NAND2X1 NAND2X1_918 ( .A(sqrto_134_), .B(u2__abc_52138_new_n4679_), .Y(u2__abc_52138_new_n4680_));
NAND2X1 NAND2X1_919 ( .A(u2__abc_52138_new_n4678_), .B(u2__abc_52138_new_n4680_), .Y(u2__abc_52138_new_n4681_));
NAND2X1 NAND2X1_92 ( .A(aNan), .B(\a[91] ), .Y(_abc_65734_new_n1104_));
NAND2X1 NAND2X1_920 ( .A(u2_remHi_135_), .B(u2__abc_52138_new_n4682_), .Y(u2__abc_52138_new_n4683_));
NAND2X1 NAND2X1_921 ( .A(sqrto_135_), .B(u2__abc_52138_new_n4684_), .Y(u2__abc_52138_new_n4685_));
NAND2X1 NAND2X1_922 ( .A(u2__abc_52138_new_n4683_), .B(u2__abc_52138_new_n4685_), .Y(u2__abc_52138_new_n4686_));
NAND2X1 NAND2X1_923 ( .A(u2_remHi_140_), .B(u2__abc_52138_new_n4689_), .Y(u2__abc_52138_new_n4690_));
NAND2X1 NAND2X1_924 ( .A(sqrto_140_), .B(u2__abc_52138_new_n4691_), .Y(u2__abc_52138_new_n4692_));
NAND2X1 NAND2X1_925 ( .A(u2__abc_52138_new_n4690_), .B(u2__abc_52138_new_n4692_), .Y(u2__abc_52138_new_n4693_));
NAND2X1 NAND2X1_926 ( .A(u2_remHi_141_), .B(u2__abc_52138_new_n4694_), .Y(u2__abc_52138_new_n4695_));
NAND2X1 NAND2X1_927 ( .A(sqrto_141_), .B(u2__abc_52138_new_n4696_), .Y(u2__abc_52138_new_n4697_));
NAND2X1 NAND2X1_928 ( .A(u2__abc_52138_new_n4695_), .B(u2__abc_52138_new_n4697_), .Y(u2__abc_52138_new_n4698_));
NAND2X1 NAND2X1_929 ( .A(u2_remHi_139_), .B(u2__abc_52138_new_n4700_), .Y(u2__abc_52138_new_n4701_));
NAND2X1 NAND2X1_93 ( .A(aNan), .B(\a[92] ), .Y(_abc_65734_new_n1107_));
NAND2X1 NAND2X1_930 ( .A(sqrto_139_), .B(u2__abc_52138_new_n4702_), .Y(u2__abc_52138_new_n4703_));
NAND2X1 NAND2X1_931 ( .A(u2__abc_52138_new_n4701_), .B(u2__abc_52138_new_n4703_), .Y(u2__abc_52138_new_n4704_));
NAND2X1 NAND2X1_932 ( .A(u2_remHi_138_), .B(u2__abc_52138_new_n4705_), .Y(u2__abc_52138_new_n4706_));
NAND2X1 NAND2X1_933 ( .A(sqrto_138_), .B(u2__abc_52138_new_n4707_), .Y(u2__abc_52138_new_n4708_));
NAND2X1 NAND2X1_934 ( .A(u2__abc_52138_new_n4706_), .B(u2__abc_52138_new_n4708_), .Y(u2__abc_52138_new_n4709_));
NAND2X1 NAND2X1_935 ( .A(u2__abc_52138_new_n4688_), .B(u2__abc_52138_new_n4711_), .Y(u2__abc_52138_new_n4712_));
NAND2X1 NAND2X1_936 ( .A(u2_remHi_126_), .B(u2__abc_52138_new_n4713_), .Y(u2__abc_52138_new_n4714_));
NAND2X1 NAND2X1_937 ( .A(sqrto_126_), .B(u2__abc_52138_new_n4715_), .Y(u2__abc_52138_new_n4716_));
NAND2X1 NAND2X1_938 ( .A(u2__abc_52138_new_n4714_), .B(u2__abc_52138_new_n4716_), .Y(u2__abc_52138_new_n4717_));
NAND2X1 NAND2X1_939 ( .A(u2_remHi_127_), .B(u2__abc_52138_new_n4719_), .Y(u2__abc_52138_new_n4720_));
NAND2X1 NAND2X1_94 ( .A(aNan), .B(\a[93] ), .Y(_abc_65734_new_n1110_));
NAND2X1 NAND2X1_940 ( .A(sqrto_127_), .B(u2__abc_52138_new_n4721_), .Y(u2__abc_52138_new_n4722_));
NAND2X1 NAND2X1_941 ( .A(u2__abc_52138_new_n4720_), .B(u2__abc_52138_new_n4722_), .Y(u2__abc_52138_new_n4723_));
NAND2X1 NAND2X1_942 ( .A(u2__abc_52138_new_n4718_), .B(u2__abc_52138_new_n4724_), .Y(u2__abc_52138_new_n4725_));
NAND2X1 NAND2X1_943 ( .A(u2_remHi_129_), .B(u2__abc_52138_new_n4727_), .Y(u2__abc_52138_new_n4728_));
NAND2X1 NAND2X1_944 ( .A(sqrto_129_), .B(u2__abc_52138_new_n4729_), .Y(u2__abc_52138_new_n4730_));
NAND2X1 NAND2X1_945 ( .A(u2_remHi_132_), .B(u2__abc_52138_new_n4733_), .Y(u2__abc_52138_new_n4734_));
NAND2X1 NAND2X1_946 ( .A(sqrto_132_), .B(u2__abc_52138_new_n4735_), .Y(u2__abc_52138_new_n4736_));
NAND2X1 NAND2X1_947 ( .A(u2__abc_52138_new_n4734_), .B(u2__abc_52138_new_n4736_), .Y(u2__abc_52138_new_n4737_));
NAND2X1 NAND2X1_948 ( .A(u2_remHi_133_), .B(u2__abc_52138_new_n4738_), .Y(u2__abc_52138_new_n4739_));
NAND2X1 NAND2X1_949 ( .A(sqrto_133_), .B(u2__abc_52138_new_n4740_), .Y(u2__abc_52138_new_n4741_));
NAND2X1 NAND2X1_95 ( .A(aNan), .B(\a[94] ), .Y(_abc_65734_new_n1113_));
NAND2X1 NAND2X1_950 ( .A(u2__abc_52138_new_n4739_), .B(u2__abc_52138_new_n4741_), .Y(u2__abc_52138_new_n4742_));
NAND2X1 NAND2X1_951 ( .A(u2_remHi_131_), .B(u2__abc_52138_new_n4744_), .Y(u2__abc_52138_new_n4745_));
NAND2X1 NAND2X1_952 ( .A(sqrto_131_), .B(u2__abc_52138_new_n4746_), .Y(u2__abc_52138_new_n4747_));
NAND2X1 NAND2X1_953 ( .A(u2__abc_52138_new_n4570_), .B(u2__abc_52138_new_n4547_), .Y(u2__abc_52138_new_n4757_));
NAND2X1 NAND2X1_954 ( .A(u2__abc_52138_new_n4754_), .B(u2__abc_52138_new_n4758_), .Y(u2__abc_52138_new_n4759_));
NAND2X1 NAND2X1_955 ( .A(u2__abc_52138_new_n4641_), .B(u2__abc_52138_new_n4664_), .Y(u2__abc_52138_new_n4761_));
NAND2X1 NAND2X1_956 ( .A(u2__abc_52138_new_n4749_), .B(u2__abc_52138_new_n4748_), .Y(u2__abc_52138_new_n4765_));
NAND2X1 NAND2X1_957 ( .A(sqrto_130_), .B(u2__abc_52138_new_n4776_), .Y(u2__abc_52138_new_n4777_));
NAND2X1 NAND2X1_958 ( .A(u2__abc_52138_new_n4794_), .B(u2__abc_52138_new_n4699_), .Y(u2__abc_52138_new_n4795_));
NAND2X1 NAND2X1_959 ( .A(u2__abc_52138_new_n4797_), .B(u2__abc_52138_new_n4795_), .Y(u2__abc_52138_new_n4798_));
NAND2X1 NAND2X1_96 ( .A(aNan), .B(\a[95] ), .Y(_abc_65734_new_n1116_));
NAND2X1 NAND2X1_960 ( .A(u2__abc_52138_new_n4817_), .B(u2__abc_52138_new_n4583_), .Y(u2__abc_52138_new_n4818_));
NAND2X1 NAND2X1_961 ( .A(u2__abc_52138_new_n4820_), .B(u2__abc_52138_new_n4818_), .Y(u2__abc_52138_new_n4821_));
NAND2X1 NAND2X1_962 ( .A(u2__abc_52138_new_n4606_), .B(u2__abc_52138_new_n4823_), .Y(u2__abc_52138_new_n4824_));
NAND2X1 NAND2X1_963 ( .A(u2__abc_52138_new_n4826_), .B(u2__abc_52138_new_n4824_), .Y(u2__abc_52138_new_n4827_));
NAND2X1 NAND2X1_964 ( .A(u2__abc_52138_new_n4511_), .B(u2__abc_52138_new_n4846_), .Y(u2__abc_52138_new_n4847_));
NAND2X1 NAND2X1_965 ( .A(u2__abc_52138_new_n4849_), .B(u2__abc_52138_new_n4847_), .Y(u2__abc_52138_new_n4850_));
NAND2X1 NAND2X1_966 ( .A(u2__abc_52138_new_n4488_), .B(u2__abc_52138_new_n4851_), .Y(u2__abc_52138_new_n4852_));
NAND2X1 NAND2X1_967 ( .A(u2__abc_52138_new_n4428_), .B(u2__abc_52138_new_n4866_), .Y(u2__abc_52138_new_n4867_));
NAND2X1 NAND2X1_968 ( .A(u2__abc_52138_new_n4876_), .B(u2__abc_52138_new_n4867_), .Y(u2__abc_52138_new_n4877_));
NAND2X1 NAND2X1_969 ( .A(u2__abc_52138_new_n4880_), .B(u2__abc_52138_new_n4883_), .Y(u2__abc_52138_new_n4884_));
NAND2X1 NAND2X1_97 ( .A(aNan), .B(\a[96] ), .Y(_abc_65734_new_n1119_));
NAND2X1 NAND2X1_970 ( .A(u2__abc_52138_new_n4899_), .B(u2__abc_52138_new_n4299_), .Y(u2__abc_52138_new_n4900_));
NAND2X1 NAND2X1_971 ( .A(u2__abc_52138_new_n4902_), .B(u2__abc_52138_new_n4900_), .Y(u2__abc_52138_new_n4903_));
NAND2X1 NAND2X1_972 ( .A(sqrto_202_), .B(u2__abc_52138_new_n4905_), .Y(u2__abc_52138_new_n4906_));
NAND2X1 NAND2X1_973 ( .A(u2__abc_52138_new_n4907_), .B(u2__abc_52138_new_n4322_), .Y(u2__abc_52138_new_n4908_));
NAND2X1 NAND2X1_974 ( .A(u2__abc_52138_new_n4928_), .B(u2__abc_52138_new_n4929_), .Y(u2__abc_52138_new_n4930_));
NAND2X1 NAND2X1_975 ( .A(u2__abc_52138_new_n4932_), .B(u2__abc_52138_new_n4930_), .Y(u2__abc_52138_new_n4933_));
NAND2X1 NAND2X1_976 ( .A(u2__abc_52138_new_n4946_), .B(u2__abc_52138_new_n4156_), .Y(u2__abc_52138_new_n4947_));
NAND2X1 NAND2X1_977 ( .A(u2__abc_52138_new_n4949_), .B(u2__abc_52138_new_n4947_), .Y(u2__abc_52138_new_n4950_));
NAND2X1 NAND2X1_978 ( .A(u2__abc_52138_new_n4179_), .B(u2__abc_52138_new_n4952_), .Y(u2__abc_52138_new_n4953_));
NAND2X1 NAND2X1_979 ( .A(u2__abc_52138_new_n4956_), .B(u2__abc_52138_new_n4953_), .Y(u2__abc_52138_new_n4957_));
NAND2X1 NAND2X1_98 ( .A(aNan), .B(\a[97] ), .Y(_abc_65734_new_n1122_));
NAND2X1 NAND2X1_980 ( .A(u2__abc_52138_new_n4024_), .B(u2__abc_52138_new_n4972_), .Y(u2__abc_52138_new_n4973_));
NAND2X1 NAND2X1_981 ( .A(u2__abc_52138_new_n4975_), .B(u2__abc_52138_new_n4973_), .Y(u2__abc_52138_new_n4976_));
NAND2X1 NAND2X1_982 ( .A(u2__abc_52138_new_n4084_), .B(u2__abc_52138_new_n4095_), .Y(u2__abc_52138_new_n4983_));
NAND2X1 NAND2X1_983 ( .A(u2__abc_52138_new_n4982_), .B(u2__abc_52138_new_n4992_), .Y(u2__abc_52138_new_n4993_));
NAND2X1 NAND2X1_984 ( .A(u2__abc_52138_new_n4981_), .B(u2__abc_52138_new_n4993_), .Y(u2__abc_52138_new_n4994_));
NAND2X1 NAND2X1_985 ( .A(u2__abc_52138_new_n5003_), .B(u2__abc_52138_new_n5008_), .Y(u2__abc_52138_new_n5009_));
NAND2X1 NAND2X1_986 ( .A(u2__abc_52138_new_n5010_), .B(u2__abc_52138_new_n5015_), .Y(u2__abc_52138_new_n5016_));
NAND2X1 NAND2X1_987 ( .A(u2_o_375_), .B(u2__abc_52138_new_n5023_), .Y(u2__abc_52138_new_n5024_));
NAND2X1 NAND2X1_988 ( .A(u2_remHi_375_), .B(u2__abc_52138_new_n5025_), .Y(u2__abc_52138_new_n5026_));
NAND2X1 NAND2X1_989 ( .A(u2__abc_52138_new_n5024_), .B(u2__abc_52138_new_n5026_), .Y(u2__abc_52138_new_n5027_));
NAND2X1 NAND2X1_99 ( .A(aNan), .B(\a[98] ), .Y(_abc_65734_new_n1125_));
NAND2X1 NAND2X1_990 ( .A(u2__abc_52138_new_n5022_), .B(u2__abc_52138_new_n5028_), .Y(u2__abc_52138_new_n5029_));
NAND2X1 NAND2X1_991 ( .A(u2__abc_52138_new_n5037_), .B(u2__abc_52138_new_n5040_), .Y(u2__abc_52138_new_n5041_));
NAND2X1 NAND2X1_992 ( .A(u2__abc_52138_new_n5017_), .B(u2__abc_52138_new_n5043_), .Y(u2__abc_52138_new_n5044_));
NAND2X1 NAND2X1_993 ( .A(u2__abc_52138_new_n5050_), .B(u2__abc_52138_new_n5049_), .Y(u2__abc_52138_new_n5051_));
NAND2X1 NAND2X1_994 ( .A(u2_o_366_), .B(u2__abc_52138_new_n5052_), .Y(u2__abc_52138_new_n5055_));
NAND2X1 NAND2X1_995 ( .A(u2_remHi_367_), .B(u2__abc_52138_new_n5057_), .Y(u2__abc_52138_new_n5058_));
NAND2X1 NAND2X1_996 ( .A(u2_o_367_), .B(u2__abc_52138_new_n5059_), .Y(u2__abc_52138_new_n5060_));
NAND2X1 NAND2X1_997 ( .A(u2__abc_52138_new_n5058_), .B(u2__abc_52138_new_n5060_), .Y(u2__abc_52138_new_n5061_));
NAND2X1 NAND2X1_998 ( .A(u2__abc_52138_new_n5062_), .B(u2__abc_52138_new_n5056_), .Y(u2__abc_52138_new_n5063_));
NAND2X1 NAND2X1_999 ( .A(u2__abc_52138_new_n5069_), .B(u2__abc_52138_new_n5074_), .Y(u2__abc_52138_new_n5075_));
NAND3X1 NAND3X1_1 ( .A(_abc_65734_new_n1458_), .B(_abc_65734_new_n1463_), .C(_abc_65734_new_n1453_), .Y(_abc_65734_new_n1464_));
NAND3X1 NAND3X1_10 ( .A(_abc_65734_new_n1533_), .B(_abc_65734_new_n1535_), .C(_abc_65734_new_n1524_), .Y(_abc_65734_new_n1536_));
NAND3X1 NAND3X1_100 ( .A(u2__abc_52138_new_n6785_), .B(u2__abc_52138_new_n6786_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6787_));
NAND3X1 NAND3X1_101 ( .A(u2__abc_52138_new_n6807_), .B(u2__abc_52138_new_n6809_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6810_));
NAND3X1 NAND3X1_102 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n6865_), .C(u2__abc_52138_new_n6864_), .Y(u2__abc_52138_new_n6866_));
NAND3X1 NAND3X1_103 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n6907_), .C(u2__abc_52138_new_n6908_), .Y(u2__abc_52138_new_n6909_));
NAND3X1 NAND3X1_104 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n6972_), .C(u2__abc_52138_new_n6973_), .Y(u2__abc_52138_new_n6974_));
NAND3X1 NAND3X1_105 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n7033_), .C(u2__abc_52138_new_n7036_), .Y(u2__abc_52138_new_n7037_));
NAND3X1 NAND3X1_106 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n7057_), .C(u2__abc_52138_new_n7058_), .Y(u2__abc_52138_new_n7059_));
NAND3X1 NAND3X1_107 ( .A(u2__abc_52138_new_n3312_), .B(u2__abc_52138_new_n3314_), .C(u2__abc_52138_new_n7076_), .Y(u2__abc_52138_new_n7084_));
NAND3X1 NAND3X1_108 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n7101_), .C(u2__abc_52138_new_n7102_), .Y(u2__abc_52138_new_n7103_));
NAND3X1 NAND3X1_109 ( .A(u2__abc_52138_new_n3241_), .B(u2__abc_52138_new_n3243_), .C(u2__abc_52138_new_n7118_), .Y(u2__abc_52138_new_n7126_));
NAND3X1 NAND3X1_11 ( .A(_abc_65734_new_n1529_), .B(_abc_65734_new_n1540_), .C(_abc_65734_new_n1515_), .Y(_abc_65734_new_n1544_));
NAND3X1 NAND3X1_110 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n7187_), .C(u2__abc_52138_new_n7188_), .Y(u2__abc_52138_new_n7189_));
NAND3X1 NAND3X1_111 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n7273_), .C(u2__abc_52138_new_n7272_), .Y(u2__abc_52138_new_n7274_));
NAND3X1 NAND3X1_112 ( .A(u2__abc_52138_new_n3790_), .B(u2__abc_52138_new_n3795_), .C(u2__abc_52138_new_n7309_), .Y(u2__abc_52138_new_n7310_));
NAND3X1 NAND3X1_113 ( .A(u2__abc_52138_new_n3823_), .B(u2__abc_52138_new_n3828_), .C(u2__abc_52138_new_n7354_), .Y(u2__abc_52138_new_n7355_));
NAND3X1 NAND3X1_114 ( .A(u2__abc_52138_new_n7532_), .B(u2__abc_52138_new_n7538_), .C(u2__abc_52138_new_n7531_), .Y(u2__abc_52138_new_n7539_));
NAND3X1 NAND3X1_115 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n7544_), .C(u2__abc_52138_new_n7542_), .Y(u2__abc_52138_new_n7545_));
NAND3X1 NAND3X1_116 ( .A(u2__abc_52138_new_n7684_), .B(u2__abc_52138_new_n3638_), .C(u2__abc_52138_new_n3962_), .Y(u2__abc_52138_new_n7714_));
NAND3X1 NAND3X1_117 ( .A(u2__abc_52138_new_n7805_), .B(u2__abc_52138_new_n7807_), .C(u2__abc_52138_new_n7801_), .Y(u2__abc_52138_new_n7808_));
NAND3X1 NAND3X1_118 ( .A(u2__abc_52138_new_n6499_), .B(u2__abc_52138_new_n7900_), .C(u2__abc_52138_new_n7902_), .Y(u2__abc_52138_new_n7903_));
NAND3X1 NAND3X1_119 ( .A(u2__abc_52138_new_n8688_), .B(u2__abc_52138_new_n8689_), .C(u2__abc_52138_new_n8686_), .Y(u2__abc_52138_new_n8690_));
NAND3X1 NAND3X1_12 ( .A(\a[119] ), .B(_abc_65734_new_n1535_), .C(_abc_65734_new_n1511_), .Y(_abc_65734_new_n1546_));
NAND3X1 NAND3X1_120 ( .A(u2__abc_52138_new_n4242_), .B(u2__abc_52138_new_n4244_), .C(u2__abc_52138_new_n8794_), .Y(u2__abc_52138_new_n8802_));
NAND3X1 NAND3X1_121 ( .A(u2__abc_52138_new_n8937_), .B(u2__abc_52138_new_n8941_), .C(u2__abc_52138_new_n8936_), .Y(u2__abc_52138_new_n8942_));
NAND3X1 NAND3X1_122 ( .A(u2__abc_52138_new_n4288_), .B(u2__abc_52138_new_n4379_), .C(u2__abc_52138_new_n9267_), .Y(u2__abc_52138_new_n9268_));
NAND3X1 NAND3X1_123 ( .A(u2__abc_52138_new_n9593_), .B(u2__abc_52138_new_n9594_), .C(u2__abc_52138_new_n5774_), .Y(u2__abc_52138_new_n9614_));
NAND3X1 NAND3X1_124 ( .A(u2__abc_52138_new_n9767_), .B(u2__abc_52138_new_n9768_), .C(u2__abc_52138_new_n5801_), .Y(u2__abc_52138_new_n9789_));
NAND3X1 NAND3X1_125 ( .A(u2__abc_52138_new_n9789_), .B(u2__abc_52138_new_n9790_), .C(u2__abc_52138_new_n9788_), .Y(u2__abc_52138_new_n9791_));
NAND3X1 NAND3X1_126 ( .A(u2__abc_52138_new_n9958_), .B(u2__abc_52138_new_n9964_), .C(u2__abc_52138_new_n9957_), .Y(u2__abc_52138_new_n9965_));
NAND3X1 NAND3X1_127 ( .A(u2__abc_52138_new_n10111_), .B(u2__abc_52138_new_n10112_), .C(u2__abc_52138_new_n5854_), .Y(u2__abc_52138_new_n10132_));
NAND3X1 NAND3X1_128 ( .A(u2__abc_52138_new_n10132_), .B(u2__abc_52138_new_n10133_), .C(u2__abc_52138_new_n10134_), .Y(u2__abc_52138_new_n10135_));
NAND3X1 NAND3X1_129 ( .A(u2__abc_52138_new_n10461_), .B(u2__abc_52138_new_n5912_), .C(u2__abc_52138_new_n5909_), .Y(u2__abc_52138_new_n10480_));
NAND3X1 NAND3X1_13 ( .A(\a[122] ), .B(\a[123] ), .C(_abc_65734_new_n1548_), .Y(_abc_65734_new_n1549_));
NAND3X1 NAND3X1_130 ( .A(u2__abc_52138_new_n10658_), .B(u2__abc_52138_new_n10650_), .C(u2__abc_52138_new_n10649_), .Y(u2__abc_52138_new_n10659_));
NAND3X1 NAND3X1_131 ( .A(u2__abc_52138_new_n6346_), .B(u2__abc_52138_new_n10811_), .C(u2__abc_52138_new_n6345_), .Y(u2__abc_52138_new_n10830_));
NAND3X1 NAND3X1_132 ( .A(u2__abc_52138_new_n10830_), .B(u2__abc_52138_new_n10831_), .C(u2__abc_52138_new_n10832_), .Y(u2__abc_52138_new_n10833_));
NAND3X1 NAND3X1_133 ( .A(u2__abc_52138_new_n6365_), .B(u2__abc_52138_new_n10983_), .C(u2__abc_52138_new_n6364_), .Y(u2__abc_52138_new_n11003_));
NAND3X1 NAND3X1_134 ( .A(u2_remLo_0_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11418_));
NAND3X1 NAND3X1_135 ( .A(u2_remLo_1_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11421_));
NAND3X1 NAND3X1_136 ( .A(u2_remLo_2_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11424_));
NAND3X1 NAND3X1_137 ( .A(u2_remLo_3_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11427_));
NAND3X1 NAND3X1_138 ( .A(u2_remLo_4_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11430_));
NAND3X1 NAND3X1_139 ( .A(u2_remLo_5_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11433_));
NAND3X1 NAND3X1_14 ( .A(_abc_65734_new_n1550_), .B(_abc_65734_new_n1556_), .C(_abc_65734_new_n1539_), .Y(_abc_65734_new_n1557_));
NAND3X1 NAND3X1_140 ( .A(u2_remLo_6_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11436_));
NAND3X1 NAND3X1_141 ( .A(u2_remLo_7_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11439_));
NAND3X1 NAND3X1_142 ( .A(u2_remLo_8_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11442_));
NAND3X1 NAND3X1_143 ( .A(u2_remLo_9_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11445_));
NAND3X1 NAND3X1_144 ( .A(u2_remLo_10_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11448_));
NAND3X1 NAND3X1_145 ( .A(u2_remLo_11_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11451_));
NAND3X1 NAND3X1_146 ( .A(u2_remLo_12_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11454_));
NAND3X1 NAND3X1_147 ( .A(u2_remLo_13_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11457_));
NAND3X1 NAND3X1_148 ( .A(u2_remLo_14_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11460_));
NAND3X1 NAND3X1_149 ( .A(u2_remLo_15_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11463_));
NAND3X1 NAND3X1_15 ( .A(\a[124] ), .B(\a[125] ), .C(_abc_65734_new_n1565_), .Y(_abc_65734_new_n1566_));
NAND3X1 NAND3X1_150 ( .A(u2_remLo_16_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11466_));
NAND3X1 NAND3X1_151 ( .A(u2_remLo_17_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11469_));
NAND3X1 NAND3X1_152 ( .A(u2_remLo_18_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11472_));
NAND3X1 NAND3X1_153 ( .A(u2_remLo_19_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11475_));
NAND3X1 NAND3X1_154 ( .A(u2_remLo_20_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11478_));
NAND3X1 NAND3X1_155 ( .A(u2_remLo_21_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11481_));
NAND3X1 NAND3X1_156 ( .A(u2_remLo_22_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11484_));
NAND3X1 NAND3X1_157 ( .A(u2_remLo_23_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11487_));
NAND3X1 NAND3X1_158 ( .A(u2_remLo_24_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11490_));
NAND3X1 NAND3X1_159 ( .A(u2_remLo_25_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11493_));
NAND3X1 NAND3X1_16 ( .A(_abc_65734_new_n1567_), .B(_abc_65734_new_n1575_), .C(_abc_65734_new_n1574_), .Y(_abc_65734_new_n1576_));
NAND3X1 NAND3X1_160 ( .A(u2_remLo_26_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11496_));
NAND3X1 NAND3X1_161 ( .A(u2_remLo_27_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11499_));
NAND3X1 NAND3X1_162 ( .A(u2_remLo_28_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11502_));
NAND3X1 NAND3X1_163 ( .A(u2_remLo_29_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n11505_));
NAND3X1 NAND3X1_164 ( .A(u2_remLo_256_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12235_));
NAND3X1 NAND3X1_165 ( .A(u2_remLo_257_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12238_));
NAND3X1 NAND3X1_166 ( .A(u2_remLo_258_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12241_));
NAND3X1 NAND3X1_167 ( .A(u2_remLo_259_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12244_));
NAND3X1 NAND3X1_168 ( .A(u2_remLo_260_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12247_));
NAND3X1 NAND3X1_169 ( .A(u2_remLo_261_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12250_));
NAND3X1 NAND3X1_17 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1573_), .C(_abc_65734_new_n1576_), .Y(_abc_65734_new_n1577_));
NAND3X1 NAND3X1_170 ( .A(u2_remLo_262_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12253_));
NAND3X1 NAND3X1_171 ( .A(u2_remLo_263_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12256_));
NAND3X1 NAND3X1_172 ( .A(u2_remLo_264_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12259_));
NAND3X1 NAND3X1_173 ( .A(u2_remLo_265_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12262_));
NAND3X1 NAND3X1_174 ( .A(u2_remLo_266_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12265_));
NAND3X1 NAND3X1_175 ( .A(u2_remLo_267_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12268_));
NAND3X1 NAND3X1_176 ( .A(u2_remLo_268_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12271_));
NAND3X1 NAND3X1_177 ( .A(u2_remLo_269_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12274_));
NAND3X1 NAND3X1_178 ( .A(u2_remLo_270_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12277_));
NAND3X1 NAND3X1_179 ( .A(u2_remLo_271_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12280_));
NAND3X1 NAND3X1_18 ( .A(\a[123] ), .B(\a[124] ), .C(_abc_65734_new_n1581_), .Y(_abc_65734_new_n1582_));
NAND3X1 NAND3X1_180 ( .A(u2_remLo_272_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12283_));
NAND3X1 NAND3X1_181 ( .A(u2_remLo_273_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12286_));
NAND3X1 NAND3X1_182 ( .A(u2_remLo_274_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12289_));
NAND3X1 NAND3X1_183 ( .A(u2_remLo_275_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12292_));
NAND3X1 NAND3X1_184 ( .A(u2_remLo_276_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12295_));
NAND3X1 NAND3X1_185 ( .A(u2_remLo_277_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12298_));
NAND3X1 NAND3X1_186 ( .A(u2_remLo_278_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12301_));
NAND3X1 NAND3X1_187 ( .A(u2_remLo_279_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12304_));
NAND3X1 NAND3X1_188 ( .A(u2_remLo_280_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12307_));
NAND3X1 NAND3X1_189 ( .A(u2_remLo_281_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12310_));
NAND3X1 NAND3X1_19 ( .A(\a[112] ), .B(u1__abc_51895_new_n160_), .C(u1__abc_51895_new_n163_), .Y(u1__abc_51895_new_n164_));
NAND3X1 NAND3X1_190 ( .A(u2_remLo_282_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12313_));
NAND3X1 NAND3X1_191 ( .A(u2_remLo_283_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12316_));
NAND3X1 NAND3X1_192 ( .A(u2_remLo_284_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12319_));
NAND3X1 NAND3X1_193 ( .A(u2_remLo_285_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12322_));
NAND3X1 NAND3X1_194 ( .A(u2_remLo_286_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12325_));
NAND3X1 NAND3X1_195 ( .A(u2_remLo_287_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12328_));
NAND3X1 NAND3X1_196 ( .A(u2_remLo_288_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12331_));
NAND3X1 NAND3X1_197 ( .A(u2_remLo_289_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12334_));
NAND3X1 NAND3X1_198 ( .A(u2_remLo_290_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12337_));
NAND3X1 NAND3X1_199 ( .A(u2_remLo_291_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12340_));
NAND3X1 NAND3X1_2 ( .A(\a[116] ), .B(_abc_65734_new_n1452_), .C(_abc_65734_new_n1470_), .Y(_abc_65734_new_n1472_));
NAND3X1 NAND3X1_20 ( .A(u2__abc_52138_new_n3018_), .B(u2__abc_52138_new_n3020_), .C(u2__abc_52138_new_n3016_), .Y(u2__abc_52138_new_n3021_));
NAND3X1 NAND3X1_200 ( .A(u2_remLo_292_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12343_));
NAND3X1 NAND3X1_201 ( .A(u2_remLo_293_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12346_));
NAND3X1 NAND3X1_202 ( .A(u2_remLo_294_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12349_));
NAND3X1 NAND3X1_203 ( .A(u2_remLo_295_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12352_));
NAND3X1 NAND3X1_204 ( .A(u2_remLo_296_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12355_));
NAND3X1 NAND3X1_205 ( .A(u2_remLo_297_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12358_));
NAND3X1 NAND3X1_206 ( .A(u2_remLo_298_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12361_));
NAND3X1 NAND3X1_207 ( .A(u2_remLo_299_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12364_));
NAND3X1 NAND3X1_208 ( .A(u2_remLo_300_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12367_));
NAND3X1 NAND3X1_209 ( .A(u2_remLo_301_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12370_));
NAND3X1 NAND3X1_21 ( .A(u2__abc_52138_new_n3036_), .B(u2__abc_52138_new_n3038_), .C(u2__abc_52138_new_n3034_), .Y(u2__abc_52138_new_n3039_));
NAND3X1 NAND3X1_210 ( .A(u2_remLo_302_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12373_));
NAND3X1 NAND3X1_211 ( .A(u2_remLo_303_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12376_));
NAND3X1 NAND3X1_212 ( .A(u2_remLo_304_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12379_));
NAND3X1 NAND3X1_213 ( .A(u2_remLo_305_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12382_));
NAND3X1 NAND3X1_214 ( .A(u2_remLo_306_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12385_));
NAND3X1 NAND3X1_215 ( .A(u2_remLo_307_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12388_));
NAND3X1 NAND3X1_216 ( .A(u2_remLo_308_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12391_));
NAND3X1 NAND3X1_217 ( .A(u2_remLo_309_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12394_));
NAND3X1 NAND3X1_218 ( .A(u2_remLo_310_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12397_));
NAND3X1 NAND3X1_219 ( .A(u2_remLo_311_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12400_));
NAND3X1 NAND3X1_22 ( .A(u2__abc_52138_new_n3055_), .B(u2__abc_52138_new_n3057_), .C(u2__abc_52138_new_n3053_), .Y(u2__abc_52138_new_n3058_));
NAND3X1 NAND3X1_220 ( .A(u2_remLo_312_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12403_));
NAND3X1 NAND3X1_221 ( .A(u2_remLo_313_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12406_));
NAND3X1 NAND3X1_222 ( .A(u2_remLo_314_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12409_));
NAND3X1 NAND3X1_223 ( .A(u2_remLo_315_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12412_));
NAND3X1 NAND3X1_224 ( .A(u2_remLo_316_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12415_));
NAND3X1 NAND3X1_225 ( .A(u2_remLo_317_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12418_));
NAND3X1 NAND3X1_226 ( .A(u2_remLo_318_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12421_));
NAND3X1 NAND3X1_227 ( .A(u2_remLo_319_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12424_));
NAND3X1 NAND3X1_228 ( .A(u2_remLo_320_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12427_));
NAND3X1 NAND3X1_229 ( .A(u2_remLo_321_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12430_));
NAND3X1 NAND3X1_23 ( .A(u2__abc_52138_new_n3061_), .B(u2__abc_52138_new_n3063_), .C(u2__abc_52138_new_n3059_), .Y(u2__abc_52138_new_n3064_));
NAND3X1 NAND3X1_230 ( .A(u2_remLo_322_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12433_));
NAND3X1 NAND3X1_231 ( .A(u2_remLo_323_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12436_));
NAND3X1 NAND3X1_232 ( .A(u2_remLo_324_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12439_));
NAND3X1 NAND3X1_233 ( .A(u2_remLo_325_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12442_));
NAND3X1 NAND3X1_234 ( .A(u2_remLo_326_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12445_));
NAND3X1 NAND3X1_235 ( .A(u2_remLo_327_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12448_));
NAND3X1 NAND3X1_236 ( .A(u2_remLo_328_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12451_));
NAND3X1 NAND3X1_237 ( .A(u2_remLo_329_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12454_));
NAND3X1 NAND3X1_238 ( .A(u2_remLo_330_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12457_));
NAND3X1 NAND3X1_239 ( .A(u2_remLo_331_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12460_));
NAND3X1 NAND3X1_24 ( .A(u2__abc_52138_new_n3184_), .B(u2__abc_52138_new_n3186_), .C(u2__abc_52138_new_n3182_), .Y(u2__abc_52138_new_n3187_));
NAND3X1 NAND3X1_240 ( .A(u2_remLo_332_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12463_));
NAND3X1 NAND3X1_241 ( .A(u2_remLo_333_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12466_));
NAND3X1 NAND3X1_242 ( .A(u2_remLo_334_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12469_));
NAND3X1 NAND3X1_243 ( .A(u2_remLo_335_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12472_));
NAND3X1 NAND3X1_244 ( .A(u2_remLo_336_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12475_));
NAND3X1 NAND3X1_245 ( .A(u2_remLo_337_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12478_));
NAND3X1 NAND3X1_246 ( .A(u2_remLo_338_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12481_));
NAND3X1 NAND3X1_247 ( .A(u2_remLo_339_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12484_));
NAND3X1 NAND3X1_248 ( .A(u2_remLo_340_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12487_));
NAND3X1 NAND3X1_249 ( .A(u2_remLo_341_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12490_));
NAND3X1 NAND3X1_25 ( .A(u2__abc_52138_new_n3190_), .B(u2__abc_52138_new_n3192_), .C(u2__abc_52138_new_n3188_), .Y(u2__abc_52138_new_n3193_));
NAND3X1 NAND3X1_250 ( .A(u2_remLo_342_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12493_));
NAND3X1 NAND3X1_251 ( .A(u2_remLo_343_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12496_));
NAND3X1 NAND3X1_252 ( .A(u2_remLo_344_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12499_));
NAND3X1 NAND3X1_253 ( .A(u2_remLo_345_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12502_));
NAND3X1 NAND3X1_254 ( .A(u2_remLo_346_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12505_));
NAND3X1 NAND3X1_255 ( .A(u2_remLo_347_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12508_));
NAND3X1 NAND3X1_256 ( .A(u2_remLo_348_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12511_));
NAND3X1 NAND3X1_257 ( .A(u2_remLo_349_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12514_));
NAND3X1 NAND3X1_258 ( .A(u2_remLo_350_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12517_));
NAND3X1 NAND3X1_259 ( .A(u2_remLo_351_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12520_));
NAND3X1 NAND3X1_26 ( .A(u2__abc_52138_new_n3165_), .B(u2__abc_52138_new_n3167_), .C(u2__abc_52138_new_n3197_), .Y(u2__abc_52138_new_n3198_));
NAND3X1 NAND3X1_260 ( .A(u2_remLo_352_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12523_));
NAND3X1 NAND3X1_261 ( .A(u2_remLo_353_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12526_));
NAND3X1 NAND3X1_262 ( .A(u2_remLo_354_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12529_));
NAND3X1 NAND3X1_263 ( .A(u2_remLo_355_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12532_));
NAND3X1 NAND3X1_264 ( .A(u2_remLo_356_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12535_));
NAND3X1 NAND3X1_265 ( .A(u2_remLo_357_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12538_));
NAND3X1 NAND3X1_266 ( .A(u2_remLo_358_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12541_));
NAND3X1 NAND3X1_267 ( .A(u2_remLo_359_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12544_));
NAND3X1 NAND3X1_268 ( .A(u2_remLo_360_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12547_));
NAND3X1 NAND3X1_269 ( .A(u2_remLo_361_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12550_));
NAND3X1 NAND3X1_27 ( .A(u2__abc_52138_new_n3310_), .B(u2__abc_52138_new_n3333_), .C(u2__abc_52138_new_n3286_), .Y(u2__abc_52138_new_n3334_));
NAND3X1 NAND3X1_270 ( .A(u2_remLo_362_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12553_));
NAND3X1 NAND3X1_271 ( .A(u2_remLo_363_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12556_));
NAND3X1 NAND3X1_272 ( .A(u2_remLo_364_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12559_));
NAND3X1 NAND3X1_273 ( .A(u2_remLo_365_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12562_));
NAND3X1 NAND3X1_274 ( .A(u2_remLo_366_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12565_));
NAND3X1 NAND3X1_275 ( .A(u2_remLo_367_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12568_));
NAND3X1 NAND3X1_276 ( .A(u2_remLo_368_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12571_));
NAND3X1 NAND3X1_277 ( .A(u2_remLo_369_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12574_));
NAND3X1 NAND3X1_278 ( .A(u2_remLo_370_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12577_));
NAND3X1 NAND3X1_279 ( .A(u2_remLo_371_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12580_));
NAND3X1 NAND3X1_28 ( .A(u2__abc_52138_new_n3416_), .B(u2__abc_52138_new_n3417_), .C(u2__abc_52138_new_n3411_), .Y(u2__abc_52138_new_n3418_));
NAND3X1 NAND3X1_280 ( .A(u2_remLo_372_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12583_));
NAND3X1 NAND3X1_281 ( .A(u2_remLo_373_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12586_));
NAND3X1 NAND3X1_282 ( .A(u2_remLo_374_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12589_));
NAND3X1 NAND3X1_283 ( .A(u2_remLo_375_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12592_));
NAND3X1 NAND3X1_284 ( .A(u2_remLo_376_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12595_));
NAND3X1 NAND3X1_285 ( .A(u2_remLo_377_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12598_));
NAND3X1 NAND3X1_286 ( .A(u2_remLo_378_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12601_));
NAND3X1 NAND3X1_287 ( .A(u2_remLo_379_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12604_));
NAND3X1 NAND3X1_288 ( .A(u2_remLo_380_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12607_));
NAND3X1 NAND3X1_289 ( .A(u2_remLo_381_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12610_));
NAND3X1 NAND3X1_29 ( .A(u2__abc_52138_new_n3407_), .B(u2__abc_52138_new_n3409_), .C(u2__abc_52138_new_n3428_), .Y(u2__abc_52138_new_n3429_));
NAND3X1 NAND3X1_290 ( .A(u2_remLo_382_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12613_));
NAND3X1 NAND3X1_291 ( .A(u2_remLo_383_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12616_));
NAND3X1 NAND3X1_292 ( .A(u2_remLo_384_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12619_));
NAND3X1 NAND3X1_293 ( .A(u2_remLo_385_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12622_));
NAND3X1 NAND3X1_294 ( .A(u2_remLo_386_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12625_));
NAND3X1 NAND3X1_295 ( .A(u2_remLo_387_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12628_));
NAND3X1 NAND3X1_296 ( .A(u2_remLo_388_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12631_));
NAND3X1 NAND3X1_297 ( .A(u2_remLo_389_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12634_));
NAND3X1 NAND3X1_298 ( .A(u2_remLo_390_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12637_));
NAND3X1 NAND3X1_299 ( .A(u2_remLo_391_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12640_));
NAND3X1 NAND3X1_3 ( .A(\a[117] ), .B(\a[118] ), .C(_abc_65734_new_n1486_), .Y(_abc_65734_new_n1492_));
NAND3X1 NAND3X1_30 ( .A(u2__abc_52138_new_n3384_), .B(u2__abc_52138_new_n3386_), .C(u2__abc_52138_new_n3432_), .Y(u2__abc_52138_new_n3433_));
NAND3X1 NAND3X1_300 ( .A(u2_remLo_392_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12643_));
NAND3X1 NAND3X1_301 ( .A(u2_remLo_393_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12646_));
NAND3X1 NAND3X1_302 ( .A(u2_remLo_394_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12649_));
NAND3X1 NAND3X1_303 ( .A(u2_remLo_395_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12652_));
NAND3X1 NAND3X1_304 ( .A(u2_remLo_396_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12655_));
NAND3X1 NAND3X1_305 ( .A(u2_remLo_397_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12658_));
NAND3X1 NAND3X1_306 ( .A(u2_remLo_398_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12661_));
NAND3X1 NAND3X1_307 ( .A(u2_remLo_399_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12664_));
NAND3X1 NAND3X1_308 ( .A(u2_remLo_400_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12667_));
NAND3X1 NAND3X1_309 ( .A(u2_remLo_401_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12670_));
NAND3X1 NAND3X1_31 ( .A(u2__abc_52138_new_n3269_), .B(u2__abc_52138_new_n3497_), .C(u2__abc_52138_new_n3496_), .Y(u2__abc_52138_new_n3498_));
NAND3X1 NAND3X1_310 ( .A(u2_remLo_402_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12673_));
NAND3X1 NAND3X1_311 ( .A(u2_remLo_403_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12676_));
NAND3X1 NAND3X1_312 ( .A(u2_remLo_404_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12679_));
NAND3X1 NAND3X1_313 ( .A(u2_remLo_405_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12682_));
NAND3X1 NAND3X1_314 ( .A(u2_remLo_406_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12685_));
NAND3X1 NAND3X1_315 ( .A(u2_remLo_407_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12688_));
NAND3X1 NAND3X1_316 ( .A(u2_remLo_408_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12691_));
NAND3X1 NAND3X1_317 ( .A(u2_remLo_409_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12694_));
NAND3X1 NAND3X1_318 ( .A(u2_remLo_410_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12697_));
NAND3X1 NAND3X1_319 ( .A(u2_remLo_411_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12700_));
NAND3X1 NAND3X1_32 ( .A(u2__abc_52138_new_n3539_), .B(u2__abc_52138_new_n3541_), .C(u2__abc_52138_new_n3546_), .Y(u2__abc_52138_new_n3547_));
NAND3X1 NAND3X1_320 ( .A(u2_remLo_412_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12703_));
NAND3X1 NAND3X1_321 ( .A(u2_remLo_413_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12706_));
NAND3X1 NAND3X1_322 ( .A(u2_remLo_414_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12709_));
NAND3X1 NAND3X1_323 ( .A(u2_remLo_415_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12712_));
NAND3X1 NAND3X1_324 ( .A(u2_remLo_416_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12715_));
NAND3X1 NAND3X1_325 ( .A(u2_remLo_417_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12718_));
NAND3X1 NAND3X1_326 ( .A(u2_remLo_418_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12721_));
NAND3X1 NAND3X1_327 ( .A(u2_remLo_419_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12724_));
NAND3X1 NAND3X1_328 ( .A(u2_remLo_420_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12727_));
NAND3X1 NAND3X1_329 ( .A(u2_remLo_421_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12730_));
NAND3X1 NAND3X1_33 ( .A(u2__abc_52138_new_n3515_), .B(u2__abc_52138_new_n3526_), .C(u2__abc_52138_new_n3548_), .Y(u2__abc_52138_new_n3549_));
NAND3X1 NAND3X1_330 ( .A(u2_remLo_422_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12733_));
NAND3X1 NAND3X1_331 ( .A(u2_remLo_423_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12736_));
NAND3X1 NAND3X1_332 ( .A(u2_remLo_424_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12739_));
NAND3X1 NAND3X1_333 ( .A(u2_remLo_425_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12742_));
NAND3X1 NAND3X1_334 ( .A(u2_remLo_426_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12745_));
NAND3X1 NAND3X1_335 ( .A(u2_remLo_427_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12748_));
NAND3X1 NAND3X1_336 ( .A(u2_remLo_428_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12751_));
NAND3X1 NAND3X1_337 ( .A(u2_remLo_429_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12754_));
NAND3X1 NAND3X1_338 ( .A(u2_remLo_430_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12757_));
NAND3X1 NAND3X1_339 ( .A(u2_remLo_431_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12760_));
NAND3X1 NAND3X1_34 ( .A(u2__abc_52138_new_n3579_), .B(u2__abc_52138_new_n3581_), .C(u2__abc_52138_new_n3577_), .Y(u2__abc_52138_new_n3582_));
NAND3X1 NAND3X1_340 ( .A(u2_remLo_432_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12763_));
NAND3X1 NAND3X1_341 ( .A(u2_remLo_433_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12766_));
NAND3X1 NAND3X1_342 ( .A(u2_remLo_434_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12769_));
NAND3X1 NAND3X1_343 ( .A(u2_remLo_435_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12772_));
NAND3X1 NAND3X1_344 ( .A(u2_remLo_436_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12775_));
NAND3X1 NAND3X1_345 ( .A(u2_remLo_437_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12778_));
NAND3X1 NAND3X1_346 ( .A(u2_remLo_438_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12781_));
NAND3X1 NAND3X1_347 ( .A(u2_remLo_439_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12784_));
NAND3X1 NAND3X1_348 ( .A(u2_remLo_440_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12787_));
NAND3X1 NAND3X1_349 ( .A(u2_remLo_441_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12790_));
NAND3X1 NAND3X1_35 ( .A(u2__abc_52138_new_n3609_), .B(u2__abc_52138_new_n3611_), .C(u2__abc_52138_new_n3616_), .Y(u2__abc_52138_new_n3617_));
NAND3X1 NAND3X1_350 ( .A(u2_remLo_442_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12793_));
NAND3X1 NAND3X1_351 ( .A(u2_remLo_443_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12796_));
NAND3X1 NAND3X1_352 ( .A(u2_remLo_444_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12799_));
NAND3X1 NAND3X1_353 ( .A(u2_remLo_445_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12802_));
NAND3X1 NAND3X1_354 ( .A(u2_remLo_446_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12805_));
NAND3X1 NAND3X1_355 ( .A(u2_remLo_447_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12808_));
NAND3X1 NAND3X1_356 ( .A(u2_remLo_448_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12811_));
NAND3X1 NAND3X1_357 ( .A(u2_remLo_449_), .B(u2__abc_52138_new_n6504_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n12814_));
NAND3X1 NAND3X1_358 ( .A(u2__abc_52138_new_n3026_), .B(u2__abc_52138_new_n3031_), .C(u2__abc_52138_new_n6668_), .Y(u2__abc_52138_new_n12819_));
NAND3X1 NAND3X1_359 ( .A(u2__abc_52138_new_n3044_), .B(u2__abc_52138_new_n3049_), .C(u2__abc_52138_new_n12820_), .Y(u2__abc_52138_new_n12821_));
NAND3X1 NAND3X1_36 ( .A(u2__abc_52138_new_n3631_), .B(u2__abc_52138_new_n3633_), .C(u2__abc_52138_new_n3638_), .Y(u2__abc_52138_new_n3639_));
NAND3X1 NAND3X1_360 ( .A(u2__abc_52138_new_n3070_), .B(u2__abc_52138_new_n3066_), .C(u2__abc_52138_new_n3067_), .Y(u2__abc_52138_new_n12823_));
NAND3X1 NAND3X1_361 ( .A(u2__abc_52138_new_n3181_), .B(u2__abc_52138_new_n3194_), .C(u2__abc_52138_new_n12838_), .Y(u2__abc_52138_new_n12839_));
NAND3X1 NAND3X1_362 ( .A(u2__abc_52138_new_n5928_), .B(u2__abc_52138_new_n13036_), .C(u2__abc_52138_new_n13035_), .Y(u2__abc_52138_new_n13037_));
NAND3X1 NAND3X1_363 ( .A(sqrto_2_), .B(sqrto_1_), .C(u2__abc_52138_new_n13051_), .Y(u2__abc_52138_new_n13067_));
NAND3X1 NAND3X1_364 ( .A(sqrto_1_), .B(sqrto_0_), .C(u2__abc_52138_new_n13044_), .Y(u2__abc_52138_new_n13075_));
NAND3X1 NAND3X1_365 ( .A(sqrto_3_), .B(sqrto_2_), .C(u2__abc_52138_new_n13060_), .Y(u2__abc_52138_new_n13090_));
NAND3X1 NAND3X1_366 ( .A(sqrto_6_), .B(sqrto_5_), .C(u2__abc_52138_new_n13083_), .Y(u2__abc_52138_new_n13098_));
NAND3X1 NAND3X1_367 ( .A(sqrto_5_), .B(sqrto_4_), .C(u2__abc_52138_new_n13076_), .Y(u2__abc_52138_new_n13106_));
NAND3X1 NAND3X1_368 ( .A(sqrto_7_), .B(sqrto_6_), .C(u2__abc_52138_new_n13091_), .Y(u2__abc_52138_new_n13121_));
NAND3X1 NAND3X1_369 ( .A(sqrto_10_), .B(sqrto_9_), .C(u2__abc_52138_new_n13114_), .Y(u2__abc_52138_new_n13129_));
NAND3X1 NAND3X1_37 ( .A(u2__abc_52138_new_n3703_), .B(u2__abc_52138_new_n3705_), .C(u2__abc_52138_new_n3710_), .Y(u2__abc_52138_new_n3711_));
NAND3X1 NAND3X1_370 ( .A(sqrto_9_), .B(sqrto_8_), .C(u2__abc_52138_new_n13107_), .Y(u2__abc_52138_new_n13137_));
NAND3X1 NAND3X1_371 ( .A(sqrto_11_), .B(sqrto_10_), .C(u2__abc_52138_new_n13122_), .Y(u2__abc_52138_new_n13152_));
NAND3X1 NAND3X1_372 ( .A(sqrto_14_), .B(sqrto_13_), .C(u2__abc_52138_new_n13145_), .Y(u2__abc_52138_new_n13160_));
NAND3X1 NAND3X1_373 ( .A(sqrto_13_), .B(sqrto_12_), .C(u2__abc_52138_new_n13138_), .Y(u2__abc_52138_new_n13168_));
NAND3X1 NAND3X1_374 ( .A(sqrto_15_), .B(sqrto_14_), .C(u2__abc_52138_new_n13153_), .Y(u2__abc_52138_new_n13183_));
NAND3X1 NAND3X1_375 ( .A(sqrto_18_), .B(sqrto_17_), .C(u2__abc_52138_new_n13176_), .Y(u2__abc_52138_new_n13191_));
NAND3X1 NAND3X1_376 ( .A(sqrto_17_), .B(sqrto_16_), .C(u2__abc_52138_new_n13169_), .Y(u2__abc_52138_new_n13199_));
NAND3X1 NAND3X1_377 ( .A(sqrto_19_), .B(sqrto_18_), .C(u2__abc_52138_new_n13184_), .Y(u2__abc_52138_new_n13214_));
NAND3X1 NAND3X1_378 ( .A(sqrto_22_), .B(sqrto_21_), .C(u2__abc_52138_new_n13207_), .Y(u2__abc_52138_new_n13222_));
NAND3X1 NAND3X1_379 ( .A(sqrto_21_), .B(sqrto_20_), .C(u2__abc_52138_new_n13200_), .Y(u2__abc_52138_new_n13230_));
NAND3X1 NAND3X1_38 ( .A(u2__abc_52138_new_n3726_), .B(u2__abc_52138_new_n3729_), .C(u2__abc_52138_new_n3734_), .Y(u2__abc_52138_new_n3735_));
NAND3X1 NAND3X1_380 ( .A(sqrto_23_), .B(sqrto_22_), .C(u2__abc_52138_new_n13215_), .Y(u2__abc_52138_new_n13245_));
NAND3X1 NAND3X1_381 ( .A(sqrto_26_), .B(sqrto_25_), .C(u2__abc_52138_new_n13238_), .Y(u2__abc_52138_new_n13253_));
NAND3X1 NAND3X1_382 ( .A(sqrto_25_), .B(sqrto_24_), .C(u2__abc_52138_new_n13231_), .Y(u2__abc_52138_new_n13261_));
NAND3X1 NAND3X1_383 ( .A(sqrto_27_), .B(sqrto_26_), .C(u2__abc_52138_new_n13246_), .Y(u2__abc_52138_new_n13276_));
NAND3X1 NAND3X1_384 ( .A(sqrto_30_), .B(sqrto_29_), .C(u2__abc_52138_new_n13269_), .Y(u2__abc_52138_new_n13284_));
NAND3X1 NAND3X1_385 ( .A(sqrto_29_), .B(sqrto_28_), .C(u2__abc_52138_new_n13262_), .Y(u2__abc_52138_new_n13292_));
NAND3X1 NAND3X1_386 ( .A(sqrto_31_), .B(sqrto_30_), .C(u2__abc_52138_new_n13277_), .Y(u2__abc_52138_new_n13307_));
NAND3X1 NAND3X1_387 ( .A(sqrto_34_), .B(sqrto_33_), .C(u2__abc_52138_new_n13300_), .Y(u2__abc_52138_new_n13316_));
NAND3X1 NAND3X1_388 ( .A(sqrto_33_), .B(sqrto_32_), .C(u2__abc_52138_new_n13293_), .Y(u2__abc_52138_new_n13324_));
NAND3X1 NAND3X1_389 ( .A(sqrto_35_), .B(sqrto_34_), .C(u2__abc_52138_new_n13308_), .Y(u2__abc_52138_new_n13339_));
NAND3X1 NAND3X1_39 ( .A(u2__abc_52138_new_n3803_), .B(u2__abc_52138_new_n3805_), .C(u2__abc_52138_new_n3801_), .Y(u2__abc_52138_new_n3806_));
NAND3X1 NAND3X1_390 ( .A(sqrto_38_), .B(sqrto_37_), .C(u2__abc_52138_new_n13332_), .Y(u2__abc_52138_new_n13347_));
NAND3X1 NAND3X1_391 ( .A(sqrto_37_), .B(sqrto_36_), .C(u2__abc_52138_new_n13325_), .Y(u2__abc_52138_new_n13355_));
NAND3X1 NAND3X1_392 ( .A(sqrto_39_), .B(sqrto_38_), .C(u2__abc_52138_new_n13340_), .Y(u2__abc_52138_new_n13370_));
NAND3X1 NAND3X1_393 ( .A(sqrto_42_), .B(sqrto_41_), .C(u2__abc_52138_new_n13363_), .Y(u2__abc_52138_new_n13378_));
NAND3X1 NAND3X1_394 ( .A(sqrto_41_), .B(sqrto_40_), .C(u2__abc_52138_new_n13356_), .Y(u2__abc_52138_new_n13386_));
NAND3X1 NAND3X1_395 ( .A(sqrto_43_), .B(sqrto_42_), .C(u2__abc_52138_new_n13371_), .Y(u2__abc_52138_new_n13401_));
NAND3X1 NAND3X1_396 ( .A(sqrto_46_), .B(sqrto_45_), .C(u2__abc_52138_new_n13394_), .Y(u2__abc_52138_new_n13409_));
NAND3X1 NAND3X1_397 ( .A(sqrto_45_), .B(sqrto_44_), .C(u2__abc_52138_new_n13387_), .Y(u2__abc_52138_new_n13417_));
NAND3X1 NAND3X1_398 ( .A(sqrto_47_), .B(sqrto_46_), .C(u2__abc_52138_new_n13402_), .Y(u2__abc_52138_new_n13432_));
NAND3X1 NAND3X1_399 ( .A(sqrto_50_), .B(sqrto_49_), .C(u2__abc_52138_new_n13425_), .Y(u2__abc_52138_new_n13440_));
NAND3X1 NAND3X1_4 ( .A(\a[118] ), .B(\a[119] ), .C(_abc_65734_new_n1482_), .Y(_abc_65734_new_n1502_));
NAND3X1 NAND3X1_40 ( .A(u2__abc_52138_new_n3857_), .B(u2__abc_52138_new_n3859_), .C(u2__abc_52138_new_n3855_), .Y(u2__abc_52138_new_n3860_));
NAND3X1 NAND3X1_400 ( .A(sqrto_49_), .B(sqrto_48_), .C(u2__abc_52138_new_n13418_), .Y(u2__abc_52138_new_n13448_));
NAND3X1 NAND3X1_401 ( .A(sqrto_51_), .B(sqrto_50_), .C(u2__abc_52138_new_n13433_), .Y(u2__abc_52138_new_n13463_));
NAND3X1 NAND3X1_402 ( .A(sqrto_54_), .B(sqrto_53_), .C(u2__abc_52138_new_n13456_), .Y(u2__abc_52138_new_n13471_));
NAND3X1 NAND3X1_403 ( .A(sqrto_53_), .B(sqrto_52_), .C(u2__abc_52138_new_n13449_), .Y(u2__abc_52138_new_n13479_));
NAND3X1 NAND3X1_404 ( .A(sqrto_55_), .B(sqrto_54_), .C(u2__abc_52138_new_n13464_), .Y(u2__abc_52138_new_n13494_));
NAND3X1 NAND3X1_405 ( .A(sqrto_58_), .B(sqrto_57_), .C(u2__abc_52138_new_n13487_), .Y(u2__abc_52138_new_n13502_));
NAND3X1 NAND3X1_406 ( .A(sqrto_57_), .B(sqrto_56_), .C(u2__abc_52138_new_n13480_), .Y(u2__abc_52138_new_n13510_));
NAND3X1 NAND3X1_407 ( .A(sqrto_59_), .B(sqrto_58_), .C(u2__abc_52138_new_n13495_), .Y(u2__abc_52138_new_n13525_));
NAND3X1 NAND3X1_408 ( .A(sqrto_62_), .B(sqrto_61_), .C(u2__abc_52138_new_n13518_), .Y(u2__abc_52138_new_n13533_));
NAND3X1 NAND3X1_409 ( .A(sqrto_61_), .B(sqrto_60_), .C(u2__abc_52138_new_n13511_), .Y(u2__abc_52138_new_n13541_));
NAND3X1 NAND3X1_41 ( .A(u2__abc_52138_new_n3863_), .B(u2__abc_52138_new_n3865_), .C(u2__abc_52138_new_n3861_), .Y(u2__abc_52138_new_n3866_));
NAND3X1 NAND3X1_410 ( .A(sqrto_63_), .B(sqrto_62_), .C(u2__abc_52138_new_n13526_), .Y(u2__abc_52138_new_n13556_));
NAND3X1 NAND3X1_411 ( .A(sqrto_66_), .B(sqrto_65_), .C(u2__abc_52138_new_n13549_), .Y(u2__abc_52138_new_n13564_));
NAND3X1 NAND3X1_412 ( .A(sqrto_65_), .B(sqrto_64_), .C(u2__abc_52138_new_n13542_), .Y(u2__abc_52138_new_n13572_));
NAND3X1 NAND3X1_413 ( .A(sqrto_67_), .B(sqrto_66_), .C(u2__abc_52138_new_n13557_), .Y(u2__abc_52138_new_n13587_));
NAND3X1 NAND3X1_414 ( .A(sqrto_70_), .B(sqrto_69_), .C(u2__abc_52138_new_n13580_), .Y(u2__abc_52138_new_n13595_));
NAND3X1 NAND3X1_415 ( .A(sqrto_69_), .B(sqrto_68_), .C(u2__abc_52138_new_n13573_), .Y(u2__abc_52138_new_n13603_));
NAND3X1 NAND3X1_416 ( .A(sqrto_71_), .B(sqrto_70_), .C(u2__abc_52138_new_n13588_), .Y(u2__abc_52138_new_n13618_));
NAND3X1 NAND3X1_417 ( .A(sqrto_74_), .B(sqrto_73_), .C(u2__abc_52138_new_n13611_), .Y(u2__abc_52138_new_n13626_));
NAND3X1 NAND3X1_418 ( .A(sqrto_73_), .B(sqrto_72_), .C(u2__abc_52138_new_n13604_), .Y(u2__abc_52138_new_n13634_));
NAND3X1 NAND3X1_419 ( .A(sqrto_75_), .B(sqrto_74_), .C(u2__abc_52138_new_n13619_), .Y(u2__abc_52138_new_n13649_));
NAND3X1 NAND3X1_42 ( .A(u2__abc_52138_new_n3849_), .B(u2__abc_52138_new_n3851_), .C(u2__abc_52138_new_n3872_), .Y(u2__abc_52138_new_n3873_));
NAND3X1 NAND3X1_420 ( .A(sqrto_78_), .B(sqrto_77_), .C(u2__abc_52138_new_n13642_), .Y(u2__abc_52138_new_n13657_));
NAND3X1 NAND3X1_421 ( .A(sqrto_77_), .B(sqrto_76_), .C(u2__abc_52138_new_n13635_), .Y(u2__abc_52138_new_n13664_));
NAND3X1 NAND3X1_422 ( .A(sqrto_79_), .B(sqrto_78_), .C(u2__abc_52138_new_n13650_), .Y(u2__abc_52138_new_n13680_));
NAND3X1 NAND3X1_423 ( .A(sqrto_82_), .B(sqrto_81_), .C(u2__abc_52138_new_n13673_), .Y(u2__abc_52138_new_n13688_));
NAND3X1 NAND3X1_424 ( .A(sqrto_81_), .B(sqrto_80_), .C(u2__abc_52138_new_n13665_), .Y(u2__abc_52138_new_n13696_));
NAND3X1 NAND3X1_425 ( .A(sqrto_83_), .B(sqrto_82_), .C(u2__abc_52138_new_n13681_), .Y(u2__abc_52138_new_n13711_));
NAND3X1 NAND3X1_426 ( .A(sqrto_86_), .B(sqrto_85_), .C(u2__abc_52138_new_n13704_), .Y(u2__abc_52138_new_n13719_));
NAND3X1 NAND3X1_427 ( .A(sqrto_85_), .B(sqrto_84_), .C(u2__abc_52138_new_n13697_), .Y(u2__abc_52138_new_n13726_));
NAND3X1 NAND3X1_428 ( .A(sqrto_87_), .B(sqrto_86_), .C(u2__abc_52138_new_n13712_), .Y(u2__abc_52138_new_n13742_));
NAND3X1 NAND3X1_429 ( .A(sqrto_90_), .B(sqrto_89_), .C(u2__abc_52138_new_n13735_), .Y(u2__abc_52138_new_n13750_));
NAND3X1 NAND3X1_43 ( .A(sqrto_82_), .B(u2__abc_52138_new_n3779_), .C(u2__abc_52138_new_n3773_), .Y(u2__abc_52138_new_n3916_));
NAND3X1 NAND3X1_430 ( .A(sqrto_89_), .B(sqrto_88_), .C(u2__abc_52138_new_n13727_), .Y(u2__abc_52138_new_n13757_));
NAND3X1 NAND3X1_431 ( .A(sqrto_91_), .B(sqrto_90_), .C(u2__abc_52138_new_n13743_), .Y(u2__abc_52138_new_n13772_));
NAND3X1 NAND3X1_432 ( .A(sqrto_94_), .B(sqrto_93_), .C(u2__abc_52138_new_n13766_), .Y(u2__abc_52138_new_n13781_));
NAND3X1 NAND3X1_433 ( .A(sqrto_93_), .B(sqrto_92_), .C(u2__abc_52138_new_n13758_), .Y(u2__abc_52138_new_n13789_));
NAND3X1 NAND3X1_434 ( .A(sqrto_95_), .B(sqrto_94_), .C(u2__abc_52138_new_n13773_), .Y(u2__abc_52138_new_n13804_));
NAND3X1 NAND3X1_435 ( .A(sqrto_98_), .B(sqrto_97_), .C(u2__abc_52138_new_n13797_), .Y(u2__abc_52138_new_n13812_));
NAND3X1 NAND3X1_436 ( .A(sqrto_97_), .B(sqrto_96_), .C(u2__abc_52138_new_n13790_), .Y(u2__abc_52138_new_n13820_));
NAND3X1 NAND3X1_437 ( .A(sqrto_99_), .B(sqrto_98_), .C(u2__abc_52138_new_n13805_), .Y(u2__abc_52138_new_n13835_));
NAND3X1 NAND3X1_438 ( .A(sqrto_102_), .B(sqrto_101_), .C(u2__abc_52138_new_n13828_), .Y(u2__abc_52138_new_n13843_));
NAND3X1 NAND3X1_439 ( .A(sqrto_101_), .B(sqrto_100_), .C(u2__abc_52138_new_n13821_), .Y(u2__abc_52138_new_n13850_));
NAND3X1 NAND3X1_44 ( .A(sqrto_88_), .B(u2__abc_52138_new_n3715_), .C(u2__abc_52138_new_n3719_), .Y(u2__abc_52138_new_n3924_));
NAND3X1 NAND3X1_440 ( .A(sqrto_103_), .B(sqrto_102_), .C(u2__abc_52138_new_n13836_), .Y(u2__abc_52138_new_n13866_));
NAND3X1 NAND3X1_441 ( .A(sqrto_106_), .B(sqrto_105_), .C(u2__abc_52138_new_n13859_), .Y(u2__abc_52138_new_n13874_));
NAND3X1 NAND3X1_442 ( .A(sqrto_105_), .B(sqrto_104_), .C(u2__abc_52138_new_n13851_), .Y(u2__abc_52138_new_n13881_));
NAND3X1 NAND3X1_443 ( .A(sqrto_107_), .B(sqrto_106_), .C(u2__abc_52138_new_n13867_), .Y(u2__abc_52138_new_n13896_));
NAND3X1 NAND3X1_444 ( .A(sqrto_110_), .B(sqrto_109_), .C(u2__abc_52138_new_n13890_), .Y(u2__abc_52138_new_n13905_));
NAND3X1 NAND3X1_445 ( .A(sqrto_109_), .B(sqrto_108_), .C(u2__abc_52138_new_n13882_), .Y(u2__abc_52138_new_n13913_));
NAND3X1 NAND3X1_446 ( .A(sqrto_111_), .B(sqrto_110_), .C(u2__abc_52138_new_n13897_), .Y(u2__abc_52138_new_n13928_));
NAND3X1 NAND3X1_447 ( .A(sqrto_114_), .B(sqrto_113_), .C(u2__abc_52138_new_n13921_), .Y(u2__abc_52138_new_n13936_));
NAND3X1 NAND3X1_448 ( .A(sqrto_113_), .B(sqrto_112_), .C(u2__abc_52138_new_n13914_), .Y(u2__abc_52138_new_n13943_));
NAND3X1 NAND3X1_449 ( .A(sqrto_115_), .B(sqrto_114_), .C(u2__abc_52138_new_n13929_), .Y(u2__abc_52138_new_n13958_));
NAND3X1 NAND3X1_45 ( .A(u2__abc_52138_new_n3627_), .B(u2__abc_52138_new_n3967_), .C(u2__abc_52138_new_n3965_), .Y(u2__abc_52138_new_n3968_));
NAND3X1 NAND3X1_450 ( .A(sqrto_118_), .B(sqrto_117_), .C(u2__abc_52138_new_n13952_), .Y(u2__abc_52138_new_n13968_));
NAND3X1 NAND3X1_451 ( .A(sqrto_117_), .B(sqrto_116_), .C(u2__abc_52138_new_n13944_), .Y(u2__abc_52138_new_n13976_));
NAND3X1 NAND3X1_452 ( .A(sqrto_119_), .B(sqrto_118_), .C(u2__abc_52138_new_n13959_), .Y(u2__abc_52138_new_n13990_));
NAND3X1 NAND3X1_453 ( .A(sqrto_122_), .B(sqrto_121_), .C(u2__abc_52138_new_n13984_), .Y(u2__abc_52138_new_n13999_));
NAND3X1 NAND3X1_454 ( .A(sqrto_121_), .B(sqrto_120_), .C(u2__abc_52138_new_n13977_), .Y(u2__abc_52138_new_n14007_));
NAND3X1 NAND3X1_455 ( .A(sqrto_123_), .B(sqrto_122_), .C(u2__abc_52138_new_n13991_), .Y(u2__abc_52138_new_n14021_));
NAND3X1 NAND3X1_456 ( .A(sqrto_126_), .B(sqrto_125_), .C(u2__abc_52138_new_n14015_), .Y(u2__abc_52138_new_n14030_));
NAND3X1 NAND3X1_457 ( .A(sqrto_125_), .B(sqrto_124_), .C(u2__abc_52138_new_n14008_), .Y(u2__abc_52138_new_n14038_));
NAND3X1 NAND3X1_458 ( .A(sqrto_127_), .B(sqrto_126_), .C(u2__abc_52138_new_n14022_), .Y(u2__abc_52138_new_n14053_));
NAND3X1 NAND3X1_459 ( .A(sqrto_130_), .B(sqrto_129_), .C(u2__abc_52138_new_n14046_), .Y(u2__abc_52138_new_n14062_));
NAND3X1 NAND3X1_46 ( .A(u2__abc_52138_new_n3524_), .B(u2__abc_52138_new_n3989_), .C(u2__abc_52138_new_n3988_), .Y(u2__abc_52138_new_n3990_));
NAND3X1 NAND3X1_460 ( .A(sqrto_129_), .B(sqrto_128_), .C(u2__abc_52138_new_n14039_), .Y(u2__abc_52138_new_n14070_));
NAND3X1 NAND3X1_461 ( .A(sqrto_131_), .B(sqrto_130_), .C(u2__abc_52138_new_n14054_), .Y(u2__abc_52138_new_n14085_));
NAND3X1 NAND3X1_462 ( .A(sqrto_134_), .B(sqrto_133_), .C(u2__abc_52138_new_n14078_), .Y(u2__abc_52138_new_n14093_));
NAND3X1 NAND3X1_463 ( .A(sqrto_133_), .B(sqrto_132_), .C(u2__abc_52138_new_n14071_), .Y(u2__abc_52138_new_n14100_));
NAND3X1 NAND3X1_464 ( .A(sqrto_135_), .B(sqrto_134_), .C(u2__abc_52138_new_n14086_), .Y(u2__abc_52138_new_n14116_));
NAND3X1 NAND3X1_465 ( .A(sqrto_138_), .B(sqrto_137_), .C(u2__abc_52138_new_n14109_), .Y(u2__abc_52138_new_n14124_));
NAND3X1 NAND3X1_466 ( .A(sqrto_137_), .B(sqrto_136_), .C(u2__abc_52138_new_n14101_), .Y(u2__abc_52138_new_n14131_));
NAND3X1 NAND3X1_467 ( .A(sqrto_139_), .B(sqrto_138_), .C(u2__abc_52138_new_n14117_), .Y(u2__abc_52138_new_n14146_));
NAND3X1 NAND3X1_468 ( .A(sqrto_142_), .B(sqrto_141_), .C(u2__abc_52138_new_n14140_), .Y(u2__abc_52138_new_n14155_));
NAND3X1 NAND3X1_469 ( .A(sqrto_141_), .B(sqrto_140_), .C(u2__abc_52138_new_n14132_), .Y(u2__abc_52138_new_n14163_));
NAND3X1 NAND3X1_47 ( .A(u2__abc_52138_new_n4136_), .B(u2__abc_52138_new_n4137_), .C(u2__abc_52138_new_n4142_), .Y(u2__abc_52138_new_n4143_));
NAND3X1 NAND3X1_470 ( .A(sqrto_143_), .B(sqrto_142_), .C(u2__abc_52138_new_n14147_), .Y(u2__abc_52138_new_n14178_));
NAND3X1 NAND3X1_471 ( .A(sqrto_146_), .B(sqrto_145_), .C(u2__abc_52138_new_n14171_), .Y(u2__abc_52138_new_n14186_));
NAND3X1 NAND3X1_472 ( .A(sqrto_145_), .B(sqrto_144_), .C(u2__abc_52138_new_n14164_), .Y(u2__abc_52138_new_n14193_));
NAND3X1 NAND3X1_473 ( .A(sqrto_147_), .B(sqrto_146_), .C(u2__abc_52138_new_n14179_), .Y(u2__abc_52138_new_n14208_));
NAND3X1 NAND3X1_474 ( .A(sqrto_150_), .B(sqrto_149_), .C(u2__abc_52138_new_n14202_), .Y(u2__abc_52138_new_n14217_));
NAND3X1 NAND3X1_475 ( .A(sqrto_149_), .B(sqrto_148_), .C(u2__abc_52138_new_n14194_), .Y(u2__abc_52138_new_n14225_));
NAND3X1 NAND3X1_476 ( .A(sqrto_151_), .B(sqrto_150_), .C(u2__abc_52138_new_n14209_), .Y(u2__abc_52138_new_n14239_));
NAND3X1 NAND3X1_477 ( .A(sqrto_154_), .B(sqrto_153_), .C(u2__abc_52138_new_n14233_), .Y(u2__abc_52138_new_n14248_));
NAND3X1 NAND3X1_478 ( .A(sqrto_153_), .B(sqrto_152_), .C(u2__abc_52138_new_n14226_), .Y(u2__abc_52138_new_n14256_));
NAND3X1 NAND3X1_479 ( .A(sqrto_155_), .B(sqrto_154_), .C(u2__abc_52138_new_n14240_), .Y(u2__abc_52138_new_n14270_));
NAND3X1 NAND3X1_48 ( .A(u2__abc_52138_new_n4184_), .B(u2__abc_52138_new_n4189_), .C(u2__abc_52138_new_n4179_), .Y(u2__abc_52138_new_n4190_));
NAND3X1 NAND3X1_480 ( .A(sqrto_158_), .B(sqrto_157_), .C(u2__abc_52138_new_n14264_), .Y(u2__abc_52138_new_n14279_));
NAND3X1 NAND3X1_481 ( .A(sqrto_157_), .B(sqrto_156_), .C(u2__abc_52138_new_n14257_), .Y(u2__abc_52138_new_n14287_));
NAND3X1 NAND3X1_482 ( .A(sqrto_159_), .B(sqrto_158_), .C(u2__abc_52138_new_n14271_), .Y(u2__abc_52138_new_n14302_));
NAND3X1 NAND3X1_483 ( .A(sqrto_162_), .B(sqrto_161_), .C(u2__abc_52138_new_n14295_), .Y(u2__abc_52138_new_n14310_));
NAND3X1 NAND3X1_484 ( .A(sqrto_161_), .B(sqrto_160_), .C(u2__abc_52138_new_n14288_), .Y(u2__abc_52138_new_n14317_));
NAND3X1 NAND3X1_485 ( .A(sqrto_163_), .B(sqrto_162_), .C(u2__abc_52138_new_n14303_), .Y(u2__abc_52138_new_n14332_));
NAND3X1 NAND3X1_486 ( .A(sqrto_166_), .B(sqrto_165_), .C(u2__abc_52138_new_n14326_), .Y(u2__abc_52138_new_n14341_));
NAND3X1 NAND3X1_487 ( .A(sqrto_165_), .B(sqrto_164_), .C(u2__abc_52138_new_n14318_), .Y(u2__abc_52138_new_n14349_));
NAND3X1 NAND3X1_488 ( .A(sqrto_167_), .B(sqrto_166_), .C(u2__abc_52138_new_n14333_), .Y(u2__abc_52138_new_n14363_));
NAND3X1 NAND3X1_489 ( .A(sqrto_170_), .B(sqrto_169_), .C(u2__abc_52138_new_n14357_), .Y(u2__abc_52138_new_n14372_));
NAND3X1 NAND3X1_49 ( .A(u2__abc_52138_new_n4327_), .B(u2__abc_52138_new_n4328_), .C(u2__abc_52138_new_n4322_), .Y(u2__abc_52138_new_n4329_));
NAND3X1 NAND3X1_490 ( .A(sqrto_169_), .B(sqrto_168_), .C(u2__abc_52138_new_n14350_), .Y(u2__abc_52138_new_n14380_));
NAND3X1 NAND3X1_491 ( .A(sqrto_171_), .B(sqrto_170_), .C(u2__abc_52138_new_n14364_), .Y(u2__abc_52138_new_n14394_));
NAND3X1 NAND3X1_492 ( .A(sqrto_174_), .B(sqrto_173_), .C(u2__abc_52138_new_n14388_), .Y(u2__abc_52138_new_n14403_));
NAND3X1 NAND3X1_493 ( .A(sqrto_173_), .B(sqrto_172_), .C(u2__abc_52138_new_n14381_), .Y(u2__abc_52138_new_n14411_));
NAND3X1 NAND3X1_494 ( .A(sqrto_175_), .B(sqrto_174_), .C(u2__abc_52138_new_n14395_), .Y(u2__abc_52138_new_n14425_));
NAND3X1 NAND3X1_495 ( .A(sqrto_178_), .B(sqrto_177_), .C(u2__abc_52138_new_n14419_), .Y(u2__abc_52138_new_n14434_));
NAND3X1 NAND3X1_496 ( .A(sqrto_177_), .B(sqrto_176_), .C(u2__abc_52138_new_n14412_), .Y(u2__abc_52138_new_n14442_));
NAND3X1 NAND3X1_497 ( .A(sqrto_179_), .B(sqrto_178_), .C(u2__abc_52138_new_n14426_), .Y(u2__abc_52138_new_n14456_));
NAND3X1 NAND3X1_498 ( .A(sqrto_182_), .B(sqrto_181_), .C(u2__abc_52138_new_n14450_), .Y(u2__abc_52138_new_n14465_));
NAND3X1 NAND3X1_499 ( .A(sqrto_181_), .B(sqrto_180_), .C(u2__abc_52138_new_n14443_), .Y(u2__abc_52138_new_n14473_));
NAND3X1 NAND3X1_5 ( .A(_abc_65734_new_n1475_), .B(_abc_65734_new_n1488_), .C(_abc_65734_new_n1496_), .Y(_abc_65734_new_n1505_));
NAND3X1 NAND3X1_50 ( .A(u2__abc_52138_new_n4468_), .B(u2__abc_52138_new_n4474_), .C(u2__abc_52138_new_n4462_), .Y(u2__abc_52138_new_n4475_));
NAND3X1 NAND3X1_500 ( .A(sqrto_183_), .B(sqrto_182_), .C(u2__abc_52138_new_n14457_), .Y(u2__abc_52138_new_n14487_));
NAND3X1 NAND3X1_501 ( .A(sqrto_186_), .B(sqrto_185_), .C(u2__abc_52138_new_n14481_), .Y(u2__abc_52138_new_n14496_));
NAND3X1 NAND3X1_502 ( .A(sqrto_185_), .B(sqrto_184_), .C(u2__abc_52138_new_n14474_), .Y(u2__abc_52138_new_n14504_));
NAND3X1 NAND3X1_503 ( .A(sqrto_187_), .B(sqrto_186_), .C(u2__abc_52138_new_n14488_), .Y(u2__abc_52138_new_n14518_));
NAND3X1 NAND3X1_504 ( .A(sqrto_190_), .B(sqrto_189_), .C(u2__abc_52138_new_n14512_), .Y(u2__abc_52138_new_n14527_));
NAND3X1 NAND3X1_505 ( .A(sqrto_189_), .B(sqrto_188_), .C(u2__abc_52138_new_n14505_), .Y(u2__abc_52138_new_n14534_));
NAND3X1 NAND3X1_506 ( .A(sqrto_191_), .B(sqrto_190_), .C(u2__abc_52138_new_n14519_), .Y(u2__abc_52138_new_n14550_));
NAND3X1 NAND3X1_507 ( .A(sqrto_194_), .B(sqrto_193_), .C(u2__abc_52138_new_n14543_), .Y(u2__abc_52138_new_n14558_));
NAND3X1 NAND3X1_508 ( .A(sqrto_193_), .B(sqrto_192_), .C(u2__abc_52138_new_n14535_), .Y(u2__abc_52138_new_n14565_));
NAND3X1 NAND3X1_509 ( .A(sqrto_195_), .B(sqrto_194_), .C(u2__abc_52138_new_n14551_), .Y(u2__abc_52138_new_n14580_));
NAND3X1 NAND3X1_51 ( .A(u2__abc_52138_new_n4547_), .B(u2__abc_52138_new_n4570_), .C(u2__abc_52138_new_n4524_), .Y(u2__abc_52138_new_n4571_));
NAND3X1 NAND3X1_510 ( .A(sqrto_198_), .B(sqrto_197_), .C(u2__abc_52138_new_n14574_), .Y(u2__abc_52138_new_n14589_));
NAND3X1 NAND3X1_511 ( .A(sqrto_197_), .B(sqrto_196_), .C(u2__abc_52138_new_n14566_), .Y(u2__abc_52138_new_n14597_));
NAND3X1 NAND3X1_512 ( .A(sqrto_199_), .B(sqrto_198_), .C(u2__abc_52138_new_n14581_), .Y(u2__abc_52138_new_n14611_));
NAND3X1 NAND3X1_513 ( .A(sqrto_202_), .B(sqrto_201_), .C(u2__abc_52138_new_n14605_), .Y(u2__abc_52138_new_n14621_));
NAND3X1 NAND3X1_514 ( .A(sqrto_201_), .B(sqrto_200_), .C(u2__abc_52138_new_n14598_), .Y(u2__abc_52138_new_n14629_));
NAND3X1 NAND3X1_515 ( .A(sqrto_203_), .B(sqrto_202_), .C(u2__abc_52138_new_n14612_), .Y(u2__abc_52138_new_n14643_));
NAND3X1 NAND3X1_516 ( .A(sqrto_206_), .B(sqrto_205_), .C(u2__abc_52138_new_n14637_), .Y(u2__abc_52138_new_n14652_));
NAND3X1 NAND3X1_517 ( .A(sqrto_205_), .B(sqrto_204_), .C(u2__abc_52138_new_n14630_), .Y(u2__abc_52138_new_n14660_));
NAND3X1 NAND3X1_518 ( .A(sqrto_207_), .B(sqrto_206_), .C(u2__abc_52138_new_n14644_), .Y(u2__abc_52138_new_n14674_));
NAND3X1 NAND3X1_519 ( .A(sqrto_210_), .B(sqrto_209_), .C(u2__abc_52138_new_n14668_), .Y(u2__abc_52138_new_n14683_));
NAND3X1 NAND3X1_52 ( .A(u2__abc_52138_new_n4611_), .B(u2__abc_52138_new_n4616_), .C(u2__abc_52138_new_n4606_), .Y(u2__abc_52138_new_n4617_));
NAND3X1 NAND3X1_520 ( .A(sqrto_209_), .B(sqrto_208_), .C(u2__abc_52138_new_n14661_), .Y(u2__abc_52138_new_n14691_));
NAND3X1 NAND3X1_521 ( .A(sqrto_211_), .B(sqrto_210_), .C(u2__abc_52138_new_n14675_), .Y(u2__abc_52138_new_n14705_));
NAND3X1 NAND3X1_522 ( .A(sqrto_214_), .B(sqrto_213_), .C(u2__abc_52138_new_n14699_), .Y(u2__abc_52138_new_n14714_));
NAND3X1 NAND3X1_523 ( .A(sqrto_213_), .B(sqrto_212_), .C(u2__abc_52138_new_n14692_), .Y(u2__abc_52138_new_n14722_));
NAND3X1 NAND3X1_524 ( .A(sqrto_215_), .B(sqrto_214_), .C(u2__abc_52138_new_n14706_), .Y(u2__abc_52138_new_n14736_));
NAND3X1 NAND3X1_525 ( .A(sqrto_218_), .B(sqrto_217_), .C(u2__abc_52138_new_n14730_), .Y(u2__abc_52138_new_n14745_));
NAND3X1 NAND3X1_526 ( .A(sqrto_217_), .B(sqrto_216_), .C(u2__abc_52138_new_n14723_), .Y(u2__abc_52138_new_n14753_));
NAND3X1 NAND3X1_527 ( .A(sqrto_219_), .B(sqrto_218_), .C(u2__abc_52138_new_n14737_), .Y(u2__abc_52138_new_n14767_));
NAND3X1 NAND3X1_528 ( .A(sqrto_222_), .B(sqrto_221_), .C(u2__abc_52138_new_n14761_), .Y(u2__abc_52138_new_n14776_));
NAND3X1 NAND3X1_529 ( .A(sqrto_221_), .B(sqrto_220_), .C(u2__abc_52138_new_n14754_), .Y(u2__abc_52138_new_n14783_));
NAND3X1 NAND3X1_53 ( .A(u2__abc_52138_new_n4648_), .B(u2__abc_52138_new_n4650_), .C(u2__abc_52138_new_n4646_), .Y(u2__abc_52138_new_n4651_));
NAND3X1 NAND3X1_530 ( .A(sqrto_223_), .B(sqrto_222_), .C(u2__abc_52138_new_n14768_), .Y(u2__abc_52138_new_n14798_));
NAND3X1 NAND3X1_531 ( .A(u2_o_226_), .B(sqrto_225_), .C(u2__abc_52138_new_n14792_), .Y(u2__abc_52138_new_n14807_));
NAND3X1 NAND3X1_532 ( .A(sqrto_225_), .B(sqrto_224_), .C(u2__abc_52138_new_n14784_), .Y(u2__abc_52138_new_n14815_));
NAND3X1 NAND3X1_533 ( .A(u2_o_227_), .B(u2_o_226_), .C(u2__abc_52138_new_n14799_), .Y(u2__abc_52138_new_n14829_));
NAND3X1 NAND3X1_534 ( .A(u2_o_230_), .B(u2_o_229_), .C(u2__abc_52138_new_n14823_), .Y(u2__abc_52138_new_n14838_));
NAND3X1 NAND3X1_535 ( .A(u2_o_229_), .B(u2_o_228_), .C(u2__abc_52138_new_n14816_), .Y(u2__abc_52138_new_n14846_));
NAND3X1 NAND3X1_536 ( .A(u2_o_231_), .B(u2_o_230_), .C(u2__abc_52138_new_n14830_), .Y(u2__abc_52138_new_n14860_));
NAND3X1 NAND3X1_537 ( .A(u2_o_234_), .B(u2_o_233_), .C(u2__abc_52138_new_n14854_), .Y(u2__abc_52138_new_n14869_));
NAND3X1 NAND3X1_538 ( .A(u2_o_233_), .B(u2_o_232_), .C(u2__abc_52138_new_n14847_), .Y(u2__abc_52138_new_n14877_));
NAND3X1 NAND3X1_539 ( .A(u2_o_235_), .B(u2_o_234_), .C(u2__abc_52138_new_n14861_), .Y(u2__abc_52138_new_n14891_));
NAND3X1 NAND3X1_54 ( .A(u2__abc_52138_new_n4654_), .B(u2__abc_52138_new_n4657_), .C(u2__abc_52138_new_n4662_), .Y(u2__abc_52138_new_n4663_));
NAND3X1 NAND3X1_540 ( .A(u2_o_238_), .B(u2_o_237_), .C(u2__abc_52138_new_n14885_), .Y(u2__abc_52138_new_n14900_));
NAND3X1 NAND3X1_541 ( .A(u2_o_237_), .B(u2_o_236_), .C(u2__abc_52138_new_n14878_), .Y(u2__abc_52138_new_n14907_));
NAND3X1 NAND3X1_542 ( .A(u2_o_239_), .B(u2_o_238_), .C(u2__abc_52138_new_n14892_), .Y(u2__abc_52138_new_n14922_));
NAND3X1 NAND3X1_543 ( .A(u2_o_242_), .B(u2_o_241_), .C(u2__abc_52138_new_n14916_), .Y(u2__abc_52138_new_n14931_));
NAND3X1 NAND3X1_544 ( .A(u2_o_241_), .B(u2_o_240_), .C(u2__abc_52138_new_n14908_), .Y(u2__abc_52138_new_n14939_));
NAND3X1 NAND3X1_545 ( .A(u2_o_243_), .B(u2_o_242_), .C(u2__abc_52138_new_n14923_), .Y(u2__abc_52138_new_n14953_));
NAND3X1 NAND3X1_546 ( .A(u2_o_246_), .B(u2_o_245_), .C(u2__abc_52138_new_n14947_), .Y(u2__abc_52138_new_n14962_));
NAND3X1 NAND3X1_547 ( .A(u2_o_245_), .B(u2_o_244_), .C(u2__abc_52138_new_n14940_), .Y(u2__abc_52138_new_n14969_));
NAND3X1 NAND3X1_548 ( .A(u2_o_247_), .B(u2_o_246_), .C(u2__abc_52138_new_n14954_), .Y(u2__abc_52138_new_n14984_));
NAND3X1 NAND3X1_549 ( .A(u2_o_250_), .B(u2_o_249_), .C(u2__abc_52138_new_n14978_), .Y(u2__abc_52138_new_n14993_));
NAND3X1 NAND3X1_55 ( .A(u2__abc_52138_new_n4641_), .B(u2__abc_52138_new_n4664_), .C(u2__abc_52138_new_n4618_), .Y(u2__abc_52138_new_n4665_));
NAND3X1 NAND3X1_550 ( .A(u2_o_249_), .B(u2_o_248_), .C(u2__abc_52138_new_n14970_), .Y(u2__abc_52138_new_n15000_));
NAND3X1 NAND3X1_551 ( .A(u2_o_251_), .B(u2_o_250_), .C(u2__abc_52138_new_n14985_), .Y(u2__abc_52138_new_n15015_));
NAND3X1 NAND3X1_552 ( .A(u2_o_254_), .B(u2_o_253_), .C(u2__abc_52138_new_n15009_), .Y(u2__abc_52138_new_n15024_));
NAND3X1 NAND3X1_553 ( .A(u2_o_253_), .B(u2_o_252_), .C(u2__abc_52138_new_n15001_), .Y(u2__abc_52138_new_n15031_));
NAND3X1 NAND3X1_554 ( .A(u2_o_255_), .B(u2_o_254_), .C(u2__abc_52138_new_n15016_), .Y(u2__abc_52138_new_n15047_));
NAND3X1 NAND3X1_555 ( .A(u2_o_258_), .B(u2_o_257_), .C(u2__abc_52138_new_n15040_), .Y(u2__abc_52138_new_n15055_));
NAND3X1 NAND3X1_556 ( .A(u2_o_257_), .B(u2_o_256_), .C(u2__abc_52138_new_n15032_), .Y(u2__abc_52138_new_n15062_));
NAND3X1 NAND3X1_557 ( .A(u2_o_259_), .B(u2_o_258_), .C(u2__abc_52138_new_n15048_), .Y(u2__abc_52138_new_n15077_));
NAND3X1 NAND3X1_558 ( .A(u2_o_262_), .B(u2_o_261_), .C(u2__abc_52138_new_n15071_), .Y(u2__abc_52138_new_n15086_));
NAND3X1 NAND3X1_559 ( .A(u2_o_261_), .B(u2_o_260_), .C(u2__abc_52138_new_n15063_), .Y(u2__abc_52138_new_n15094_));
NAND3X1 NAND3X1_56 ( .A(u2__abc_52138_new_n4728_), .B(u2__abc_52138_new_n4730_), .C(u2__abc_52138_new_n4726_), .Y(u2__abc_52138_new_n4731_));
NAND3X1 NAND3X1_560 ( .A(u2_o_263_), .B(u2_o_262_), .C(u2__abc_52138_new_n15078_), .Y(u2__abc_52138_new_n15108_));
NAND3X1 NAND3X1_561 ( .A(u2_o_266_), .B(u2_o_265_), .C(u2__abc_52138_new_n15102_), .Y(u2__abc_52138_new_n15117_));
NAND3X1 NAND3X1_562 ( .A(u2_o_265_), .B(u2_o_264_), .C(u2__abc_52138_new_n15095_), .Y(u2__abc_52138_new_n15125_));
NAND3X1 NAND3X1_563 ( .A(u2_o_267_), .B(u2_o_266_), .C(u2__abc_52138_new_n15109_), .Y(u2__abc_52138_new_n15139_));
NAND3X1 NAND3X1_564 ( .A(u2_o_270_), .B(u2_o_269_), .C(u2__abc_52138_new_n15133_), .Y(u2__abc_52138_new_n15148_));
NAND3X1 NAND3X1_565 ( .A(u2_o_269_), .B(u2_o_268_), .C(u2__abc_52138_new_n15126_), .Y(u2__abc_52138_new_n15156_));
NAND3X1 NAND3X1_566 ( .A(u2_o_271_), .B(u2_o_270_), .C(u2__abc_52138_new_n15140_), .Y(u2__abc_52138_new_n15170_));
NAND3X1 NAND3X1_567 ( .A(u2_o_274_), .B(u2_o_273_), .C(u2__abc_52138_new_n15164_), .Y(u2__abc_52138_new_n15179_));
NAND3X1 NAND3X1_568 ( .A(u2_o_273_), .B(u2_o_272_), .C(u2__abc_52138_new_n15157_), .Y(u2__abc_52138_new_n15187_));
NAND3X1 NAND3X1_569 ( .A(u2_o_275_), .B(u2_o_274_), .C(u2__abc_52138_new_n15171_), .Y(u2__abc_52138_new_n15201_));
NAND3X1 NAND3X1_57 ( .A(u2__abc_52138_new_n4748_), .B(u2__abc_52138_new_n4749_), .C(u2__abc_52138_new_n4743_), .Y(u2__abc_52138_new_n4750_));
NAND3X1 NAND3X1_570 ( .A(u2_o_278_), .B(u2_o_277_), .C(u2__abc_52138_new_n15195_), .Y(u2__abc_52138_new_n15210_));
NAND3X1 NAND3X1_571 ( .A(u2_o_277_), .B(u2_o_276_), .C(u2__abc_52138_new_n15188_), .Y(u2__abc_52138_new_n15218_));
NAND3X1 NAND3X1_572 ( .A(u2_o_279_), .B(u2_o_278_), .C(u2__abc_52138_new_n15202_), .Y(u2__abc_52138_new_n15232_));
NAND3X1 NAND3X1_573 ( .A(u2_o_282_), .B(u2_o_281_), .C(u2__abc_52138_new_n15226_), .Y(u2__abc_52138_new_n15241_));
NAND3X1 NAND3X1_574 ( .A(u2_o_281_), .B(u2_o_280_), .C(u2__abc_52138_new_n15219_), .Y(u2__abc_52138_new_n15249_));
NAND3X1 NAND3X1_575 ( .A(u2_o_283_), .B(u2_o_282_), .C(u2__abc_52138_new_n15233_), .Y(u2__abc_52138_new_n15263_));
NAND3X1 NAND3X1_576 ( .A(u2_o_286_), .B(u2_o_285_), .C(u2__abc_52138_new_n15257_), .Y(u2__abc_52138_new_n15272_));
NAND3X1 NAND3X1_577 ( .A(u2_o_285_), .B(u2_o_284_), .C(u2__abc_52138_new_n15250_), .Y(u2__abc_52138_new_n15279_));
NAND3X1 NAND3X1_578 ( .A(u2_o_287_), .B(u2_o_286_), .C(u2__abc_52138_new_n15264_), .Y(u2__abc_52138_new_n15294_));
NAND3X1 NAND3X1_579 ( .A(u2_o_290_), .B(u2_o_289_), .C(u2__abc_52138_new_n15288_), .Y(u2__abc_52138_new_n15303_));
NAND3X1 NAND3X1_58 ( .A(u2__abc_52138_new_n4572_), .B(u2__abc_52138_new_n4752_), .C(u2__abc_52138_new_n4381_), .Y(u2__abc_52138_new_n4753_));
NAND3X1 NAND3X1_580 ( .A(u2_o_289_), .B(u2_o_288_), .C(u2__abc_52138_new_n15280_), .Y(u2__abc_52138_new_n15311_));
NAND3X1 NAND3X1_581 ( .A(u2_o_291_), .B(u2_o_290_), .C(u2__abc_52138_new_n15295_), .Y(u2__abc_52138_new_n15325_));
NAND3X1 NAND3X1_582 ( .A(u2_o_294_), .B(u2_o_293_), .C(u2__abc_52138_new_n15319_), .Y(u2__abc_52138_new_n15334_));
NAND3X1 NAND3X1_583 ( .A(u2_o_293_), .B(u2_o_292_), .C(u2__abc_52138_new_n15312_), .Y(u2__abc_52138_new_n15342_));
NAND3X1 NAND3X1_584 ( .A(u2_o_295_), .B(u2_o_294_), .C(u2__abc_52138_new_n15326_), .Y(u2__abc_52138_new_n15356_));
NAND3X1 NAND3X1_585 ( .A(u2_o_298_), .B(u2_o_297_), .C(u2__abc_52138_new_n15350_), .Y(u2__abc_52138_new_n15365_));
NAND3X1 NAND3X1_586 ( .A(u2_o_297_), .B(u2_o_296_), .C(u2__abc_52138_new_n15343_), .Y(u2__abc_52138_new_n15373_));
NAND3X1 NAND3X1_587 ( .A(u2_o_299_), .B(u2_o_298_), .C(u2__abc_52138_new_n15357_), .Y(u2__abc_52138_new_n15387_));
NAND3X1 NAND3X1_588 ( .A(u2_o_302_), .B(u2_o_301_), .C(u2__abc_52138_new_n15381_), .Y(u2__abc_52138_new_n15396_));
NAND3X1 NAND3X1_589 ( .A(u2_o_301_), .B(u2_o_300_), .C(u2__abc_52138_new_n15374_), .Y(u2__abc_52138_new_n15403_));
NAND3X1 NAND3X1_59 ( .A(u2__abc_52138_new_n4511_), .B(u2__abc_52138_new_n4522_), .C(u2__abc_52138_new_n4755_), .Y(u2__abc_52138_new_n4756_));
NAND3X1 NAND3X1_590 ( .A(u2_o_303_), .B(u2_o_302_), .C(u2__abc_52138_new_n15388_), .Y(u2__abc_52138_new_n15418_));
NAND3X1 NAND3X1_591 ( .A(u2_o_306_), .B(u2_o_305_), .C(u2__abc_52138_new_n15412_), .Y(u2__abc_52138_new_n15427_));
NAND3X1 NAND3X1_592 ( .A(u2_o_305_), .B(u2_o_304_), .C(u2__abc_52138_new_n15404_), .Y(u2__abc_52138_new_n15435_));
NAND3X1 NAND3X1_593 ( .A(u2_o_307_), .B(u2_o_306_), .C(u2__abc_52138_new_n15419_), .Y(u2__abc_52138_new_n15449_));
NAND3X1 NAND3X1_594 ( .A(u2_o_310_), .B(u2_o_309_), .C(u2__abc_52138_new_n15443_), .Y(u2__abc_52138_new_n15458_));
NAND3X1 NAND3X1_595 ( .A(u2_o_309_), .B(u2_o_308_), .C(u2__abc_52138_new_n15436_), .Y(u2__abc_52138_new_n15465_));
NAND3X1 NAND3X1_596 ( .A(u2_o_311_), .B(u2_o_310_), .C(u2__abc_52138_new_n15450_), .Y(u2__abc_52138_new_n15480_));
NAND3X1 NAND3X1_597 ( .A(u2_o_314_), .B(u2_o_313_), .C(u2__abc_52138_new_n15474_), .Y(u2__abc_52138_new_n15490_));
NAND3X1 NAND3X1_598 ( .A(u2_o_313_), .B(u2_o_312_), .C(u2__abc_52138_new_n15466_), .Y(u2__abc_52138_new_n15497_));
NAND3X1 NAND3X1_599 ( .A(u2_o_315_), .B(u2_o_314_), .C(u2__abc_52138_new_n15481_), .Y(u2__abc_52138_new_n15512_));
NAND3X1 NAND3X1_6 ( .A(\a[119] ), .B(_abc_65734_new_n1510_), .C(_abc_65734_new_n1511_), .Y(_abc_65734_new_n1512_));
NAND3X1 NAND3X1_60 ( .A(u2__abc_52138_new_n4739_), .B(u2__abc_52138_new_n4741_), .C(u2__abc_52138_new_n4763_), .Y(u2__abc_52138_new_n4764_));
NAND3X1 NAND3X1_600 ( .A(u2_o_318_), .B(u2_o_317_), .C(u2__abc_52138_new_n15506_), .Y(u2__abc_52138_new_n15521_));
NAND3X1 NAND3X1_601 ( .A(u2_o_317_), .B(u2_o_316_), .C(u2__abc_52138_new_n15498_), .Y(u2__abc_52138_new_n15528_));
NAND3X1 NAND3X1_602 ( .A(u2_o_319_), .B(u2_o_318_), .C(u2__abc_52138_new_n15513_), .Y(u2__abc_52138_new_n15543_));
NAND3X1 NAND3X1_603 ( .A(u2_o_322_), .B(u2_o_321_), .C(u2__abc_52138_new_n15537_), .Y(u2__abc_52138_new_n15552_));
NAND3X1 NAND3X1_604 ( .A(u2_o_321_), .B(u2_o_320_), .C(u2__abc_52138_new_n15529_), .Y(u2__abc_52138_new_n15560_));
NAND3X1 NAND3X1_605 ( .A(u2_o_323_), .B(u2_o_322_), .C(u2__abc_52138_new_n15544_), .Y(u2__abc_52138_new_n15574_));
NAND3X1 NAND3X1_606 ( .A(u2_o_326_), .B(u2_o_325_), .C(u2__abc_52138_new_n15568_), .Y(u2__abc_52138_new_n15583_));
NAND3X1 NAND3X1_607 ( .A(u2_o_325_), .B(u2_o_324_), .C(u2__abc_52138_new_n15561_), .Y(u2__abc_52138_new_n15591_));
NAND3X1 NAND3X1_608 ( .A(u2_o_327_), .B(u2_o_326_), .C(u2__abc_52138_new_n15575_), .Y(u2__abc_52138_new_n15605_));
NAND3X1 NAND3X1_609 ( .A(u2_o_330_), .B(u2_o_329_), .C(u2__abc_52138_new_n15599_), .Y(u2__abc_52138_new_n15614_));
NAND3X1 NAND3X1_61 ( .A(u2__abc_52138_new_n4486_), .B(u2__abc_52138_new_n4854_), .C(u2__abc_52138_new_n4852_), .Y(u2__abc_52138_new_n4855_));
NAND3X1 NAND3X1_610 ( .A(u2_o_329_), .B(u2_o_328_), .C(u2__abc_52138_new_n15592_), .Y(u2__abc_52138_new_n15622_));
NAND3X1 NAND3X1_611 ( .A(u2_o_331_), .B(u2_o_330_), .C(u2__abc_52138_new_n15606_), .Y(u2__abc_52138_new_n15636_));
NAND3X1 NAND3X1_612 ( .A(u2_o_334_), .B(u2_o_333_), .C(u2__abc_52138_new_n15630_), .Y(u2__abc_52138_new_n15646_));
NAND3X1 NAND3X1_613 ( .A(u2_o_333_), .B(u2_o_332_), .C(u2__abc_52138_new_n15623_), .Y(u2__abc_52138_new_n15653_));
NAND3X1 NAND3X1_614 ( .A(u2_o_335_), .B(u2_o_334_), .C(u2__abc_52138_new_n15637_), .Y(u2__abc_52138_new_n15668_));
NAND3X1 NAND3X1_615 ( .A(u2_o_338_), .B(u2_o_337_), .C(u2__abc_52138_new_n15662_), .Y(u2__abc_52138_new_n15678_));
NAND3X1 NAND3X1_616 ( .A(u2_o_337_), .B(u2_o_336_), .C(u2__abc_52138_new_n15654_), .Y(u2__abc_52138_new_n15686_));
NAND3X1 NAND3X1_617 ( .A(u2_o_339_), .B(u2_o_338_), .C(u2__abc_52138_new_n15669_), .Y(u2__abc_52138_new_n15700_));
NAND3X1 NAND3X1_618 ( .A(u2_o_342_), .B(u2_o_341_), .C(u2__abc_52138_new_n15694_), .Y(u2__abc_52138_new_n15709_));
NAND3X1 NAND3X1_619 ( .A(u2_o_341_), .B(u2_o_340_), .C(u2__abc_52138_new_n15687_), .Y(u2__abc_52138_new_n15716_));
NAND3X1 NAND3X1_62 ( .A(u2__abc_52138_new_n4320_), .B(u2__abc_52138_new_n4910_), .C(u2__abc_52138_new_n4908_), .Y(u2__abc_52138_new_n4911_));
NAND3X1 NAND3X1_620 ( .A(u2_o_343_), .B(u2_o_342_), .C(u2__abc_52138_new_n15701_), .Y(u2__abc_52138_new_n15731_));
NAND3X1 NAND3X1_621 ( .A(u2_o_346_), .B(u2_o_345_), .C(u2__abc_52138_new_n15725_), .Y(u2__abc_52138_new_n15740_));
NAND3X1 NAND3X1_622 ( .A(u2_o_345_), .B(u2_o_344_), .C(u2__abc_52138_new_n15717_), .Y(u2__abc_52138_new_n15747_));
NAND3X1 NAND3X1_623 ( .A(u2_o_347_), .B(u2_o_346_), .C(u2__abc_52138_new_n15732_), .Y(u2__abc_52138_new_n15762_));
NAND3X1 NAND3X1_624 ( .A(u2_o_350_), .B(u2_o_349_), .C(u2__abc_52138_new_n15756_), .Y(u2__abc_52138_new_n15771_));
NAND3X1 NAND3X1_625 ( .A(u2_o_349_), .B(u2_o_348_), .C(u2__abc_52138_new_n15748_), .Y(u2__abc_52138_new_n15778_));
NAND3X1 NAND3X1_626 ( .A(u2_o_351_), .B(u2_o_350_), .C(u2__abc_52138_new_n15763_), .Y(u2__abc_52138_new_n15793_));
NAND3X1 NAND3X1_627 ( .A(u2_o_354_), .B(u2_o_353_), .C(u2__abc_52138_new_n15787_), .Y(u2__abc_52138_new_n15802_));
NAND3X1 NAND3X1_628 ( .A(u2_o_353_), .B(u2_o_352_), .C(u2__abc_52138_new_n15779_), .Y(u2__abc_52138_new_n15810_));
NAND3X1 NAND3X1_629 ( .A(u2_o_355_), .B(u2_o_354_), .C(u2__abc_52138_new_n15794_), .Y(u2__abc_52138_new_n15824_));
NAND3X1 NAND3X1_63 ( .A(u2__abc_52138_new_n5199_), .B(u2__abc_52138_new_n5204_), .C(u2__abc_52138_new_n5194_), .Y(u2__abc_52138_new_n5205_));
NAND3X1 NAND3X1_630 ( .A(u2_o_358_), .B(u2_o_357_), .C(u2__abc_52138_new_n15818_), .Y(u2__abc_52138_new_n15833_));
NAND3X1 NAND3X1_631 ( .A(u2_o_357_), .B(u2_o_356_), .C(u2__abc_52138_new_n15811_), .Y(u2__abc_52138_new_n15840_));
NAND3X1 NAND3X1_632 ( .A(u2_o_359_), .B(u2_o_358_), .C(u2__abc_52138_new_n15825_), .Y(u2__abc_52138_new_n15855_));
NAND3X1 NAND3X1_633 ( .A(u2_o_362_), .B(u2_o_361_), .C(u2__abc_52138_new_n15849_), .Y(u2__abc_52138_new_n15864_));
NAND3X1 NAND3X1_634 ( .A(u2_o_361_), .B(u2_o_360_), .C(u2__abc_52138_new_n15841_), .Y(u2__abc_52138_new_n15871_));
NAND3X1 NAND3X1_635 ( .A(u2_o_363_), .B(u2_o_362_), .C(u2__abc_52138_new_n15856_), .Y(u2__abc_52138_new_n15886_));
NAND3X1 NAND3X1_636 ( .A(u2_o_366_), .B(u2_o_365_), .C(u2__abc_52138_new_n15880_), .Y(u2__abc_52138_new_n15895_));
NAND3X1 NAND3X1_637 ( .A(u2_o_365_), .B(u2_o_364_), .C(u2__abc_52138_new_n15872_), .Y(u2__abc_52138_new_n15902_));
NAND3X1 NAND3X1_638 ( .A(u2_o_367_), .B(u2_o_366_), .C(u2__abc_52138_new_n15887_), .Y(u2__abc_52138_new_n15918_));
NAND3X1 NAND3X1_639 ( .A(u2_o_370_), .B(u2_o_369_), .C(u2__abc_52138_new_n15911_), .Y(u2__abc_52138_new_n15927_));
NAND3X1 NAND3X1_64 ( .A(u2__abc_52138_new_n5207_), .B(u2__abc_52138_new_n5209_), .C(u2__abc_52138_new_n5214_), .Y(u2__abc_52138_new_n5215_));
NAND3X1 NAND3X1_640 ( .A(u2_o_369_), .B(u2_o_368_), .C(u2__abc_52138_new_n15903_), .Y(u2__abc_52138_new_n15934_));
NAND3X1 NAND3X1_641 ( .A(u2_o_371_), .B(u2_o_370_), .C(u2__abc_52138_new_n15919_), .Y(u2__abc_52138_new_n15949_));
NAND3X1 NAND3X1_642 ( .A(u2_o_374_), .B(u2_o_373_), .C(u2__abc_52138_new_n15943_), .Y(u2__abc_52138_new_n15958_));
NAND3X1 NAND3X1_643 ( .A(u2_o_373_), .B(u2_o_372_), .C(u2__abc_52138_new_n15935_), .Y(u2__abc_52138_new_n15965_));
NAND3X1 NAND3X1_644 ( .A(u2_o_375_), .B(u2_o_374_), .C(u2__abc_52138_new_n15950_), .Y(u2__abc_52138_new_n15980_));
NAND3X1 NAND3X1_645 ( .A(u2_o_378_), .B(u2_o_377_), .C(u2__abc_52138_new_n15974_), .Y(u2__abc_52138_new_n15989_));
NAND3X1 NAND3X1_646 ( .A(u2_o_377_), .B(u2_o_376_), .C(u2__abc_52138_new_n15966_), .Y(u2__abc_52138_new_n15996_));
NAND3X1 NAND3X1_647 ( .A(u2_o_379_), .B(u2_o_378_), .C(u2__abc_52138_new_n15981_), .Y(u2__abc_52138_new_n16011_));
NAND3X1 NAND3X1_648 ( .A(u2_o_382_), .B(u2_o_381_), .C(u2__abc_52138_new_n16005_), .Y(u2__abc_52138_new_n16020_));
NAND3X1 NAND3X1_649 ( .A(u2_o_381_), .B(u2_o_380_), .C(u2__abc_52138_new_n15997_), .Y(u2__abc_52138_new_n16027_));
NAND3X1 NAND3X1_65 ( .A(u2__abc_52138_new_n5241_), .B(u2__abc_52138_new_n5247_), .C(u2__abc_52138_new_n5240_), .Y(u2__abc_52138_new_n5248_));
NAND3X1 NAND3X1_650 ( .A(u2_o_383_), .B(u2_o_382_), .C(u2__abc_52138_new_n16012_), .Y(u2__abc_52138_new_n16042_));
NAND3X1 NAND3X1_651 ( .A(u2_o_386_), .B(u2_o_385_), .C(u2__abc_52138_new_n16036_), .Y(u2__abc_52138_new_n16051_));
NAND3X1 NAND3X1_652 ( .A(u2_o_385_), .B(u2_o_384_), .C(u2__abc_52138_new_n16028_), .Y(u2__abc_52138_new_n16059_));
NAND3X1 NAND3X1_653 ( .A(u2_o_387_), .B(u2_o_386_), .C(u2__abc_52138_new_n16043_), .Y(u2__abc_52138_new_n16073_));
NAND3X1 NAND3X1_654 ( .A(u2_o_390_), .B(u2_o_389_), .C(u2__abc_52138_new_n16067_), .Y(u2__abc_52138_new_n16083_));
NAND3X1 NAND3X1_655 ( .A(u2_o_389_), .B(u2_o_388_), .C(u2__abc_52138_new_n16060_), .Y(u2__abc_52138_new_n16092_));
NAND3X1 NAND3X1_656 ( .A(u2_o_391_), .B(u2_o_390_), .C(u2__abc_52138_new_n16074_), .Y(u2__abc_52138_new_n16106_));
NAND3X1 NAND3X1_657 ( .A(u2_o_394_), .B(u2_o_393_), .C(u2__abc_52138_new_n16100_), .Y(u2__abc_52138_new_n16116_));
NAND3X1 NAND3X1_658 ( .A(u2_o_393_), .B(u2_o_392_), .C(u2__abc_52138_new_n16093_), .Y(u2__abc_52138_new_n16124_));
NAND3X1 NAND3X1_659 ( .A(u2_o_395_), .B(u2_o_394_), .C(u2__abc_52138_new_n16107_), .Y(u2__abc_52138_new_n16138_));
NAND3X1 NAND3X1_66 ( .A(u2__abc_52138_new_n5265_), .B(u2__abc_52138_new_n5270_), .C(u2__abc_52138_new_n5260_), .Y(u2__abc_52138_new_n5271_));
NAND3X1 NAND3X1_660 ( .A(u2_o_398_), .B(u2_o_397_), .C(u2__abc_52138_new_n16132_), .Y(u2__abc_52138_new_n16147_));
NAND3X1 NAND3X1_661 ( .A(u2_o_397_), .B(u2_o_396_), .C(u2__abc_52138_new_n16125_), .Y(u2__abc_52138_new_n16154_));
NAND3X1 NAND3X1_662 ( .A(u2_o_399_), .B(u2_o_398_), .C(u2__abc_52138_new_n16139_), .Y(u2__abc_52138_new_n16169_));
NAND3X1 NAND3X1_663 ( .A(u2_o_402_), .B(u2_o_401_), .C(u2__abc_52138_new_n16163_), .Y(u2__abc_52138_new_n16178_));
NAND3X1 NAND3X1_664 ( .A(u2_o_401_), .B(u2_o_400_), .C(u2__abc_52138_new_n16155_), .Y(u2__abc_52138_new_n16186_));
NAND3X1 NAND3X1_665 ( .A(u2_o_403_), .B(u2_o_402_), .C(u2__abc_52138_new_n16170_), .Y(u2__abc_52138_new_n16200_));
NAND3X1 NAND3X1_666 ( .A(u2_o_406_), .B(u2_o_405_), .C(u2__abc_52138_new_n16194_), .Y(u2__abc_52138_new_n16209_));
NAND3X1 NAND3X1_667 ( .A(u2_o_405_), .B(u2_o_404_), .C(u2__abc_52138_new_n16187_), .Y(u2__abc_52138_new_n16216_));
NAND3X1 NAND3X1_668 ( .A(u2_o_407_), .B(u2_o_406_), .C(u2__abc_52138_new_n16201_), .Y(u2__abc_52138_new_n16231_));
NAND3X1 NAND3X1_669 ( .A(u2_o_410_), .B(u2_o_409_), .C(u2__abc_52138_new_n16225_), .Y(u2__abc_52138_new_n16240_));
NAND3X1 NAND3X1_67 ( .A(u2__abc_52138_new_n5751_), .B(u2__abc_52138_new_n5753_), .C(u2__abc_52138_new_n5750_), .Y(u2__abc_52138_new_n5754_));
NAND3X1 NAND3X1_670 ( .A(u2_o_409_), .B(u2_o_408_), .C(u2__abc_52138_new_n16217_), .Y(u2__abc_52138_new_n16247_));
NAND3X1 NAND3X1_671 ( .A(u2_o_411_), .B(u2_o_410_), .C(u2__abc_52138_new_n16232_), .Y(u2__abc_52138_new_n16262_));
NAND3X1 NAND3X1_672 ( .A(u2_o_414_), .B(u2_o_413_), .C(u2__abc_52138_new_n16256_), .Y(u2__abc_52138_new_n16271_));
NAND3X1 NAND3X1_673 ( .A(u2_o_413_), .B(u2_o_412_), .C(u2__abc_52138_new_n16248_), .Y(u2__abc_52138_new_n16278_));
NAND3X1 NAND3X1_674 ( .A(u2_o_415_), .B(u2_o_414_), .C(u2__abc_52138_new_n16263_), .Y(u2__abc_52138_new_n16293_));
NAND3X1 NAND3X1_675 ( .A(u2_o_418_), .B(u2_o_417_), .C(u2__abc_52138_new_n16287_), .Y(u2__abc_52138_new_n16302_));
NAND3X1 NAND3X1_676 ( .A(u2_o_417_), .B(u2_o_416_), .C(u2__abc_52138_new_n16279_), .Y(u2__abc_52138_new_n16310_));
NAND3X1 NAND3X1_677 ( .A(u2_o_419_), .B(u2_o_418_), .C(u2__abc_52138_new_n16294_), .Y(u2__abc_52138_new_n16324_));
NAND3X1 NAND3X1_678 ( .A(u2_o_422_), .B(u2_o_421_), .C(u2__abc_52138_new_n16318_), .Y(u2__abc_52138_new_n16333_));
NAND3X1 NAND3X1_679 ( .A(u2_o_421_), .B(u2_o_420_), .C(u2__abc_52138_new_n16311_), .Y(u2__abc_52138_new_n16340_));
NAND3X1 NAND3X1_68 ( .A(u2__abc_52138_new_n5776_), .B(u2__abc_52138_new_n5778_), .C(u2__abc_52138_new_n5773_), .Y(u2__abc_52138_new_n5779_));
NAND3X1 NAND3X1_680 ( .A(u2_o_423_), .B(u2_o_422_), .C(u2__abc_52138_new_n16325_), .Y(u2__abc_52138_new_n16355_));
NAND3X1 NAND3X1_681 ( .A(u2_o_426_), .B(u2_o_425_), .C(u2__abc_52138_new_n16349_), .Y(u2__abc_52138_new_n16364_));
NAND3X1 NAND3X1_682 ( .A(u2_o_425_), .B(u2_o_424_), .C(u2__abc_52138_new_n16341_), .Y(u2__abc_52138_new_n16371_));
NAND3X1 NAND3X1_683 ( .A(u2_o_427_), .B(u2_o_426_), .C(u2__abc_52138_new_n16356_), .Y(u2__abc_52138_new_n16386_));
NAND3X1 NAND3X1_684 ( .A(u2_o_430_), .B(u2_o_429_), .C(u2__abc_52138_new_n16380_), .Y(u2__abc_52138_new_n16395_));
NAND3X1 NAND3X1_685 ( .A(u2_o_429_), .B(u2_o_428_), .C(u2__abc_52138_new_n16372_), .Y(u2__abc_52138_new_n16402_));
NAND3X1 NAND3X1_686 ( .A(u2_o_431_), .B(u2_o_430_), .C(u2__abc_52138_new_n16387_), .Y(u2__abc_52138_new_n16417_));
NAND3X1 NAND3X1_687 ( .A(u2_o_434_), .B(u2_o_433_), .C(u2__abc_52138_new_n16411_), .Y(u2__abc_52138_new_n16426_));
NAND3X1 NAND3X1_688 ( .A(u2_o_433_), .B(u2_o_432_), .C(u2__abc_52138_new_n16403_), .Y(u2__abc_52138_new_n16433_));
NAND3X1 NAND3X1_689 ( .A(u2_o_435_), .B(u2_o_434_), .C(u2__abc_52138_new_n16418_), .Y(u2__abc_52138_new_n16448_));
NAND3X1 NAND3X1_69 ( .A(u2__abc_52138_new_n5804_), .B(u2__abc_52138_new_n5805_), .C(u2__abc_52138_new_n5800_), .Y(u2__abc_52138_new_n5806_));
NAND3X1 NAND3X1_690 ( .A(u2_o_438_), .B(u2_o_437_), .C(u2__abc_52138_new_n16442_), .Y(u2__abc_52138_new_n16457_));
NAND3X1 NAND3X1_691 ( .A(u2_o_437_), .B(u2_o_436_), .C(u2__abc_52138_new_n16434_), .Y(u2__abc_52138_new_n16464_));
NAND3X1 NAND3X1_692 ( .A(u2_o_439_), .B(u2_o_438_), .C(u2__abc_52138_new_n16449_), .Y(u2__abc_52138_new_n16479_));
NAND3X1 NAND3X1_693 ( .A(u2_o_442_), .B(u2_o_441_), .C(u2__abc_52138_new_n16473_), .Y(u2__abc_52138_new_n16488_));
NAND3X1 NAND3X1_694 ( .A(u2_o_441_), .B(u2_o_440_), .C(u2__abc_52138_new_n16465_), .Y(u2__abc_52138_new_n16495_));
NAND3X1 NAND3X1_695 ( .A(u2_o_443_), .B(u2_o_442_), .C(u2__abc_52138_new_n16480_), .Y(u2__abc_52138_new_n16510_));
NAND3X1 NAND3X1_696 ( .A(u2_o_446_), .B(u2_o_445_), .C(u2__abc_52138_new_n16504_), .Y(u2__abc_52138_new_n16519_));
NAND3X1 NAND3X1_697 ( .A(u2_o_445_), .B(u2_o_444_), .C(u2__abc_52138_new_n16496_), .Y(u2__abc_52138_new_n16527_));
NAND3X1 NAND3X1_7 ( .A(\a[119] ), .B(\a[120] ), .C(_abc_65734_new_n1511_), .Y(_abc_65734_new_n1516_));
NAND3X1 NAND3X1_70 ( .A(u2__abc_52138_new_n5809_), .B(u2__abc_52138_new_n5822_), .C(u2__abc_52138_new_n5817_), .Y(u2__abc_52138_new_n5823_));
NAND3X1 NAND3X1_71 ( .A(u2__abc_52138_new_n5334_), .B(u2__abc_52138_new_n5845_), .C(u2__abc_52138_new_n5843_), .Y(u2__abc_52138_new_n5846_));
NAND3X1 NAND3X1_72 ( .A(u2__abc_52138_new_n5842_), .B(u2__abc_52138_new_n5846_), .C(u2__abc_52138_new_n5841_), .Y(u2__abc_52138_new_n5847_));
NAND3X1 NAND3X1_73 ( .A(u2__abc_52138_new_n5856_), .B(u2__abc_52138_new_n5857_), .C(u2__abc_52138_new_n5853_), .Y(u2__abc_52138_new_n5858_));
NAND3X1 NAND3X1_74 ( .A(u2__abc_52138_new_n5894_), .B(u2__abc_52138_new_n5898_), .C(u2__abc_52138_new_n5897_), .Y(u2__abc_52138_new_n5899_));
NAND3X1 NAND3X1_75 ( .A(u2__abc_52138_new_n5910_), .B(u2__abc_52138_new_n5913_), .C(u2__abc_52138_new_n5909_), .Y(u2__abc_52138_new_n5914_));
NAND3X1 NAND3X1_76 ( .A(u2__abc_52138_new_n5914_), .B(u2__abc_52138_new_n5916_), .C(u2__abc_52138_new_n5908_), .Y(u2__abc_52138_new_n5917_));
NAND3X1 NAND3X1_77 ( .A(u2__abc_52138_new_n5901_), .B(u2__abc_52138_new_n5939_), .C(u2__abc_52138_new_n5928_), .Y(u2__abc_52138_new_n5940_));
NAND3X1 NAND3X1_78 ( .A(u2__abc_52138_new_n6051_), .B(u2__abc_52138_new_n6056_), .C(u2__abc_52138_new_n6046_), .Y(u2__abc_52138_new_n6057_));
NAND3X1 NAND3X1_79 ( .A(u2__abc_52138_new_n6348_), .B(u2__abc_52138_new_n6349_), .C(u2__abc_52138_new_n6355_), .Y(u2__abc_52138_new_n6356_));
NAND3X1 NAND3X1_8 ( .A(_abc_65734_new_n1503_), .B(_abc_65734_new_n1518_), .C(_abc_65734_new_n1495_), .Y(_abc_65734_new_n1522_));
NAND3X1 NAND3X1_80 ( .A(u2__abc_52138_new_n6423_), .B(u2__abc_52138_new_n6425_), .C(u2__abc_52138_new_n6421_), .Y(u2__abc_52138_new_n6426_));
NAND3X1 NAND3X1_81 ( .A(u2__abc_52138_new_n4192_), .B(u2__abc_52138_new_n4754_), .C(u2__abc_52138_new_n6451_), .Y(u2__abc_52138_new_n6452_));
NAND3X1 NAND3X1_82 ( .A(u2__abc_52138_new_n6107_), .B(u2__abc_52138_new_n6131_), .C(u2__abc_52138_new_n4377_), .Y(u2__abc_52138_new_n6453_));
NAND3X1 NAND3X1_83 ( .A(u2__abc_52138_new_n6457_), .B(u2__abc_52138_new_n6468_), .C(u2__abc_52138_new_n3015_), .Y(u2__abc_52138_new_n6469_));
NAND3X1 NAND3X1_84 ( .A(u2__abc_52138_new_n3196_), .B(u2__abc_52138_new_n3424_), .C(u2__abc_52138_new_n6470_), .Y(u2__abc_52138_new_n6471_));
NAND3X1 NAND3X1_85 ( .A(u2__abc_52138_new_n5228_), .B(u2__abc_52138_new_n5272_), .C(u2__abc_52138_new_n5181_), .Y(u2__abc_52138_new_n6476_));
NAND3X1 NAND3X1_86 ( .A(u2__abc_52138_new_n4752_), .B(u2__abc_52138_new_n6481_), .C(u2__abc_52138_new_n6330_), .Y(u2__abc_52138_new_n6482_));
NAND3X1 NAND3X1_87 ( .A(u2__abc_52138_new_n6483_), .B(u2__abc_52138_new_n6484_), .C(u2__abc_52138_new_n6485_), .Y(u2__abc_52138_new_n6486_));
NAND3X1 NAND3X1_88 ( .A(u2__abc_52138_new_n3419_), .B(u2__abc_52138_new_n6489_), .C(u2__abc_52138_new_n6490_), .Y(u2__abc_52138_new_n6491_));
NAND3X1 NAND3X1_89 ( .A(u2__abc_52138_new_n6495_), .B(u2__abc_52138_new_n5547_), .C(u2__abc_52138_new_n6492_), .Y(u2__abc_52138_new_n6496_));
NAND3X1 NAND3X1_9 ( .A(\a[120] ), .B(_abc_65734_new_n1523_), .C(_abc_65734_new_n1524_), .Y(_abc_65734_new_n1525_));
NAND3X1 NAND3X1_90 ( .A(u2__abc_52138_new_n6521_), .B(u2__abc_52138_new_n6522_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6523_));
NAND3X1 NAND3X1_91 ( .A(u2__abc_52138_new_n6530_), .B(u2__abc_52138_new_n6531_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6532_));
NAND3X1 NAND3X1_92 ( .A(u2__abc_52138_new_n6605_), .B(u2__abc_52138_new_n6607_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6608_));
NAND3X1 NAND3X1_93 ( .A(u2__abc_52138_new_n6627_), .B(u2__abc_52138_new_n6628_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6629_));
NAND3X1 NAND3X1_94 ( .A(u2__abc_52138_new_n6675_), .B(u2__abc_52138_new_n6676_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6677_));
NAND3X1 NAND3X1_95 ( .A(u2__abc_52138_new_n6694_), .B(u2__abc_52138_new_n6695_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6696_));
NAND3X1 NAND3X1_96 ( .A(u2__abc_52138_new_n6717_), .B(u2__abc_52138_new_n6718_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6719_));
NAND3X1 NAND3X1_97 ( .A(u2__abc_52138_new_n6739_), .B(u2__abc_52138_new_n6740_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6741_));
NAND3X1 NAND3X1_98 ( .A(u2__abc_52138_new_n6759_), .B(u2__abc_52138_new_n6761_), .C(u2__abc_52138_new_n6757_), .Y(u2__abc_52138_new_n6762_));
NAND3X1 NAND3X1_99 ( .A(u2__abc_52138_new_n6764_), .B(u2__abc_52138_new_n6766_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6767_));
NOR2X1 NOR2X1_1 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1169_), .Y(fracta1_0_));
NOR2X1 NOR2X1_10 ( .A(_abc_65734_new_n1496_), .B(_abc_65734_new_n1484_), .Y(_abc_65734_new_n1497_));
NOR2X1 NOR2X1_100 ( .A(\a[79] ), .B(\a[76] ), .Y(u1__abc_51895_new_n368_));
NOR2X1 NOR2X1_1000 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7301_), .Y(u2__abc_52138_new_n7302_));
NOR2X1 NOR2X1_1001 ( .A(u2__abc_52138_new_n7308_), .B(u2__abc_52138_new_n7298_), .Y(u2__abc_52138_new_n7309_));
NOR2X1 NOR2X1_1002 ( .A(u2__abc_52138_new_n3828_), .B(u2__abc_52138_new_n7314_), .Y(u2__abc_52138_new_n7317_));
NOR2X1 NOR2X1_1003 ( .A(u2__abc_52138_new_n7328_), .B(u2__abc_52138_new_n7326_), .Y(u2__abc_52138_new_n7329_));
NOR2X1 NOR2X1_1004 ( .A(u2__abc_52138_new_n3820_), .B(u2__abc_52138_new_n7326_), .Y(u2__abc_52138_new_n7336_));
NOR2X1 NOR2X1_1005 ( .A(u2__abc_52138_new_n7355_), .B(u2__abc_52138_new_n7313_), .Y(u2__abc_52138_new_n7356_));
NOR2X1 NOR2X1_1006 ( .A(u2__abc_52138_new_n7360_), .B(u2__abc_52138_new_n7356_), .Y(u2__abc_52138_new_n7361_));
NOR2X1 NOR2X1_1007 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7383_), .Y(u2__abc_52138_new_n7384_));
NOR2X1 NOR2X1_1008 ( .A(u2__abc_52138_new_n7401_), .B(u2__abc_52138_new_n7402_), .Y(u2__abc_52138_new_n7403_));
NOR2X1 NOR2X1_1009 ( .A(u2__abc_52138_new_n7399_), .B(u2__abc_52138_new_n7406_), .Y(u2__abc_52138_new_n7409_));
NOR2X1 NOR2X1_101 ( .A(\a[67] ), .B(\a[64] ), .Y(u1__abc_51895_new_n370_));
NOR2X1 NOR2X1_1010 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7418_), .Y(u2__abc_52138_new_n7419_));
NOR2X1 NOR2X1_1011 ( .A(u2__abc_52138_new_n3765_), .B(u2__abc_52138_new_n7426_), .Y(u2__abc_52138_new_n7427_));
NOR2X1 NOR2X1_1012 ( .A(u2__abc_52138_new_n7427_), .B(u2__abc_52138_new_n7429_), .Y(u2__abc_52138_new_n7430_));
NOR2X1 NOR2X1_1013 ( .A(u2_remHi_85_), .B(u2__abc_52138_new_n3766_), .Y(u2__abc_52138_new_n7436_));
NOR2X1 NOR2X1_1014 ( .A(u2__abc_52138_new_n3918_), .B(u2__abc_52138_new_n7436_), .Y(u2__abc_52138_new_n7437_));
NOR2X1 NOR2X1_1015 ( .A(u2__abc_52138_new_n7446_), .B(u2__abc_52138_new_n7449_), .Y(u2__abc_52138_new_n7450_));
NOR2X1 NOR2X1_1016 ( .A(u2__abc_52138_new_n3734_), .B(u2__abc_52138_new_n7451_), .Y(u2__abc_52138_new_n7454_));
NOR2X1 NOR2X1_1017 ( .A(u2__abc_52138_new_n7476_), .B(u2__abc_52138_new_n7475_), .Y(u2__abc_52138_new_n7477_));
NOR2X1 NOR2X1_1018 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7484_), .Y(u2__abc_52138_new_n7485_));
NOR2X1 NOR2X1_1019 ( .A(u2__abc_52138_new_n7491_), .B(u2__abc_52138_new_n7493_), .Y(u2__abc_52138_new_n7494_));
NOR2X1 NOR2X1_102 ( .A(\a[70] ), .B(\a[69] ), .Y(u1__abc_51895_new_n371_));
NOR2X1 NOR2X1_1020 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7505_), .Y(u2__abc_52138_new_n7506_));
NOR2X1 NOR2X1_1021 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7515_), .Y(u2__abc_52138_new_n7516_));
NOR2X1 NOR2X1_1022 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7524_), .Y(u2__abc_52138_new_n7525_));
NOR2X1 NOR2X1_1023 ( .A(u2__abc_52138_new_n3870_), .B(u2__abc_52138_new_n7186_), .Y(u2__abc_52138_new_n7540_));
NOR2X1 NOR2X1_1024 ( .A(u2__abc_52138_new_n7539_), .B(u2__abc_52138_new_n7540_), .Y(u2__abc_52138_new_n7541_));
NOR2X1 NOR2X1_1025 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7552_), .Y(u2__abc_52138_new_n7553_));
NOR2X1 NOR2X1_1026 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7562_), .Y(u2__abc_52138_new_n7563_));
NOR2X1 NOR2X1_1027 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7572_), .Y(u2__abc_52138_new_n7573_));
NOR2X1 NOR2X1_1028 ( .A(u2__abc_52138_new_n7579_), .B(u2__abc_52138_new_n7586_), .Y(u2__abc_52138_new_n7589_));
NOR2X1 NOR2X1_1029 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7598_), .Y(u2__abc_52138_new_n7599_));
NOR2X1 NOR2X1_103 ( .A(u1__abc_51895_new_n369_), .B(u1__abc_51895_new_n372_), .Y(u1__abc_51895_new_n373_));
NOR2X1 NOR2X1_1030 ( .A(u2__abc_52138_new_n3669_), .B(u2__abc_52138_new_n7606_), .Y(u2__abc_52138_new_n7607_));
NOR2X1 NOR2X1_1031 ( .A(u2__abc_52138_new_n7607_), .B(u2__abc_52138_new_n7609_), .Y(u2__abc_52138_new_n7610_));
NOR2X1 NOR2X1_1032 ( .A(u2__abc_52138_new_n3948_), .B(u2__abc_52138_new_n3947_), .Y(u2__abc_52138_new_n7626_));
NOR2X1 NOR2X1_1033 ( .A(u2__abc_52138_new_n3616_), .B(u2__abc_52138_new_n7631_), .Y(u2__abc_52138_new_n7634_));
NOR2X1 NOR2X1_1034 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7644_), .Y(u2__abc_52138_new_n7645_));
NOR2X1 NOR2X1_1035 ( .A(u2__abc_52138_new_n3601_), .B(u2__abc_52138_new_n7652_), .Y(u2__abc_52138_new_n7653_));
NOR2X1 NOR2X1_1036 ( .A(u2__abc_52138_new_n7653_), .B(u2__abc_52138_new_n7655_), .Y(u2__abc_52138_new_n7656_));
NOR2X1 NOR2X1_1037 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7663_), .Y(u2__abc_52138_new_n7664_));
NOR2X1 NOR2X1_1038 ( .A(u2__abc_52138_new_n3598_), .B(u2__abc_52138_new_n3606_), .Y(u2__abc_52138_new_n7671_));
NOR2X1 NOR2X1_1039 ( .A(u2__abc_52138_new_n3958_), .B(u2__abc_52138_new_n7671_), .Y(u2__abc_52138_new_n7672_));
NOR2X1 NOR2X1_104 ( .A(u2__abc_52138_new_n2962_), .B(u2__abc_52138_new_n2963_), .Y(u2__abc_52138_new_n2964_));
NOR2X1 NOR2X1_1040 ( .A(u2__abc_52138_new_n7673_), .B(u2__abc_52138_new_n7674_), .Y(u2__abc_52138_new_n7676_));
NOR2X1 NOR2X1_1041 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7686_), .Y(u2__abc_52138_new_n7687_));
NOR2X1 NOR2X1_1042 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7696_), .Y(u2__abc_52138_new_n7697_));
NOR2X1 NOR2X1_1043 ( .A(u2__abc_52138_new_n3966_), .B(u2__abc_52138_new_n7703_), .Y(u2__abc_52138_new_n7704_));
NOR2X1 NOR2X1_1044 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7722_), .Y(u2__abc_52138_new_n7723_));
NOR2X1 NOR2X1_1045 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7731_), .Y(u2__abc_52138_new_n7732_));
NOR2X1 NOR2X1_1046 ( .A(u2__abc_52138_new_n3565_), .B(u2__abc_52138_new_n7739_), .Y(u2__abc_52138_new_n7740_));
NOR2X1 NOR2X1_1047 ( .A(u2__abc_52138_new_n7740_), .B(u2__abc_52138_new_n7742_), .Y(u2__abc_52138_new_n7743_));
NOR2X1 NOR2X1_1048 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7750_), .Y(u2__abc_52138_new_n7751_));
NOR2X1 NOR2X1_1049 ( .A(u2__abc_52138_new_n3562_), .B(u2__abc_52138_new_n3570_), .Y(u2__abc_52138_new_n7758_));
NOR2X1 NOR2X1_105 ( .A(u2__abc_52138_new_n2968_), .B(u2__abc_52138_new_n2970_), .Y(u2__abc_52138_new_n2971_));
NOR2X1 NOR2X1_1050 ( .A(u2__abc_52138_new_n3975_), .B(u2__abc_52138_new_n7758_), .Y(u2__abc_52138_new_n7759_));
NOR2X1 NOR2X1_1051 ( .A(u2__abc_52138_new_n3592_), .B(u2__abc_52138_new_n7761_), .Y(u2__abc_52138_new_n7762_));
NOR2X1 NOR2X1_1052 ( .A(u2__abc_52138_new_n7762_), .B(u2__abc_52138_new_n7764_), .Y(u2__abc_52138_new_n7765_));
NOR2X1 NOR2X1_1053 ( .A(u2__abc_52138_new_n3577_), .B(u2__abc_52138_new_n7782_), .Y(u2__abc_52138_new_n7784_));
NOR2X1 NOR2X1_1054 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7784_), .Y(u2__abc_52138_new_n7785_));
NOR2X1 NOR2X1_1055 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7794_), .Y(u2__abc_52138_new_n7795_));
NOR2X1 NOR2X1_1056 ( .A(u2__abc_52138_new_n7792_), .B(u2__abc_52138_new_n7802_), .Y(u2__abc_52138_new_n7803_));
NOR2X1 NOR2X1_1057 ( .A(u2__abc_52138_new_n3595_), .B(u2__abc_52138_new_n7729_), .Y(u2__abc_52138_new_n7809_));
NOR2X1 NOR2X1_1058 ( .A(u2__abc_52138_new_n7808_), .B(u2__abc_52138_new_n7809_), .Y(u2__abc_52138_new_n7810_));
NOR2X1 NOR2X1_1059 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7842_), .Y(u2__abc_52138_new_n7843_));
NOR2X1 NOR2X1_106 ( .A(u2_cnt_3_), .B(u2_cnt_2_), .Y(u2__abc_52138_new_n2972_));
NOR2X1 NOR2X1_1060 ( .A(u2__abc_52138_new_n7854_), .B(u2__abc_52138_new_n7853_), .Y(u2__abc_52138_new_n7855_));
NOR2X1 NOR2X1_1061 ( .A(u2__abc_52138_new_n7856_), .B(u2__abc_52138_new_n7855_), .Y(u2__abc_52138_new_n7857_));
NOR2X1 NOR2X1_1062 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7864_), .Y(u2__abc_52138_new_n7865_));
NOR2X1 NOR2X1_1063 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7873_), .Y(u2__abc_52138_new_n7874_));
NOR2X1 NOR2X1_1064 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7881_), .Y(u2__abc_52138_new_n7882_));
NOR2X1 NOR2X1_1065 ( .A(u2__abc_52138_new_n7888_), .B(u2__abc_52138_new_n7186_), .Y(u2__abc_52138_new_n7889_));
NOR2X1 NOR2X1_1066 ( .A(u2__abc_52138_new_n7899_), .B(u2__abc_52138_new_n7889_), .Y(u2__abc_52138_new_n7901_));
NOR2X1 NOR2X1_1067 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7921_), .Y(u2__abc_52138_new_n7922_));
NOR2X1 NOR2X1_1068 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7931_), .Y(u2__abc_52138_new_n7932_));
NOR2X1 NOR2X1_1069 ( .A(u2__abc_52138_new_n7938_), .B(u2__abc_52138_new_n7928_), .Y(u2__abc_52138_new_n7939_));
NOR2X1 NOR2X1_107 ( .A(u2_cnt_0_), .B(u2__abc_52138_new_n2974_), .Y(u2__abc_52138_new_n2975_));
NOR2X1 NOR2X1_1070 ( .A(u2__abc_52138_new_n4749_), .B(u2__abc_52138_new_n7943_), .Y(u2__abc_52138_new_n7946_));
NOR2X1 NOR2X1_1071 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7955_), .Y(u2__abc_52138_new_n7956_));
NOR2X1 NOR2X1_1072 ( .A(u2__abc_52138_new_n4737_), .B(u2__abc_52138_new_n7963_), .Y(u2__abc_52138_new_n7964_));
NOR2X1 NOR2X1_1073 ( .A(u2__abc_52138_new_n7964_), .B(u2__abc_52138_new_n7966_), .Y(u2__abc_52138_new_n7967_));
NOR2X1 NOR2X1_1074 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7974_), .Y(u2__abc_52138_new_n7975_));
NOR2X1 NOR2X1_1075 ( .A(u2__abc_52138_new_n4750_), .B(u2__abc_52138_new_n7942_), .Y(u2__abc_52138_new_n7982_));
NOR2X1 NOR2X1_1076 ( .A(u2__abc_52138_new_n7986_), .B(u2__abc_52138_new_n7982_), .Y(u2__abc_52138_new_n7987_));
NOR2X1 NOR2X1_1077 ( .A(u2__abc_52138_new_n7981_), .B(u2__abc_52138_new_n7988_), .Y(u2__abc_52138_new_n7991_));
NOR2X1 NOR2X1_1078 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8000_), .Y(u2__abc_52138_new_n8001_));
NOR2X1 NOR2X1_1079 ( .A(u2__abc_52138_new_n4670_), .B(u2__abc_52138_new_n8008_), .Y(u2__abc_52138_new_n8009_));
NOR2X1 NOR2X1_108 ( .A(u2__abc_52138_new_n2973_), .B(u2__abc_52138_new_n2976_), .Y(u2__abc_52138_new_n2977_));
NOR2X1 NOR2X1_1080 ( .A(sqrto_136_), .B(u2__abc_52138_new_n4668_), .Y(u2__abc_52138_new_n8010_));
NOR2X1 NOR2X1_1081 ( .A(u2_remHi_136_), .B(u2__abc_52138_new_n4666_), .Y(u2__abc_52138_new_n8011_));
NOR2X1 NOR2X1_1082 ( .A(u2__abc_52138_new_n8009_), .B(u2__abc_52138_new_n8013_), .Y(u2__abc_52138_new_n8014_));
NOR2X1 NOR2X1_1083 ( .A(u2_remHi_137_), .B(u2__abc_52138_new_n4671_), .Y(u2__abc_52138_new_n8020_));
NOR2X1 NOR2X1_1084 ( .A(u2__abc_52138_new_n4789_), .B(u2__abc_52138_new_n8020_), .Y(u2__abc_52138_new_n8021_));
NOR2X1 NOR2X1_1085 ( .A(u2__abc_52138_new_n4709_), .B(u2__abc_52138_new_n8034_), .Y(u2__abc_52138_new_n8035_));
NOR2X1 NOR2X1_1086 ( .A(u2__abc_52138_new_n8035_), .B(u2__abc_52138_new_n8037_), .Y(u2__abc_52138_new_n8038_));
NOR2X1 NOR2X1_1087 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8045_), .Y(u2__abc_52138_new_n8046_));
NOR2X1 NOR2X1_1088 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8054_), .Y(u2__abc_52138_new_n8055_));
NOR2X1 NOR2X1_1089 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8062_), .Y(u2__abc_52138_new_n8063_));
NOR2X1 NOR2X1_109 ( .A(rst), .B(u2__abc_52138_new_n2966_), .Y(u2__abc_52138_new_n2981_));
NOR2X1 NOR2X1_1090 ( .A(u2__abc_52138_new_n8069_), .B(u2__abc_52138_new_n8070_), .Y(u2__abc_52138_new_n8071_));
NOR2X1 NOR2X1_1091 ( .A(u2__abc_52138_new_n4712_), .B(u2__abc_52138_new_n4751_), .Y(u2__abc_52138_new_n8079_));
NOR2X1 NOR2X1_1092 ( .A(u2__abc_52138_new_n4662_), .B(u2__abc_52138_new_n8081_), .Y(u2__abc_52138_new_n8084_));
NOR2X1 NOR2X1_1093 ( .A(u2__abc_52138_new_n4653_), .B(u2__abc_52138_new_n4656_), .Y(u2__abc_52138_new_n8092_));
NOR2X1 NOR2X1_1094 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8094_), .Y(u2__abc_52138_new_n8095_));
NOR2X1 NOR2X1_1095 ( .A(u2__abc_52138_new_n8101_), .B(u2__abc_52138_new_n8102_), .Y(u2__abc_52138_new_n8103_));
NOR2X1 NOR2X1_1096 ( .A(u2__abc_52138_new_n8103_), .B(u2__abc_52138_new_n8105_), .Y(u2__abc_52138_new_n8106_));
NOR2X1 NOR2X1_1097 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8114_), .Y(u2__abc_52138_new_n8115_));
NOR2X1 NOR2X1_1098 ( .A(u2__abc_52138_new_n4639_), .B(u2__abc_52138_new_n8122_), .Y(u2__abc_52138_new_n8123_));
NOR2X1 NOR2X1_1099 ( .A(u2__abc_52138_new_n8123_), .B(u2__abc_52138_new_n8125_), .Y(u2__abc_52138_new_n8126_));
NOR2X1 NOR2X1_11 ( .A(_abc_65734_new_n1503_), .B(_abc_65734_new_n1495_), .Y(_abc_65734_new_n1504_));
NOR2X1 NOR2X1_110 ( .A(rst), .B(ce), .Y(u2__abc_52138_new_n2982_));
NOR2X1 NOR2X1_1100 ( .A(sqrto_148_), .B(u2__abc_52138_new_n4621_), .Y(u2__abc_52138_new_n8141_));
NOR2X1 NOR2X1_1101 ( .A(u2__abc_52138_new_n8141_), .B(u2__abc_52138_new_n4810_), .Y(u2__abc_52138_new_n8142_));
NOR2X1 NOR2X1_1102 ( .A(u2__abc_52138_new_n8142_), .B(u2__abc_52138_new_n8144_), .Y(u2__abc_52138_new_n8146_));
NOR2X1 NOR2X1_1103 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8146_), .Y(u2__abc_52138_new_n8147_));
NOR2X1 NOR2X1_1104 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8155_), .Y(u2__abc_52138_new_n8156_));
NOR2X1 NOR2X1_1105 ( .A(u2__abc_52138_new_n4636_), .B(u2__abc_52138_new_n4634_), .Y(u2__abc_52138_new_n8163_));
NOR2X1 NOR2X1_1106 ( .A(u2__abc_52138_new_n8170_), .B(u2__abc_52138_new_n8171_), .Y(u2__abc_52138_new_n8173_));
NOR2X1 NOR2X1_1107 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8182_), .Y(u2__abc_52138_new_n8183_));
NOR2X1 NOR2X1_1108 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8192_), .Y(u2__abc_52138_new_n8193_));
NOR2X1 NOR2X1_1109 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8200_), .Y(u2__abc_52138_new_n8201_));
NOR2X1 NOR2X1_111 ( .A(ld), .B(u2__abc_52138_new_n2963_), .Y(u2__abc_52138_new_n2983_));
NOR2X1 NOR2X1_1110 ( .A(u2__abc_52138_new_n8213_), .B(u2__abc_52138_new_n8212_), .Y(u2__abc_52138_new_n8214_));
NOR2X1 NOR2X1_1111 ( .A(u2__abc_52138_new_n8215_), .B(u2__abc_52138_new_n8214_), .Y(u2__abc_52138_new_n8216_));
NOR2X1 NOR2X1_1112 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8222_), .Y(u2__abc_52138_new_n8223_));
NOR2X1 NOR2X1_1113 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8232_), .Y(u2__abc_52138_new_n8233_));
NOR2X1 NOR2X1_1114 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8240_), .Y(u2__abc_52138_new_n8241_));
NOR2X1 NOR2X1_1115 ( .A(u2__abc_52138_new_n4665_), .B(u2__abc_52138_new_n8078_), .Y(u2__abc_52138_new_n8248_));
NOR2X1 NOR2X1_1116 ( .A(u2__abc_52138_new_n4545_), .B(u2__abc_52138_new_n8257_), .Y(u2__abc_52138_new_n8258_));
NOR2X1 NOR2X1_1117 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8261_), .Y(u2__abc_52138_new_n8262_));
NOR2X1 NOR2X1_1118 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8269_), .Y(u2__abc_52138_new_n8270_));
NOR2X1 NOR2X1_1119 ( .A(u2__abc_52138_new_n4529_), .B(u2__abc_52138_new_n8277_), .Y(u2__abc_52138_new_n8278_));
NOR2X1 NOR2X1_112 ( .A(done), .B(u2__abc_52138_new_n2983_), .Y(u2__abc_52138_new_n2984_));
NOR2X1 NOR2X1_1120 ( .A(sqrto_160_), .B(u2__abc_52138_new_n4527_), .Y(u2__abc_52138_new_n8279_));
NOR2X1 NOR2X1_1121 ( .A(u2_remHi_160_), .B(u2__abc_52138_new_n4525_), .Y(u2__abc_52138_new_n8280_));
NOR2X1 NOR2X1_1122 ( .A(u2__abc_52138_new_n8278_), .B(u2__abc_52138_new_n8282_), .Y(u2__abc_52138_new_n8283_));
NOR2X1 NOR2X1_1123 ( .A(u2_remHi_161_), .B(u2__abc_52138_new_n4530_), .Y(u2__abc_52138_new_n8289_));
NOR2X1 NOR2X1_1124 ( .A(u2__abc_52138_new_n4833_), .B(u2__abc_52138_new_n8289_), .Y(u2__abc_52138_new_n8290_));
NOR2X1 NOR2X1_1125 ( .A(u2__abc_52138_new_n4568_), .B(u2__abc_52138_new_n8302_), .Y(u2__abc_52138_new_n8303_));
NOR2X1 NOR2X1_1126 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8324_), .Y(u2__abc_52138_new_n8325_));
NOR2X1 NOR2X1_1127 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8333_), .Y(u2__abc_52138_new_n8334_));
NOR2X1 NOR2X1_1128 ( .A(u2__abc_52138_new_n4521_), .B(u2__abc_52138_new_n8345_), .Y(u2__abc_52138_new_n8346_));
NOR2X1 NOR2X1_1129 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8356_), .Y(u2__abc_52138_new_n8357_));
NOR2X1 NOR2X1_113 ( .A(u2__abc_52138_new_n2968_), .B(u2__abc_52138_new_n2973_), .Y(u2__abc_52138_new_n2988_));
NOR2X1 NOR2X1_1130 ( .A(u2__abc_52138_new_n4505_), .B(u2__abc_52138_new_n8364_), .Y(u2__abc_52138_new_n8365_));
NOR2X1 NOR2X1_1131 ( .A(u2__abc_52138_new_n8365_), .B(u2__abc_52138_new_n8367_), .Y(u2__abc_52138_new_n8368_));
NOR2X1 NOR2X1_1132 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8375_), .Y(u2__abc_52138_new_n8376_));
NOR2X1 NOR2X1_1133 ( .A(u2__abc_52138_new_n4498_), .B(u2__abc_52138_new_n8383_), .Y(u2__abc_52138_new_n8384_));
NOR2X1 NOR2X1_1134 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8394_), .Y(u2__abc_52138_new_n8395_));
NOR2X1 NOR2X1_1135 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8403_), .Y(u2__abc_52138_new_n8404_));
NOR2X1 NOR2X1_1136 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8411_), .Y(u2__abc_52138_new_n8412_));
NOR2X1 NOR2X1_1137 ( .A(u2__abc_52138_new_n4571_), .B(u2__abc_52138_new_n8257_), .Y(u2__abc_52138_new_n8430_));
NOR2X1 NOR2X1_1138 ( .A(u2__abc_52138_new_n8429_), .B(u2__abc_52138_new_n8430_), .Y(u2__abc_52138_new_n8432_));
NOR2X1 NOR2X1_1139 ( .A(u2__abc_52138_new_n8448_), .B(u2__abc_52138_new_n8453_), .Y(u2__abc_52138_new_n8455_));
NOR2X1 NOR2X1_114 ( .A(u2__abc_52138_new_n2970_), .B(u2__abc_52138_new_n2976_), .Y(u2__abc_52138_new_n2989_));
NOR2X1 NOR2X1_1140 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8455_), .Y(u2__abc_52138_new_n8456_));
NOR2X1 NOR2X1_1141 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8464_), .Y(u2__abc_52138_new_n8465_));
NOR2X1 NOR2X1_1142 ( .A(u2__abc_52138_new_n4449_), .B(u2__abc_52138_new_n8474_), .Y(u2__abc_52138_new_n8475_));
NOR2X1 NOR2X1_1143 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8485_), .Y(u2__abc_52138_new_n8486_));
NOR2X1 NOR2X1_1144 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8494_), .Y(u2__abc_52138_new_n8495_));
NOR2X1 NOR2X1_1145 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8502_), .Y(u2__abc_52138_new_n8503_));
NOR2X1 NOR2X1_1146 ( .A(u2__abc_52138_new_n4430_), .B(u2__abc_52138_new_n4438_), .Y(u2__abc_52138_new_n8510_));
NOR2X1 NOR2X1_1147 ( .A(u2__abc_52138_new_n4862_), .B(u2__abc_52138_new_n8510_), .Y(u2__abc_52138_new_n8511_));
NOR2X1 NOR2X1_1148 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8525_), .Y(u2__abc_52138_new_n8526_));
NOR2X1 NOR2X1_1149 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8536_), .Y(u2__abc_52138_new_n8537_));
NOR2X1 NOR2X1_115 ( .A(u2_remHi_448_), .B(u2__abc_52138_new_n2997_), .Y(u2__abc_52138_new_n2998_));
NOR2X1 NOR2X1_1150 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8545_), .Y(u2__abc_52138_new_n8546_));
NOR2X1 NOR2X1_1151 ( .A(u2__abc_52138_new_n4425_), .B(u2__abc_52138_new_n8555_), .Y(u2__abc_52138_new_n8556_));
NOR2X1 NOR2X1_1152 ( .A(u2__abc_52138_new_n8556_), .B(u2__abc_52138_new_n8558_), .Y(u2__abc_52138_new_n8559_));
NOR2X1 NOR2X1_1153 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8566_), .Y(u2__abc_52138_new_n8567_));
NOR2X1 NOR2X1_1154 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8575_), .Y(u2__abc_52138_new_n8576_));
NOR2X1 NOR2X1_1155 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8583_), .Y(u2__abc_52138_new_n8584_));
NOR2X1 NOR2X1_1156 ( .A(u2__abc_52138_new_n8591_), .B(u2__abc_52138_new_n8513_), .Y(u2__abc_52138_new_n8592_));
NOR2X1 NOR2X1_1157 ( .A(u2__abc_52138_new_n4427_), .B(u2__abc_52138_new_n8553_), .Y(u2__abc_52138_new_n8593_));
NOR2X1 NOR2X1_1158 ( .A(u2__abc_52138_new_n8592_), .B(u2__abc_52138_new_n8601_), .Y(u2__abc_52138_new_n8602_));
NOR2X1 NOR2X1_1159 ( .A(u2__abc_52138_new_n4368_), .B(u2__abc_52138_new_n8604_), .Y(u2__abc_52138_new_n8605_));
NOR2X1 NOR2X1_116 ( .A(u2__abc_52138_new_n2998_), .B(u2__abc_52138_new_n3001_), .Y(u2__abc_52138_new_n3002_));
NOR2X1 NOR2X1_1160 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8608_), .Y(u2__abc_52138_new_n8609_));
NOR2X1 NOR2X1_1161 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8616_), .Y(u2__abc_52138_new_n8617_));
NOR2X1 NOR2X1_1162 ( .A(u2__abc_52138_new_n4351_), .B(u2__abc_52138_new_n8644_), .Y(u2__abc_52138_new_n8645_));
NOR2X1 NOR2X1_1163 ( .A(u2__abc_52138_new_n8645_), .B(u2__abc_52138_new_n8647_), .Y(u2__abc_52138_new_n8648_));
NOR2X1 NOR2X1_1164 ( .A(sqrto_196_), .B(u2__abc_52138_new_n4333_), .Y(u2__abc_52138_new_n8663_));
NOR2X1 NOR2X1_1165 ( .A(u2_remHi_196_), .B(u2__abc_52138_new_n4331_), .Y(u2__abc_52138_new_n8664_));
NOR2X1 NOR2X1_1166 ( .A(u2__abc_52138_new_n8663_), .B(u2__abc_52138_new_n8664_), .Y(u2__abc_52138_new_n8665_));
NOR2X1 NOR2X1_1167 ( .A(u2__abc_52138_new_n8665_), .B(u2__abc_52138_new_n8667_), .Y(u2__abc_52138_new_n8669_));
NOR2X1 NOR2X1_1168 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8669_), .Y(u2__abc_52138_new_n8670_));
NOR2X1 NOR2X1_1169 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8678_), .Y(u2__abc_52138_new_n8679_));
NOR2X1 NOR2X1_117 ( .A(u2_o_447_), .B(u2__abc_52138_new_n3003_), .Y(u2__abc_52138_new_n3004_));
NOR2X1 NOR2X1_1170 ( .A(u2__abc_52138_new_n4378_), .B(u2__abc_52138_new_n8604_), .Y(u2__abc_52138_new_n8691_));
NOR2X1 NOR2X1_1171 ( .A(u2__abc_52138_new_n8690_), .B(u2__abc_52138_new_n8691_), .Y(u2__abc_52138_new_n8693_));
NOR2X1 NOR2X1_1172 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8702_), .Y(u2__abc_52138_new_n8703_));
NOR2X1 NOR2X1_1173 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8712_), .Y(u2__abc_52138_new_n8713_));
NOR2X1 NOR2X1_1174 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8720_), .Y(u2__abc_52138_new_n8721_));
NOR2X1 NOR2X1_1175 ( .A(u2__abc_52138_new_n8733_), .B(u2__abc_52138_new_n8732_), .Y(u2__abc_52138_new_n8734_));
NOR2X1 NOR2X1_1176 ( .A(u2__abc_52138_new_n8735_), .B(u2__abc_52138_new_n8734_), .Y(u2__abc_52138_new_n8736_));
NOR2X1 NOR2X1_1177 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8742_), .Y(u2__abc_52138_new_n8743_));
NOR2X1 NOR2X1_1178 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8752_), .Y(u2__abc_52138_new_n8753_));
NOR2X1 NOR2X1_1179 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8760_), .Y(u2__abc_52138_new_n8761_));
NOR2X1 NOR2X1_118 ( .A(u2_remHi_447_), .B(u2__abc_52138_new_n3005_), .Y(u2__abc_52138_new_n3006_));
NOR2X1 NOR2X1_1180 ( .A(u2__abc_52138_new_n4311_), .B(u2__abc_52138_new_n4329_), .Y(u2__abc_52138_new_n8768_));
NOR2X1 NOR2X1_1181 ( .A(u2__abc_52138_new_n8774_), .B(u2__abc_52138_new_n8775_), .Y(u2__abc_52138_new_n8777_));
NOR2X1 NOR2X1_1182 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8786_), .Y(u2__abc_52138_new_n8787_));
NOR2X1 NOR2X1_1183 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8795_), .Y(u2__abc_52138_new_n8796_));
NOR2X1 NOR2X1_1184 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8804_), .Y(u2__abc_52138_new_n8805_));
NOR2X1 NOR2X1_1185 ( .A(u2__abc_52138_new_n4245_), .B(u2__abc_52138_new_n4250_), .Y(u2__abc_52138_new_n8811_));
NOR2X1 NOR2X1_1186 ( .A(u2__abc_52138_new_n4284_), .B(u2__abc_52138_new_n8816_), .Y(u2__abc_52138_new_n8818_));
NOR2X1 NOR2X1_1187 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8818_), .Y(u2__abc_52138_new_n8819_));
NOR2X1 NOR2X1_1188 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8844_), .Y(u2__abc_52138_new_n8845_));
NOR2X1 NOR2X1_1189 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8868_), .Y(u2__abc_52138_new_n8869_));
NOR2X1 NOR2X1_119 ( .A(u2__abc_52138_new_n3004_), .B(u2__abc_52138_new_n3006_), .Y(u2__abc_52138_new_n3007_));
NOR2X1 NOR2X1_1190 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8878_), .Y(u2__abc_52138_new_n8879_));
NOR2X1 NOR2X1_1191 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8887_), .Y(u2__abc_52138_new_n8888_));
NOR2X1 NOR2X1_1192 ( .A(u2__abc_52138_new_n8894_), .B(u2__abc_52138_new_n8899_), .Y(u2__abc_52138_new_n8900_));
NOR2X1 NOR2X1_1193 ( .A(u2__abc_52138_new_n8901_), .B(u2__abc_52138_new_n8900_), .Y(u2__abc_52138_new_n8902_));
NOR2X1 NOR2X1_1194 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8909_), .Y(u2__abc_52138_new_n8910_));
NOR2X1 NOR2X1_1195 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8919_), .Y(u2__abc_52138_new_n8920_));
NOR2X1 NOR2X1_1196 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8928_), .Y(u2__abc_52138_new_n8929_));
NOR2X1 NOR2X1_1197 ( .A(u2__abc_52138_new_n4240_), .B(u2__abc_52138_new_n8857_), .Y(u2__abc_52138_new_n8938_));
NOR2X1 NOR2X1_1198 ( .A(u2__abc_52138_new_n8940_), .B(u2__abc_52138_new_n8938_), .Y(u2__abc_52138_new_n8941_));
NOR2X1 NOR2X1_1199 ( .A(u2__abc_52138_new_n4380_), .B(u2__abc_52138_new_n8604_), .Y(u2__abc_52138_new_n8943_));
NOR2X1 NOR2X1_12 ( .A(_abc_65734_new_n1505_), .B(_abc_65734_new_n1506_), .Y(_abc_65734_new_n1507_));
NOR2X1 NOR2X1_120 ( .A(u2_o_446_), .B(u2__abc_52138_new_n3008_), .Y(u2__abc_52138_new_n3009_));
NOR2X1 NOR2X1_1200 ( .A(u2__abc_52138_new_n8942_), .B(u2__abc_52138_new_n8943_), .Y(u2__abc_52138_new_n8946_));
NOR2X1 NOR2X1_1201 ( .A(u2__abc_52138_new_n8945_), .B(u2__abc_52138_new_n8948_), .Y(u2__abc_52138_new_n8949_));
NOR2X1 NOR2X1_1202 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8956_), .Y(u2__abc_52138_new_n8957_));
NOR2X1 NOR2X1_1203 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8965_), .Y(u2__abc_52138_new_n8966_));
NOR2X1 NOR2X1_1204 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8973_), .Y(u2__abc_52138_new_n8974_));
NOR2X1 NOR2X1_1205 ( .A(u2__abc_52138_new_n8985_), .B(u2__abc_52138_new_n8984_), .Y(u2__abc_52138_new_n8986_));
NOR2X1 NOR2X1_1206 ( .A(u2__abc_52138_new_n8987_), .B(u2__abc_52138_new_n8986_), .Y(u2__abc_52138_new_n8988_));
NOR2X1 NOR2X1_1207 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n8994_), .Y(u2__abc_52138_new_n8995_));
NOR2X1 NOR2X1_1208 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9004_), .Y(u2__abc_52138_new_n9005_));
NOR2X1 NOR2X1_1209 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9012_), .Y(u2__abc_52138_new_n9013_));
NOR2X1 NOR2X1_121 ( .A(u2_remHi_446_), .B(u2__abc_52138_new_n3010_), .Y(u2__abc_52138_new_n3011_));
NOR2X1 NOR2X1_1210 ( .A(u2__abc_52138_new_n4142_), .B(u2__abc_52138_new_n9024_), .Y(u2__abc_52138_new_n9026_));
NOR2X1 NOR2X1_1211 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9026_), .Y(u2__abc_52138_new_n9027_));
NOR2X1 NOR2X1_1212 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9036_), .Y(u2__abc_52138_new_n9037_));
NOR2X1 NOR2X1_1213 ( .A(u2__abc_52138_new_n4127_), .B(u2__abc_52138_new_n9043_), .Y(u2__abc_52138_new_n9044_));
NOR2X1 NOR2X1_1214 ( .A(u2__abc_52138_new_n9044_), .B(u2__abc_52138_new_n9046_), .Y(u2__abc_52138_new_n9047_));
NOR2X1 NOR2X1_1215 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9054_), .Y(u2__abc_52138_new_n9055_));
NOR2X1 NOR2X1_1216 ( .A(u2__abc_52138_new_n4119_), .B(u2__abc_52138_new_n9062_), .Y(u2__abc_52138_new_n9063_));
NOR2X1 NOR2X1_1217 ( .A(u2__abc_52138_new_n9063_), .B(u2__abc_52138_new_n9065_), .Y(u2__abc_52138_new_n9066_));
NOR2X1 NOR2X1_1218 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9073_), .Y(u2__abc_52138_new_n9074_));
NOR2X1 NOR2X1_1219 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9082_), .Y(u2__abc_52138_new_n9083_));
NOR2X1 NOR2X1_122 ( .A(u2__abc_52138_new_n3009_), .B(u2__abc_52138_new_n3011_), .Y(u2__abc_52138_new_n3012_));
NOR2X1 NOR2X1_1220 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9090_), .Y(u2__abc_52138_new_n9091_));
NOR2X1 NOR2X1_1221 ( .A(u2__abc_52138_new_n9097_), .B(u2__abc_52138_new_n9104_), .Y(u2__abc_52138_new_n9105_));
NOR2X1 NOR2X1_1222 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9108_), .Y(u2__abc_52138_new_n9109_));
NOR2X1 NOR2X1_1223 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9117_), .Y(u2__abc_52138_new_n9118_));
NOR2X1 NOR2X1_1224 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9127_), .Y(u2__abc_52138_new_n9128_));
NOR2X1 NOR2X1_1225 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9136_), .Y(u2__abc_52138_new_n9137_));
NOR2X1 NOR2X1_1226 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9148_), .Y(u2__abc_52138_new_n9149_));
NOR2X1 NOR2X1_1227 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9175_), .Y(u2__abc_52138_new_n9176_));
NOR2X1 NOR2X1_1228 ( .A(u2__abc_52138_new_n4097_), .B(u2__abc_52138_new_n9115_), .Y(u2__abc_52138_new_n9187_));
NOR2X1 NOR2X1_1229 ( .A(u2__abc_52138_new_n9186_), .B(u2__abc_52138_new_n9187_), .Y(u2__abc_52138_new_n9188_));
NOR2X1 NOR2X1_123 ( .A(u2__abc_52138_new_n3021_), .B(u2__abc_52138_new_n3032_), .Y(u2__abc_52138_new_n3033_));
NOR2X1 NOR2X1_1230 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9198_), .Y(u2__abc_52138_new_n9199_));
NOR2X1 NOR2X1_1231 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9219_), .Y(u2__abc_52138_new_n9220_));
NOR2X1 NOR2X1_1232 ( .A(u2__abc_52138_new_n9232_), .B(u2__abc_52138_new_n9231_), .Y(u2__abc_52138_new_n9233_));
NOR2X1 NOR2X1_1233 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9240_), .Y(u2__abc_52138_new_n9241_));
NOR2X1 NOR2X1_1234 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9257_), .Y(u2__abc_52138_new_n9258_));
NOR2X1 NOR2X1_1235 ( .A(u2_remHi_254_), .B(u2__abc_52138_new_n5687_), .Y(u2__abc_52138_new_n9264_));
NOR2X1 NOR2X1_1236 ( .A(u2_o_254_), .B(u2__abc_52138_new_n5691_), .Y(u2__abc_52138_new_n9265_));
NOR2X1 NOR2X1_1237 ( .A(u2__abc_52138_new_n9264_), .B(u2__abc_52138_new_n9265_), .Y(u2__abc_52138_new_n9266_));
NOR2X1 NOR2X1_1238 ( .A(u2__abc_52138_new_n9324_), .B(u2__abc_52138_new_n9323_), .Y(u2__abc_52138_new_n9325_));
NOR2X1 NOR2X1_1239 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9332_), .Y(u2__abc_52138_new_n9333_));
NOR2X1 NOR2X1_124 ( .A(u2__abc_52138_new_n3039_), .B(u2__abc_52138_new_n3050_), .Y(u2__abc_52138_new_n3051_));
NOR2X1 NOR2X1_1240 ( .A(u2__abc_52138_new_n9343_), .B(u2__abc_52138_new_n9344_), .Y(u2__abc_52138_new_n9345_));
NOR2X1 NOR2X1_1241 ( .A(u2__abc_52138_new_n5710_), .B(u2__abc_52138_new_n9343_), .Y(u2__abc_52138_new_n9351_));
NOR2X1 NOR2X1_1242 ( .A(u2__abc_52138_new_n5664_), .B(u2__abc_52138_new_n5669_), .Y(u2__abc_52138_new_n9400_));
NOR2X1 NOR2X1_1243 ( .A(u2__abc_52138_new_n9402_), .B(u2__abc_52138_new_n9403_), .Y(u2__abc_52138_new_n9404_));
NOR2X1 NOR2X1_1244 ( .A(u2__abc_52138_new_n5652_), .B(u2__abc_52138_new_n9402_), .Y(u2__abc_52138_new_n9410_));
NOR2X1 NOR2X1_1245 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9411_), .Y(u2__abc_52138_new_n9412_));
NOR2X1 NOR2X1_1246 ( .A(u2__abc_52138_new_n5733_), .B(u2__abc_52138_new_n9288_), .Y(u2__abc_52138_new_n9445_));
NOR2X1 NOR2X1_1247 ( .A(u2__abc_52138_new_n9444_), .B(u2__abc_52138_new_n9445_), .Y(u2__abc_52138_new_n9448_));
NOR2X1 NOR2X1_1248 ( .A(u2__abc_52138_new_n9447_), .B(u2__abc_52138_new_n9450_), .Y(u2__abc_52138_new_n9451_));
NOR2X1 NOR2X1_1249 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9458_), .Y(u2__abc_52138_new_n9459_));
NOR2X1 NOR2X1_125 ( .A(u2__abc_52138_new_n3058_), .B(u2__abc_52138_new_n3064_), .Y(u2__abc_52138_new_n3065_));
NOR2X1 NOR2X1_1250 ( .A(u2__abc_52138_new_n9493_), .B(u2__abc_52138_new_n9492_), .Y(u2__abc_52138_new_n9494_));
NOR2X1 NOR2X1_1251 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9501_), .Y(u2__abc_52138_new_n9502_));
NOR2X1 NOR2X1_1252 ( .A(u2__abc_52138_new_n9535_), .B(u2__abc_52138_new_n9534_), .Y(u2__abc_52138_new_n9536_));
NOR2X1 NOR2X1_1253 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9543_), .Y(u2__abc_52138_new_n9544_));
NOR2X1 NOR2X1_1254 ( .A(u2__abc_52138_new_n9577_), .B(u2__abc_52138_new_n9576_), .Y(u2__abc_52138_new_n9578_));
NOR2X1 NOR2X1_1255 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9586_), .Y(u2__abc_52138_new_n9587_));
NOR2X1 NOR2X1_1256 ( .A(u2__abc_52138_new_n9619_), .B(u2__abc_52138_new_n9620_), .Y(u2__abc_52138_new_n9623_));
NOR2X1 NOR2X1_1257 ( .A(u2__abc_52138_new_n9622_), .B(u2__abc_52138_new_n9625_), .Y(u2__abc_52138_new_n9626_));
NOR2X1 NOR2X1_1258 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9633_), .Y(u2__abc_52138_new_n9634_));
NOR2X1 NOR2X1_1259 ( .A(u2__abc_52138_new_n9669_), .B(u2__abc_52138_new_n9668_), .Y(u2__abc_52138_new_n9670_));
NOR2X1 NOR2X1_126 ( .A(u2_remHi_0_), .B(u2__abc_52138_new_n3072_), .Y(u2__abc_52138_new_n3073_));
NOR2X1 NOR2X1_1260 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9677_), .Y(u2__abc_52138_new_n9678_));
NOR2X1 NOR2X1_1261 ( .A(u2__abc_52138_new_n9751_), .B(u2__abc_52138_new_n9750_), .Y(u2__abc_52138_new_n9752_));
NOR2X1 NOR2X1_1262 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9759_), .Y(u2__abc_52138_new_n9760_));
NOR2X1 NOR2X1_1263 ( .A(u2__abc_52138_new_n5501_), .B(u2__abc_52138_new_n9707_), .Y(u2__abc_52138_new_n9787_));
NOR2X1 NOR2X1_1264 ( .A(u2__abc_52138_new_n9791_), .B(u2__abc_52138_new_n9787_), .Y(u2__abc_52138_new_n9792_));
NOR2X1 NOR2X1_1265 ( .A(u2__abc_52138_new_n9837_), .B(u2__abc_52138_new_n9836_), .Y(u2__abc_52138_new_n9838_));
NOR2X1 NOR2X1_1266 ( .A(u2__abc_52138_new_n9847_), .B(u2__abc_52138_new_n9845_), .Y(u2__abc_52138_new_n9848_));
NOR2X1 NOR2X1_1267 ( .A(u2__abc_52138_new_n9879_), .B(u2__abc_52138_new_n9878_), .Y(u2__abc_52138_new_n9880_));
NOR2X1 NOR2X1_1268 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9887_), .Y(u2__abc_52138_new_n9888_));
NOR2X1 NOR2X1_1269 ( .A(u2__abc_52138_new_n9922_), .B(u2__abc_52138_new_n9921_), .Y(u2__abc_52138_new_n9923_));
NOR2X1 NOR2X1_127 ( .A(u2_remHi_1_), .B(u2__abc_52138_new_n3074_), .Y(u2__abc_52138_new_n3075_));
NOR2X1 NOR2X1_1270 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n9930_), .Y(u2__abc_52138_new_n9931_));
NOR2X1 NOR2X1_1271 ( .A(u2__abc_52138_new_n5402_), .B(u2__abc_52138_new_n5397_), .Y(u2__abc_52138_new_n9960_));
NOR2X1 NOR2X1_1272 ( .A(u2__abc_52138_new_n5735_), .B(u2__abc_52138_new_n9288_), .Y(u2__abc_52138_new_n9966_));
NOR2X1 NOR2X1_1273 ( .A(u2__abc_52138_new_n9965_), .B(u2__abc_52138_new_n9966_), .Y(u2__abc_52138_new_n9967_));
NOR2X1 NOR2X1_1274 ( .A(u2__abc_52138_new_n10012_), .B(u2__abc_52138_new_n10011_), .Y(u2__abc_52138_new_n10013_));
NOR2X1 NOR2X1_1275 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10020_), .Y(u2__abc_52138_new_n10021_));
NOR2X1 NOR2X1_1276 ( .A(u2__abc_52138_new_n5340_), .B(u2__abc_52138_new_n10008_), .Y(u2__abc_52138_new_n10046_));
NOR2X1 NOR2X1_1277 ( .A(u2__abc_52138_new_n10049_), .B(u2__abc_52138_new_n10046_), .Y(u2__abc_52138_new_n10050_));
NOR2X1 NOR2X1_1278 ( .A(u2__abc_52138_new_n10095_), .B(u2__abc_52138_new_n10094_), .Y(u2__abc_52138_new_n10096_));
NOR2X1 NOR2X1_1279 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10104_), .Y(u2__abc_52138_new_n10105_));
NOR2X1 NOR2X1_128 ( .A(u2_remHi_8_), .B(u2__abc_52138_new_n3096_), .Y(u2__abc_52138_new_n3097_));
NOR2X1 NOR2X1_1280 ( .A(u2__abc_52138_new_n10140_), .B(u2__abc_52138_new_n10139_), .Y(u2__abc_52138_new_n10141_));
NOR2X1 NOR2X1_1281 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10148_), .Y(u2__abc_52138_new_n10149_));
NOR2X1 NOR2X1_1282 ( .A(u2__abc_52138_new_n10183_), .B(u2__abc_52138_new_n10182_), .Y(u2__abc_52138_new_n10184_));
NOR2X1 NOR2X1_1283 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10191_), .Y(u2__abc_52138_new_n10192_));
NOR2X1 NOR2X1_1284 ( .A(u2_remHi_340_), .B(u2__abc_52138_new_n5249_), .Y(u2__abc_52138_new_n10208_));
NOR2X1 NOR2X1_1285 ( .A(u2__abc_52138_new_n5269_), .B(u2__abc_52138_new_n5259_), .Y(u2__abc_52138_new_n10217_));
NOR2X1 NOR2X1_1286 ( .A(u2__abc_52138_new_n10226_), .B(u2__abc_52138_new_n10225_), .Y(u2__abc_52138_new_n10227_));
NOR2X1 NOR2X1_1287 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10235_), .Y(u2__abc_52138_new_n10236_));
NOR2X1 NOR2X1_1288 ( .A(u2_remHi_344_), .B(u2__abc_52138_new_n5183_), .Y(u2__abc_52138_new_n10253_));
NOR2X1 NOR2X1_1289 ( .A(u2__abc_52138_new_n10270_), .B(u2__abc_52138_new_n10269_), .Y(u2__abc_52138_new_n10271_));
NOR2X1 NOR2X1_129 ( .A(u2__abc_52138_new_n3116_), .B(u2__abc_52138_new_n3121_), .Y(u2__abc_52138_new_n3122_));
NOR2X1 NOR2X1_1290 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10278_), .Y(u2__abc_52138_new_n10279_));
NOR2X1 NOR2X1_1291 ( .A(u2__abc_52138_new_n10285_), .B(u2__abc_52138_new_n10287_), .Y(u2__abc_52138_new_n10288_));
NOR2X1 NOR2X1_1292 ( .A(u2__abc_52138_new_n10288_), .B(u2__abc_52138_new_n10290_), .Y(u2__abc_52138_new_n10291_));
NOR2X1 NOR2X1_1293 ( .A(u2__abc_52138_new_n5227_), .B(u2__abc_52138_new_n10266_), .Y(u2__abc_52138_new_n10305_));
NOR2X1 NOR2X1_1294 ( .A(u2__abc_52138_new_n10305_), .B(u2__abc_52138_new_n10310_), .Y(u2__abc_52138_new_n10311_));
NOR2X1 NOR2X1_1295 ( .A(u2__abc_52138_new_n10316_), .B(u2__abc_52138_new_n10315_), .Y(u2__abc_52138_new_n10317_));
NOR2X1 NOR2X1_1296 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10324_), .Y(u2__abc_52138_new_n10325_));
NOR2X1 NOR2X1_1297 ( .A(u2__abc_52138_new_n10358_), .B(u2__abc_52138_new_n10357_), .Y(u2__abc_52138_new_n10359_));
NOR2X1 NOR2X1_1298 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10367_), .Y(u2__abc_52138_new_n10368_));
NOR2X1 NOR2X1_1299 ( .A(u2__abc_52138_new_n10398_), .B(u2__abc_52138_new_n10399_), .Y(u2__abc_52138_new_n10400_));
NOR2X1 NOR2X1_13 ( .A(_abc_65734_new_n1518_), .B(_abc_65734_new_n1507_), .Y(_abc_65734_new_n1519_));
NOR2X1 NOR2X1_130 ( .A(u2__abc_52138_new_n3127_), .B(u2__abc_52138_new_n3132_), .Y(u2__abc_52138_new_n3133_));
NOR2X1 NOR2X1_1300 ( .A(u2__abc_52138_new_n5112_), .B(u2__abc_52138_new_n10420_), .Y(u2__abc_52138_new_n10439_));
NOR2X1 NOR2X1_1301 ( .A(u2__abc_52138_new_n10441_), .B(u2__abc_52138_new_n10439_), .Y(u2__abc_52138_new_n10442_));
NOR2X1 NOR2X1_1302 ( .A(u2__abc_52138_new_n10446_), .B(u2__abc_52138_new_n10445_), .Y(u2__abc_52138_new_n10447_));
NOR2X1 NOR2X1_1303 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10454_), .Y(u2__abc_52138_new_n10455_));
NOR2X1 NOR2X1_1304 ( .A(u2__abc_52138_new_n10481_), .B(u2__abc_52138_new_n10482_), .Y(u2__abc_52138_new_n10483_));
NOR2X1 NOR2X1_1305 ( .A(u2__abc_52138_new_n10484_), .B(u2__abc_52138_new_n10485_), .Y(u2__abc_52138_new_n10488_));
NOR2X1 NOR2X1_1306 ( .A(u2__abc_52138_new_n10487_), .B(u2__abc_52138_new_n10490_), .Y(u2__abc_52138_new_n10491_));
NOR2X1 NOR2X1_1307 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10498_), .Y(u2__abc_52138_new_n10499_));
NOR2X1 NOR2X1_1308 ( .A(u2__abc_52138_new_n10611_), .B(u2__abc_52138_new_n10610_), .Y(u2__abc_52138_new_n10612_));
NOR2X1 NOR2X1_1309 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10619_), .Y(u2__abc_52138_new_n10620_));
NOR2X1 NOR2X1_131 ( .A(u2__abc_52138_new_n3139_), .B(u2__abc_52138_new_n3144_), .Y(u2__abc_52138_new_n3145_));
NOR2X1 NOR2X1_1310 ( .A(u2__abc_52138_new_n10646_), .B(u2__abc_52138_new_n9288_), .Y(u2__abc_52138_new_n10647_));
NOR2X1 NOR2X1_1311 ( .A(u2__abc_52138_new_n10659_), .B(u2__abc_52138_new_n10647_), .Y(u2__abc_52138_new_n10662_));
NOR2X1 NOR2X1_1312 ( .A(u2__abc_52138_new_n10661_), .B(u2__abc_52138_new_n10664_), .Y(u2__abc_52138_new_n10665_));
NOR2X1 NOR2X1_1313 ( .A(u2__abc_52138_new_n10707_), .B(u2__abc_52138_new_n10706_), .Y(u2__abc_52138_new_n10708_));
NOR2X1 NOR2X1_1314 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10715_), .Y(u2__abc_52138_new_n10716_));
NOR2X1 NOR2X1_1315 ( .A(u2__abc_52138_new_n10722_), .B(u2__abc_52138_new_n10725_), .Y(u2__abc_52138_new_n10726_));
NOR2X1 NOR2X1_1316 ( .A(u2__abc_52138_new_n10726_), .B(u2__abc_52138_new_n10728_), .Y(u2__abc_52138_new_n10729_));
NOR2X1 NOR2X1_1317 ( .A(u2__abc_52138_new_n6148_), .B(u2__abc_52138_new_n6146_), .Y(u2__abc_52138_new_n10744_));
NOR2X1 NOR2X1_1318 ( .A(u2__abc_52138_new_n10796_), .B(u2__abc_52138_new_n10795_), .Y(u2__abc_52138_new_n10797_));
NOR2X1 NOR2X1_1319 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10804_), .Y(u2__abc_52138_new_n10805_));
NOR2X1 NOR2X1_132 ( .A(u2__abc_52138_new_n3150_), .B(u2__abc_52138_new_n3155_), .Y(u2__abc_52138_new_n3156_));
NOR2X1 NOR2X1_1320 ( .A(u2__abc_52138_new_n10833_), .B(u2__abc_52138_new_n10834_), .Y(u2__abc_52138_new_n10835_));
NOR2X1 NOR2X1_1321 ( .A(u2__abc_52138_new_n10880_), .B(u2__abc_52138_new_n10879_), .Y(u2__abc_52138_new_n10881_));
NOR2X1 NOR2X1_1322 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10888_), .Y(u2__abc_52138_new_n10889_));
NOR2X1 NOR2X1_1323 ( .A(u2__abc_52138_new_n10915_), .B(u2__abc_52138_new_n10876_), .Y(u2__abc_52138_new_n10916_));
NOR2X1 NOR2X1_1324 ( .A(u2__abc_52138_new_n10919_), .B(u2__abc_52138_new_n10916_), .Y(u2__abc_52138_new_n10920_));
NOR2X1 NOR2X1_1325 ( .A(u2__abc_52138_new_n10924_), .B(u2__abc_52138_new_n10923_), .Y(u2__abc_52138_new_n10925_));
NOR2X1 NOR2X1_1326 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10932_), .Y(u2__abc_52138_new_n10933_));
NOR2X1 NOR2X1_1327 ( .A(u2__abc_52138_new_n10967_), .B(u2__abc_52138_new_n10966_), .Y(u2__abc_52138_new_n10968_));
NOR2X1 NOR2X1_1328 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n10976_), .Y(u2__abc_52138_new_n10977_));
NOR2X1 NOR2X1_1329 ( .A(u2__abc_52138_new_n11007_), .B(u2__abc_52138_new_n11009_), .Y(u2__abc_52138_new_n11010_));
NOR2X1 NOR2X1_133 ( .A(u2__abc_52138_new_n3163_), .B(u2__abc_52138_new_n3168_), .Y(u2__abc_52138_new_n3169_));
NOR2X1 NOR2X1_1330 ( .A(u2__abc_52138_new_n11014_), .B(u2__abc_52138_new_n11013_), .Y(u2__abc_52138_new_n11015_));
NOR2X1 NOR2X1_1331 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n11022_), .Y(u2__abc_52138_new_n11023_));
NOR2X1 NOR2X1_1332 ( .A(u2__abc_52138_new_n6112_), .B(u2__abc_52138_new_n11031_), .Y(u2__abc_52138_new_n11032_));
NOR2X1 NOR2X1_1333 ( .A(u2__abc_52138_new_n11032_), .B(u2__abc_52138_new_n11034_), .Y(u2__abc_52138_new_n11035_));
NOR2X1 NOR2X1_1334 ( .A(u2__abc_52138_new_n11058_), .B(u2__abc_52138_new_n11057_), .Y(u2__abc_52138_new_n11059_));
NOR2X1 NOR2X1_1335 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n11067_), .Y(u2__abc_52138_new_n11068_));
NOR2X1 NOR2X1_1336 ( .A(u2__abc_52138_new_n6088_), .B(u2__abc_52138_new_n11075_), .Y(u2__abc_52138_new_n11076_));
NOR2X1 NOR2X1_1337 ( .A(u2__abc_52138_new_n11076_), .B(u2__abc_52138_new_n11078_), .Y(u2__abc_52138_new_n11079_));
NOR2X1 NOR2X1_1338 ( .A(u2__abc_52138_new_n6097_), .B(u2__abc_52138_new_n6095_), .Y(u2__abc_52138_new_n11095_));
NOR2X1 NOR2X1_1339 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n11110_), .Y(u2__abc_52138_new_n11111_));
NOR2X1 NOR2X1_134 ( .A(u2__abc_52138_new_n3174_), .B(u2__abc_52138_new_n3179_), .Y(u2__abc_52138_new_n3180_));
NOR2X1 NOR2X1_1340 ( .A(u2__abc_52138_new_n6040_), .B(u2__abc_52138_new_n11118_), .Y(u2__abc_52138_new_n11119_));
NOR2X1 NOR2X1_1341 ( .A(u2__abc_52138_new_n11119_), .B(u2__abc_52138_new_n11121_), .Y(u2__abc_52138_new_n11122_));
NOR2X1 NOR2X1_1342 ( .A(u2__abc_52138_new_n11143_), .B(u2__abc_52138_new_n11142_), .Y(u2__abc_52138_new_n11144_));
NOR2X1 NOR2X1_1343 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n11151_), .Y(u2__abc_52138_new_n11152_));
NOR2X1 NOR2X1_1344 ( .A(u2__abc_52138_new_n6073_), .B(u2__abc_52138_new_n6076_), .Y(u2__abc_52138_new_n11158_));
NOR2X1 NOR2X1_1345 ( .A(u2__abc_52138_new_n6062_), .B(u2__abc_52138_new_n11160_), .Y(u2__abc_52138_new_n11161_));
NOR2X1 NOR2X1_1346 ( .A(u2__abc_52138_new_n11161_), .B(u2__abc_52138_new_n11163_), .Y(u2__abc_52138_new_n11164_));
NOR2X1 NOR2X1_1347 ( .A(u2__abc_52138_new_n6071_), .B(u2__abc_52138_new_n11158_), .Y(u2__abc_52138_new_n11180_));
NOR2X1 NOR2X1_1348 ( .A(u2__abc_52138_new_n11208_), .B(u2__abc_52138_new_n11207_), .Y(u2__abc_52138_new_n11209_));
NOR2X1 NOR2X1_1349 ( .A(u2__abc_52138_new_n11238_), .B(u2__abc_52138_new_n11237_), .Y(u2__abc_52138_new_n11239_));
NOR2X1 NOR2X1_135 ( .A(u2__abc_52138_new_n3187_), .B(u2__abc_52138_new_n3193_), .Y(u2__abc_52138_new_n3194_));
NOR2X1 NOR2X1_1350 ( .A(u2__abc_52138_new_n5991_), .B(u2__abc_52138_new_n11246_), .Y(u2__abc_52138_new_n11247_));
NOR2X1 NOR2X1_1351 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n11247_), .Y(u2__abc_52138_new_n11248_));
NOR2X1 NOR2X1_1352 ( .A(u2__abc_52138_new_n11286_), .B(u2__abc_52138_new_n11290_), .Y(u2__abc_52138_new_n11291_));
NOR2X1 NOR2X1_1353 ( .A(u2__abc_52138_new_n11291_), .B(u2__abc_52138_new_n11293_), .Y(u2__abc_52138_new_n11294_));
NOR2X1 NOR2X1_1354 ( .A(u2__abc_52138_new_n11316_), .B(u2__abc_52138_new_n11315_), .Y(u2__abc_52138_new_n11317_));
NOR2X1 NOR2X1_1355 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n11324_), .Y(u2__abc_52138_new_n11325_));
NOR2X1 NOR2X1_1356 ( .A(u2__abc_52138_new_n5958_), .B(u2__abc_52138_new_n5961_), .Y(u2__abc_52138_new_n11332_));
NOR2X1 NOR2X1_1357 ( .A(u2__abc_52138_new_n5986_), .B(u2__abc_52138_new_n11268_), .Y(u2__abc_52138_new_n11352_));
NOR2X1 NOR2X1_1358 ( .A(u2__abc_52138_new_n5956_), .B(u2__abc_52138_new_n5954_), .Y(u2__abc_52138_new_n11355_));
NOR2X1 NOR2X1_1359 ( .A(u2__abc_52138_new_n11357_), .B(u2__abc_52138_new_n11352_), .Y(u2__abc_52138_new_n11358_));
NOR2X1 NOR2X1_136 ( .A(u2__abc_52138_new_n3195_), .B(u2__abc_52138_new_n3158_), .Y(u2__abc_52138_new_n3196_));
NOR2X1 NOR2X1_1360 ( .A(u2__abc_52138_new_n11377_), .B(u2__abc_52138_new_n2974_), .Y(u2__abc_52138_new_n11382_));
NOR2X1 NOR2X1_1361 ( .A(u2__abc_52138_new_n11382_), .B(u2__abc_52138_new_n11378_), .Y(u2__abc_52138_new_n11383_));
NOR2X1 NOR2X1_1362 ( .A(u2__abc_52138_new_n2966_), .B(u2__abc_52138_new_n11388_), .Y(u2__abc_52138_new_n11391_));
NOR2X1 NOR2X1_1363 ( .A(rst), .B(u2__abc_52138_new_n11394_), .Y(u2__abc_52138_new_n11395_));
NOR2X1 NOR2X1_1364 ( .A(u2__abc_52138_new_n11393_), .B(u2__abc_52138_new_n11396_), .Y(u2__0cnt_7_0__3_));
NOR2X1 NOR2X1_1365 ( .A(u2__abc_52138_new_n2967_), .B(u2__abc_52138_new_n11392_), .Y(u2__abc_52138_new_n11398_));
NOR2X1 NOR2X1_1366 ( .A(u2__abc_52138_new_n11398_), .B(u2__abc_52138_new_n11399_), .Y(u2__0cnt_7_0__4_));
NOR2X1 NOR2X1_1367 ( .A(u2__abc_52138_new_n11403_), .B(u2__abc_52138_new_n11402_), .Y(u2__0cnt_7_0__5_));
NOR2X1 NOR2X1_1368 ( .A(u2_cnt_6_), .B(u2__abc_52138_new_n11402_), .Y(u2__abc_52138_new_n11405_));
NOR2X1 NOR2X1_1369 ( .A(u2__abc_52138_new_n11406_), .B(u2__abc_52138_new_n11401_), .Y(u2__abc_52138_new_n11409_));
NOR2X1 NOR2X1_137 ( .A(u2_remHi_19_), .B(u2__abc_52138_new_n3206_), .Y(u2__abc_52138_new_n3208_));
NOR2X1 NOR2X1_1370 ( .A(rst), .B(u2__abc_52138_new_n11413_), .Y(u2__0remLo_451_0__0_));
NOR2X1 NOR2X1_1371 ( .A(rst), .B(u2__abc_52138_new_n11415_), .Y(u2__0remLo_451_0__1_));
NOR2X1 NOR2X1_1372 ( .A(u2__abc_52138_new_n6503_), .B(u2__abc_52138_new_n2991_), .Y(u2__abc_52138_new_n11509_));
NOR2X1 NOR2X1_1373 ( .A(rst), .B(u2__abc_52138_new_n2965_), .Y(u2__abc_52138_new_n11717_));
NOR2X1 NOR2X1_1374 ( .A(u2__abc_52138_new_n11710_), .B(u2__abc_52138_new_n2986_), .Y(u2__abc_52138_new_n11718_));
NOR2X1 NOR2X1_1375 ( .A(u2__abc_52138_new_n11716_), .B(u2__abc_52138_new_n2986_), .Y(u2__abc_52138_new_n11725_));
NOR2X1 NOR2X1_1376 ( .A(u2__abc_52138_new_n11830_), .B(u2__abc_52138_new_n2986_), .Y(u2__abc_52138_new_n11840_));
NOR2X1 NOR2X1_1377 ( .A(u2__abc_52138_new_n11960_), .B(u2__abc_52138_new_n2986_), .Y(u2__abc_52138_new_n11967_));
NOR2X1 NOR2X1_1378 ( .A(u2__abc_52138_new_n12060_), .B(u2__abc_52138_new_n2986_), .Y(u2__abc_52138_new_n12070_));
NOR2X1 NOR2X1_1379 ( .A(u2__abc_52138_new_n12154_), .B(u2__abc_52138_new_n2986_), .Y(u2__abc_52138_new_n12161_));
NOR2X1 NOR2X1_138 ( .A(sqrto_21_), .B(u2__abc_52138_new_n3185_), .Y(u2__abc_52138_new_n3213_));
NOR2X1 NOR2X1_1380 ( .A(u2__abc_52138_new_n12221_), .B(u2__abc_52138_new_n2986_), .Y(u2__abc_52138_new_n12228_));
NOR2X1 NOR2X1_1381 ( .A(rst), .B(u2__abc_52138_new_n12816_), .Y(u2__0root_452_0__0_));
NOR2X1 NOR2X1_1382 ( .A(u2__abc_52138_new_n6599_), .B(u2__abc_52138_new_n6614_), .Y(u2__abc_52138_new_n12820_));
NOR2X1 NOR2X1_1383 ( .A(u2__abc_52138_new_n12821_), .B(u2__abc_52138_new_n12819_), .Y(u2__abc_52138_new_n12822_));
NOR2X1 NOR2X1_1384 ( .A(u2__abc_52138_new_n3134_), .B(u2__abc_52138_new_n3157_), .Y(u2__abc_52138_new_n12838_));
NOR2X1 NOR2X1_1385 ( .A(u2__abc_52138_new_n3420_), .B(u2__abc_52138_new_n3334_), .Y(u2__abc_52138_new_n12857_));
NOR2X1 NOR2X1_1386 ( .A(u2__abc_52138_new_n7035_), .B(u2__abc_52138_new_n12872_), .Y(u2__abc_52138_new_n12873_));
NOR2X1 NOR2X1_1387 ( .A(u2__abc_52138_new_n7447_), .B(u2__abc_52138_new_n7400_), .Y(u2__abc_52138_new_n12887_));
NOR2X1 NOR2X1_1388 ( .A(u2__abc_52138_new_n7310_), .B(u2__abc_52138_new_n7355_), .Y(u2__abc_52138_new_n12889_));
NOR2X1 NOR2X1_1389 ( .A(u2__abc_52138_new_n12894_), .B(u2__abc_52138_new_n7252_), .Y(u2__abc_52138_new_n12895_));
NOR2X1 NOR2X1_139 ( .A(sqrto_25_), .B(u2__abc_52138_new_n3119_), .Y(u2__abc_52138_new_n3225_));
NOR2X1 NOR2X1_1390 ( .A(u2__abc_52138_new_n7503_), .B(u2__abc_52138_new_n7491_), .Y(u2__abc_52138_new_n12916_));
NOR2X1 NOR2X1_1391 ( .A(u2__abc_52138_new_n3717_), .B(u2__abc_52138_new_n3722_), .Y(u2__abc_52138_new_n12918_));
NOR2X1 NOR2X1_1392 ( .A(u2__abc_52138_new_n12926_), .B(u2__abc_52138_new_n7570_), .Y(u2__abc_52138_new_n12927_));
NOR2X1 NOR2X1_1393 ( .A(u2__abc_52138_new_n3601_), .B(u2__abc_52138_new_n3606_), .Y(u2__abc_52138_new_n12934_));
NOR2X1 NOR2X1_1394 ( .A(u2__abc_52138_new_n3587_), .B(u2__abc_52138_new_n3592_), .Y(u2__abc_52138_new_n12941_));
NOR2X1 NOR2X1_1395 ( .A(u2__abc_52138_new_n8590_), .B(u2__abc_52138_new_n9268_), .Y(u2__abc_52138_new_n12954_));
NOR2X1 NOR2X1_1396 ( .A(u2__abc_52138_new_n8101_), .B(u2__abc_52138_new_n8112_), .Y(u2__abc_52138_new_n12968_));
NOR2X1 NOR2X1_1397 ( .A(u2__abc_52138_new_n8939_), .B(u2__abc_52138_new_n8895_), .Y(u2__abc_52138_new_n13006_));
NOR2X1 NOR2X1_1398 ( .A(u2_root_0_), .B(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n13045_));
NOR2X1 NOR2X1_1399 ( .A(sqrto_0_), .B(u2__abc_52138_new_n13044_), .Y(u2__abc_52138_new_n13052_));
NOR2X1 NOR2X1_14 ( .A(_abc_65734_new_n1500_), .B(_abc_65734_new_n1492_), .Y(_abc_65734_new_n1524_));
NOR2X1 NOR2X1_140 ( .A(u2_remHi_29_), .B(u2__abc_52138_new_n3142_), .Y(u2__abc_52138_new_n3231_));
NOR2X1 NOR2X1_1400 ( .A(sqrto_1_), .B(u2__abc_52138_new_n13051_), .Y(u2__abc_52138_new_n13058_));
NOR2X1 NOR2X1_1401 ( .A(sqrto_2_), .B(u2__abc_52138_new_n13060_), .Y(u2__abc_52138_new_n13066_));
NOR2X1 NOR2X1_1402 ( .A(sqrto_3_), .B(u2__abc_52138_new_n13068_), .Y(u2__abc_52138_new_n13074_));
NOR2X1 NOR2X1_1403 ( .A(sqrto_4_), .B(u2__abc_52138_new_n13076_), .Y(u2__abc_52138_new_n13082_));
NOR2X1 NOR2X1_1404 ( .A(sqrto_5_), .B(u2__abc_52138_new_n13083_), .Y(u2__abc_52138_new_n13089_));
NOR2X1 NOR2X1_1405 ( .A(sqrto_6_), .B(u2__abc_52138_new_n13091_), .Y(u2__abc_52138_new_n13097_));
NOR2X1 NOR2X1_1406 ( .A(sqrto_7_), .B(u2__abc_52138_new_n13099_), .Y(u2__abc_52138_new_n13105_));
NOR2X1 NOR2X1_1407 ( .A(sqrto_8_), .B(u2__abc_52138_new_n13107_), .Y(u2__abc_52138_new_n13113_));
NOR2X1 NOR2X1_1408 ( .A(sqrto_9_), .B(u2__abc_52138_new_n13114_), .Y(u2__abc_52138_new_n13120_));
NOR2X1 NOR2X1_1409 ( .A(sqrto_10_), .B(u2__abc_52138_new_n13122_), .Y(u2__abc_52138_new_n13128_));
NOR2X1 NOR2X1_141 ( .A(u2__abc_52138_new_n3244_), .B(u2__abc_52138_new_n3249_), .Y(u2__abc_52138_new_n3250_));
NOR2X1 NOR2X1_1410 ( .A(sqrto_11_), .B(u2__abc_52138_new_n13130_), .Y(u2__abc_52138_new_n13136_));
NOR2X1 NOR2X1_1411 ( .A(sqrto_12_), .B(u2__abc_52138_new_n13138_), .Y(u2__abc_52138_new_n13144_));
NOR2X1 NOR2X1_1412 ( .A(sqrto_13_), .B(u2__abc_52138_new_n13145_), .Y(u2__abc_52138_new_n13151_));
NOR2X1 NOR2X1_1413 ( .A(sqrto_14_), .B(u2__abc_52138_new_n13153_), .Y(u2__abc_52138_new_n13159_));
NOR2X1 NOR2X1_1414 ( .A(sqrto_15_), .B(u2__abc_52138_new_n13161_), .Y(u2__abc_52138_new_n13167_));
NOR2X1 NOR2X1_1415 ( .A(sqrto_16_), .B(u2__abc_52138_new_n13169_), .Y(u2__abc_52138_new_n13175_));
NOR2X1 NOR2X1_1416 ( .A(sqrto_17_), .B(u2__abc_52138_new_n13176_), .Y(u2__abc_52138_new_n13182_));
NOR2X1 NOR2X1_1417 ( .A(sqrto_18_), .B(u2__abc_52138_new_n13184_), .Y(u2__abc_52138_new_n13190_));
NOR2X1 NOR2X1_1418 ( .A(sqrto_19_), .B(u2__abc_52138_new_n13192_), .Y(u2__abc_52138_new_n13198_));
NOR2X1 NOR2X1_1419 ( .A(sqrto_20_), .B(u2__abc_52138_new_n13200_), .Y(u2__abc_52138_new_n13206_));
NOR2X1 NOR2X1_142 ( .A(u2__abc_52138_new_n3255_), .B(u2__abc_52138_new_n3260_), .Y(u2__abc_52138_new_n3261_));
NOR2X1 NOR2X1_1420 ( .A(sqrto_21_), .B(u2__abc_52138_new_n13207_), .Y(u2__abc_52138_new_n13213_));
NOR2X1 NOR2X1_1421 ( .A(sqrto_22_), .B(u2__abc_52138_new_n13215_), .Y(u2__abc_52138_new_n13221_));
NOR2X1 NOR2X1_1422 ( .A(sqrto_23_), .B(u2__abc_52138_new_n13223_), .Y(u2__abc_52138_new_n13229_));
NOR2X1 NOR2X1_1423 ( .A(sqrto_24_), .B(u2__abc_52138_new_n13231_), .Y(u2__abc_52138_new_n13237_));
NOR2X1 NOR2X1_1424 ( .A(sqrto_25_), .B(u2__abc_52138_new_n13238_), .Y(u2__abc_52138_new_n13244_));
NOR2X1 NOR2X1_1425 ( .A(sqrto_26_), .B(u2__abc_52138_new_n13246_), .Y(u2__abc_52138_new_n13252_));
NOR2X1 NOR2X1_1426 ( .A(sqrto_27_), .B(u2__abc_52138_new_n13254_), .Y(u2__abc_52138_new_n13260_));
NOR2X1 NOR2X1_1427 ( .A(sqrto_28_), .B(u2__abc_52138_new_n13262_), .Y(u2__abc_52138_new_n13268_));
NOR2X1 NOR2X1_1428 ( .A(sqrto_29_), .B(u2__abc_52138_new_n13269_), .Y(u2__abc_52138_new_n13275_));
NOR2X1 NOR2X1_1429 ( .A(sqrto_30_), .B(u2__abc_52138_new_n13277_), .Y(u2__abc_52138_new_n13283_));
NOR2X1 NOR2X1_143 ( .A(u2__abc_52138_new_n3267_), .B(u2__abc_52138_new_n3272_), .Y(u2__abc_52138_new_n3273_));
NOR2X1 NOR2X1_1430 ( .A(sqrto_31_), .B(u2__abc_52138_new_n13285_), .Y(u2__abc_52138_new_n13291_));
NOR2X1 NOR2X1_1431 ( .A(sqrto_32_), .B(u2__abc_52138_new_n13293_), .Y(u2__abc_52138_new_n13299_));
NOR2X1 NOR2X1_1432 ( .A(sqrto_33_), .B(u2__abc_52138_new_n13300_), .Y(u2__abc_52138_new_n13306_));
NOR2X1 NOR2X1_1433 ( .A(sqrto_34_), .B(u2__abc_52138_new_n13308_), .Y(u2__abc_52138_new_n13315_));
NOR2X1 NOR2X1_1434 ( .A(sqrto_35_), .B(u2__abc_52138_new_n13317_), .Y(u2__abc_52138_new_n13323_));
NOR2X1 NOR2X1_1435 ( .A(sqrto_36_), .B(u2__abc_52138_new_n13325_), .Y(u2__abc_52138_new_n13331_));
NOR2X1 NOR2X1_1436 ( .A(sqrto_37_), .B(u2__abc_52138_new_n13332_), .Y(u2__abc_52138_new_n13338_));
NOR2X1 NOR2X1_1437 ( .A(sqrto_38_), .B(u2__abc_52138_new_n13340_), .Y(u2__abc_52138_new_n13346_));
NOR2X1 NOR2X1_1438 ( .A(sqrto_39_), .B(u2__abc_52138_new_n13348_), .Y(u2__abc_52138_new_n13354_));
NOR2X1 NOR2X1_1439 ( .A(sqrto_40_), .B(u2__abc_52138_new_n13356_), .Y(u2__abc_52138_new_n13362_));
NOR2X1 NOR2X1_144 ( .A(u2__abc_52138_new_n3278_), .B(u2__abc_52138_new_n3283_), .Y(u2__abc_52138_new_n3284_));
NOR2X1 NOR2X1_1440 ( .A(sqrto_41_), .B(u2__abc_52138_new_n13363_), .Y(u2__abc_52138_new_n13369_));
NOR2X1 NOR2X1_1441 ( .A(sqrto_42_), .B(u2__abc_52138_new_n13371_), .Y(u2__abc_52138_new_n13377_));
NOR2X1 NOR2X1_1442 ( .A(sqrto_43_), .B(u2__abc_52138_new_n13379_), .Y(u2__abc_52138_new_n13385_));
NOR2X1 NOR2X1_1443 ( .A(sqrto_44_), .B(u2__abc_52138_new_n13387_), .Y(u2__abc_52138_new_n13393_));
NOR2X1 NOR2X1_1444 ( .A(sqrto_45_), .B(u2__abc_52138_new_n13394_), .Y(u2__abc_52138_new_n13400_));
NOR2X1 NOR2X1_1445 ( .A(sqrto_46_), .B(u2__abc_52138_new_n13402_), .Y(u2__abc_52138_new_n13408_));
NOR2X1 NOR2X1_1446 ( .A(sqrto_47_), .B(u2__abc_52138_new_n13410_), .Y(u2__abc_52138_new_n13416_));
NOR2X1 NOR2X1_1447 ( .A(sqrto_48_), .B(u2__abc_52138_new_n13418_), .Y(u2__abc_52138_new_n13424_));
NOR2X1 NOR2X1_1448 ( .A(sqrto_49_), .B(u2__abc_52138_new_n13425_), .Y(u2__abc_52138_new_n13431_));
NOR2X1 NOR2X1_1449 ( .A(sqrto_50_), .B(u2__abc_52138_new_n13433_), .Y(u2__abc_52138_new_n13439_));
NOR2X1 NOR2X1_145 ( .A(u2__abc_52138_new_n3262_), .B(u2__abc_52138_new_n3285_), .Y(u2__abc_52138_new_n3286_));
NOR2X1 NOR2X1_1450 ( .A(sqrto_51_), .B(u2__abc_52138_new_n13441_), .Y(u2__abc_52138_new_n13447_));
NOR2X1 NOR2X1_1451 ( .A(sqrto_52_), .B(u2__abc_52138_new_n13449_), .Y(u2__abc_52138_new_n13455_));
NOR2X1 NOR2X1_1452 ( .A(sqrto_53_), .B(u2__abc_52138_new_n13456_), .Y(u2__abc_52138_new_n13462_));
NOR2X1 NOR2X1_1453 ( .A(sqrto_54_), .B(u2__abc_52138_new_n13464_), .Y(u2__abc_52138_new_n13470_));
NOR2X1 NOR2X1_1454 ( .A(sqrto_55_), .B(u2__abc_52138_new_n13472_), .Y(u2__abc_52138_new_n13478_));
NOR2X1 NOR2X1_1455 ( .A(sqrto_56_), .B(u2__abc_52138_new_n13480_), .Y(u2__abc_52138_new_n13486_));
NOR2X1 NOR2X1_1456 ( .A(sqrto_57_), .B(u2__abc_52138_new_n13487_), .Y(u2__abc_52138_new_n13493_));
NOR2X1 NOR2X1_1457 ( .A(sqrto_58_), .B(u2__abc_52138_new_n13495_), .Y(u2__abc_52138_new_n13501_));
NOR2X1 NOR2X1_1458 ( .A(sqrto_59_), .B(u2__abc_52138_new_n13503_), .Y(u2__abc_52138_new_n13509_));
NOR2X1 NOR2X1_1459 ( .A(sqrto_60_), .B(u2__abc_52138_new_n13511_), .Y(u2__abc_52138_new_n13517_));
NOR2X1 NOR2X1_146 ( .A(sqrto_48_), .B(u2__abc_52138_new_n3287_), .Y(u2__abc_52138_new_n3288_));
NOR2X1 NOR2X1_1460 ( .A(sqrto_61_), .B(u2__abc_52138_new_n13518_), .Y(u2__abc_52138_new_n13524_));
NOR2X1 NOR2X1_1461 ( .A(sqrto_62_), .B(u2__abc_52138_new_n13526_), .Y(u2__abc_52138_new_n13532_));
NOR2X1 NOR2X1_1462 ( .A(sqrto_63_), .B(u2__abc_52138_new_n13534_), .Y(u2__abc_52138_new_n13540_));
NOR2X1 NOR2X1_1463 ( .A(sqrto_64_), .B(u2__abc_52138_new_n13542_), .Y(u2__abc_52138_new_n13548_));
NOR2X1 NOR2X1_1464 ( .A(sqrto_65_), .B(u2__abc_52138_new_n13549_), .Y(u2__abc_52138_new_n13555_));
NOR2X1 NOR2X1_1465 ( .A(sqrto_66_), .B(u2__abc_52138_new_n13557_), .Y(u2__abc_52138_new_n13563_));
NOR2X1 NOR2X1_1466 ( .A(sqrto_67_), .B(u2__abc_52138_new_n13565_), .Y(u2__abc_52138_new_n13571_));
NOR2X1 NOR2X1_1467 ( .A(sqrto_68_), .B(u2__abc_52138_new_n13573_), .Y(u2__abc_52138_new_n13579_));
NOR2X1 NOR2X1_1468 ( .A(sqrto_69_), .B(u2__abc_52138_new_n13580_), .Y(u2__abc_52138_new_n13586_));
NOR2X1 NOR2X1_1469 ( .A(sqrto_70_), .B(u2__abc_52138_new_n13588_), .Y(u2__abc_52138_new_n13594_));
NOR2X1 NOR2X1_147 ( .A(u2_remHi_48_), .B(u2__abc_52138_new_n3289_), .Y(u2__abc_52138_new_n3290_));
NOR2X1 NOR2X1_1470 ( .A(sqrto_71_), .B(u2__abc_52138_new_n13596_), .Y(u2__abc_52138_new_n13602_));
NOR2X1 NOR2X1_1471 ( .A(sqrto_72_), .B(u2__abc_52138_new_n13604_), .Y(u2__abc_52138_new_n13610_));
NOR2X1 NOR2X1_1472 ( .A(sqrto_73_), .B(u2__abc_52138_new_n13611_), .Y(u2__abc_52138_new_n13617_));
NOR2X1 NOR2X1_1473 ( .A(sqrto_74_), .B(u2__abc_52138_new_n13619_), .Y(u2__abc_52138_new_n13625_));
NOR2X1 NOR2X1_1474 ( .A(sqrto_75_), .B(u2__abc_52138_new_n13627_), .Y(u2__abc_52138_new_n13633_));
NOR2X1 NOR2X1_1475 ( .A(sqrto_76_), .B(u2__abc_52138_new_n13635_), .Y(u2__abc_52138_new_n13641_));
NOR2X1 NOR2X1_1476 ( .A(sqrto_77_), .B(u2__abc_52138_new_n13642_), .Y(u2__abc_52138_new_n13648_));
NOR2X1 NOR2X1_1477 ( .A(sqrto_78_), .B(u2__abc_52138_new_n13650_), .Y(u2__abc_52138_new_n13656_));
NOR2X1 NOR2X1_1478 ( .A(sqrto_79_), .B(u2__abc_52138_new_n13658_), .Y(u2__abc_52138_new_n13666_));
NOR2X1 NOR2X1_1479 ( .A(sqrto_80_), .B(u2__abc_52138_new_n13665_), .Y(u2__abc_52138_new_n13672_));
NOR2X1 NOR2X1_148 ( .A(u2__abc_52138_new_n3288_), .B(u2__abc_52138_new_n3290_), .Y(u2__abc_52138_new_n3291_));
NOR2X1 NOR2X1_1480 ( .A(sqrto_81_), .B(u2__abc_52138_new_n13673_), .Y(u2__abc_52138_new_n13679_));
NOR2X1 NOR2X1_1481 ( .A(sqrto_82_), .B(u2__abc_52138_new_n13681_), .Y(u2__abc_52138_new_n13687_));
NOR2X1 NOR2X1_1482 ( .A(sqrto_83_), .B(u2__abc_52138_new_n13689_), .Y(u2__abc_52138_new_n13695_));
NOR2X1 NOR2X1_1483 ( .A(sqrto_84_), .B(u2__abc_52138_new_n13697_), .Y(u2__abc_52138_new_n13703_));
NOR2X1 NOR2X1_1484 ( .A(sqrto_85_), .B(u2__abc_52138_new_n13704_), .Y(u2__abc_52138_new_n13710_));
NOR2X1 NOR2X1_1485 ( .A(sqrto_86_), .B(u2__abc_52138_new_n13712_), .Y(u2__abc_52138_new_n13718_));
NOR2X1 NOR2X1_1486 ( .A(sqrto_87_), .B(u2__abc_52138_new_n13720_), .Y(u2__abc_52138_new_n13728_));
NOR2X1 NOR2X1_1487 ( .A(sqrto_88_), .B(u2__abc_52138_new_n13727_), .Y(u2__abc_52138_new_n13734_));
NOR2X1 NOR2X1_1488 ( .A(sqrto_89_), .B(u2__abc_52138_new_n13735_), .Y(u2__abc_52138_new_n13741_));
NOR2X1 NOR2X1_1489 ( .A(sqrto_90_), .B(u2__abc_52138_new_n13743_), .Y(u2__abc_52138_new_n13749_));
NOR2X1 NOR2X1_149 ( .A(sqrto_49_), .B(u2__abc_52138_new_n3292_), .Y(u2__abc_52138_new_n3293_));
NOR2X1 NOR2X1_1490 ( .A(sqrto_91_), .B(u2__abc_52138_new_n13751_), .Y(u2__abc_52138_new_n13759_));
NOR2X1 NOR2X1_1491 ( .A(sqrto_92_), .B(u2__abc_52138_new_n13758_), .Y(u2__abc_52138_new_n13765_));
NOR2X1 NOR2X1_1492 ( .A(sqrto_93_), .B(u2__abc_52138_new_n13766_), .Y(u2__abc_52138_new_n13774_));
NOR2X1 NOR2X1_1493 ( .A(sqrto_94_), .B(u2__abc_52138_new_n13773_), .Y(u2__abc_52138_new_n13780_));
NOR2X1 NOR2X1_1494 ( .A(sqrto_95_), .B(u2__abc_52138_new_n13782_), .Y(u2__abc_52138_new_n13788_));
NOR2X1 NOR2X1_1495 ( .A(sqrto_96_), .B(u2__abc_52138_new_n13790_), .Y(u2__abc_52138_new_n13796_));
NOR2X1 NOR2X1_1496 ( .A(sqrto_97_), .B(u2__abc_52138_new_n13797_), .Y(u2__abc_52138_new_n13803_));
NOR2X1 NOR2X1_1497 ( .A(sqrto_98_), .B(u2__abc_52138_new_n13805_), .Y(u2__abc_52138_new_n13811_));
NOR2X1 NOR2X1_1498 ( .A(sqrto_99_), .B(u2__abc_52138_new_n13813_), .Y(u2__abc_52138_new_n13819_));
NOR2X1 NOR2X1_1499 ( .A(sqrto_100_), .B(u2__abc_52138_new_n13821_), .Y(u2__abc_52138_new_n13827_));
NOR2X1 NOR2X1_15 ( .A(_abc_65734_new_n1527_), .B(_abc_65734_new_n1522_), .Y(_abc_65734_new_n1528_));
NOR2X1 NOR2X1_150 ( .A(u2_remHi_49_), .B(u2__abc_52138_new_n3294_), .Y(u2__abc_52138_new_n3295_));
NOR2X1 NOR2X1_1500 ( .A(sqrto_101_), .B(u2__abc_52138_new_n13828_), .Y(u2__abc_52138_new_n13834_));
NOR2X1 NOR2X1_1501 ( .A(sqrto_102_), .B(u2__abc_52138_new_n13836_), .Y(u2__abc_52138_new_n13842_));
NOR2X1 NOR2X1_1502 ( .A(sqrto_103_), .B(u2__abc_52138_new_n13844_), .Y(u2__abc_52138_new_n13852_));
NOR2X1 NOR2X1_1503 ( .A(sqrto_104_), .B(u2__abc_52138_new_n13851_), .Y(u2__abc_52138_new_n13858_));
NOR2X1 NOR2X1_1504 ( .A(sqrto_105_), .B(u2__abc_52138_new_n13859_), .Y(u2__abc_52138_new_n13865_));
NOR2X1 NOR2X1_1505 ( .A(sqrto_106_), .B(u2__abc_52138_new_n13867_), .Y(u2__abc_52138_new_n13873_));
NOR2X1 NOR2X1_1506 ( .A(sqrto_107_), .B(u2__abc_52138_new_n13875_), .Y(u2__abc_52138_new_n13883_));
NOR2X1 NOR2X1_1507 ( .A(sqrto_108_), .B(u2__abc_52138_new_n13882_), .Y(u2__abc_52138_new_n13889_));
NOR2X1 NOR2X1_1508 ( .A(sqrto_109_), .B(u2__abc_52138_new_n13890_), .Y(u2__abc_52138_new_n13898_));
NOR2X1 NOR2X1_1509 ( .A(sqrto_110_), .B(u2__abc_52138_new_n13897_), .Y(u2__abc_52138_new_n13904_));
NOR2X1 NOR2X1_151 ( .A(u2__abc_52138_new_n3293_), .B(u2__abc_52138_new_n3295_), .Y(u2__abc_52138_new_n3296_));
NOR2X1 NOR2X1_1510 ( .A(sqrto_111_), .B(u2__abc_52138_new_n13906_), .Y(u2__abc_52138_new_n13912_));
NOR2X1 NOR2X1_1511 ( .A(sqrto_112_), .B(u2__abc_52138_new_n13914_), .Y(u2__abc_52138_new_n13920_));
NOR2X1 NOR2X1_1512 ( .A(sqrto_113_), .B(u2__abc_52138_new_n13921_), .Y(u2__abc_52138_new_n13927_));
NOR2X1 NOR2X1_1513 ( .A(sqrto_114_), .B(u2__abc_52138_new_n13929_), .Y(u2__abc_52138_new_n13935_));
NOR2X1 NOR2X1_1514 ( .A(sqrto_115_), .B(u2__abc_52138_new_n13937_), .Y(u2__abc_52138_new_n13945_));
NOR2X1 NOR2X1_1515 ( .A(sqrto_116_), .B(u2__abc_52138_new_n13944_), .Y(u2__abc_52138_new_n13951_));
NOR2X1 NOR2X1_1516 ( .A(sqrto_117_), .B(u2__abc_52138_new_n13952_), .Y(u2__abc_52138_new_n13960_));
NOR2X1 NOR2X1_1517 ( .A(sqrto_118_), .B(u2__abc_52138_new_n13959_), .Y(u2__abc_52138_new_n13967_));
NOR2X1 NOR2X1_1518 ( .A(sqrto_119_), .B(u2__abc_52138_new_n13969_), .Y(u2__abc_52138_new_n13975_));
NOR2X1 NOR2X1_1519 ( .A(sqrto_120_), .B(u2__abc_52138_new_n13977_), .Y(u2__abc_52138_new_n13983_));
NOR2X1 NOR2X1_152 ( .A(sqrto_47_), .B(u2__abc_52138_new_n3298_), .Y(u2__abc_52138_new_n3299_));
NOR2X1 NOR2X1_1520 ( .A(sqrto_121_), .B(u2__abc_52138_new_n13984_), .Y(u2__abc_52138_new_n13992_));
NOR2X1 NOR2X1_1521 ( .A(sqrto_122_), .B(u2__abc_52138_new_n13991_), .Y(u2__abc_52138_new_n13998_));
NOR2X1 NOR2X1_1522 ( .A(sqrto_123_), .B(u2__abc_52138_new_n14000_), .Y(u2__abc_52138_new_n14006_));
NOR2X1 NOR2X1_1523 ( .A(sqrto_124_), .B(u2__abc_52138_new_n14008_), .Y(u2__abc_52138_new_n14014_));
NOR2X1 NOR2X1_1524 ( .A(sqrto_125_), .B(u2__abc_52138_new_n14015_), .Y(u2__abc_52138_new_n14023_));
NOR2X1 NOR2X1_1525 ( .A(sqrto_126_), .B(u2__abc_52138_new_n14022_), .Y(u2__abc_52138_new_n14029_));
NOR2X1 NOR2X1_1526 ( .A(sqrto_127_), .B(u2__abc_52138_new_n14031_), .Y(u2__abc_52138_new_n14037_));
NOR2X1 NOR2X1_1527 ( .A(sqrto_128_), .B(u2__abc_52138_new_n14039_), .Y(u2__abc_52138_new_n14045_));
NOR2X1 NOR2X1_1528 ( .A(sqrto_129_), .B(u2__abc_52138_new_n14046_), .Y(u2__abc_52138_new_n14052_));
NOR2X1 NOR2X1_1529 ( .A(sqrto_130_), .B(u2__abc_52138_new_n14054_), .Y(u2__abc_52138_new_n14061_));
NOR2X1 NOR2X1_153 ( .A(u2_remHi_47_), .B(u2__abc_52138_new_n3300_), .Y(u2__abc_52138_new_n3301_));
NOR2X1 NOR2X1_1530 ( .A(sqrto_131_), .B(u2__abc_52138_new_n14063_), .Y(u2__abc_52138_new_n14069_));
NOR2X1 NOR2X1_1531 ( .A(sqrto_132_), .B(u2__abc_52138_new_n14071_), .Y(u2__abc_52138_new_n14077_));
NOR2X1 NOR2X1_1532 ( .A(sqrto_133_), .B(u2__abc_52138_new_n14078_), .Y(u2__abc_52138_new_n14084_));
NOR2X1 NOR2X1_1533 ( .A(sqrto_134_), .B(u2__abc_52138_new_n14086_), .Y(u2__abc_52138_new_n14092_));
NOR2X1 NOR2X1_1534 ( .A(sqrto_135_), .B(u2__abc_52138_new_n14094_), .Y(u2__abc_52138_new_n14102_));
NOR2X1 NOR2X1_1535 ( .A(sqrto_136_), .B(u2__abc_52138_new_n14101_), .Y(u2__abc_52138_new_n14108_));
NOR2X1 NOR2X1_1536 ( .A(sqrto_137_), .B(u2__abc_52138_new_n14109_), .Y(u2__abc_52138_new_n14115_));
NOR2X1 NOR2X1_1537 ( .A(sqrto_138_), .B(u2__abc_52138_new_n14117_), .Y(u2__abc_52138_new_n14123_));
NOR2X1 NOR2X1_1538 ( .A(sqrto_139_), .B(u2__abc_52138_new_n14125_), .Y(u2__abc_52138_new_n14133_));
NOR2X1 NOR2X1_1539 ( .A(sqrto_140_), .B(u2__abc_52138_new_n14132_), .Y(u2__abc_52138_new_n14139_));
NOR2X1 NOR2X1_154 ( .A(u2__abc_52138_new_n3299_), .B(u2__abc_52138_new_n3301_), .Y(u2__abc_52138_new_n3302_));
NOR2X1 NOR2X1_1540 ( .A(sqrto_141_), .B(u2__abc_52138_new_n14140_), .Y(u2__abc_52138_new_n14148_));
NOR2X1 NOR2X1_1541 ( .A(sqrto_142_), .B(u2__abc_52138_new_n14147_), .Y(u2__abc_52138_new_n14154_));
NOR2X1 NOR2X1_1542 ( .A(sqrto_143_), .B(u2__abc_52138_new_n14156_), .Y(u2__abc_52138_new_n14162_));
NOR2X1 NOR2X1_1543 ( .A(sqrto_144_), .B(u2__abc_52138_new_n14164_), .Y(u2__abc_52138_new_n14170_));
NOR2X1 NOR2X1_1544 ( .A(sqrto_145_), .B(u2__abc_52138_new_n14171_), .Y(u2__abc_52138_new_n14177_));
NOR2X1 NOR2X1_1545 ( .A(sqrto_146_), .B(u2__abc_52138_new_n14179_), .Y(u2__abc_52138_new_n14185_));
NOR2X1 NOR2X1_1546 ( .A(sqrto_147_), .B(u2__abc_52138_new_n14187_), .Y(u2__abc_52138_new_n14195_));
NOR2X1 NOR2X1_1547 ( .A(sqrto_148_), .B(u2__abc_52138_new_n14194_), .Y(u2__abc_52138_new_n14201_));
NOR2X1 NOR2X1_1548 ( .A(sqrto_149_), .B(u2__abc_52138_new_n14202_), .Y(u2__abc_52138_new_n14210_));
NOR2X1 NOR2X1_1549 ( .A(sqrto_150_), .B(u2__abc_52138_new_n14209_), .Y(u2__abc_52138_new_n14216_));
NOR2X1 NOR2X1_155 ( .A(u2__abc_52138_new_n3297_), .B(u2__abc_52138_new_n3309_), .Y(u2__abc_52138_new_n3310_));
NOR2X1 NOR2X1_1550 ( .A(sqrto_151_), .B(u2__abc_52138_new_n14218_), .Y(u2__abc_52138_new_n14224_));
NOR2X1 NOR2X1_1551 ( .A(sqrto_152_), .B(u2__abc_52138_new_n14226_), .Y(u2__abc_52138_new_n14232_));
NOR2X1 NOR2X1_1552 ( .A(sqrto_153_), .B(u2__abc_52138_new_n14233_), .Y(u2__abc_52138_new_n14241_));
NOR2X1 NOR2X1_1553 ( .A(sqrto_154_), .B(u2__abc_52138_new_n14240_), .Y(u2__abc_52138_new_n14247_));
NOR2X1 NOR2X1_1554 ( .A(sqrto_155_), .B(u2__abc_52138_new_n14249_), .Y(u2__abc_52138_new_n14255_));
NOR2X1 NOR2X1_1555 ( .A(sqrto_156_), .B(u2__abc_52138_new_n14257_), .Y(u2__abc_52138_new_n14263_));
NOR2X1 NOR2X1_1556 ( .A(sqrto_157_), .B(u2__abc_52138_new_n14264_), .Y(u2__abc_52138_new_n14272_));
NOR2X1 NOR2X1_1557 ( .A(sqrto_158_), .B(u2__abc_52138_new_n14271_), .Y(u2__abc_52138_new_n14278_));
NOR2X1 NOR2X1_1558 ( .A(sqrto_159_), .B(u2__abc_52138_new_n14280_), .Y(u2__abc_52138_new_n14286_));
NOR2X1 NOR2X1_1559 ( .A(sqrto_160_), .B(u2__abc_52138_new_n14288_), .Y(u2__abc_52138_new_n14294_));
NOR2X1 NOR2X1_156 ( .A(u2__abc_52138_new_n3315_), .B(u2__abc_52138_new_n3320_), .Y(u2__abc_52138_new_n3321_));
NOR2X1 NOR2X1_1560 ( .A(sqrto_161_), .B(u2__abc_52138_new_n14295_), .Y(u2__abc_52138_new_n14301_));
NOR2X1 NOR2X1_1561 ( .A(sqrto_162_), .B(u2__abc_52138_new_n14303_), .Y(u2__abc_52138_new_n14309_));
NOR2X1 NOR2X1_1562 ( .A(sqrto_163_), .B(u2__abc_52138_new_n14311_), .Y(u2__abc_52138_new_n14319_));
NOR2X1 NOR2X1_1563 ( .A(sqrto_164_), .B(u2__abc_52138_new_n14318_), .Y(u2__abc_52138_new_n14325_));
NOR2X1 NOR2X1_1564 ( .A(sqrto_165_), .B(u2__abc_52138_new_n14326_), .Y(u2__abc_52138_new_n14334_));
NOR2X1 NOR2X1_1565 ( .A(sqrto_166_), .B(u2__abc_52138_new_n14333_), .Y(u2__abc_52138_new_n14340_));
NOR2X1 NOR2X1_1566 ( .A(sqrto_167_), .B(u2__abc_52138_new_n14342_), .Y(u2__abc_52138_new_n14348_));
NOR2X1 NOR2X1_1567 ( .A(sqrto_168_), .B(u2__abc_52138_new_n14350_), .Y(u2__abc_52138_new_n14356_));
NOR2X1 NOR2X1_1568 ( .A(sqrto_169_), .B(u2__abc_52138_new_n14357_), .Y(u2__abc_52138_new_n14365_));
NOR2X1 NOR2X1_1569 ( .A(sqrto_170_), .B(u2__abc_52138_new_n14364_), .Y(u2__abc_52138_new_n14371_));
NOR2X1 NOR2X1_157 ( .A(u2__abc_52138_new_n3326_), .B(u2__abc_52138_new_n3331_), .Y(u2__abc_52138_new_n3332_));
NOR2X1 NOR2X1_1570 ( .A(sqrto_171_), .B(u2__abc_52138_new_n14373_), .Y(u2__abc_52138_new_n14379_));
NOR2X1 NOR2X1_1571 ( .A(sqrto_172_), .B(u2__abc_52138_new_n14381_), .Y(u2__abc_52138_new_n14387_));
NOR2X1 NOR2X1_1572 ( .A(sqrto_173_), .B(u2__abc_52138_new_n14388_), .Y(u2__abc_52138_new_n14396_));
NOR2X1 NOR2X1_1573 ( .A(sqrto_174_), .B(u2__abc_52138_new_n14395_), .Y(u2__abc_52138_new_n14402_));
NOR2X1 NOR2X1_1574 ( .A(sqrto_175_), .B(u2__abc_52138_new_n14404_), .Y(u2__abc_52138_new_n14410_));
NOR2X1 NOR2X1_1575 ( .A(sqrto_176_), .B(u2__abc_52138_new_n14412_), .Y(u2__abc_52138_new_n14418_));
NOR2X1 NOR2X1_1576 ( .A(sqrto_177_), .B(u2__abc_52138_new_n14419_), .Y(u2__abc_52138_new_n14427_));
NOR2X1 NOR2X1_1577 ( .A(sqrto_178_), .B(u2__abc_52138_new_n14426_), .Y(u2__abc_52138_new_n14433_));
NOR2X1 NOR2X1_1578 ( .A(sqrto_179_), .B(u2__abc_52138_new_n14435_), .Y(u2__abc_52138_new_n14441_));
NOR2X1 NOR2X1_1579 ( .A(sqrto_180_), .B(u2__abc_52138_new_n14443_), .Y(u2__abc_52138_new_n14449_));
NOR2X1 NOR2X1_158 ( .A(u2__abc_52138_new_n3339_), .B(u2__abc_52138_new_n3344_), .Y(u2__abc_52138_new_n3345_));
NOR2X1 NOR2X1_1580 ( .A(sqrto_181_), .B(u2__abc_52138_new_n14450_), .Y(u2__abc_52138_new_n14458_));
NOR2X1 NOR2X1_1581 ( .A(sqrto_182_), .B(u2__abc_52138_new_n14457_), .Y(u2__abc_52138_new_n14464_));
NOR2X1 NOR2X1_1582 ( .A(sqrto_183_), .B(u2__abc_52138_new_n14466_), .Y(u2__abc_52138_new_n14472_));
NOR2X1 NOR2X1_1583 ( .A(sqrto_184_), .B(u2__abc_52138_new_n14474_), .Y(u2__abc_52138_new_n14480_));
NOR2X1 NOR2X1_1584 ( .A(sqrto_185_), .B(u2__abc_52138_new_n14481_), .Y(u2__abc_52138_new_n14489_));
NOR2X1 NOR2X1_1585 ( .A(sqrto_186_), .B(u2__abc_52138_new_n14488_), .Y(u2__abc_52138_new_n14495_));
NOR2X1 NOR2X1_1586 ( .A(sqrto_187_), .B(u2__abc_52138_new_n14497_), .Y(u2__abc_52138_new_n14503_));
NOR2X1 NOR2X1_1587 ( .A(sqrto_188_), .B(u2__abc_52138_new_n14505_), .Y(u2__abc_52138_new_n14511_));
NOR2X1 NOR2X1_1588 ( .A(sqrto_189_), .B(u2__abc_52138_new_n14512_), .Y(u2__abc_52138_new_n14520_));
NOR2X1 NOR2X1_1589 ( .A(sqrto_190_), .B(u2__abc_52138_new_n14519_), .Y(u2__abc_52138_new_n14526_));
NOR2X1 NOR2X1_159 ( .A(u2__abc_52138_new_n3350_), .B(u2__abc_52138_new_n3355_), .Y(u2__abc_52138_new_n3356_));
NOR2X1 NOR2X1_1590 ( .A(sqrto_191_), .B(u2__abc_52138_new_n14528_), .Y(u2__abc_52138_new_n14536_));
NOR2X1 NOR2X1_1591 ( .A(sqrto_192_), .B(u2__abc_52138_new_n14535_), .Y(u2__abc_52138_new_n14542_));
NOR2X1 NOR2X1_1592 ( .A(sqrto_193_), .B(u2__abc_52138_new_n14543_), .Y(u2__abc_52138_new_n14549_));
NOR2X1 NOR2X1_1593 ( .A(sqrto_194_), .B(u2__abc_52138_new_n14551_), .Y(u2__abc_52138_new_n14557_));
NOR2X1 NOR2X1_1594 ( .A(sqrto_195_), .B(u2__abc_52138_new_n14559_), .Y(u2__abc_52138_new_n14567_));
NOR2X1 NOR2X1_1595 ( .A(sqrto_196_), .B(u2__abc_52138_new_n14566_), .Y(u2__abc_52138_new_n14573_));
NOR2X1 NOR2X1_1596 ( .A(sqrto_197_), .B(u2__abc_52138_new_n14574_), .Y(u2__abc_52138_new_n14582_));
NOR2X1 NOR2X1_1597 ( .A(sqrto_198_), .B(u2__abc_52138_new_n14581_), .Y(u2__abc_52138_new_n14588_));
NOR2X1 NOR2X1_1598 ( .A(sqrto_199_), .B(u2__abc_52138_new_n14590_), .Y(u2__abc_52138_new_n14596_));
NOR2X1 NOR2X1_1599 ( .A(sqrto_200_), .B(u2__abc_52138_new_n14598_), .Y(u2__abc_52138_new_n14604_));
NOR2X1 NOR2X1_16 ( .A(_abc_65734_new_n1529_), .B(_abc_65734_new_n1515_), .Y(_abc_65734_new_n1530_));
NOR2X1 NOR2X1_160 ( .A(u2__abc_52138_new_n3362_), .B(u2__abc_52138_new_n3367_), .Y(u2__abc_52138_new_n3368_));
NOR2X1 NOR2X1_1600 ( .A(sqrto_201_), .B(u2__abc_52138_new_n14605_), .Y(u2__abc_52138_new_n14613_));
NOR2X1 NOR2X1_1601 ( .A(sqrto_202_), .B(u2__abc_52138_new_n14612_), .Y(u2__abc_52138_new_n14620_));
NOR2X1 NOR2X1_1602 ( .A(sqrto_203_), .B(u2__abc_52138_new_n14622_), .Y(u2__abc_52138_new_n14628_));
NOR2X1 NOR2X1_1603 ( .A(sqrto_204_), .B(u2__abc_52138_new_n14630_), .Y(u2__abc_52138_new_n14636_));
NOR2X1 NOR2X1_1604 ( .A(sqrto_205_), .B(u2__abc_52138_new_n14637_), .Y(u2__abc_52138_new_n14645_));
NOR2X1 NOR2X1_1605 ( .A(sqrto_206_), .B(u2__abc_52138_new_n14644_), .Y(u2__abc_52138_new_n14651_));
NOR2X1 NOR2X1_1606 ( .A(sqrto_207_), .B(u2__abc_52138_new_n14653_), .Y(u2__abc_52138_new_n14659_));
NOR2X1 NOR2X1_1607 ( .A(sqrto_208_), .B(u2__abc_52138_new_n14661_), .Y(u2__abc_52138_new_n14667_));
NOR2X1 NOR2X1_1608 ( .A(sqrto_209_), .B(u2__abc_52138_new_n14668_), .Y(u2__abc_52138_new_n14676_));
NOR2X1 NOR2X1_1609 ( .A(sqrto_210_), .B(u2__abc_52138_new_n14675_), .Y(u2__abc_52138_new_n14682_));
NOR2X1 NOR2X1_161 ( .A(u2__abc_52138_new_n3373_), .B(u2__abc_52138_new_n3378_), .Y(u2__abc_52138_new_n3379_));
NOR2X1 NOR2X1_1610 ( .A(sqrto_211_), .B(u2__abc_52138_new_n14684_), .Y(u2__abc_52138_new_n14690_));
NOR2X1 NOR2X1_1611 ( .A(sqrto_212_), .B(u2__abc_52138_new_n14692_), .Y(u2__abc_52138_new_n14698_));
NOR2X1 NOR2X1_1612 ( .A(sqrto_213_), .B(u2__abc_52138_new_n14699_), .Y(u2__abc_52138_new_n14707_));
NOR2X1 NOR2X1_1613 ( .A(sqrto_214_), .B(u2__abc_52138_new_n14706_), .Y(u2__abc_52138_new_n14713_));
NOR2X1 NOR2X1_1614 ( .A(sqrto_215_), .B(u2__abc_52138_new_n14715_), .Y(u2__abc_52138_new_n14721_));
NOR2X1 NOR2X1_1615 ( .A(sqrto_216_), .B(u2__abc_52138_new_n14723_), .Y(u2__abc_52138_new_n14729_));
NOR2X1 NOR2X1_1616 ( .A(sqrto_217_), .B(u2__abc_52138_new_n14730_), .Y(u2__abc_52138_new_n14738_));
NOR2X1 NOR2X1_1617 ( .A(sqrto_218_), .B(u2__abc_52138_new_n14737_), .Y(u2__abc_52138_new_n14744_));
NOR2X1 NOR2X1_1618 ( .A(sqrto_219_), .B(u2__abc_52138_new_n14746_), .Y(u2__abc_52138_new_n14752_));
NOR2X1 NOR2X1_1619 ( .A(sqrto_220_), .B(u2__abc_52138_new_n14754_), .Y(u2__abc_52138_new_n14760_));
NOR2X1 NOR2X1_162 ( .A(u2__abc_52138_new_n3357_), .B(u2__abc_52138_new_n3380_), .Y(u2__abc_52138_new_n3381_));
NOR2X1 NOR2X1_1620 ( .A(sqrto_221_), .B(u2__abc_52138_new_n14761_), .Y(u2__abc_52138_new_n14769_));
NOR2X1 NOR2X1_1621 ( .A(sqrto_222_), .B(u2__abc_52138_new_n14768_), .Y(u2__abc_52138_new_n14775_));
NOR2X1 NOR2X1_1622 ( .A(sqrto_223_), .B(u2__abc_52138_new_n14777_), .Y(u2__abc_52138_new_n14785_));
NOR2X1 NOR2X1_1623 ( .A(sqrto_224_), .B(u2__abc_52138_new_n14784_), .Y(u2__abc_52138_new_n14791_));
NOR2X1 NOR2X1_1624 ( .A(sqrto_225_), .B(u2__abc_52138_new_n14792_), .Y(u2__abc_52138_new_n14800_));
NOR2X1 NOR2X1_1625 ( .A(u2_o_226_), .B(u2__abc_52138_new_n14799_), .Y(u2__abc_52138_new_n14806_));
NOR2X1 NOR2X1_1626 ( .A(u2_o_227_), .B(u2__abc_52138_new_n14808_), .Y(u2__abc_52138_new_n14814_));
NOR2X1 NOR2X1_1627 ( .A(u2_o_228_), .B(u2__abc_52138_new_n14816_), .Y(u2__abc_52138_new_n14822_));
NOR2X1 NOR2X1_1628 ( .A(u2_o_229_), .B(u2__abc_52138_new_n14823_), .Y(u2__abc_52138_new_n14831_));
NOR2X1 NOR2X1_1629 ( .A(u2_o_230_), .B(u2__abc_52138_new_n14830_), .Y(u2__abc_52138_new_n14837_));
NOR2X1 NOR2X1_163 ( .A(u2__abc_52138_new_n3382_), .B(u2__abc_52138_new_n3387_), .Y(u2__abc_52138_new_n3388_));
NOR2X1 NOR2X1_1630 ( .A(u2_o_231_), .B(u2__abc_52138_new_n14839_), .Y(u2__abc_52138_new_n14845_));
NOR2X1 NOR2X1_1631 ( .A(u2_o_232_), .B(u2__abc_52138_new_n14847_), .Y(u2__abc_52138_new_n14853_));
NOR2X1 NOR2X1_1632 ( .A(u2_o_233_), .B(u2__abc_52138_new_n14854_), .Y(u2__abc_52138_new_n14862_));
NOR2X1 NOR2X1_1633 ( .A(u2_o_234_), .B(u2__abc_52138_new_n14861_), .Y(u2__abc_52138_new_n14868_));
NOR2X1 NOR2X1_1634 ( .A(u2_o_235_), .B(u2__abc_52138_new_n14870_), .Y(u2__abc_52138_new_n14876_));
NOR2X1 NOR2X1_1635 ( .A(u2_o_236_), .B(u2__abc_52138_new_n14878_), .Y(u2__abc_52138_new_n14884_));
NOR2X1 NOR2X1_1636 ( .A(u2_o_237_), .B(u2__abc_52138_new_n14885_), .Y(u2__abc_52138_new_n14893_));
NOR2X1 NOR2X1_1637 ( .A(u2_o_238_), .B(u2__abc_52138_new_n14892_), .Y(u2__abc_52138_new_n14899_));
NOR2X1 NOR2X1_1638 ( .A(u2_o_239_), .B(u2__abc_52138_new_n14901_), .Y(u2__abc_52138_new_n14909_));
NOR2X1 NOR2X1_1639 ( .A(u2_o_240_), .B(u2__abc_52138_new_n14908_), .Y(u2__abc_52138_new_n14915_));
NOR2X1 NOR2X1_164 ( .A(u2__abc_52138_new_n3393_), .B(u2__abc_52138_new_n3398_), .Y(u2__abc_52138_new_n3399_));
NOR2X1 NOR2X1_1640 ( .A(u2_o_241_), .B(u2__abc_52138_new_n14916_), .Y(u2__abc_52138_new_n14924_));
NOR2X1 NOR2X1_1641 ( .A(u2_o_242_), .B(u2__abc_52138_new_n14923_), .Y(u2__abc_52138_new_n14930_));
NOR2X1 NOR2X1_1642 ( .A(u2_o_243_), .B(u2__abc_52138_new_n14932_), .Y(u2__abc_52138_new_n14938_));
NOR2X1 NOR2X1_1643 ( .A(u2_o_244_), .B(u2__abc_52138_new_n14940_), .Y(u2__abc_52138_new_n14946_));
NOR2X1 NOR2X1_1644 ( .A(u2_o_245_), .B(u2__abc_52138_new_n14947_), .Y(u2__abc_52138_new_n14955_));
NOR2X1 NOR2X1_1645 ( .A(u2_o_246_), .B(u2__abc_52138_new_n14954_), .Y(u2__abc_52138_new_n14961_));
NOR2X1 NOR2X1_1646 ( .A(u2_o_247_), .B(u2__abc_52138_new_n14963_), .Y(u2__abc_52138_new_n14971_));
NOR2X1 NOR2X1_1647 ( .A(u2_o_248_), .B(u2__abc_52138_new_n14970_), .Y(u2__abc_52138_new_n14977_));
NOR2X1 NOR2X1_1648 ( .A(u2_o_249_), .B(u2__abc_52138_new_n14978_), .Y(u2__abc_52138_new_n14986_));
NOR2X1 NOR2X1_1649 ( .A(u2_o_250_), .B(u2__abc_52138_new_n14985_), .Y(u2__abc_52138_new_n14992_));
NOR2X1 NOR2X1_165 ( .A(u2__abc_52138_new_n3405_), .B(u2__abc_52138_new_n3410_), .Y(u2__abc_52138_new_n3411_));
NOR2X1 NOR2X1_1650 ( .A(u2_o_251_), .B(u2__abc_52138_new_n14994_), .Y(u2__abc_52138_new_n15002_));
NOR2X1 NOR2X1_1651 ( .A(u2_o_252_), .B(u2__abc_52138_new_n15001_), .Y(u2__abc_52138_new_n15008_));
NOR2X1 NOR2X1_1652 ( .A(u2_o_253_), .B(u2__abc_52138_new_n15009_), .Y(u2__abc_52138_new_n15017_));
NOR2X1 NOR2X1_1653 ( .A(u2_o_254_), .B(u2__abc_52138_new_n15016_), .Y(u2__abc_52138_new_n15023_));
NOR2X1 NOR2X1_1654 ( .A(u2_o_255_), .B(u2__abc_52138_new_n15025_), .Y(u2__abc_52138_new_n15033_));
NOR2X1 NOR2X1_1655 ( .A(u2_o_256_), .B(u2__abc_52138_new_n15032_), .Y(u2__abc_52138_new_n15039_));
NOR2X1 NOR2X1_1656 ( .A(u2_o_257_), .B(u2__abc_52138_new_n15040_), .Y(u2__abc_52138_new_n15046_));
NOR2X1 NOR2X1_1657 ( .A(u2_o_258_), .B(u2__abc_52138_new_n15048_), .Y(u2__abc_52138_new_n15054_));
NOR2X1 NOR2X1_1658 ( .A(u2_o_259_), .B(u2__abc_52138_new_n15056_), .Y(u2__abc_52138_new_n15064_));
NOR2X1 NOR2X1_1659 ( .A(u2_o_260_), .B(u2__abc_52138_new_n15063_), .Y(u2__abc_52138_new_n15070_));
NOR2X1 NOR2X1_166 ( .A(u2__abc_52138_new_n3400_), .B(u2__abc_52138_new_n3418_), .Y(u2__abc_52138_new_n3419_));
NOR2X1 NOR2X1_1660 ( .A(u2_o_261_), .B(u2__abc_52138_new_n15071_), .Y(u2__abc_52138_new_n15079_));
NOR2X1 NOR2X1_1661 ( .A(u2_o_262_), .B(u2__abc_52138_new_n15078_), .Y(u2__abc_52138_new_n15085_));
NOR2X1 NOR2X1_1662 ( .A(u2_o_263_), .B(u2__abc_52138_new_n15087_), .Y(u2__abc_52138_new_n15093_));
NOR2X1 NOR2X1_1663 ( .A(u2_o_264_), .B(u2__abc_52138_new_n15095_), .Y(u2__abc_52138_new_n15101_));
NOR2X1 NOR2X1_1664 ( .A(u2_o_265_), .B(u2__abc_52138_new_n15102_), .Y(u2__abc_52138_new_n15110_));
NOR2X1 NOR2X1_1665 ( .A(u2_o_266_), .B(u2__abc_52138_new_n15109_), .Y(u2__abc_52138_new_n15116_));
NOR2X1 NOR2X1_1666 ( .A(u2_o_267_), .B(u2__abc_52138_new_n15118_), .Y(u2__abc_52138_new_n15124_));
NOR2X1 NOR2X1_1667 ( .A(u2_o_268_), .B(u2__abc_52138_new_n15126_), .Y(u2__abc_52138_new_n15132_));
NOR2X1 NOR2X1_1668 ( .A(u2_o_269_), .B(u2__abc_52138_new_n15133_), .Y(u2__abc_52138_new_n15141_));
NOR2X1 NOR2X1_1669 ( .A(u2_o_270_), .B(u2__abc_52138_new_n15140_), .Y(u2__abc_52138_new_n15147_));
NOR2X1 NOR2X1_167 ( .A(u2__abc_52138_new_n3423_), .B(u2__abc_52138_new_n3422_), .Y(u2__abc_52138_new_n3424_));
NOR2X1 NOR2X1_1670 ( .A(u2_o_271_), .B(u2__abc_52138_new_n15149_), .Y(u2__abc_52138_new_n15155_));
NOR2X1 NOR2X1_1671 ( .A(u2_o_272_), .B(u2__abc_52138_new_n15157_), .Y(u2__abc_52138_new_n15163_));
NOR2X1 NOR2X1_1672 ( .A(u2_o_273_), .B(u2__abc_52138_new_n15164_), .Y(u2__abc_52138_new_n15172_));
NOR2X1 NOR2X1_1673 ( .A(u2_o_274_), .B(u2__abc_52138_new_n15171_), .Y(u2__abc_52138_new_n15178_));
NOR2X1 NOR2X1_1674 ( .A(u2_o_275_), .B(u2__abc_52138_new_n15180_), .Y(u2__abc_52138_new_n15186_));
NOR2X1 NOR2X1_1675 ( .A(u2_o_276_), .B(u2__abc_52138_new_n15188_), .Y(u2__abc_52138_new_n15194_));
NOR2X1 NOR2X1_1676 ( .A(u2_o_277_), .B(u2__abc_52138_new_n15195_), .Y(u2__abc_52138_new_n15203_));
NOR2X1 NOR2X1_1677 ( .A(u2_o_278_), .B(u2__abc_52138_new_n15202_), .Y(u2__abc_52138_new_n15209_));
NOR2X1 NOR2X1_1678 ( .A(u2_o_279_), .B(u2__abc_52138_new_n15211_), .Y(u2__abc_52138_new_n15217_));
NOR2X1 NOR2X1_1679 ( .A(u2_o_280_), .B(u2__abc_52138_new_n15219_), .Y(u2__abc_52138_new_n15225_));
NOR2X1 NOR2X1_168 ( .A(u2__abc_52138_new_n3429_), .B(u2__abc_52138_new_n3430_), .Y(u2__abc_52138_new_n3431_));
NOR2X1 NOR2X1_1680 ( .A(u2_o_281_), .B(u2__abc_52138_new_n15226_), .Y(u2__abc_52138_new_n15234_));
NOR2X1 NOR2X1_1681 ( .A(u2_o_282_), .B(u2__abc_52138_new_n15233_), .Y(u2__abc_52138_new_n15240_));
NOR2X1 NOR2X1_1682 ( .A(u2_o_283_), .B(u2__abc_52138_new_n15242_), .Y(u2__abc_52138_new_n15248_));
NOR2X1 NOR2X1_1683 ( .A(u2_o_284_), .B(u2__abc_52138_new_n15250_), .Y(u2__abc_52138_new_n15256_));
NOR2X1 NOR2X1_1684 ( .A(u2_o_285_), .B(u2__abc_52138_new_n15257_), .Y(u2__abc_52138_new_n15265_));
NOR2X1 NOR2X1_1685 ( .A(u2_o_286_), .B(u2__abc_52138_new_n15264_), .Y(u2__abc_52138_new_n15271_));
NOR2X1 NOR2X1_1686 ( .A(u2_o_287_), .B(u2__abc_52138_new_n15273_), .Y(u2__abc_52138_new_n15281_));
NOR2X1 NOR2X1_1687 ( .A(u2_o_288_), .B(u2__abc_52138_new_n15280_), .Y(u2__abc_52138_new_n15287_));
NOR2X1 NOR2X1_1688 ( .A(u2_o_289_), .B(u2__abc_52138_new_n15288_), .Y(u2__abc_52138_new_n15296_));
NOR2X1 NOR2X1_1689 ( .A(u2_o_290_), .B(u2__abc_52138_new_n15295_), .Y(u2__abc_52138_new_n15302_));
NOR2X1 NOR2X1_169 ( .A(u2_remHi_32_), .B(u2__abc_52138_new_n3437_), .Y(u2__abc_52138_new_n3438_));
NOR2X1 NOR2X1_1690 ( .A(u2_o_291_), .B(u2__abc_52138_new_n15304_), .Y(u2__abc_52138_new_n15310_));
NOR2X1 NOR2X1_1691 ( .A(u2_o_292_), .B(u2__abc_52138_new_n15312_), .Y(u2__abc_52138_new_n15318_));
NOR2X1 NOR2X1_1692 ( .A(u2_o_293_), .B(u2__abc_52138_new_n15319_), .Y(u2__abc_52138_new_n15327_));
NOR2X1 NOR2X1_1693 ( .A(u2_o_294_), .B(u2__abc_52138_new_n15326_), .Y(u2__abc_52138_new_n15333_));
NOR2X1 NOR2X1_1694 ( .A(u2_o_295_), .B(u2__abc_52138_new_n15335_), .Y(u2__abc_52138_new_n15341_));
NOR2X1 NOR2X1_1695 ( .A(u2_o_296_), .B(u2__abc_52138_new_n15343_), .Y(u2__abc_52138_new_n15349_));
NOR2X1 NOR2X1_1696 ( .A(u2_o_297_), .B(u2__abc_52138_new_n15350_), .Y(u2__abc_52138_new_n15358_));
NOR2X1 NOR2X1_1697 ( .A(u2_o_298_), .B(u2__abc_52138_new_n15357_), .Y(u2__abc_52138_new_n15364_));
NOR2X1 NOR2X1_1698 ( .A(u2_o_299_), .B(u2__abc_52138_new_n15366_), .Y(u2__abc_52138_new_n15372_));
NOR2X1 NOR2X1_1699 ( .A(u2_o_300_), .B(u2__abc_52138_new_n15374_), .Y(u2__abc_52138_new_n15380_));
NOR2X1 NOR2X1_17 ( .A(_abc_65734_new_n1540_), .B(_abc_65734_new_n1528_), .Y(_abc_65734_new_n1541_));
NOR2X1 NOR2X1_170 ( .A(sqrto_41_), .B(u2__abc_52138_new_n3342_), .Y(u2__abc_52138_new_n3456_));
NOR2X1 NOR2X1_1700 ( .A(u2_o_301_), .B(u2__abc_52138_new_n15381_), .Y(u2__abc_52138_new_n15389_));
NOR2X1 NOR2X1_1701 ( .A(u2_o_302_), .B(u2__abc_52138_new_n15388_), .Y(u2__abc_52138_new_n15395_));
NOR2X1 NOR2X1_1702 ( .A(u2_o_303_), .B(u2__abc_52138_new_n15397_), .Y(u2__abc_52138_new_n15405_));
NOR2X1 NOR2X1_1703 ( .A(u2_o_304_), .B(u2__abc_52138_new_n15404_), .Y(u2__abc_52138_new_n15411_));
NOR2X1 NOR2X1_1704 ( .A(u2_o_305_), .B(u2__abc_52138_new_n15412_), .Y(u2__abc_52138_new_n15420_));
NOR2X1 NOR2X1_1705 ( .A(u2_o_306_), .B(u2__abc_52138_new_n15419_), .Y(u2__abc_52138_new_n15426_));
NOR2X1 NOR2X1_1706 ( .A(u2_o_307_), .B(u2__abc_52138_new_n15428_), .Y(u2__abc_52138_new_n15434_));
NOR2X1 NOR2X1_1707 ( .A(u2_o_308_), .B(u2__abc_52138_new_n15436_), .Y(u2__abc_52138_new_n15442_));
NOR2X1 NOR2X1_1708 ( .A(u2_o_309_), .B(u2__abc_52138_new_n15443_), .Y(u2__abc_52138_new_n15451_));
NOR2X1 NOR2X1_1709 ( .A(u2_o_310_), .B(u2__abc_52138_new_n15450_), .Y(u2__abc_52138_new_n15457_));
NOR2X1 NOR2X1_171 ( .A(sqrto_51_), .B(u2__abc_52138_new_n3324_), .Y(u2__abc_52138_new_n3478_));
NOR2X1 NOR2X1_1710 ( .A(u2_o_311_), .B(u2__abc_52138_new_n15459_), .Y(u2__abc_52138_new_n15467_));
NOR2X1 NOR2X1_1711 ( .A(u2_o_312_), .B(u2__abc_52138_new_n15466_), .Y(u2__abc_52138_new_n15473_));
NOR2X1 NOR2X1_1712 ( .A(u2_o_313_), .B(u2__abc_52138_new_n15474_), .Y(u2__abc_52138_new_n15482_));
NOR2X1 NOR2X1_1713 ( .A(u2_o_314_), .B(u2__abc_52138_new_n15481_), .Y(u2__abc_52138_new_n15489_));
NOR2X1 NOR2X1_1714 ( .A(u2_o_315_), .B(u2__abc_52138_new_n15491_), .Y(u2__abc_52138_new_n15499_));
NOR2X1 NOR2X1_1715 ( .A(u2_o_316_), .B(u2__abc_52138_new_n15498_), .Y(u2__abc_52138_new_n15505_));
NOR2X1 NOR2X1_1716 ( .A(u2_o_317_), .B(u2__abc_52138_new_n15506_), .Y(u2__abc_52138_new_n15514_));
NOR2X1 NOR2X1_1717 ( .A(u2_o_318_), .B(u2__abc_52138_new_n15513_), .Y(u2__abc_52138_new_n15520_));
NOR2X1 NOR2X1_1718 ( .A(u2_o_319_), .B(u2__abc_52138_new_n15522_), .Y(u2__abc_52138_new_n15530_));
NOR2X1 NOR2X1_1719 ( .A(u2_o_320_), .B(u2__abc_52138_new_n15529_), .Y(u2__abc_52138_new_n15536_));
NOR2X1 NOR2X1_172 ( .A(sqrto_118_), .B(u2__abc_52138_new_n3503_), .Y(u2__abc_52138_new_n3504_));
NOR2X1 NOR2X1_1720 ( .A(u2_o_321_), .B(u2__abc_52138_new_n15537_), .Y(u2__abc_52138_new_n15545_));
NOR2X1 NOR2X1_1721 ( .A(u2_o_322_), .B(u2__abc_52138_new_n15544_), .Y(u2__abc_52138_new_n15551_));
NOR2X1 NOR2X1_1722 ( .A(u2_o_323_), .B(u2__abc_52138_new_n15553_), .Y(u2__abc_52138_new_n15559_));
NOR2X1 NOR2X1_1723 ( .A(u2_o_324_), .B(u2__abc_52138_new_n15561_), .Y(u2__abc_52138_new_n15567_));
NOR2X1 NOR2X1_1724 ( .A(u2_o_325_), .B(u2__abc_52138_new_n15568_), .Y(u2__abc_52138_new_n15576_));
NOR2X1 NOR2X1_1725 ( .A(u2_o_326_), .B(u2__abc_52138_new_n15575_), .Y(u2__abc_52138_new_n15582_));
NOR2X1 NOR2X1_1726 ( .A(u2_o_327_), .B(u2__abc_52138_new_n15584_), .Y(u2__abc_52138_new_n15590_));
NOR2X1 NOR2X1_1727 ( .A(u2_o_328_), .B(u2__abc_52138_new_n15592_), .Y(u2__abc_52138_new_n15598_));
NOR2X1 NOR2X1_1728 ( .A(u2_o_329_), .B(u2__abc_52138_new_n15599_), .Y(u2__abc_52138_new_n15607_));
NOR2X1 NOR2X1_1729 ( .A(u2_o_330_), .B(u2__abc_52138_new_n15606_), .Y(u2__abc_52138_new_n15613_));
NOR2X1 NOR2X1_173 ( .A(sqrto_119_), .B(u2__abc_52138_new_n3508_), .Y(u2__abc_52138_new_n3509_));
NOR2X1 NOR2X1_1730 ( .A(u2_o_331_), .B(u2__abc_52138_new_n15615_), .Y(u2__abc_52138_new_n15621_));
NOR2X1 NOR2X1_1731 ( .A(u2_o_332_), .B(u2__abc_52138_new_n15623_), .Y(u2__abc_52138_new_n15629_));
NOR2X1 NOR2X1_1732 ( .A(u2_o_333_), .B(u2__abc_52138_new_n15630_), .Y(u2__abc_52138_new_n15638_));
NOR2X1 NOR2X1_1733 ( .A(u2_o_334_), .B(u2__abc_52138_new_n15637_), .Y(u2__abc_52138_new_n15645_));
NOR2X1 NOR2X1_1734 ( .A(u2_o_335_), .B(u2__abc_52138_new_n15647_), .Y(u2__abc_52138_new_n15655_));
NOR2X1 NOR2X1_1735 ( .A(u2_o_336_), .B(u2__abc_52138_new_n15654_), .Y(u2__abc_52138_new_n15661_));
NOR2X1 NOR2X1_1736 ( .A(u2_o_337_), .B(u2__abc_52138_new_n15662_), .Y(u2__abc_52138_new_n15670_));
NOR2X1 NOR2X1_1737 ( .A(u2_o_338_), .B(u2__abc_52138_new_n15669_), .Y(u2__abc_52138_new_n15677_));
NOR2X1 NOR2X1_1738 ( .A(u2_o_339_), .B(u2__abc_52138_new_n15679_), .Y(u2__abc_52138_new_n15685_));
NOR2X1 NOR2X1_1739 ( .A(u2_o_340_), .B(u2__abc_52138_new_n15687_), .Y(u2__abc_52138_new_n15693_));
NOR2X1 NOR2X1_174 ( .A(u2_remHi_119_), .B(u2__abc_52138_new_n3511_), .Y(u2__abc_52138_new_n3512_));
NOR2X1 NOR2X1_1740 ( .A(u2_o_341_), .B(u2__abc_52138_new_n15694_), .Y(u2__abc_52138_new_n15702_));
NOR2X1 NOR2X1_1741 ( .A(u2_o_342_), .B(u2__abc_52138_new_n15701_), .Y(u2__abc_52138_new_n15708_));
NOR2X1 NOR2X1_1742 ( .A(u2_o_343_), .B(u2__abc_52138_new_n15710_), .Y(u2__abc_52138_new_n15718_));
NOR2X1 NOR2X1_1743 ( .A(u2_o_344_), .B(u2__abc_52138_new_n15717_), .Y(u2__abc_52138_new_n15724_));
NOR2X1 NOR2X1_1744 ( .A(u2_o_345_), .B(u2__abc_52138_new_n15725_), .Y(u2__abc_52138_new_n15733_));
NOR2X1 NOR2X1_1745 ( .A(u2_o_346_), .B(u2__abc_52138_new_n15732_), .Y(u2__abc_52138_new_n15739_));
NOR2X1 NOR2X1_1746 ( .A(u2_o_347_), .B(u2__abc_52138_new_n15741_), .Y(u2__abc_52138_new_n15749_));
NOR2X1 NOR2X1_1747 ( .A(u2_o_348_), .B(u2__abc_52138_new_n15748_), .Y(u2__abc_52138_new_n15755_));
NOR2X1 NOR2X1_1748 ( .A(u2_o_349_), .B(u2__abc_52138_new_n15756_), .Y(u2__abc_52138_new_n15764_));
NOR2X1 NOR2X1_1749 ( .A(u2_o_350_), .B(u2__abc_52138_new_n15763_), .Y(u2__abc_52138_new_n15770_));
NOR2X1 NOR2X1_175 ( .A(u2__abc_52138_new_n3507_), .B(u2__abc_52138_new_n3514_), .Y(u2__abc_52138_new_n3515_));
NOR2X1 NOR2X1_1750 ( .A(u2_o_351_), .B(u2__abc_52138_new_n15772_), .Y(u2__abc_52138_new_n15780_));
NOR2X1 NOR2X1_1751 ( .A(u2_o_352_), .B(u2__abc_52138_new_n15779_), .Y(u2__abc_52138_new_n15786_));
NOR2X1 NOR2X1_1752 ( .A(u2_o_353_), .B(u2__abc_52138_new_n15787_), .Y(u2__abc_52138_new_n15795_));
NOR2X1 NOR2X1_1753 ( .A(u2_o_354_), .B(u2__abc_52138_new_n15794_), .Y(u2__abc_52138_new_n15801_));
NOR2X1 NOR2X1_1754 ( .A(u2_o_355_), .B(u2__abc_52138_new_n15803_), .Y(u2__abc_52138_new_n15809_));
NOR2X1 NOR2X1_1755 ( .A(u2_o_356_), .B(u2__abc_52138_new_n15811_), .Y(u2__abc_52138_new_n15817_));
NOR2X1 NOR2X1_1756 ( .A(u2_o_357_), .B(u2__abc_52138_new_n15818_), .Y(u2__abc_52138_new_n15826_));
NOR2X1 NOR2X1_1757 ( .A(u2_o_358_), .B(u2__abc_52138_new_n15825_), .Y(u2__abc_52138_new_n15832_));
NOR2X1 NOR2X1_1758 ( .A(u2_o_359_), .B(u2__abc_52138_new_n15834_), .Y(u2__abc_52138_new_n15842_));
NOR2X1 NOR2X1_1759 ( .A(u2_o_360_), .B(u2__abc_52138_new_n15841_), .Y(u2__abc_52138_new_n15848_));
NOR2X1 NOR2X1_176 ( .A(u2__abc_52138_new_n3520_), .B(u2__abc_52138_new_n3525_), .Y(u2__abc_52138_new_n3526_));
NOR2X1 NOR2X1_1760 ( .A(u2_o_361_), .B(u2__abc_52138_new_n15849_), .Y(u2__abc_52138_new_n15857_));
NOR2X1 NOR2X1_1761 ( .A(u2_o_362_), .B(u2__abc_52138_new_n15856_), .Y(u2__abc_52138_new_n15863_));
NOR2X1 NOR2X1_1762 ( .A(u2_o_363_), .B(u2__abc_52138_new_n15865_), .Y(u2__abc_52138_new_n15873_));
NOR2X1 NOR2X1_1763 ( .A(u2_o_364_), .B(u2__abc_52138_new_n15872_), .Y(u2__abc_52138_new_n15879_));
NOR2X1 NOR2X1_1764 ( .A(u2_o_365_), .B(u2__abc_52138_new_n15880_), .Y(u2__abc_52138_new_n15888_));
NOR2X1 NOR2X1_1765 ( .A(u2_o_366_), .B(u2__abc_52138_new_n15887_), .Y(u2__abc_52138_new_n15894_));
NOR2X1 NOR2X1_1766 ( .A(u2_o_367_), .B(u2__abc_52138_new_n15896_), .Y(u2__abc_52138_new_n15904_));
NOR2X1 NOR2X1_1767 ( .A(u2_o_368_), .B(u2__abc_52138_new_n15903_), .Y(u2__abc_52138_new_n15910_));
NOR2X1 NOR2X1_1768 ( .A(u2_o_369_), .B(u2__abc_52138_new_n15911_), .Y(u2__abc_52138_new_n15920_));
NOR2X1 NOR2X1_1769 ( .A(u2_o_370_), .B(u2__abc_52138_new_n15919_), .Y(u2__abc_52138_new_n15926_));
NOR2X1 NOR2X1_177 ( .A(sqrto_122_), .B(u2__abc_52138_new_n3542_), .Y(u2__abc_52138_new_n3543_));
NOR2X1 NOR2X1_1770 ( .A(u2_o_371_), .B(u2__abc_52138_new_n15928_), .Y(u2__abc_52138_new_n15936_));
NOR2X1 NOR2X1_1771 ( .A(u2_o_372_), .B(u2__abc_52138_new_n15935_), .Y(u2__abc_52138_new_n15942_));
NOR2X1 NOR2X1_1772 ( .A(u2_o_373_), .B(u2__abc_52138_new_n15943_), .Y(u2__abc_52138_new_n15951_));
NOR2X1 NOR2X1_1773 ( .A(u2_o_374_), .B(u2__abc_52138_new_n15950_), .Y(u2__abc_52138_new_n15957_));
NOR2X1 NOR2X1_1774 ( .A(u2_o_375_), .B(u2__abc_52138_new_n15959_), .Y(u2__abc_52138_new_n15967_));
NOR2X1 NOR2X1_1775 ( .A(u2_o_376_), .B(u2__abc_52138_new_n15966_), .Y(u2__abc_52138_new_n15973_));
NOR2X1 NOR2X1_1776 ( .A(u2_o_377_), .B(u2__abc_52138_new_n15974_), .Y(u2__abc_52138_new_n15982_));
NOR2X1 NOR2X1_1777 ( .A(u2_o_378_), .B(u2__abc_52138_new_n15981_), .Y(u2__abc_52138_new_n15988_));
NOR2X1 NOR2X1_1778 ( .A(u2_o_379_), .B(u2__abc_52138_new_n15990_), .Y(u2__abc_52138_new_n15998_));
NOR2X1 NOR2X1_1779 ( .A(u2_o_380_), .B(u2__abc_52138_new_n15997_), .Y(u2__abc_52138_new_n16004_));
NOR2X1 NOR2X1_178 ( .A(u2_remHi_122_), .B(u2__abc_52138_new_n3544_), .Y(u2__abc_52138_new_n3545_));
NOR2X1 NOR2X1_1780 ( .A(u2_o_381_), .B(u2__abc_52138_new_n16005_), .Y(u2__abc_52138_new_n16013_));
NOR2X1 NOR2X1_1781 ( .A(u2_o_382_), .B(u2__abc_52138_new_n16012_), .Y(u2__abc_52138_new_n16019_));
NOR2X1 NOR2X1_1782 ( .A(u2_o_383_), .B(u2__abc_52138_new_n16021_), .Y(u2__abc_52138_new_n16029_));
NOR2X1 NOR2X1_1783 ( .A(u2_o_384_), .B(u2__abc_52138_new_n16028_), .Y(u2__abc_52138_new_n16035_));
NOR2X1 NOR2X1_1784 ( .A(u2_o_385_), .B(u2__abc_52138_new_n16036_), .Y(u2__abc_52138_new_n16044_));
NOR2X1 NOR2X1_1785 ( .A(u2_o_386_), .B(u2__abc_52138_new_n16043_), .Y(u2__abc_52138_new_n16050_));
NOR2X1 NOR2X1_1786 ( .A(u2_o_387_), .B(u2__abc_52138_new_n16052_), .Y(u2__abc_52138_new_n16058_));
NOR2X1 NOR2X1_1787 ( .A(u2_o_388_), .B(u2__abc_52138_new_n16060_), .Y(u2__abc_52138_new_n16066_));
NOR2X1 NOR2X1_1788 ( .A(u2_o_389_), .B(u2__abc_52138_new_n16067_), .Y(u2__abc_52138_new_n16075_));
NOR2X1 NOR2X1_1789 ( .A(u2_o_390_), .B(u2__abc_52138_new_n16074_), .Y(u2__abc_52138_new_n16082_));
NOR2X1 NOR2X1_179 ( .A(u2__abc_52138_new_n3543_), .B(u2__abc_52138_new_n3545_), .Y(u2__abc_52138_new_n3546_));
NOR2X1 NOR2X1_1790 ( .A(u2_o_391_), .B(u2__abc_52138_new_n16084_), .Y(u2__abc_52138_new_n16091_));
NOR2X1 NOR2X1_1791 ( .A(u2_o_392_), .B(u2__abc_52138_new_n16093_), .Y(u2__abc_52138_new_n16099_));
NOR2X1 NOR2X1_1792 ( .A(u2_o_393_), .B(u2__abc_52138_new_n16100_), .Y(u2__abc_52138_new_n16108_));
NOR2X1 NOR2X1_1793 ( .A(u2_o_394_), .B(u2__abc_52138_new_n16107_), .Y(u2__abc_52138_new_n16115_));
NOR2X1 NOR2X1_1794 ( .A(u2_o_395_), .B(u2__abc_52138_new_n16117_), .Y(u2__abc_52138_new_n16123_));
NOR2X1 NOR2X1_1795 ( .A(u2_o_396_), .B(u2__abc_52138_new_n16125_), .Y(u2__abc_52138_new_n16131_));
NOR2X1 NOR2X1_1796 ( .A(u2_o_397_), .B(u2__abc_52138_new_n16132_), .Y(u2__abc_52138_new_n16140_));
NOR2X1 NOR2X1_1797 ( .A(u2_o_398_), .B(u2__abc_52138_new_n16139_), .Y(u2__abc_52138_new_n16146_));
NOR2X1 NOR2X1_1798 ( .A(u2_o_399_), .B(u2__abc_52138_new_n16148_), .Y(u2__abc_52138_new_n16156_));
NOR2X1 NOR2X1_1799 ( .A(u2_o_400_), .B(u2__abc_52138_new_n16155_), .Y(u2__abc_52138_new_n16162_));
NOR2X1 NOR2X1_18 ( .A(_abc_65734_new_n1523_), .B(_abc_65734_new_n1516_), .Y(_abc_65734_new_n1580_));
NOR2X1 NOR2X1_180 ( .A(u2__abc_52138_new_n3537_), .B(u2__abc_52138_new_n3547_), .Y(u2__abc_52138_new_n3548_));
NOR2X1 NOR2X1_1800 ( .A(u2_o_401_), .B(u2__abc_52138_new_n16163_), .Y(u2__abc_52138_new_n16171_));
NOR2X1 NOR2X1_1801 ( .A(u2_o_402_), .B(u2__abc_52138_new_n16170_), .Y(u2__abc_52138_new_n16177_));
NOR2X1 NOR2X1_1802 ( .A(u2_o_403_), .B(u2__abc_52138_new_n16179_), .Y(u2__abc_52138_new_n16185_));
NOR2X1 NOR2X1_1803 ( .A(u2_o_404_), .B(u2__abc_52138_new_n16187_), .Y(u2__abc_52138_new_n16193_));
NOR2X1 NOR2X1_1804 ( .A(u2_o_405_), .B(u2__abc_52138_new_n16194_), .Y(u2__abc_52138_new_n16202_));
NOR2X1 NOR2X1_1805 ( .A(u2_o_406_), .B(u2__abc_52138_new_n16201_), .Y(u2__abc_52138_new_n16208_));
NOR2X1 NOR2X1_1806 ( .A(u2_o_407_), .B(u2__abc_52138_new_n16210_), .Y(u2__abc_52138_new_n16218_));
NOR2X1 NOR2X1_1807 ( .A(u2_o_408_), .B(u2__abc_52138_new_n16217_), .Y(u2__abc_52138_new_n16224_));
NOR2X1 NOR2X1_1808 ( .A(u2_o_409_), .B(u2__abc_52138_new_n16225_), .Y(u2__abc_52138_new_n16233_));
NOR2X1 NOR2X1_1809 ( .A(u2_o_410_), .B(u2__abc_52138_new_n16232_), .Y(u2__abc_52138_new_n16239_));
NOR2X1 NOR2X1_181 ( .A(u2__abc_52138_new_n3554_), .B(u2__abc_52138_new_n3559_), .Y(u2__abc_52138_new_n3560_));
NOR2X1 NOR2X1_1810 ( .A(u2_o_411_), .B(u2__abc_52138_new_n16241_), .Y(u2__abc_52138_new_n16249_));
NOR2X1 NOR2X1_1811 ( .A(u2_o_412_), .B(u2__abc_52138_new_n16248_), .Y(u2__abc_52138_new_n16255_));
NOR2X1 NOR2X1_1812 ( .A(u2_o_413_), .B(u2__abc_52138_new_n16256_), .Y(u2__abc_52138_new_n16264_));
NOR2X1 NOR2X1_1813 ( .A(u2_o_414_), .B(u2__abc_52138_new_n16263_), .Y(u2__abc_52138_new_n16270_));
NOR2X1 NOR2X1_1814 ( .A(u2_o_415_), .B(u2__abc_52138_new_n16272_), .Y(u2__abc_52138_new_n16280_));
NOR2X1 NOR2X1_1815 ( .A(u2_o_416_), .B(u2__abc_52138_new_n16279_), .Y(u2__abc_52138_new_n16286_));
NOR2X1 NOR2X1_1816 ( .A(u2_o_417_), .B(u2__abc_52138_new_n16287_), .Y(u2__abc_52138_new_n16295_));
NOR2X1 NOR2X1_1817 ( .A(u2_o_418_), .B(u2__abc_52138_new_n16294_), .Y(u2__abc_52138_new_n16301_));
NOR2X1 NOR2X1_1818 ( .A(u2_o_419_), .B(u2__abc_52138_new_n16303_), .Y(u2__abc_52138_new_n16309_));
NOR2X1 NOR2X1_1819 ( .A(u2_o_420_), .B(u2__abc_52138_new_n16311_), .Y(u2__abc_52138_new_n16317_));
NOR2X1 NOR2X1_182 ( .A(u2__abc_52138_new_n3565_), .B(u2__abc_52138_new_n3570_), .Y(u2__abc_52138_new_n3571_));
NOR2X1 NOR2X1_1820 ( .A(u2_o_421_), .B(u2__abc_52138_new_n16318_), .Y(u2__abc_52138_new_n16326_));
NOR2X1 NOR2X1_1821 ( .A(u2_o_422_), .B(u2__abc_52138_new_n16325_), .Y(u2__abc_52138_new_n16332_));
NOR2X1 NOR2X1_1822 ( .A(u2_o_423_), .B(u2__abc_52138_new_n16334_), .Y(u2__abc_52138_new_n16342_));
NOR2X1 NOR2X1_1823 ( .A(u2_o_424_), .B(u2__abc_52138_new_n16341_), .Y(u2__abc_52138_new_n16348_));
NOR2X1 NOR2X1_1824 ( .A(u2_o_425_), .B(u2__abc_52138_new_n16349_), .Y(u2__abc_52138_new_n16357_));
NOR2X1 NOR2X1_1825 ( .A(u2_o_426_), .B(u2__abc_52138_new_n16356_), .Y(u2__abc_52138_new_n16363_));
NOR2X1 NOR2X1_1826 ( .A(u2_o_427_), .B(u2__abc_52138_new_n16365_), .Y(u2__abc_52138_new_n16373_));
NOR2X1 NOR2X1_1827 ( .A(u2_o_428_), .B(u2__abc_52138_new_n16372_), .Y(u2__abc_52138_new_n16379_));
NOR2X1 NOR2X1_1828 ( .A(u2_o_429_), .B(u2__abc_52138_new_n16380_), .Y(u2__abc_52138_new_n16388_));
NOR2X1 NOR2X1_1829 ( .A(u2_o_430_), .B(u2__abc_52138_new_n16387_), .Y(u2__abc_52138_new_n16394_));
NOR2X1 NOR2X1_183 ( .A(sqrto_116_), .B(u2__abc_52138_new_n3573_), .Y(u2__abc_52138_new_n3574_));
NOR2X1 NOR2X1_1830 ( .A(u2_o_431_), .B(u2__abc_52138_new_n16396_), .Y(u2__abc_52138_new_n16404_));
NOR2X1 NOR2X1_1831 ( .A(u2_o_432_), .B(u2__abc_52138_new_n16403_), .Y(u2__abc_52138_new_n16410_));
NOR2X1 NOR2X1_1832 ( .A(u2_o_433_), .B(u2__abc_52138_new_n16411_), .Y(u2__abc_52138_new_n16419_));
NOR2X1 NOR2X1_1833 ( .A(u2_o_434_), .B(u2__abc_52138_new_n16418_), .Y(u2__abc_52138_new_n16425_));
NOR2X1 NOR2X1_1834 ( .A(u2_o_435_), .B(u2__abc_52138_new_n16427_), .Y(u2__abc_52138_new_n16435_));
NOR2X1 NOR2X1_1835 ( .A(u2_o_436_), .B(u2__abc_52138_new_n16434_), .Y(u2__abc_52138_new_n16441_));
NOR2X1 NOR2X1_1836 ( .A(u2_o_437_), .B(u2__abc_52138_new_n16442_), .Y(u2__abc_52138_new_n16450_));
NOR2X1 NOR2X1_1837 ( .A(u2_o_438_), .B(u2__abc_52138_new_n16449_), .Y(u2__abc_52138_new_n16456_));
NOR2X1 NOR2X1_1838 ( .A(u2_o_439_), .B(u2__abc_52138_new_n16458_), .Y(u2__abc_52138_new_n16466_));
NOR2X1 NOR2X1_1839 ( .A(u2_o_440_), .B(u2__abc_52138_new_n16465_), .Y(u2__abc_52138_new_n16472_));
NOR2X1 NOR2X1_184 ( .A(u2_remHi_116_), .B(u2__abc_52138_new_n3575_), .Y(u2__abc_52138_new_n3576_));
NOR2X1 NOR2X1_1840 ( .A(u2_o_441_), .B(u2__abc_52138_new_n16473_), .Y(u2__abc_52138_new_n16481_));
NOR2X1 NOR2X1_1841 ( .A(u2_o_442_), .B(u2__abc_52138_new_n16480_), .Y(u2__abc_52138_new_n16487_));
NOR2X1 NOR2X1_1842 ( .A(u2_o_443_), .B(u2__abc_52138_new_n16489_), .Y(u2__abc_52138_new_n16497_));
NOR2X1 NOR2X1_1843 ( .A(u2_o_444_), .B(u2__abc_52138_new_n16496_), .Y(u2__abc_52138_new_n16503_));
NOR2X1 NOR2X1_1844 ( .A(u2_o_445_), .B(u2__abc_52138_new_n16504_), .Y(u2__abc_52138_new_n16512_));
NOR2X1 NOR2X1_1845 ( .A(u2_o_446_), .B(u2__abc_52138_new_n16511_), .Y(u2__abc_52138_new_n16518_));
NOR2X1 NOR2X1_1846 ( .A(u2_o_447_), .B(u2__abc_52138_new_n16520_), .Y(u2__abc_52138_new_n16526_));
NOR2X1 NOR2X1_1847 ( .A(u2_o_448_), .B(u2__abc_52138_new_n16528_), .Y(u2__abc_52138_new_n16534_));
NOR2X1 NOR2X1_185 ( .A(u2__abc_52138_new_n3574_), .B(u2__abc_52138_new_n3576_), .Y(u2__abc_52138_new_n3577_));
NOR2X1 NOR2X1_186 ( .A(u2__abc_52138_new_n3593_), .B(u2__abc_52138_new_n3582_), .Y(u2__abc_52138_new_n3594_));
NOR2X1 NOR2X1_187 ( .A(u2__abc_52138_new_n3595_), .B(u2__abc_52138_new_n3549_), .Y(u2__abc_52138_new_n3596_));
NOR2X1 NOR2X1_188 ( .A(sqrto_102_), .B(u2__abc_52138_new_n3612_), .Y(u2__abc_52138_new_n3613_));
NOR2X1 NOR2X1_189 ( .A(u2_remHi_102_), .B(u2__abc_52138_new_n3614_), .Y(u2__abc_52138_new_n3615_));
NOR2X1 NOR2X1_19 ( .A(\a[121] ), .B(\a[122] ), .Y(u1__abc_51895_new_n137_));
NOR2X1 NOR2X1_190 ( .A(u2__abc_52138_new_n3613_), .B(u2__abc_52138_new_n3615_), .Y(u2__abc_52138_new_n3616_));
NOR2X1 NOR2X1_191 ( .A(u2__abc_52138_new_n3607_), .B(u2__abc_52138_new_n3617_), .Y(u2__abc_52138_new_n3618_));
NOR2X1 NOR2X1_192 ( .A(sqrto_106_), .B(u2__abc_52138_new_n3634_), .Y(u2__abc_52138_new_n3635_));
NOR2X1 NOR2X1_193 ( .A(u2_remHi_106_), .B(u2__abc_52138_new_n3636_), .Y(u2__abc_52138_new_n3637_));
NOR2X1 NOR2X1_194 ( .A(u2__abc_52138_new_n3635_), .B(u2__abc_52138_new_n3637_), .Y(u2__abc_52138_new_n3638_));
NOR2X1 NOR2X1_195 ( .A(u2__abc_52138_new_n3629_), .B(u2__abc_52138_new_n3639_), .Y(u2__abc_52138_new_n3640_));
NOR2X1 NOR2X1_196 ( .A(sqrto_96_), .B(u2__abc_52138_new_n3642_), .Y(u2__abc_52138_new_n3643_));
NOR2X1 NOR2X1_197 ( .A(u2_remHi_96_), .B(u2__abc_52138_new_n3644_), .Y(u2__abc_52138_new_n3645_));
NOR2X1 NOR2X1_198 ( .A(u2__abc_52138_new_n3643_), .B(u2__abc_52138_new_n3645_), .Y(u2__abc_52138_new_n3646_));
NOR2X1 NOR2X1_199 ( .A(sqrto_97_), .B(u2__abc_52138_new_n3647_), .Y(u2__abc_52138_new_n3648_));
NOR2X1 NOR2X1_2 ( .A(\a[112] ), .B(_abc_65734_new_n1448_), .Y(fracta1_113_));
NOR2X1 NOR2X1_20 ( .A(\a[119] ), .B(\a[120] ), .Y(u1__abc_51895_new_n138_));
NOR2X1 NOR2X1_200 ( .A(u2_remHi_97_), .B(u2__abc_52138_new_n3649_), .Y(u2__abc_52138_new_n3650_));
NOR2X1 NOR2X1_201 ( .A(u2__abc_52138_new_n3648_), .B(u2__abc_52138_new_n3650_), .Y(u2__abc_52138_new_n3651_));
NOR2X1 NOR2X1_202 ( .A(u2__abc_52138_new_n3652_), .B(u2__abc_52138_new_n3663_), .Y(u2__abc_52138_new_n3664_));
NOR2X1 NOR2X1_203 ( .A(u2__abc_52138_new_n3669_), .B(u2__abc_52138_new_n3674_), .Y(u2__abc_52138_new_n3675_));
NOR2X1 NOR2X1_204 ( .A(u2__abc_52138_new_n3680_), .B(u2__abc_52138_new_n3685_), .Y(u2__abc_52138_new_n3686_));
NOR2X1 NOR2X1_205 ( .A(u2__abc_52138_new_n3688_), .B(u2__abc_52138_new_n3641_), .Y(u2__abc_52138_new_n3689_));
NOR2X1 NOR2X1_206 ( .A(sqrto_90_), .B(u2__abc_52138_new_n3706_), .Y(u2__abc_52138_new_n3707_));
NOR2X1 NOR2X1_207 ( .A(u2_remHi_90_), .B(u2__abc_52138_new_n3708_), .Y(u2__abc_52138_new_n3709_));
NOR2X1 NOR2X1_208 ( .A(u2__abc_52138_new_n3707_), .B(u2__abc_52138_new_n3709_), .Y(u2__abc_52138_new_n3710_));
NOR2X1 NOR2X1_209 ( .A(u2__abc_52138_new_n3701_), .B(u2__abc_52138_new_n3711_), .Y(u2__abc_52138_new_n3712_));
NOR2X1 NOR2X1_21 ( .A(\a[125] ), .B(\a[126] ), .Y(u1__abc_51895_new_n140_));
NOR2X1 NOR2X1_210 ( .A(sqrto_87_), .B(u2__abc_52138_new_n3724_), .Y(u2__abc_52138_new_n3725_));
NOR2X1 NOR2X1_211 ( .A(u2_remHi_87_), .B(u2__abc_52138_new_n3727_), .Y(u2__abc_52138_new_n3728_));
NOR2X1 NOR2X1_212 ( .A(sqrto_86_), .B(u2__abc_52138_new_n3730_), .Y(u2__abc_52138_new_n3731_));
NOR2X1 NOR2X1_213 ( .A(u2_remHi_86_), .B(u2__abc_52138_new_n3732_), .Y(u2__abc_52138_new_n3733_));
NOR2X1 NOR2X1_214 ( .A(u2__abc_52138_new_n3731_), .B(u2__abc_52138_new_n3733_), .Y(u2__abc_52138_new_n3734_));
NOR2X1 NOR2X1_215 ( .A(u2__abc_52138_new_n3723_), .B(u2__abc_52138_new_n3735_), .Y(u2__abc_52138_new_n3736_));
NOR2X1 NOR2X1_216 ( .A(u2__abc_52138_new_n3759_), .B(u2__abc_52138_new_n3748_), .Y(u2__abc_52138_new_n3760_));
NOR2X1 NOR2X1_217 ( .A(u2__abc_52138_new_n3765_), .B(u2__abc_52138_new_n3770_), .Y(u2__abc_52138_new_n3771_));
NOR2X1 NOR2X1_218 ( .A(u2__abc_52138_new_n3776_), .B(u2__abc_52138_new_n3781_), .Y(u2__abc_52138_new_n3782_));
NOR2X1 NOR2X1_219 ( .A(u2__abc_52138_new_n3784_), .B(u2__abc_52138_new_n3737_), .Y(u2__abc_52138_new_n3785_));
NOR2X1 NOR2X1_22 ( .A(\a[123] ), .B(\a[124] ), .Y(u1__abc_51895_new_n141_));
NOR2X1 NOR2X1_220 ( .A(sqrto_70_), .B(u2__abc_52138_new_n3786_), .Y(u2__abc_52138_new_n3787_));
NOR2X1 NOR2X1_221 ( .A(u2_remHi_70_), .B(u2__abc_52138_new_n3788_), .Y(u2__abc_52138_new_n3789_));
NOR2X1 NOR2X1_222 ( .A(u2__abc_52138_new_n3787_), .B(u2__abc_52138_new_n3789_), .Y(u2__abc_52138_new_n3790_));
NOR2X1 NOR2X1_223 ( .A(sqrto_71_), .B(u2__abc_52138_new_n3791_), .Y(u2__abc_52138_new_n3792_));
NOR2X1 NOR2X1_224 ( .A(u2_remHi_71_), .B(u2__abc_52138_new_n3793_), .Y(u2__abc_52138_new_n3794_));
NOR2X1 NOR2X1_225 ( .A(u2__abc_52138_new_n3792_), .B(u2__abc_52138_new_n3794_), .Y(u2__abc_52138_new_n3795_));
NOR2X1 NOR2X1_226 ( .A(u2__abc_52138_new_n3796_), .B(u2__abc_52138_new_n3806_), .Y(u2__abc_52138_new_n3807_));
NOR2X1 NOR2X1_227 ( .A(sqrto_76_), .B(u2__abc_52138_new_n3808_), .Y(u2__abc_52138_new_n3809_));
NOR2X1 NOR2X1_228 ( .A(u2_remHi_76_), .B(u2__abc_52138_new_n3810_), .Y(u2__abc_52138_new_n3811_));
NOR2X1 NOR2X1_229 ( .A(u2__abc_52138_new_n3809_), .B(u2__abc_52138_new_n3811_), .Y(u2__abc_52138_new_n3812_));
NOR2X1 NOR2X1_23 ( .A(u1__abc_51895_new_n139_), .B(u1__abc_51895_new_n142_), .Y(u1__abc_51895_new_n143_));
NOR2X1 NOR2X1_230 ( .A(sqrto_77_), .B(u2__abc_52138_new_n3813_), .Y(u2__abc_52138_new_n3814_));
NOR2X1 NOR2X1_231 ( .A(u2_remHi_77_), .B(u2__abc_52138_new_n3815_), .Y(u2__abc_52138_new_n3816_));
NOR2X1 NOR2X1_232 ( .A(u2__abc_52138_new_n3814_), .B(u2__abc_52138_new_n3816_), .Y(u2__abc_52138_new_n3817_));
NOR2X1 NOR2X1_233 ( .A(sqrto_75_), .B(u2__abc_52138_new_n3819_), .Y(u2__abc_52138_new_n3820_));
NOR2X1 NOR2X1_234 ( .A(u2_remHi_75_), .B(u2__abc_52138_new_n3821_), .Y(u2__abc_52138_new_n3822_));
NOR2X1 NOR2X1_235 ( .A(u2__abc_52138_new_n3820_), .B(u2__abc_52138_new_n3822_), .Y(u2__abc_52138_new_n3823_));
NOR2X1 NOR2X1_236 ( .A(sqrto_74_), .B(u2__abc_52138_new_n3824_), .Y(u2__abc_52138_new_n3825_));
NOR2X1 NOR2X1_237 ( .A(u2_remHi_74_), .B(u2__abc_52138_new_n3826_), .Y(u2__abc_52138_new_n3827_));
NOR2X1 NOR2X1_238 ( .A(u2__abc_52138_new_n3825_), .B(u2__abc_52138_new_n3827_), .Y(u2__abc_52138_new_n3828_));
NOR2X1 NOR2X1_239 ( .A(u2__abc_52138_new_n3818_), .B(u2__abc_52138_new_n3829_), .Y(u2__abc_52138_new_n3830_));
NOR2X1 NOR2X1_24 ( .A(\a[113] ), .B(\a[114] ), .Y(u1__abc_51895_new_n145_));
NOR2X1 NOR2X1_240 ( .A(u2__abc_52138_new_n3836_), .B(u2__abc_52138_new_n3841_), .Y(u2__abc_52138_new_n3842_));
NOR2X1 NOR2X1_241 ( .A(u2__abc_52138_new_n3847_), .B(u2__abc_52138_new_n3852_), .Y(u2__abc_52138_new_n3853_));
NOR2X1 NOR2X1_242 ( .A(u2__abc_52138_new_n3860_), .B(u2__abc_52138_new_n3866_), .Y(u2__abc_52138_new_n3867_));
NOR2X1 NOR2X1_243 ( .A(u2__abc_52138_new_n3868_), .B(u2__abc_52138_new_n3831_), .Y(u2__abc_52138_new_n3869_));
NOR2X1 NOR2X1_244 ( .A(u2__abc_52138_new_n3870_), .B(u2__abc_52138_new_n3690_), .Y(u2__abc_52138_new_n3871_));
NOR2X1 NOR2X1_245 ( .A(sqrto_69_), .B(u2__abc_52138_new_n3858_), .Y(u2__abc_52138_new_n3890_));
NOR2X1 NOR2X1_246 ( .A(sqrto_85_), .B(u2__abc_52138_new_n3768_), .Y(u2__abc_52138_new_n3918_));
NOR2X1 NOR2X1_247 ( .A(u2__abc_52138_new_n3695_), .B(u2__abc_52138_new_n3700_), .Y(u2__abc_52138_new_n3928_));
NOR2X1 NOR2X1_248 ( .A(u2_remHi_100_), .B(u2__abc_52138_new_n3665_), .Y(u2__abc_52138_new_n3951_));
NOR2X1 NOR2X1_249 ( .A(u2_remHi_101_), .B(u2__abc_52138_new_n3670_), .Y(u2__abc_52138_new_n3952_));
NOR2X1 NOR2X1_25 ( .A(\a[117] ), .B(\a[118] ), .Y(u1__abc_51895_new_n147_));
NOR2X1 NOR2X1_250 ( .A(u2__abc_52138_new_n3623_), .B(u2__abc_52138_new_n3628_), .Y(u2__abc_52138_new_n3962_));
NOR2X1 NOR2X1_251 ( .A(sqrto_115_), .B(u2__abc_52138_new_n3585_), .Y(u2__abc_52138_new_n3982_));
NOR2X1 NOR2X1_252 ( .A(u2__abc_52138_new_n3531_), .B(u2__abc_52138_new_n3536_), .Y(u2__abc_52138_new_n3991_));
NOR2X1 NOR2X1_253 ( .A(u2__abc_52138_new_n4007_), .B(u2__abc_52138_new_n4012_), .Y(u2__abc_52138_new_n4013_));
NOR2X1 NOR2X1_254 ( .A(u2__abc_52138_new_n4018_), .B(u2__abc_52138_new_n4023_), .Y(u2__abc_52138_new_n4024_));
NOR2X1 NOR2X1_255 ( .A(u2__abc_52138_new_n4030_), .B(u2__abc_52138_new_n4035_), .Y(u2__abc_52138_new_n4036_));
NOR2X1 NOR2X1_256 ( .A(u2__abc_52138_new_n4041_), .B(u2__abc_52138_new_n4046_), .Y(u2__abc_52138_new_n4047_));
NOR2X1 NOR2X1_257 ( .A(u2__abc_52138_new_n4065_), .B(u2__abc_52138_new_n4070_), .Y(u2__abc_52138_new_n4071_));
NOR2X1 NOR2X1_258 ( .A(u2__abc_52138_new_n4060_), .B(u2__abc_52138_new_n4072_), .Y(u2__abc_52138_new_n4073_));
NOR2X1 NOR2X1_259 ( .A(u2__abc_52138_new_n4078_), .B(u2__abc_52138_new_n4083_), .Y(u2__abc_52138_new_n4084_));
NOR2X1 NOR2X1_26 ( .A(\a[115] ), .B(\a[116] ), .Y(u1__abc_51895_new_n148_));
NOR2X1 NOR2X1_260 ( .A(u2_o_243_), .B(u2__abc_52138_new_n4085_), .Y(u2__abc_52138_new_n4086_));
NOR2X1 NOR2X1_261 ( .A(u2_remHi_243_), .B(u2__abc_52138_new_n4087_), .Y(u2__abc_52138_new_n4088_));
NOR2X1 NOR2X1_262 ( .A(u2__abc_52138_new_n4086_), .B(u2__abc_52138_new_n4088_), .Y(u2__abc_52138_new_n4089_));
NOR2X1 NOR2X1_263 ( .A(u2__abc_52138_new_n4049_), .B(u2__abc_52138_new_n4097_), .Y(u2__abc_52138_new_n4098_));
NOR2X1 NOR2X1_264 ( .A(u2__abc_52138_new_n4103_), .B(u2__abc_52138_new_n4108_), .Y(u2__abc_52138_new_n4109_));
NOR2X1 NOR2X1_265 ( .A(u2__abc_52138_new_n4114_), .B(u2__abc_52138_new_n4119_), .Y(u2__abc_52138_new_n4120_));
NOR2X1 NOR2X1_266 ( .A(u2_o_231_), .B(u2__abc_52138_new_n4134_), .Y(u2__abc_52138_new_n4135_));
NOR2X1 NOR2X1_267 ( .A(u2_o_230_), .B(u2__abc_52138_new_n4138_), .Y(u2__abc_52138_new_n4139_));
NOR2X1 NOR2X1_268 ( .A(u2_remHi_230_), .B(u2__abc_52138_new_n4140_), .Y(u2__abc_52138_new_n4141_));
NOR2X1 NOR2X1_269 ( .A(u2__abc_52138_new_n4139_), .B(u2__abc_52138_new_n4141_), .Y(u2__abc_52138_new_n4142_));
NOR2X1 NOR2X1_27 ( .A(u1__abc_51895_new_n146_), .B(u1__abc_51895_new_n149_), .Y(u1__abc_51895_new_n150_));
NOR2X1 NOR2X1_270 ( .A(u2__abc_52138_new_n4133_), .B(u2__abc_52138_new_n4143_), .Y(u2__abc_52138_new_n4144_));
NOR2X1 NOR2X1_271 ( .A(u2__abc_52138_new_n4150_), .B(u2__abc_52138_new_n4155_), .Y(u2__abc_52138_new_n4156_));
NOR2X1 NOR2X1_272 ( .A(u2__abc_52138_new_n4161_), .B(u2__abc_52138_new_n4166_), .Y(u2__abc_52138_new_n4167_));
NOR2X1 NOR2X1_273 ( .A(u2__abc_52138_new_n4173_), .B(u2__abc_52138_new_n4178_), .Y(u2__abc_52138_new_n4179_));
NOR2X1 NOR2X1_274 ( .A(u2_o_227_), .B(u2__abc_52138_new_n4180_), .Y(u2__abc_52138_new_n4181_));
NOR2X1 NOR2X1_275 ( .A(u2_remHi_227_), .B(u2__abc_52138_new_n4182_), .Y(u2__abc_52138_new_n4183_));
NOR2X1 NOR2X1_276 ( .A(u2__abc_52138_new_n4181_), .B(u2__abc_52138_new_n4183_), .Y(u2__abc_52138_new_n4184_));
NOR2X1 NOR2X1_277 ( .A(u2_o_226_), .B(u2__abc_52138_new_n4185_), .Y(u2__abc_52138_new_n4186_));
NOR2X1 NOR2X1_278 ( .A(u2_remHi_226_), .B(u2__abc_52138_new_n4187_), .Y(u2__abc_52138_new_n4188_));
NOR2X1 NOR2X1_279 ( .A(u2__abc_52138_new_n4186_), .B(u2__abc_52138_new_n4188_), .Y(u2__abc_52138_new_n4189_));
NOR2X1 NOR2X1_28 ( .A(u1__abc_51895_new_n153_), .B(u1__abc_51895_new_n154_), .Y(u1__abc_51895_new_n155_));
NOR2X1 NOR2X1_280 ( .A(u2__abc_52138_new_n4191_), .B(u2__abc_52138_new_n4145_), .Y(u2__abc_52138_new_n4192_));
NOR2X1 NOR2X1_281 ( .A(u2__abc_52138_new_n4204_), .B(u2__abc_52138_new_n4215_), .Y(u2__abc_52138_new_n4216_));
NOR2X1 NOR2X1_282 ( .A(sqrto_219_), .B(u2__abc_52138_new_n4228_), .Y(u2__abc_52138_new_n4229_));
NOR2X1 NOR2X1_283 ( .A(u2_remHi_219_), .B(u2__abc_52138_new_n4230_), .Y(u2__abc_52138_new_n4231_));
NOR2X1 NOR2X1_284 ( .A(u2__abc_52138_new_n4229_), .B(u2__abc_52138_new_n4231_), .Y(u2__abc_52138_new_n4232_));
NOR2X1 NOR2X1_285 ( .A(u2__abc_52138_new_n4238_), .B(u2__abc_52138_new_n4227_), .Y(u2__abc_52138_new_n4239_));
NOR2X1 NOR2X1_286 ( .A(u2__abc_52138_new_n4251_), .B(u2__abc_52138_new_n4262_), .Y(u2__abc_52138_new_n4263_));
NOR2X1 NOR2X1_287 ( .A(sqrto_212_), .B(u2__abc_52138_new_n4264_), .Y(u2__abc_52138_new_n4265_));
NOR2X1 NOR2X1_288 ( .A(u2_remHi_212_), .B(u2__abc_52138_new_n4266_), .Y(u2__abc_52138_new_n4267_));
NOR2X1 NOR2X1_289 ( .A(u2__abc_52138_new_n4265_), .B(u2__abc_52138_new_n4267_), .Y(u2__abc_52138_new_n4268_));
NOR2X1 NOR2X1_29 ( .A(u1__abc_51895_new_n156_), .B(u1__abc_51895_new_n157_), .Y(u1__abc_51895_new_n158_));
NOR2X1 NOR2X1_290 ( .A(sqrto_213_), .B(u2__abc_52138_new_n4269_), .Y(u2__abc_52138_new_n4270_));
NOR2X1 NOR2X1_291 ( .A(u2_remHi_213_), .B(u2__abc_52138_new_n4271_), .Y(u2__abc_52138_new_n4272_));
NOR2X1 NOR2X1_292 ( .A(u2__abc_52138_new_n4270_), .B(u2__abc_52138_new_n4272_), .Y(u2__abc_52138_new_n4273_));
NOR2X1 NOR2X1_293 ( .A(sqrto_211_), .B(u2__abc_52138_new_n4275_), .Y(u2__abc_52138_new_n4276_));
NOR2X1 NOR2X1_294 ( .A(u2_remHi_211_), .B(u2__abc_52138_new_n4277_), .Y(u2__abc_52138_new_n4278_));
NOR2X1 NOR2X1_295 ( .A(u2__abc_52138_new_n4276_), .B(u2__abc_52138_new_n4278_), .Y(u2__abc_52138_new_n4279_));
NOR2X1 NOR2X1_296 ( .A(sqrto_210_), .B(u2__abc_52138_new_n4280_), .Y(u2__abc_52138_new_n4281_));
NOR2X1 NOR2X1_297 ( .A(u2_remHi_210_), .B(u2__abc_52138_new_n4282_), .Y(u2__abc_52138_new_n4283_));
NOR2X1 NOR2X1_298 ( .A(u2__abc_52138_new_n4281_), .B(u2__abc_52138_new_n4283_), .Y(u2__abc_52138_new_n4284_));
NOR2X1 NOR2X1_299 ( .A(u2__abc_52138_new_n4285_), .B(u2__abc_52138_new_n4274_), .Y(u2__abc_52138_new_n4286_));
NOR2X1 NOR2X1_3 ( .A(\a[112] ), .B(\a[113] ), .Y(_abc_65734_new_n1453_));
NOR2X1 NOR2X1_30 ( .A(u1__abc_51895_new_n161_), .B(u1__abc_51895_new_n162_), .Y(u1__abc_51895_new_n163_));
NOR2X1 NOR2X1_300 ( .A(u2__abc_52138_new_n4240_), .B(u2__abc_52138_new_n4287_), .Y(u2__abc_52138_new_n4288_));
NOR2X1 NOR2X1_301 ( .A(u2__abc_52138_new_n4293_), .B(u2__abc_52138_new_n4298_), .Y(u2__abc_52138_new_n4299_));
NOR2X1 NOR2X1_302 ( .A(u2__abc_52138_new_n4304_), .B(u2__abc_52138_new_n4309_), .Y(u2__abc_52138_new_n4310_));
NOR2X1 NOR2X1_303 ( .A(u2__abc_52138_new_n4316_), .B(u2__abc_52138_new_n4321_), .Y(u2__abc_52138_new_n4322_));
NOR2X1 NOR2X1_304 ( .A(sqrto_203_), .B(u2__abc_52138_new_n4323_), .Y(u2__abc_52138_new_n4324_));
NOR2X1 NOR2X1_305 ( .A(u2_remHi_203_), .B(u2__abc_52138_new_n4325_), .Y(u2__abc_52138_new_n4326_));
NOR2X1 NOR2X1_306 ( .A(u2__abc_52138_new_n4324_), .B(u2__abc_52138_new_n4326_), .Y(u2__abc_52138_new_n4327_));
NOR2X1 NOR2X1_307 ( .A(u2__abc_52138_new_n4335_), .B(u2__abc_52138_new_n4340_), .Y(u2__abc_52138_new_n4341_));
NOR2X1 NOR2X1_308 ( .A(u2__abc_52138_new_n4346_), .B(u2__abc_52138_new_n4351_), .Y(u2__abc_52138_new_n4352_));
NOR2X1 NOR2X1_309 ( .A(sqrto_192_), .B(u2__abc_52138_new_n4354_), .Y(u2__abc_52138_new_n4355_));
NOR2X1 NOR2X1_31 ( .A(u1__abc_51895_new_n159_), .B(u1__abc_51895_new_n164_), .Y(u1_xinf));
NOR2X1 NOR2X1_310 ( .A(u2_remHi_192_), .B(u2__abc_52138_new_n4356_), .Y(u2__abc_52138_new_n4357_));
NOR2X1 NOR2X1_311 ( .A(sqrto_190_), .B(u2__abc_52138_new_n4364_), .Y(u2__abc_52138_new_n4365_));
NOR2X1 NOR2X1_312 ( .A(u2_remHi_190_), .B(u2__abc_52138_new_n4366_), .Y(u2__abc_52138_new_n4367_));
NOR2X1 NOR2X1_313 ( .A(sqrto_191_), .B(u2__abc_52138_new_n4369_), .Y(u2__abc_52138_new_n4370_));
NOR2X1 NOR2X1_314 ( .A(u2_remHi_191_), .B(u2__abc_52138_new_n4372_), .Y(u2__abc_52138_new_n4373_));
NOR2X1 NOR2X1_315 ( .A(u2__abc_52138_new_n4368_), .B(u2__abc_52138_new_n4375_), .Y(u2__abc_52138_new_n4376_));
NOR2X1 NOR2X1_316 ( .A(u2__abc_52138_new_n4330_), .B(u2__abc_52138_new_n4378_), .Y(u2__abc_52138_new_n4379_));
NOR2X1 NOR2X1_317 ( .A(u2__abc_52138_new_n4193_), .B(u2__abc_52138_new_n4380_), .Y(u2__abc_52138_new_n4381_));
NOR2X1 NOR2X1_318 ( .A(u2__abc_52138_new_n4386_), .B(u2__abc_52138_new_n4391_), .Y(u2__abc_52138_new_n4392_));
NOR2X1 NOR2X1_319 ( .A(u2__abc_52138_new_n4397_), .B(u2__abc_52138_new_n4402_), .Y(u2__abc_52138_new_n4403_));
NOR2X1 NOR2X1_32 ( .A(\a[10] ), .B(\a[11] ), .Y(u1__abc_51895_new_n166_));
NOR2X1 NOR2X1_320 ( .A(u2__abc_52138_new_n4409_), .B(u2__abc_52138_new_n4414_), .Y(u2__abc_52138_new_n4415_));
NOR2X1 NOR2X1_321 ( .A(u2__abc_52138_new_n4420_), .B(u2__abc_52138_new_n4425_), .Y(u2__abc_52138_new_n4426_));
NOR2X1 NOR2X1_322 ( .A(u2__abc_52138_new_n4404_), .B(u2__abc_52138_new_n4427_), .Y(u2__abc_52138_new_n4428_));
NOR2X1 NOR2X1_323 ( .A(u2__abc_52138_new_n4433_), .B(u2__abc_52138_new_n4438_), .Y(u2__abc_52138_new_n4439_));
NOR2X1 NOR2X1_324 ( .A(u2__abc_52138_new_n4444_), .B(u2__abc_52138_new_n4449_), .Y(u2__abc_52138_new_n4450_));
NOR2X1 NOR2X1_325 ( .A(u2__abc_52138_new_n4456_), .B(u2__abc_52138_new_n4461_), .Y(u2__abc_52138_new_n4462_));
NOR2X1 NOR2X1_326 ( .A(u2__abc_52138_new_n4451_), .B(u2__abc_52138_new_n4475_), .Y(u2__abc_52138_new_n4476_));
NOR2X1 NOR2X1_327 ( .A(u2__abc_52138_new_n4482_), .B(u2__abc_52138_new_n4487_), .Y(u2__abc_52138_new_n4488_));
NOR2X1 NOR2X1_328 ( .A(u2__abc_52138_new_n4493_), .B(u2__abc_52138_new_n4498_), .Y(u2__abc_52138_new_n4499_));
NOR2X1 NOR2X1_329 ( .A(u2__abc_52138_new_n4505_), .B(u2__abc_52138_new_n4510_), .Y(u2__abc_52138_new_n4511_));
NOR2X1 NOR2X1_33 ( .A(\a[8] ), .B(\a[9] ), .Y(u1__abc_51895_new_n167_));
NOR2X1 NOR2X1_330 ( .A(sqrto_166_), .B(u2__abc_52138_new_n4517_), .Y(u2__abc_52138_new_n4518_));
NOR2X1 NOR2X1_331 ( .A(u2_remHi_166_), .B(u2__abc_52138_new_n4519_), .Y(u2__abc_52138_new_n4520_));
NOR2X1 NOR2X1_332 ( .A(u2__abc_52138_new_n4516_), .B(u2__abc_52138_new_n4521_), .Y(u2__abc_52138_new_n4522_));
NOR2X1 NOR2X1_333 ( .A(u2__abc_52138_new_n4500_), .B(u2__abc_52138_new_n4523_), .Y(u2__abc_52138_new_n4524_));
NOR2X1 NOR2X1_334 ( .A(u2__abc_52138_new_n4529_), .B(u2__abc_52138_new_n4534_), .Y(u2__abc_52138_new_n4535_));
NOR2X1 NOR2X1_335 ( .A(u2_remHi_159_), .B(u2__abc_52138_new_n4536_), .Y(u2__abc_52138_new_n4538_));
NOR2X1 NOR2X1_336 ( .A(sqrto_158_), .B(u2__abc_52138_new_n4541_), .Y(u2__abc_52138_new_n4542_));
NOR2X1 NOR2X1_337 ( .A(u2_remHi_158_), .B(u2__abc_52138_new_n4543_), .Y(u2__abc_52138_new_n4544_));
NOR2X1 NOR2X1_338 ( .A(u2__abc_52138_new_n4545_), .B(u2__abc_52138_new_n4540_), .Y(u2__abc_52138_new_n4546_));
NOR2X1 NOR2X1_339 ( .A(u2__abc_52138_new_n4552_), .B(u2__abc_52138_new_n4557_), .Y(u2__abc_52138_new_n4558_));
NOR2X1 NOR2X1_34 ( .A(\a[14] ), .B(\a[15] ), .Y(u1__abc_51895_new_n169_));
NOR2X1 NOR2X1_340 ( .A(u2__abc_52138_new_n4563_), .B(u2__abc_52138_new_n4568_), .Y(u2__abc_52138_new_n4569_));
NOR2X1 NOR2X1_341 ( .A(u2__abc_52138_new_n4477_), .B(u2__abc_52138_new_n4571_), .Y(u2__abc_52138_new_n4572_));
NOR2X1 NOR2X1_342 ( .A(u2__abc_52138_new_n4577_), .B(u2__abc_52138_new_n4582_), .Y(u2__abc_52138_new_n4583_));
NOR2X1 NOR2X1_343 ( .A(u2__abc_52138_new_n4588_), .B(u2__abc_52138_new_n4593_), .Y(u2__abc_52138_new_n4594_));
NOR2X1 NOR2X1_344 ( .A(u2__abc_52138_new_n4600_), .B(u2__abc_52138_new_n4605_), .Y(u2__abc_52138_new_n4606_));
NOR2X1 NOR2X1_345 ( .A(sqrto_155_), .B(u2__abc_52138_new_n4607_), .Y(u2__abc_52138_new_n4608_));
NOR2X1 NOR2X1_346 ( .A(u2_remHi_155_), .B(u2__abc_52138_new_n4609_), .Y(u2__abc_52138_new_n4610_));
NOR2X1 NOR2X1_347 ( .A(u2__abc_52138_new_n4608_), .B(u2__abc_52138_new_n4610_), .Y(u2__abc_52138_new_n4611_));
NOR2X1 NOR2X1_348 ( .A(sqrto_154_), .B(u2__abc_52138_new_n4612_), .Y(u2__abc_52138_new_n4613_));
NOR2X1 NOR2X1_349 ( .A(u2_remHi_154_), .B(u2__abc_52138_new_n4614_), .Y(u2__abc_52138_new_n4615_));
NOR2X1 NOR2X1_35 ( .A(\a[12] ), .B(\a[13] ), .Y(u1__abc_51895_new_n170_));
NOR2X1 NOR2X1_350 ( .A(u2__abc_52138_new_n4613_), .B(u2__abc_52138_new_n4615_), .Y(u2__abc_52138_new_n4616_));
NOR2X1 NOR2X1_351 ( .A(u2__abc_52138_new_n4595_), .B(u2__abc_52138_new_n4617_), .Y(u2__abc_52138_new_n4618_));
NOR2X1 NOR2X1_352 ( .A(u2__abc_52138_new_n4623_), .B(u2__abc_52138_new_n4628_), .Y(u2__abc_52138_new_n4629_));
NOR2X1 NOR2X1_353 ( .A(u2__abc_52138_new_n4634_), .B(u2__abc_52138_new_n4639_), .Y(u2__abc_52138_new_n4640_));
NOR2X1 NOR2X1_354 ( .A(sqrto_143_), .B(u2__abc_52138_new_n4652_), .Y(u2__abc_52138_new_n4653_));
NOR2X1 NOR2X1_355 ( .A(u2_remHi_143_), .B(u2__abc_52138_new_n4655_), .Y(u2__abc_52138_new_n4656_));
NOR2X1 NOR2X1_356 ( .A(sqrto_142_), .B(u2__abc_52138_new_n4658_), .Y(u2__abc_52138_new_n4659_));
NOR2X1 NOR2X1_357 ( .A(u2_remHi_142_), .B(u2__abc_52138_new_n4660_), .Y(u2__abc_52138_new_n4661_));
NOR2X1 NOR2X1_358 ( .A(u2__abc_52138_new_n4659_), .B(u2__abc_52138_new_n4661_), .Y(u2__abc_52138_new_n4662_));
NOR2X1 NOR2X1_359 ( .A(u2__abc_52138_new_n4651_), .B(u2__abc_52138_new_n4663_), .Y(u2__abc_52138_new_n4664_));
NOR2X1 NOR2X1_36 ( .A(u1__abc_51895_new_n168_), .B(u1__abc_51895_new_n171_), .Y(u1__abc_51895_new_n172_));
NOR2X1 NOR2X1_360 ( .A(u2__abc_52138_new_n4670_), .B(u2__abc_52138_new_n4675_), .Y(u2__abc_52138_new_n4676_));
NOR2X1 NOR2X1_361 ( .A(u2__abc_52138_new_n4681_), .B(u2__abc_52138_new_n4686_), .Y(u2__abc_52138_new_n4687_));
NOR2X1 NOR2X1_362 ( .A(u2__abc_52138_new_n4693_), .B(u2__abc_52138_new_n4698_), .Y(u2__abc_52138_new_n4699_));
NOR2X1 NOR2X1_363 ( .A(u2__abc_52138_new_n4704_), .B(u2__abc_52138_new_n4709_), .Y(u2__abc_52138_new_n4710_));
NOR2X1 NOR2X1_364 ( .A(u2__abc_52138_new_n4737_), .B(u2__abc_52138_new_n4742_), .Y(u2__abc_52138_new_n4743_));
NOR2X1 NOR2X1_365 ( .A(u2__abc_52138_new_n4756_), .B(u2__abc_52138_new_n4757_), .Y(u2__abc_52138_new_n4758_));
NOR2X1 NOR2X1_366 ( .A(u2__abc_52138_new_n4761_), .B(u2__abc_52138_new_n4760_), .Y(u2__abc_52138_new_n4762_));
NOR2X1 NOR2X1_367 ( .A(u2__abc_52138_new_n4764_), .B(u2__abc_52138_new_n4765_), .Y(u2__abc_52138_new_n4766_));
NOR2X1 NOR2X1_368 ( .A(u2_remHi_128_), .B(u2__abc_52138_new_n4770_), .Y(u2__abc_52138_new_n4771_));
NOR2X1 NOR2X1_369 ( .A(sqrto_131_), .B(u2__abc_52138_new_n4746_), .Y(u2__abc_52138_new_n4775_));
NOR2X1 NOR2X1_37 ( .A(\a[2] ), .B(\a[3] ), .Y(u1__abc_51895_new_n173_));
NOR2X1 NOR2X1_370 ( .A(sqrto_133_), .B(u2__abc_52138_new_n4740_), .Y(u2__abc_52138_new_n4780_));
NOR2X1 NOR2X1_371 ( .A(sqrto_137_), .B(u2__abc_52138_new_n4673_), .Y(u2__abc_52138_new_n4789_));
NOR2X1 NOR2X1_372 ( .A(u2_remHi_144_), .B(u2__abc_52138_new_n4642_), .Y(u2__abc_52138_new_n4802_));
NOR2X1 NOR2X1_373 ( .A(sqrto_147_), .B(u2__abc_52138_new_n4632_), .Y(u2__abc_52138_new_n4807_));
NOR2X1 NOR2X1_374 ( .A(u2_remHi_148_), .B(u2__abc_52138_new_n4619_), .Y(u2__abc_52138_new_n4810_));
NOR2X1 NOR2X1_375 ( .A(u2_remHi_149_), .B(u2__abc_52138_new_n4624_), .Y(u2__abc_52138_new_n4811_));
NOR2X1 NOR2X1_376 ( .A(sqrto_161_), .B(u2__abc_52138_new_n4532_), .Y(u2__abc_52138_new_n4833_));
NOR2X1 NOR2X1_377 ( .A(sqrto_163_), .B(u2__abc_52138_new_n4561_), .Y(u2__abc_52138_new_n4838_));
NOR2X1 NOR2X1_378 ( .A(u2__abc_52138_new_n4355_), .B(u2__abc_52138_new_n4357_), .Y(u2__abc_52138_new_n4880_));
NOR2X1 NOR2X1_379 ( .A(sqrto_193_), .B(u2__abc_52138_new_n4360_), .Y(u2__abc_52138_new_n4881_));
NOR2X1 NOR2X1_38 ( .A(\a[0] ), .B(\a[1] ), .Y(u1__abc_51895_new_n174_));
NOR2X1 NOR2X1_380 ( .A(u2_remHi_193_), .B(u2__abc_52138_new_n4358_), .Y(u2__abc_52138_new_n4882_));
NOR2X1 NOR2X1_381 ( .A(u2__abc_52138_new_n4881_), .B(u2__abc_52138_new_n4882_), .Y(u2__abc_52138_new_n4883_));
NOR2X1 NOR2X1_382 ( .A(sqrto_195_), .B(u2__abc_52138_new_n4344_), .Y(u2__abc_52138_new_n4889_));
NOR2X1 NOR2X1_383 ( .A(sqrto_197_), .B(u2__abc_52138_new_n4338_), .Y(u2__abc_52138_new_n4892_));
NOR2X1 NOR2X1_384 ( .A(u2__abc_52138_new_n4198_), .B(u2__abc_52138_new_n4203_), .Y(u2__abc_52138_new_n4928_));
NOR2X1 NOR2X1_385 ( .A(u2__abc_52138_new_n4221_), .B(u2__abc_52138_new_n4226_), .Y(u2__abc_52138_new_n4934_));
NOR2X1 NOR2X1_386 ( .A(u2__abc_52138_new_n4127_), .B(u2__abc_52138_new_n4132_), .Y(u2__abc_52138_new_n4959_));
NOR2X1 NOR2X1_387 ( .A(u2__abc_52138_new_n4025_), .B(u2__abc_52138_new_n4048_), .Y(u2__abc_52138_new_n4982_));
NOR2X1 NOR2X1_388 ( .A(u2_o_380_), .B(u2__abc_52138_new_n4999_), .Y(u2__abc_52138_new_n5000_));
NOR2X1 NOR2X1_389 ( .A(u2_remHi_380_), .B(u2__abc_52138_new_n5001_), .Y(u2__abc_52138_new_n5002_));
NOR2X1 NOR2X1_39 ( .A(\a[6] ), .B(\a[7] ), .Y(u1__abc_51895_new_n176_));
NOR2X1 NOR2X1_390 ( .A(u2__abc_52138_new_n5000_), .B(u2__abc_52138_new_n5002_), .Y(u2__abc_52138_new_n5003_));
NOR2X1 NOR2X1_391 ( .A(u2_remHi_381_), .B(u2__abc_52138_new_n5004_), .Y(u2__abc_52138_new_n5005_));
NOR2X1 NOR2X1_392 ( .A(u2_o_381_), .B(u2__abc_52138_new_n5006_), .Y(u2__abc_52138_new_n5007_));
NOR2X1 NOR2X1_393 ( .A(u2__abc_52138_new_n5005_), .B(u2__abc_52138_new_n5007_), .Y(u2__abc_52138_new_n5008_));
NOR2X1 NOR2X1_394 ( .A(u2_o_379_), .B(u2__abc_52138_new_n5011_), .Y(u2__abc_52138_new_n5012_));
NOR2X1 NOR2X1_395 ( .A(u2_remHi_379_), .B(u2__abc_52138_new_n5013_), .Y(u2__abc_52138_new_n5014_));
NOR2X1 NOR2X1_396 ( .A(u2__abc_52138_new_n5012_), .B(u2__abc_52138_new_n5014_), .Y(u2__abc_52138_new_n5015_));
NOR2X1 NOR2X1_397 ( .A(u2__abc_52138_new_n5016_), .B(u2__abc_52138_new_n5009_), .Y(u2__abc_52138_new_n5017_));
NOR2X1 NOR2X1_398 ( .A(u2_remHi_374_), .B(u2__abc_52138_new_n5018_), .Y(u2__abc_52138_new_n5019_));
NOR2X1 NOR2X1_399 ( .A(u2_o_374_), .B(u2__abc_52138_new_n5020_), .Y(u2__abc_52138_new_n5021_));
NOR2X1 NOR2X1_4 ( .A(\a[114] ), .B(_abc_65734_new_n1453_), .Y(_abc_65734_new_n1457_));
NOR2X1 NOR2X1_40 ( .A(\a[4] ), .B(\a[5] ), .Y(u1__abc_51895_new_n177_));
NOR2X1 NOR2X1_400 ( .A(u2__abc_52138_new_n5019_), .B(u2__abc_52138_new_n5021_), .Y(u2__abc_52138_new_n5022_));
NOR2X1 NOR2X1_401 ( .A(u2_o_376_), .B(u2__abc_52138_new_n5030_), .Y(u2__abc_52138_new_n5031_));
NOR2X1 NOR2X1_402 ( .A(u2_remHi_376_), .B(u2__abc_52138_new_n5032_), .Y(u2__abc_52138_new_n5033_));
NOR2X1 NOR2X1_403 ( .A(u2_o_377_), .B(u2__abc_52138_new_n5035_), .Y(u2__abc_52138_new_n5036_));
NOR2X1 NOR2X1_404 ( .A(u2_remHi_377_), .B(u2__abc_52138_new_n5038_), .Y(u2__abc_52138_new_n5039_));
NOR2X1 NOR2X1_405 ( .A(u2__abc_52138_new_n5029_), .B(u2__abc_52138_new_n5042_), .Y(u2__abc_52138_new_n5043_));
NOR2X1 NOR2X1_406 ( .A(u2_o_368_), .B(u2__abc_52138_new_n5045_), .Y(u2__abc_52138_new_n5046_));
NOR2X1 NOR2X1_407 ( .A(u2_remHi_368_), .B(u2__abc_52138_new_n5047_), .Y(u2__abc_52138_new_n5048_));
NOR2X1 NOR2X1_408 ( .A(u2__abc_52138_new_n5046_), .B(u2__abc_52138_new_n5048_), .Y(u2__abc_52138_new_n5049_));
NOR2X1 NOR2X1_409 ( .A(u2_o_366_), .B(u2__abc_52138_new_n5052_), .Y(u2__abc_52138_new_n5053_));
NOR2X1 NOR2X1_41 ( .A(u1__abc_51895_new_n175_), .B(u1__abc_51895_new_n178_), .Y(u1__abc_51895_new_n179_));
NOR2X1 NOR2X1_410 ( .A(u2__abc_52138_new_n5051_), .B(u2__abc_52138_new_n5063_), .Y(u2__abc_52138_new_n5064_));
NOR2X1 NOR2X1_411 ( .A(u2_o_372_), .B(u2__abc_52138_new_n5065_), .Y(u2__abc_52138_new_n5066_));
NOR2X1 NOR2X1_412 ( .A(u2_remHi_372_), .B(u2__abc_52138_new_n5067_), .Y(u2__abc_52138_new_n5068_));
NOR2X1 NOR2X1_413 ( .A(u2__abc_52138_new_n5066_), .B(u2__abc_52138_new_n5068_), .Y(u2__abc_52138_new_n5069_));
NOR2X1 NOR2X1_414 ( .A(u2_o_373_), .B(u2__abc_52138_new_n5070_), .Y(u2__abc_52138_new_n5071_));
NOR2X1 NOR2X1_415 ( .A(u2_remHi_373_), .B(u2__abc_52138_new_n5072_), .Y(u2__abc_52138_new_n5073_));
NOR2X1 NOR2X1_416 ( .A(u2__abc_52138_new_n5071_), .B(u2__abc_52138_new_n5073_), .Y(u2__abc_52138_new_n5074_));
NOR2X1 NOR2X1_417 ( .A(u2__abc_52138_new_n5075_), .B(u2__abc_52138_new_n5087_), .Y(u2__abc_52138_new_n5088_));
NOR2X1 NOR2X1_418 ( .A(u2__abc_52138_new_n5089_), .B(u2__abc_52138_new_n5044_), .Y(u2__abc_52138_new_n5090_));
NOR2X1 NOR2X1_419 ( .A(u2_remHi_358_), .B(u2__abc_52138_new_n5091_), .Y(u2__abc_52138_new_n5092_));
NOR2X1 NOR2X1_42 ( .A(\a[27] ), .B(\a[24] ), .Y(u1__abc_51895_new_n282_));
NOR2X1 NOR2X1_420 ( .A(u2_o_358_), .B(u2__abc_52138_new_n5093_), .Y(u2__abc_52138_new_n5094_));
NOR2X1 NOR2X1_421 ( .A(u2__abc_52138_new_n5092_), .B(u2__abc_52138_new_n5094_), .Y(u2__abc_52138_new_n5095_));
NOR2X1 NOR2X1_422 ( .A(u2_o_360_), .B(u2__abc_52138_new_n5102_), .Y(u2__abc_52138_new_n5103_));
NOR2X1 NOR2X1_423 ( .A(u2_remHi_360_), .B(u2__abc_52138_new_n5104_), .Y(u2__abc_52138_new_n5105_));
NOR2X1 NOR2X1_424 ( .A(u2__abc_52138_new_n5103_), .B(u2__abc_52138_new_n5105_), .Y(u2__abc_52138_new_n5106_));
NOR2X1 NOR2X1_425 ( .A(u2_o_364_), .B(u2__abc_52138_new_n5114_), .Y(u2__abc_52138_new_n5115_));
NOR2X1 NOR2X1_426 ( .A(u2_remHi_364_), .B(u2__abc_52138_new_n5116_), .Y(u2__abc_52138_new_n5117_));
NOR2X1 NOR2X1_427 ( .A(u2__abc_52138_new_n5115_), .B(u2__abc_52138_new_n5117_), .Y(u2__abc_52138_new_n5118_));
NOR2X1 NOR2X1_428 ( .A(u2_o_365_), .B(u2__abc_52138_new_n5119_), .Y(u2__abc_52138_new_n5120_));
NOR2X1 NOR2X1_429 ( .A(u2_remHi_365_), .B(u2__abc_52138_new_n5121_), .Y(u2__abc_52138_new_n5122_));
NOR2X1 NOR2X1_43 ( .A(\a[30] ), .B(\a[29] ), .Y(u1__abc_51895_new_n283_));
NOR2X1 NOR2X1_430 ( .A(u2__abc_52138_new_n5120_), .B(u2__abc_52138_new_n5122_), .Y(u2__abc_52138_new_n5123_));
NOR2X1 NOR2X1_431 ( .A(u2_o_363_), .B(u2__abc_52138_new_n5126_), .Y(u2__abc_52138_new_n5127_));
NOR2X1 NOR2X1_432 ( .A(u2_remHi_363_), .B(u2__abc_52138_new_n5128_), .Y(u2__abc_52138_new_n5129_));
NOR2X1 NOR2X1_433 ( .A(u2__abc_52138_new_n5127_), .B(u2__abc_52138_new_n5129_), .Y(u2__abc_52138_new_n5130_));
NOR2X1 NOR2X1_434 ( .A(u2_o_352_), .B(u2__abc_52138_new_n5134_), .Y(u2__abc_52138_new_n5135_));
NOR2X1 NOR2X1_435 ( .A(u2_remHi_352_), .B(u2__abc_52138_new_n5136_), .Y(u2__abc_52138_new_n5137_));
NOR2X1 NOR2X1_436 ( .A(u2__abc_52138_new_n5135_), .B(u2__abc_52138_new_n5137_), .Y(u2__abc_52138_new_n5138_));
NOR2X1 NOR2X1_437 ( .A(u2_o_353_), .B(u2__abc_52138_new_n5139_), .Y(u2__abc_52138_new_n5140_));
NOR2X1 NOR2X1_438 ( .A(u2_remHi_353_), .B(u2__abc_52138_new_n5141_), .Y(u2__abc_52138_new_n5142_));
NOR2X1 NOR2X1_439 ( .A(u2__abc_52138_new_n5140_), .B(u2__abc_52138_new_n5142_), .Y(u2__abc_52138_new_n5143_));
NOR2X1 NOR2X1_44 ( .A(\a[18] ), .B(\a[17] ), .Y(u1__abc_51895_new_n285_));
NOR2X1 NOR2X1_440 ( .A(u2_o_350_), .B(u2__abc_52138_new_n5145_), .Y(u2__abc_52138_new_n5146_));
NOR2X1 NOR2X1_441 ( .A(u2_remHi_350_), .B(u2__abc_52138_new_n5147_), .Y(u2__abc_52138_new_n5148_));
NOR2X1 NOR2X1_442 ( .A(u2__abc_52138_new_n5146_), .B(u2__abc_52138_new_n5148_), .Y(u2__abc_52138_new_n5149_));
NOR2X1 NOR2X1_443 ( .A(u2_o_351_), .B(u2__abc_52138_new_n5150_), .Y(u2__abc_52138_new_n5151_));
NOR2X1 NOR2X1_444 ( .A(u2_remHi_351_), .B(u2__abc_52138_new_n5152_), .Y(u2__abc_52138_new_n5153_));
NOR2X1 NOR2X1_445 ( .A(u2__abc_52138_new_n5151_), .B(u2__abc_52138_new_n5153_), .Y(u2__abc_52138_new_n5154_));
NOR2X1 NOR2X1_446 ( .A(u2__abc_52138_new_n5144_), .B(u2__abc_52138_new_n5155_), .Y(u2__abc_52138_new_n5156_));
NOR2X1 NOR2X1_447 ( .A(u2_o_356_), .B(u2__abc_52138_new_n5157_), .Y(u2__abc_52138_new_n5158_));
NOR2X1 NOR2X1_448 ( .A(u2_remHi_356_), .B(u2__abc_52138_new_n5159_), .Y(u2__abc_52138_new_n5160_));
NOR2X1 NOR2X1_449 ( .A(u2__abc_52138_new_n5158_), .B(u2__abc_52138_new_n5160_), .Y(u2__abc_52138_new_n5161_));
NOR2X1 NOR2X1_45 ( .A(\a[23] ), .B(\a[20] ), .Y(u1__abc_51895_new_n286_));
NOR2X1 NOR2X1_450 ( .A(u2_o_357_), .B(u2__abc_52138_new_n5162_), .Y(u2__abc_52138_new_n5163_));
NOR2X1 NOR2X1_451 ( .A(u2_remHi_357_), .B(u2__abc_52138_new_n5164_), .Y(u2__abc_52138_new_n5165_));
NOR2X1 NOR2X1_452 ( .A(u2__abc_52138_new_n5163_), .B(u2__abc_52138_new_n5165_), .Y(u2__abc_52138_new_n5166_));
NOR2X1 NOR2X1_453 ( .A(u2_o_354_), .B(u2__abc_52138_new_n5168_), .Y(u2__abc_52138_new_n5169_));
NOR2X1 NOR2X1_454 ( .A(u2_remHi_354_), .B(u2__abc_52138_new_n5170_), .Y(u2__abc_52138_new_n5171_));
NOR2X1 NOR2X1_455 ( .A(u2__abc_52138_new_n5169_), .B(u2__abc_52138_new_n5171_), .Y(u2__abc_52138_new_n5172_));
NOR2X1 NOR2X1_456 ( .A(u2_o_355_), .B(u2__abc_52138_new_n5173_), .Y(u2__abc_52138_new_n5174_));
NOR2X1 NOR2X1_457 ( .A(u2_remHi_355_), .B(u2__abc_52138_new_n5175_), .Y(u2__abc_52138_new_n5176_));
NOR2X1 NOR2X1_458 ( .A(u2__abc_52138_new_n5174_), .B(u2__abc_52138_new_n5176_), .Y(u2__abc_52138_new_n5177_));
NOR2X1 NOR2X1_459 ( .A(u2__abc_52138_new_n5167_), .B(u2__abc_52138_new_n5178_), .Y(u2__abc_52138_new_n5179_));
NOR2X1 NOR2X1_46 ( .A(u1__abc_51895_new_n284_), .B(u1__abc_51895_new_n287_), .Y(u1__abc_51895_new_n288_));
NOR2X1 NOR2X1_460 ( .A(u2__abc_52138_new_n5180_), .B(u2__abc_52138_new_n5133_), .Y(u2__abc_52138_new_n5181_));
NOR2X1 NOR2X1_461 ( .A(u2_o_345_), .B(u2__abc_52138_new_n5188_), .Y(u2__abc_52138_new_n5189_));
NOR2X1 NOR2X1_462 ( .A(u2_remHi_345_), .B(u2__abc_52138_new_n5190_), .Y(u2__abc_52138_new_n5191_));
NOR2X1 NOR2X1_463 ( .A(u2__abc_52138_new_n5189_), .B(u2__abc_52138_new_n5191_), .Y(u2__abc_52138_new_n5192_));
NOR2X1 NOR2X1_464 ( .A(u2_o_342_), .B(u2__abc_52138_new_n5195_), .Y(u2__abc_52138_new_n5196_));
NOR2X1 NOR2X1_465 ( .A(u2_remHi_342_), .B(u2__abc_52138_new_n5197_), .Y(u2__abc_52138_new_n5198_));
NOR2X1 NOR2X1_466 ( .A(u2__abc_52138_new_n5196_), .B(u2__abc_52138_new_n5198_), .Y(u2__abc_52138_new_n5199_));
NOR2X1 NOR2X1_467 ( .A(u2_o_343_), .B(u2__abc_52138_new_n5200_), .Y(u2__abc_52138_new_n5201_));
NOR2X1 NOR2X1_468 ( .A(u2_remHi_343_), .B(u2__abc_52138_new_n5202_), .Y(u2__abc_52138_new_n5203_));
NOR2X1 NOR2X1_469 ( .A(u2__abc_52138_new_n5201_), .B(u2__abc_52138_new_n5203_), .Y(u2__abc_52138_new_n5204_));
NOR2X1 NOR2X1_47 ( .A(\a[42] ), .B(\a[41] ), .Y(u1__abc_51895_new_n289_));
NOR2X1 NOR2X1_470 ( .A(u2_o_349_), .B(u2__abc_52138_new_n5210_), .Y(u2__abc_52138_new_n5211_));
NOR2X1 NOR2X1_471 ( .A(u2_remHi_349_), .B(u2__abc_52138_new_n5212_), .Y(u2__abc_52138_new_n5213_));
NOR2X1 NOR2X1_472 ( .A(u2__abc_52138_new_n5211_), .B(u2__abc_52138_new_n5213_), .Y(u2__abc_52138_new_n5214_));
NOR2X1 NOR2X1_473 ( .A(u2_o_346_), .B(u2__abc_52138_new_n5216_), .Y(u2__abc_52138_new_n5217_));
NOR2X1 NOR2X1_474 ( .A(u2_remHi_346_), .B(u2__abc_52138_new_n5218_), .Y(u2__abc_52138_new_n5219_));
NOR2X1 NOR2X1_475 ( .A(u2__abc_52138_new_n5217_), .B(u2__abc_52138_new_n5219_), .Y(u2__abc_52138_new_n5220_));
NOR2X1 NOR2X1_476 ( .A(u2_o_347_), .B(u2__abc_52138_new_n5221_), .Y(u2__abc_52138_new_n5222_));
NOR2X1 NOR2X1_477 ( .A(u2_remHi_347_), .B(u2__abc_52138_new_n5223_), .Y(u2__abc_52138_new_n5224_));
NOR2X1 NOR2X1_478 ( .A(u2__abc_52138_new_n5222_), .B(u2__abc_52138_new_n5224_), .Y(u2__abc_52138_new_n5225_));
NOR2X1 NOR2X1_479 ( .A(u2__abc_52138_new_n5227_), .B(u2__abc_52138_new_n5205_), .Y(u2__abc_52138_new_n5228_));
NOR2X1 NOR2X1_48 ( .A(\a[47] ), .B(\a[44] ), .Y(u1__abc_51895_new_n290_));
NOR2X1 NOR2X1_480 ( .A(u2_o_336_), .B(u2__abc_52138_new_n5229_), .Y(u2__abc_52138_new_n5230_));
NOR2X1 NOR2X1_481 ( .A(u2_remHi_336_), .B(u2__abc_52138_new_n5231_), .Y(u2__abc_52138_new_n5232_));
NOR2X1 NOR2X1_482 ( .A(u2__abc_52138_new_n5230_), .B(u2__abc_52138_new_n5232_), .Y(u2__abc_52138_new_n5233_));
NOR2X1 NOR2X1_483 ( .A(u2_o_337_), .B(u2__abc_52138_new_n5234_), .Y(u2__abc_52138_new_n5235_));
NOR2X1 NOR2X1_484 ( .A(u2_remHi_337_), .B(u2__abc_52138_new_n5236_), .Y(u2__abc_52138_new_n5237_));
NOR2X1 NOR2X1_485 ( .A(u2__abc_52138_new_n5235_), .B(u2__abc_52138_new_n5237_), .Y(u2__abc_52138_new_n5238_));
NOR2X1 NOR2X1_486 ( .A(u2_o_341_), .B(u2__abc_52138_new_n5254_), .Y(u2__abc_52138_new_n5255_));
NOR2X1 NOR2X1_487 ( .A(u2_remHi_341_), .B(u2__abc_52138_new_n5256_), .Y(u2__abc_52138_new_n5257_));
NOR2X1 NOR2X1_488 ( .A(u2__abc_52138_new_n5255_), .B(u2__abc_52138_new_n5257_), .Y(u2__abc_52138_new_n5258_));
NOR2X1 NOR2X1_489 ( .A(u2_o_338_), .B(u2__abc_52138_new_n5261_), .Y(u2__abc_52138_new_n5262_));
NOR2X1 NOR2X1_49 ( .A(\a[35] ), .B(\a[32] ), .Y(u1__abc_51895_new_n292_));
NOR2X1 NOR2X1_490 ( .A(u2_o_339_), .B(u2__abc_52138_new_n5266_), .Y(u2__abc_52138_new_n5267_));
NOR2X1 NOR2X1_491 ( .A(u2_remHi_339_), .B(u2__abc_52138_new_n5268_), .Y(u2__abc_52138_new_n5269_));
NOR2X1 NOR2X1_492 ( .A(u2__abc_52138_new_n5267_), .B(u2__abc_52138_new_n5269_), .Y(u2__abc_52138_new_n5270_));
NOR2X1 NOR2X1_493 ( .A(u2__abc_52138_new_n5271_), .B(u2__abc_52138_new_n5248_), .Y(u2__abc_52138_new_n5272_));
NOR2X1 NOR2X1_494 ( .A(u2_remHi_326_), .B(u2__abc_52138_new_n5274_), .Y(u2__abc_52138_new_n5275_));
NOR2X1 NOR2X1_495 ( .A(u2_o_326_), .B(u2__abc_52138_new_n5276_), .Y(u2__abc_52138_new_n5277_));
NOR2X1 NOR2X1_496 ( .A(u2__abc_52138_new_n5275_), .B(u2__abc_52138_new_n5277_), .Y(u2__abc_52138_new_n5278_));
NOR2X1 NOR2X1_497 ( .A(u2_o_328_), .B(u2__abc_52138_new_n5285_), .Y(u2__abc_52138_new_n5286_));
NOR2X1 NOR2X1_498 ( .A(u2_remHi_328_), .B(u2__abc_52138_new_n5287_), .Y(u2__abc_52138_new_n5288_));
NOR2X1 NOR2X1_499 ( .A(u2__abc_52138_new_n5286_), .B(u2__abc_52138_new_n5288_), .Y(u2__abc_52138_new_n5289_));
NOR2X1 NOR2X1_5 ( .A(_abc_65734_new_n1463_), .B(_abc_65734_new_n1466_), .Y(_abc_65734_new_n1467_));
NOR2X1 NOR2X1_50 ( .A(\a[38] ), .B(\a[37] ), .Y(u1__abc_51895_new_n293_));
NOR2X1 NOR2X1_500 ( .A(u2_o_329_), .B(u2__abc_52138_new_n5290_), .Y(u2__abc_52138_new_n5291_));
NOR2X1 NOR2X1_501 ( .A(u2_remHi_329_), .B(u2__abc_52138_new_n5292_), .Y(u2__abc_52138_new_n5293_));
NOR2X1 NOR2X1_502 ( .A(u2__abc_52138_new_n5291_), .B(u2__abc_52138_new_n5293_), .Y(u2__abc_52138_new_n5294_));
NOR2X1 NOR2X1_503 ( .A(u2__abc_52138_new_n5284_), .B(u2__abc_52138_new_n5295_), .Y(u2__abc_52138_new_n5296_));
NOR2X1 NOR2X1_504 ( .A(u2_o_332_), .B(u2__abc_52138_new_n5297_), .Y(u2__abc_52138_new_n5298_));
NOR2X1 NOR2X1_505 ( .A(u2_remHi_332_), .B(u2__abc_52138_new_n5299_), .Y(u2__abc_52138_new_n5300_));
NOR2X1 NOR2X1_506 ( .A(u2__abc_52138_new_n5298_), .B(u2__abc_52138_new_n5300_), .Y(u2__abc_52138_new_n5301_));
NOR2X1 NOR2X1_507 ( .A(u2_o_333_), .B(u2__abc_52138_new_n5302_), .Y(u2__abc_52138_new_n5303_));
NOR2X1 NOR2X1_508 ( .A(u2_remHi_333_), .B(u2__abc_52138_new_n5304_), .Y(u2__abc_52138_new_n5305_));
NOR2X1 NOR2X1_509 ( .A(u2__abc_52138_new_n5303_), .B(u2__abc_52138_new_n5305_), .Y(u2__abc_52138_new_n5306_));
NOR2X1 NOR2X1_51 ( .A(u1__abc_51895_new_n291_), .B(u1__abc_51895_new_n294_), .Y(u1__abc_51895_new_n295_));
NOR2X1 NOR2X1_510 ( .A(u2_o_330_), .B(u2__abc_52138_new_n5308_), .Y(u2__abc_52138_new_n5309_));
NOR2X1 NOR2X1_511 ( .A(u2_remHi_330_), .B(u2__abc_52138_new_n5310_), .Y(u2__abc_52138_new_n5311_));
NOR2X1 NOR2X1_512 ( .A(u2__abc_52138_new_n5309_), .B(u2__abc_52138_new_n5311_), .Y(u2__abc_52138_new_n5312_));
NOR2X1 NOR2X1_513 ( .A(u2_o_331_), .B(u2__abc_52138_new_n5313_), .Y(u2__abc_52138_new_n5314_));
NOR2X1 NOR2X1_514 ( .A(u2_remHi_331_), .B(u2__abc_52138_new_n5315_), .Y(u2__abc_52138_new_n5316_));
NOR2X1 NOR2X1_515 ( .A(u2__abc_52138_new_n5314_), .B(u2__abc_52138_new_n5316_), .Y(u2__abc_52138_new_n5317_));
NOR2X1 NOR2X1_516 ( .A(u2__abc_52138_new_n5307_), .B(u2__abc_52138_new_n5318_), .Y(u2__abc_52138_new_n5319_));
NOR2X1 NOR2X1_517 ( .A(u2_remHi_324_), .B(u2__abc_52138_new_n5321_), .Y(u2__abc_52138_new_n5322_));
NOR2X1 NOR2X1_518 ( .A(u2_o_324_), .B(u2__abc_52138_new_n5323_), .Y(u2__abc_52138_new_n5324_));
NOR2X1 NOR2X1_519 ( .A(u2__abc_52138_new_n5322_), .B(u2__abc_52138_new_n5324_), .Y(u2__abc_52138_new_n5325_));
NOR2X1 NOR2X1_52 ( .A(u1__abc_51895_new_n180_), .B(u1__abc_51895_new_n296_), .Y(u1__abc_51895_new_n297_));
NOR2X1 NOR2X1_520 ( .A(u2_remHi_325_), .B(u2__abc_52138_new_n5326_), .Y(u2__abc_52138_new_n5327_));
NOR2X1 NOR2X1_521 ( .A(u2_o_325_), .B(u2__abc_52138_new_n5328_), .Y(u2__abc_52138_new_n5329_));
NOR2X1 NOR2X1_522 ( .A(u2__abc_52138_new_n5327_), .B(u2__abc_52138_new_n5329_), .Y(u2__abc_52138_new_n5330_));
NOR2X1 NOR2X1_523 ( .A(u2__abc_52138_new_n5338_), .B(u2__abc_52138_new_n5331_), .Y(u2__abc_52138_new_n5339_));
NOR2X1 NOR2X1_524 ( .A(u2_remHi_318_), .B(u2__abc_52138_new_n5341_), .Y(u2__abc_52138_new_n5342_));
NOR2X1 NOR2X1_525 ( .A(u2_o_318_), .B(u2__abc_52138_new_n5343_), .Y(u2__abc_52138_new_n5344_));
NOR2X1 NOR2X1_526 ( .A(u2__abc_52138_new_n5342_), .B(u2__abc_52138_new_n5344_), .Y(u2__abc_52138_new_n5345_));
NOR2X1 NOR2X1_527 ( .A(u2_o_320_), .B(u2__abc_52138_new_n5352_), .Y(u2__abc_52138_new_n5353_));
NOR2X1 NOR2X1_528 ( .A(u2_remHi_320_), .B(u2__abc_52138_new_n5354_), .Y(u2__abc_52138_new_n5355_));
NOR2X1 NOR2X1_529 ( .A(u2__abc_52138_new_n5353_), .B(u2__abc_52138_new_n5355_), .Y(u2__abc_52138_new_n5356_));
NOR2X1 NOR2X1_53 ( .A(\a[91] ), .B(\a[88] ), .Y(u1__abc_51895_new_n298_));
NOR2X1 NOR2X1_530 ( .A(u2_o_321_), .B(u2__abc_52138_new_n5357_), .Y(u2__abc_52138_new_n5358_));
NOR2X1 NOR2X1_531 ( .A(u2_remHi_321_), .B(u2__abc_52138_new_n5359_), .Y(u2__abc_52138_new_n5360_));
NOR2X1 NOR2X1_532 ( .A(u2__abc_52138_new_n5358_), .B(u2__abc_52138_new_n5360_), .Y(u2__abc_52138_new_n5361_));
NOR2X1 NOR2X1_533 ( .A(u2__abc_52138_new_n5363_), .B(u2__abc_52138_new_n5340_), .Y(u2__abc_52138_new_n5364_));
NOR2X1 NOR2X1_534 ( .A(u2__abc_52138_new_n5365_), .B(u2__abc_52138_new_n5273_), .Y(u2__abc_52138_new_n5366_));
NOR2X1 NOR2X1_535 ( .A(u2_o_312_), .B(u2__abc_52138_new_n5368_), .Y(u2__abc_52138_new_n5369_));
NOR2X1 NOR2X1_536 ( .A(u2_remHi_312_), .B(u2__abc_52138_new_n5370_), .Y(u2__abc_52138_new_n5371_));
NOR2X1 NOR2X1_537 ( .A(u2__abc_52138_new_n5369_), .B(u2__abc_52138_new_n5371_), .Y(u2__abc_52138_new_n5372_));
NOR2X1 NOR2X1_538 ( .A(u2_o_313_), .B(u2__abc_52138_new_n5373_), .Y(u2__abc_52138_new_n5374_));
NOR2X1 NOR2X1_539 ( .A(u2_remHi_313_), .B(u2__abc_52138_new_n5375_), .Y(u2__abc_52138_new_n5376_));
NOR2X1 NOR2X1_54 ( .A(\a[94] ), .B(\a[93] ), .Y(u1__abc_51895_new_n299_));
NOR2X1 NOR2X1_540 ( .A(u2__abc_52138_new_n5374_), .B(u2__abc_52138_new_n5376_), .Y(u2__abc_52138_new_n5377_));
NOR2X1 NOR2X1_541 ( .A(u2_o_311_), .B(u2__abc_52138_new_n5380_), .Y(u2__abc_52138_new_n5381_));
NOR2X1 NOR2X1_542 ( .A(u2_remHi_311_), .B(u2__abc_52138_new_n5382_), .Y(u2__abc_52138_new_n5383_));
NOR2X1 NOR2X1_543 ( .A(u2__abc_52138_new_n5381_), .B(u2__abc_52138_new_n5383_), .Y(u2__abc_52138_new_n5384_));
NOR2X1 NOR2X1_544 ( .A(u2__abc_52138_new_n5385_), .B(u2__abc_52138_new_n5378_), .Y(u2__abc_52138_new_n5386_));
NOR2X1 NOR2X1_545 ( .A(u2_o_316_), .B(u2__abc_52138_new_n5387_), .Y(u2__abc_52138_new_n5388_));
NOR2X1 NOR2X1_546 ( .A(u2_remHi_316_), .B(u2__abc_52138_new_n5389_), .Y(u2__abc_52138_new_n5390_));
NOR2X1 NOR2X1_547 ( .A(u2__abc_52138_new_n5388_), .B(u2__abc_52138_new_n5390_), .Y(u2__abc_52138_new_n5391_));
NOR2X1 NOR2X1_548 ( .A(u2_o_317_), .B(u2__abc_52138_new_n5392_), .Y(u2__abc_52138_new_n5393_));
NOR2X1 NOR2X1_549 ( .A(u2_remHi_317_), .B(u2__abc_52138_new_n5394_), .Y(u2__abc_52138_new_n5395_));
NOR2X1 NOR2X1_55 ( .A(\a[82] ), .B(\a[81] ), .Y(u1__abc_51895_new_n301_));
NOR2X1 NOR2X1_550 ( .A(u2__abc_52138_new_n5393_), .B(u2__abc_52138_new_n5395_), .Y(u2__abc_52138_new_n5396_));
NOR2X1 NOR2X1_551 ( .A(u2_o_315_), .B(u2__abc_52138_new_n5399_), .Y(u2__abc_52138_new_n5400_));
NOR2X1 NOR2X1_552 ( .A(u2_remHi_315_), .B(u2__abc_52138_new_n5401_), .Y(u2__abc_52138_new_n5402_));
NOR2X1 NOR2X1_553 ( .A(u2__abc_52138_new_n5400_), .B(u2__abc_52138_new_n5402_), .Y(u2__abc_52138_new_n5403_));
NOR2X1 NOR2X1_554 ( .A(u2__abc_52138_new_n5404_), .B(u2__abc_52138_new_n5397_), .Y(u2__abc_52138_new_n5405_));
NOR2X1 NOR2X1_555 ( .A(u2_remHi_302_), .B(u2__abc_52138_new_n5407_), .Y(u2__abc_52138_new_n5408_));
NOR2X1 NOR2X1_556 ( .A(u2_o_302_), .B(u2__abc_52138_new_n5409_), .Y(u2__abc_52138_new_n5410_));
NOR2X1 NOR2X1_557 ( .A(u2__abc_52138_new_n5408_), .B(u2__abc_52138_new_n5410_), .Y(u2__abc_52138_new_n5411_));
NOR2X1 NOR2X1_558 ( .A(u2_remHi_303_), .B(u2__abc_52138_new_n5412_), .Y(u2__abc_52138_new_n5413_));
NOR2X1 NOR2X1_559 ( .A(u2_o_303_), .B(u2__abc_52138_new_n5414_), .Y(u2__abc_52138_new_n5415_));
NOR2X1 NOR2X1_56 ( .A(\a[87] ), .B(\a[84] ), .Y(u1__abc_51895_new_n302_));
NOR2X1 NOR2X1_560 ( .A(u2__abc_52138_new_n5413_), .B(u2__abc_52138_new_n5415_), .Y(u2__abc_52138_new_n5416_));
NOR2X1 NOR2X1_561 ( .A(u2_o_304_), .B(u2__abc_52138_new_n5418_), .Y(u2__abc_52138_new_n5419_));
NOR2X1 NOR2X1_562 ( .A(u2_remHi_304_), .B(u2__abc_52138_new_n5420_), .Y(u2__abc_52138_new_n5421_));
NOR2X1 NOR2X1_563 ( .A(u2__abc_52138_new_n5419_), .B(u2__abc_52138_new_n5421_), .Y(u2__abc_52138_new_n5422_));
NOR2X1 NOR2X1_564 ( .A(u2_o_305_), .B(u2__abc_52138_new_n5423_), .Y(u2__abc_52138_new_n5424_));
NOR2X1 NOR2X1_565 ( .A(u2_remHi_305_), .B(u2__abc_52138_new_n5425_), .Y(u2__abc_52138_new_n5426_));
NOR2X1 NOR2X1_566 ( .A(u2__abc_52138_new_n5424_), .B(u2__abc_52138_new_n5426_), .Y(u2__abc_52138_new_n5427_));
NOR2X1 NOR2X1_567 ( .A(u2__abc_52138_new_n5417_), .B(u2__abc_52138_new_n5428_), .Y(u2__abc_52138_new_n5429_));
NOR2X1 NOR2X1_568 ( .A(u2_o_308_), .B(u2__abc_52138_new_n5430_), .Y(u2__abc_52138_new_n5431_));
NOR2X1 NOR2X1_569 ( .A(u2_remHi_308_), .B(u2__abc_52138_new_n5432_), .Y(u2__abc_52138_new_n5433_));
NOR2X1 NOR2X1_57 ( .A(u1__abc_51895_new_n300_), .B(u1__abc_51895_new_n303_), .Y(u1__abc_51895_new_n304_));
NOR2X1 NOR2X1_570 ( .A(u2__abc_52138_new_n5431_), .B(u2__abc_52138_new_n5433_), .Y(u2__abc_52138_new_n5434_));
NOR2X1 NOR2X1_571 ( .A(u2_o_309_), .B(u2__abc_52138_new_n5435_), .Y(u2__abc_52138_new_n5436_));
NOR2X1 NOR2X1_572 ( .A(u2_remHi_309_), .B(u2__abc_52138_new_n5437_), .Y(u2__abc_52138_new_n5438_));
NOR2X1 NOR2X1_573 ( .A(u2__abc_52138_new_n5436_), .B(u2__abc_52138_new_n5438_), .Y(u2__abc_52138_new_n5439_));
NOR2X1 NOR2X1_574 ( .A(u2_o_307_), .B(u2__abc_52138_new_n5441_), .Y(u2__abc_52138_new_n5442_));
NOR2X1 NOR2X1_575 ( .A(u2_remHi_307_), .B(u2__abc_52138_new_n5443_), .Y(u2__abc_52138_new_n5444_));
NOR2X1 NOR2X1_576 ( .A(u2__abc_52138_new_n5442_), .B(u2__abc_52138_new_n5444_), .Y(u2__abc_52138_new_n5445_));
NOR2X1 NOR2X1_577 ( .A(u2_o_306_), .B(u2__abc_52138_new_n5446_), .Y(u2__abc_52138_new_n5447_));
NOR2X1 NOR2X1_578 ( .A(u2_remHi_306_), .B(u2__abc_52138_new_n5448_), .Y(u2__abc_52138_new_n5449_));
NOR2X1 NOR2X1_579 ( .A(u2__abc_52138_new_n5447_), .B(u2__abc_52138_new_n5449_), .Y(u2__abc_52138_new_n5450_));
NOR2X1 NOR2X1_58 ( .A(\a[106] ), .B(\a[105] ), .Y(u1__abc_51895_new_n305_));
NOR2X1 NOR2X1_580 ( .A(u2__abc_52138_new_n5440_), .B(u2__abc_52138_new_n5451_), .Y(u2__abc_52138_new_n5452_));
NOR2X1 NOR2X1_581 ( .A(u2__abc_52138_new_n5406_), .B(u2__abc_52138_new_n5453_), .Y(u2__abc_52138_new_n5454_));
NOR2X1 NOR2X1_582 ( .A(u2_remHi_294_), .B(u2__abc_52138_new_n5455_), .Y(u2__abc_52138_new_n5456_));
NOR2X1 NOR2X1_583 ( .A(u2_o_294_), .B(u2__abc_52138_new_n5457_), .Y(u2__abc_52138_new_n5458_));
NOR2X1 NOR2X1_584 ( .A(u2__abc_52138_new_n5456_), .B(u2__abc_52138_new_n5458_), .Y(u2__abc_52138_new_n5459_));
NOR2X1 NOR2X1_585 ( .A(u2_o_296_), .B(u2__abc_52138_new_n5466_), .Y(u2__abc_52138_new_n5467_));
NOR2X1 NOR2X1_586 ( .A(u2_remHi_296_), .B(u2__abc_52138_new_n5468_), .Y(u2__abc_52138_new_n5469_));
NOR2X1 NOR2X1_587 ( .A(u2__abc_52138_new_n5467_), .B(u2__abc_52138_new_n5469_), .Y(u2__abc_52138_new_n5470_));
NOR2X1 NOR2X1_588 ( .A(u2_o_297_), .B(u2__abc_52138_new_n5471_), .Y(u2__abc_52138_new_n5472_));
NOR2X1 NOR2X1_589 ( .A(u2_remHi_297_), .B(u2__abc_52138_new_n5473_), .Y(u2__abc_52138_new_n5474_));
NOR2X1 NOR2X1_59 ( .A(\a[111] ), .B(\a[108] ), .Y(u1__abc_51895_new_n306_));
NOR2X1 NOR2X1_590 ( .A(u2__abc_52138_new_n5472_), .B(u2__abc_52138_new_n5474_), .Y(u2__abc_52138_new_n5475_));
NOR2X1 NOR2X1_591 ( .A(u2__abc_52138_new_n5465_), .B(u2__abc_52138_new_n5476_), .Y(u2__abc_52138_new_n5477_));
NOR2X1 NOR2X1_592 ( .A(u2_o_300_), .B(u2__abc_52138_new_n5478_), .Y(u2__abc_52138_new_n5479_));
NOR2X1 NOR2X1_593 ( .A(u2_remHi_300_), .B(u2__abc_52138_new_n5480_), .Y(u2__abc_52138_new_n5481_));
NOR2X1 NOR2X1_594 ( .A(u2__abc_52138_new_n5479_), .B(u2__abc_52138_new_n5481_), .Y(u2__abc_52138_new_n5482_));
NOR2X1 NOR2X1_595 ( .A(u2_o_301_), .B(u2__abc_52138_new_n5483_), .Y(u2__abc_52138_new_n5484_));
NOR2X1 NOR2X1_596 ( .A(u2_remHi_301_), .B(u2__abc_52138_new_n5485_), .Y(u2__abc_52138_new_n5486_));
NOR2X1 NOR2X1_597 ( .A(u2__abc_52138_new_n5484_), .B(u2__abc_52138_new_n5486_), .Y(u2__abc_52138_new_n5487_));
NOR2X1 NOR2X1_598 ( .A(u2_o_298_), .B(u2__abc_52138_new_n5489_), .Y(u2__abc_52138_new_n5490_));
NOR2X1 NOR2X1_599 ( .A(u2_remHi_298_), .B(u2__abc_52138_new_n5491_), .Y(u2__abc_52138_new_n5492_));
NOR2X1 NOR2X1_6 ( .A(_abc_65734_new_n1473_), .B(_abc_65734_new_n1465_), .Y(_abc_65734_new_n1476_));
NOR2X1 NOR2X1_60 ( .A(\a[99] ), .B(\a[96] ), .Y(u1__abc_51895_new_n308_));
NOR2X1 NOR2X1_600 ( .A(u2__abc_52138_new_n5490_), .B(u2__abc_52138_new_n5492_), .Y(u2__abc_52138_new_n5493_));
NOR2X1 NOR2X1_601 ( .A(u2_o_299_), .B(u2__abc_52138_new_n5494_), .Y(u2__abc_52138_new_n5495_));
NOR2X1 NOR2X1_602 ( .A(u2_remHi_299_), .B(u2__abc_52138_new_n5496_), .Y(u2__abc_52138_new_n5497_));
NOR2X1 NOR2X1_603 ( .A(u2__abc_52138_new_n5495_), .B(u2__abc_52138_new_n5497_), .Y(u2__abc_52138_new_n5498_));
NOR2X1 NOR2X1_604 ( .A(u2__abc_52138_new_n5488_), .B(u2__abc_52138_new_n5499_), .Y(u2__abc_52138_new_n5500_));
NOR2X1 NOR2X1_605 ( .A(u2_o_288_), .B(u2__abc_52138_new_n5502_), .Y(u2__abc_52138_new_n5503_));
NOR2X1 NOR2X1_606 ( .A(u2_remHi_288_), .B(u2__abc_52138_new_n5504_), .Y(u2__abc_52138_new_n5505_));
NOR2X1 NOR2X1_607 ( .A(u2__abc_52138_new_n5503_), .B(u2__abc_52138_new_n5505_), .Y(u2__abc_52138_new_n5506_));
NOR2X1 NOR2X1_608 ( .A(u2_o_289_), .B(u2__abc_52138_new_n5507_), .Y(u2__abc_52138_new_n5508_));
NOR2X1 NOR2X1_609 ( .A(u2_remHi_289_), .B(u2__abc_52138_new_n5509_), .Y(u2__abc_52138_new_n5510_));
NOR2X1 NOR2X1_61 ( .A(\a[102] ), .B(\a[101] ), .Y(u1__abc_51895_new_n309_));
NOR2X1 NOR2X1_610 ( .A(u2__abc_52138_new_n5508_), .B(u2__abc_52138_new_n5510_), .Y(u2__abc_52138_new_n5511_));
NOR2X1 NOR2X1_611 ( .A(u2_o_286_), .B(u2__abc_52138_new_n5513_), .Y(u2__abc_52138_new_n5514_));
NOR2X1 NOR2X1_612 ( .A(u2_remHi_286_), .B(u2__abc_52138_new_n5515_), .Y(u2__abc_52138_new_n5516_));
NOR2X1 NOR2X1_613 ( .A(u2__abc_52138_new_n5514_), .B(u2__abc_52138_new_n5516_), .Y(u2__abc_52138_new_n5517_));
NOR2X1 NOR2X1_614 ( .A(u2_o_287_), .B(u2__abc_52138_new_n5518_), .Y(u2__abc_52138_new_n5519_));
NOR2X1 NOR2X1_615 ( .A(u2_remHi_287_), .B(u2__abc_52138_new_n5520_), .Y(u2__abc_52138_new_n5521_));
NOR2X1 NOR2X1_616 ( .A(u2__abc_52138_new_n5519_), .B(u2__abc_52138_new_n5521_), .Y(u2__abc_52138_new_n5522_));
NOR2X1 NOR2X1_617 ( .A(u2__abc_52138_new_n5512_), .B(u2__abc_52138_new_n5523_), .Y(u2__abc_52138_new_n5524_));
NOR2X1 NOR2X1_618 ( .A(u2_o_292_), .B(u2__abc_52138_new_n5525_), .Y(u2__abc_52138_new_n5526_));
NOR2X1 NOR2X1_619 ( .A(u2_remHi_292_), .B(u2__abc_52138_new_n5527_), .Y(u2__abc_52138_new_n5528_));
NOR2X1 NOR2X1_62 ( .A(u1__abc_51895_new_n307_), .B(u1__abc_51895_new_n310_), .Y(u1__abc_51895_new_n311_));
NOR2X1 NOR2X1_620 ( .A(u2__abc_52138_new_n5526_), .B(u2__abc_52138_new_n5528_), .Y(u2__abc_52138_new_n5529_));
NOR2X1 NOR2X1_621 ( .A(u2_o_293_), .B(u2__abc_52138_new_n5530_), .Y(u2__abc_52138_new_n5531_));
NOR2X1 NOR2X1_622 ( .A(u2_remHi_293_), .B(u2__abc_52138_new_n5532_), .Y(u2__abc_52138_new_n5533_));
NOR2X1 NOR2X1_623 ( .A(u2__abc_52138_new_n5531_), .B(u2__abc_52138_new_n5533_), .Y(u2__abc_52138_new_n5534_));
NOR2X1 NOR2X1_624 ( .A(u2_o_291_), .B(u2__abc_52138_new_n5537_), .Y(u2__abc_52138_new_n5538_));
NOR2X1 NOR2X1_625 ( .A(u2_remHi_291_), .B(u2__abc_52138_new_n5539_), .Y(u2__abc_52138_new_n5540_));
NOR2X1 NOR2X1_626 ( .A(u2__abc_52138_new_n5538_), .B(u2__abc_52138_new_n5540_), .Y(u2__abc_52138_new_n5541_));
NOR2X1 NOR2X1_627 ( .A(u2__abc_52138_new_n5542_), .B(u2__abc_52138_new_n5535_), .Y(u2__abc_52138_new_n5543_));
NOR2X1 NOR2X1_628 ( .A(u2__abc_52138_new_n5501_), .B(u2__abc_52138_new_n5544_), .Y(u2__abc_52138_new_n5545_));
NOR2X1 NOR2X1_629 ( .A(u2_o_280_), .B(u2__abc_52138_new_n5548_), .Y(u2__abc_52138_new_n5549_));
NOR2X1 NOR2X1_63 ( .A(\a[58] ), .B(\a[57] ), .Y(u1__abc_51895_new_n313_));
NOR2X1 NOR2X1_630 ( .A(u2_remHi_280_), .B(u2__abc_52138_new_n5550_), .Y(u2__abc_52138_new_n5551_));
NOR2X1 NOR2X1_631 ( .A(u2__abc_52138_new_n5549_), .B(u2__abc_52138_new_n5551_), .Y(u2__abc_52138_new_n5552_));
NOR2X1 NOR2X1_632 ( .A(u2_o_281_), .B(u2__abc_52138_new_n5553_), .Y(u2__abc_52138_new_n5554_));
NOR2X1 NOR2X1_633 ( .A(u2_remHi_281_), .B(u2__abc_52138_new_n5555_), .Y(u2__abc_52138_new_n5556_));
NOR2X1 NOR2X1_634 ( .A(u2__abc_52138_new_n5554_), .B(u2__abc_52138_new_n5556_), .Y(u2__abc_52138_new_n5557_));
NOR2X1 NOR2X1_635 ( .A(u2_o_278_), .B(u2__abc_52138_new_n5559_), .Y(u2__abc_52138_new_n5560_));
NOR2X1 NOR2X1_636 ( .A(u2_remHi_278_), .B(u2__abc_52138_new_n5561_), .Y(u2__abc_52138_new_n5562_));
NOR2X1 NOR2X1_637 ( .A(u2__abc_52138_new_n5560_), .B(u2__abc_52138_new_n5562_), .Y(u2__abc_52138_new_n5563_));
NOR2X1 NOR2X1_638 ( .A(u2_o_279_), .B(u2__abc_52138_new_n5564_), .Y(u2__abc_52138_new_n5565_));
NOR2X1 NOR2X1_639 ( .A(u2_remHi_279_), .B(u2__abc_52138_new_n5566_), .Y(u2__abc_52138_new_n5567_));
NOR2X1 NOR2X1_64 ( .A(\a[63] ), .B(\a[60] ), .Y(u1__abc_51895_new_n314_));
NOR2X1 NOR2X1_640 ( .A(u2__abc_52138_new_n5565_), .B(u2__abc_52138_new_n5567_), .Y(u2__abc_52138_new_n5568_));
NOR2X1 NOR2X1_641 ( .A(u2__abc_52138_new_n5558_), .B(u2__abc_52138_new_n5569_), .Y(u2__abc_52138_new_n5570_));
NOR2X1 NOR2X1_642 ( .A(u2_o_284_), .B(u2__abc_52138_new_n5571_), .Y(u2__abc_52138_new_n5572_));
NOR2X1 NOR2X1_643 ( .A(u2_remHi_284_), .B(u2__abc_52138_new_n5573_), .Y(u2__abc_52138_new_n5574_));
NOR2X1 NOR2X1_644 ( .A(u2__abc_52138_new_n5572_), .B(u2__abc_52138_new_n5574_), .Y(u2__abc_52138_new_n5575_));
NOR2X1 NOR2X1_645 ( .A(u2_o_285_), .B(u2__abc_52138_new_n5576_), .Y(u2__abc_52138_new_n5577_));
NOR2X1 NOR2X1_646 ( .A(u2_remHi_285_), .B(u2__abc_52138_new_n5578_), .Y(u2__abc_52138_new_n5579_));
NOR2X1 NOR2X1_647 ( .A(u2__abc_52138_new_n5577_), .B(u2__abc_52138_new_n5579_), .Y(u2__abc_52138_new_n5580_));
NOR2X1 NOR2X1_648 ( .A(u2_o_282_), .B(u2__abc_52138_new_n5582_), .Y(u2__abc_52138_new_n5583_));
NOR2X1 NOR2X1_649 ( .A(u2_remHi_282_), .B(u2__abc_52138_new_n5584_), .Y(u2__abc_52138_new_n5585_));
NOR2X1 NOR2X1_65 ( .A(\a[51] ), .B(\a[48] ), .Y(u1__abc_51895_new_n316_));
NOR2X1 NOR2X1_650 ( .A(u2__abc_52138_new_n5583_), .B(u2__abc_52138_new_n5585_), .Y(u2__abc_52138_new_n5586_));
NOR2X1 NOR2X1_651 ( .A(u2_o_283_), .B(u2__abc_52138_new_n5587_), .Y(u2__abc_52138_new_n5588_));
NOR2X1 NOR2X1_652 ( .A(u2_remHi_283_), .B(u2__abc_52138_new_n5589_), .Y(u2__abc_52138_new_n5590_));
NOR2X1 NOR2X1_653 ( .A(u2__abc_52138_new_n5588_), .B(u2__abc_52138_new_n5590_), .Y(u2__abc_52138_new_n5591_));
NOR2X1 NOR2X1_654 ( .A(u2__abc_52138_new_n5581_), .B(u2__abc_52138_new_n5592_), .Y(u2__abc_52138_new_n5593_));
NOR2X1 NOR2X1_655 ( .A(u2_o_272_), .B(u2__abc_52138_new_n5595_), .Y(u2__abc_52138_new_n5596_));
NOR2X1 NOR2X1_656 ( .A(u2_remHi_272_), .B(u2__abc_52138_new_n5597_), .Y(u2__abc_52138_new_n5598_));
NOR2X1 NOR2X1_657 ( .A(u2__abc_52138_new_n5596_), .B(u2__abc_52138_new_n5598_), .Y(u2__abc_52138_new_n5599_));
NOR2X1 NOR2X1_658 ( .A(u2_o_273_), .B(u2__abc_52138_new_n5600_), .Y(u2__abc_52138_new_n5601_));
NOR2X1 NOR2X1_659 ( .A(u2_remHi_273_), .B(u2__abc_52138_new_n5602_), .Y(u2__abc_52138_new_n5603_));
NOR2X1 NOR2X1_66 ( .A(\a[54] ), .B(\a[53] ), .Y(u1__abc_51895_new_n317_));
NOR2X1 NOR2X1_660 ( .A(u2__abc_52138_new_n5601_), .B(u2__abc_52138_new_n5603_), .Y(u2__abc_52138_new_n5604_));
NOR2X1 NOR2X1_661 ( .A(u2_o_270_), .B(u2__abc_52138_new_n5606_), .Y(u2__abc_52138_new_n5607_));
NOR2X1 NOR2X1_662 ( .A(u2_remHi_270_), .B(u2__abc_52138_new_n5608_), .Y(u2__abc_52138_new_n5609_));
NOR2X1 NOR2X1_663 ( .A(u2__abc_52138_new_n5607_), .B(u2__abc_52138_new_n5609_), .Y(u2__abc_52138_new_n5610_));
NOR2X1 NOR2X1_664 ( .A(u2_o_271_), .B(u2__abc_52138_new_n5611_), .Y(u2__abc_52138_new_n5612_));
NOR2X1 NOR2X1_665 ( .A(u2_remHi_271_), .B(u2__abc_52138_new_n5613_), .Y(u2__abc_52138_new_n5614_));
NOR2X1 NOR2X1_666 ( .A(u2__abc_52138_new_n5612_), .B(u2__abc_52138_new_n5614_), .Y(u2__abc_52138_new_n5615_));
NOR2X1 NOR2X1_667 ( .A(u2__abc_52138_new_n5605_), .B(u2__abc_52138_new_n5616_), .Y(u2__abc_52138_new_n5617_));
NOR2X1 NOR2X1_668 ( .A(u2_o_276_), .B(u2__abc_52138_new_n5618_), .Y(u2__abc_52138_new_n5619_));
NOR2X1 NOR2X1_669 ( .A(u2_remHi_276_), .B(u2__abc_52138_new_n5620_), .Y(u2__abc_52138_new_n5621_));
NOR2X1 NOR2X1_67 ( .A(u1__abc_51895_new_n315_), .B(u1__abc_51895_new_n318_), .Y(u1__abc_51895_new_n319_));
NOR2X1 NOR2X1_670 ( .A(u2__abc_52138_new_n5619_), .B(u2__abc_52138_new_n5621_), .Y(u2__abc_52138_new_n5622_));
NOR2X1 NOR2X1_671 ( .A(u2_o_277_), .B(u2__abc_52138_new_n5623_), .Y(u2__abc_52138_new_n5624_));
NOR2X1 NOR2X1_672 ( .A(u2_remHi_277_), .B(u2__abc_52138_new_n5625_), .Y(u2__abc_52138_new_n5626_));
NOR2X1 NOR2X1_673 ( .A(u2__abc_52138_new_n5624_), .B(u2__abc_52138_new_n5626_), .Y(u2__abc_52138_new_n5627_));
NOR2X1 NOR2X1_674 ( .A(u2_o_275_), .B(u2__abc_52138_new_n5630_), .Y(u2__abc_52138_new_n5631_));
NOR2X1 NOR2X1_675 ( .A(u2_remHi_275_), .B(u2__abc_52138_new_n5632_), .Y(u2__abc_52138_new_n5633_));
NOR2X1 NOR2X1_676 ( .A(u2__abc_52138_new_n5631_), .B(u2__abc_52138_new_n5633_), .Y(u2__abc_52138_new_n5634_));
NOR2X1 NOR2X1_677 ( .A(u2__abc_52138_new_n5635_), .B(u2__abc_52138_new_n5628_), .Y(u2__abc_52138_new_n5636_));
NOR2X1 NOR2X1_678 ( .A(u2__abc_52138_new_n5637_), .B(u2__abc_52138_new_n5594_), .Y(u2__abc_52138_new_n5638_));
NOR2X1 NOR2X1_679 ( .A(u2_remHi_268_), .B(u2__abc_52138_new_n5640_), .Y(u2__abc_52138_new_n5641_));
NOR2X1 NOR2X1_68 ( .A(\a[75] ), .B(\a[72] ), .Y(u1__abc_51895_new_n320_));
NOR2X1 NOR2X1_680 ( .A(u2_o_268_), .B(u2__abc_52138_new_n5642_), .Y(u2__abc_52138_new_n5643_));
NOR2X1 NOR2X1_681 ( .A(u2__abc_52138_new_n5641_), .B(u2__abc_52138_new_n5643_), .Y(u2__abc_52138_new_n5644_));
NOR2X1 NOR2X1_682 ( .A(u2_remHi_269_), .B(u2__abc_52138_new_n5645_), .Y(u2__abc_52138_new_n5646_));
NOR2X1 NOR2X1_683 ( .A(u2_o_269_), .B(u2__abc_52138_new_n5647_), .Y(u2__abc_52138_new_n5648_));
NOR2X1 NOR2X1_684 ( .A(u2__abc_52138_new_n5646_), .B(u2__abc_52138_new_n5648_), .Y(u2__abc_52138_new_n5649_));
NOR2X1 NOR2X1_685 ( .A(u2_o_266_), .B(u2__abc_52138_new_n5651_), .Y(u2__abc_52138_new_n5652_));
NOR2X1 NOR2X1_686 ( .A(u2_remHi_266_), .B(u2__abc_52138_new_n5653_), .Y(u2__abc_52138_new_n5654_));
NOR2X1 NOR2X1_687 ( .A(u2__abc_52138_new_n5652_), .B(u2__abc_52138_new_n5654_), .Y(u2__abc_52138_new_n5655_));
NOR2X1 NOR2X1_688 ( .A(u2_o_267_), .B(u2__abc_52138_new_n5656_), .Y(u2__abc_52138_new_n5657_));
NOR2X1 NOR2X1_689 ( .A(u2_remHi_267_), .B(u2__abc_52138_new_n5658_), .Y(u2__abc_52138_new_n5659_));
NOR2X1 NOR2X1_69 ( .A(\a[78] ), .B(\a[77] ), .Y(u1__abc_51895_new_n321_));
NOR2X1 NOR2X1_690 ( .A(u2__abc_52138_new_n5657_), .B(u2__abc_52138_new_n5659_), .Y(u2__abc_52138_new_n5660_));
NOR2X1 NOR2X1_691 ( .A(u2__abc_52138_new_n5650_), .B(u2__abc_52138_new_n5661_), .Y(u2__abc_52138_new_n5662_));
NOR2X1 NOR2X1_692 ( .A(u2_o_264_), .B(u2__abc_52138_new_n5663_), .Y(u2__abc_52138_new_n5664_));
NOR2X1 NOR2X1_693 ( .A(u2_remHi_264_), .B(u2__abc_52138_new_n5665_), .Y(u2__abc_52138_new_n5666_));
NOR2X1 NOR2X1_694 ( .A(u2__abc_52138_new_n5664_), .B(u2__abc_52138_new_n5666_), .Y(u2__abc_52138_new_n5667_));
NOR2X1 NOR2X1_695 ( .A(u2_o_265_), .B(u2__abc_52138_new_n5668_), .Y(u2__abc_52138_new_n5669_));
NOR2X1 NOR2X1_696 ( .A(u2_remHi_265_), .B(u2__abc_52138_new_n5670_), .Y(u2__abc_52138_new_n5671_));
NOR2X1 NOR2X1_697 ( .A(u2__abc_52138_new_n5669_), .B(u2__abc_52138_new_n5671_), .Y(u2__abc_52138_new_n5672_));
NOR2X1 NOR2X1_698 ( .A(u2_remHi_262_), .B(u2__abc_52138_new_n5674_), .Y(u2__abc_52138_new_n5675_));
NOR2X1 NOR2X1_699 ( .A(u2_o_262_), .B(u2__abc_52138_new_n5676_), .Y(u2__abc_52138_new_n5677_));
NOR2X1 NOR2X1_7 ( .A(_abc_65734_new_n1461_), .B(_abc_65734_new_n1462_), .Y(_abc_65734_new_n1479_));
NOR2X1 NOR2X1_70 ( .A(\a[66] ), .B(\a[65] ), .Y(u1__abc_51895_new_n323_));
NOR2X1 NOR2X1_700 ( .A(u2__abc_52138_new_n5675_), .B(u2__abc_52138_new_n5677_), .Y(u2__abc_52138_new_n5678_));
NOR2X1 NOR2X1_701 ( .A(u2_remHi_263_), .B(u2__abc_52138_new_n5679_), .Y(u2__abc_52138_new_n5680_));
NOR2X1 NOR2X1_702 ( .A(u2_o_263_), .B(u2__abc_52138_new_n5681_), .Y(u2__abc_52138_new_n5682_));
NOR2X1 NOR2X1_703 ( .A(u2__abc_52138_new_n5680_), .B(u2__abc_52138_new_n5682_), .Y(u2__abc_52138_new_n5683_));
NOR2X1 NOR2X1_704 ( .A(u2__abc_52138_new_n5673_), .B(u2__abc_52138_new_n5684_), .Y(u2__abc_52138_new_n5685_));
NOR2X1 NOR2X1_705 ( .A(u2__abc_52138_new_n5690_), .B(u2__abc_52138_new_n5694_), .Y(u2__abc_52138_new_n5695_));
NOR2X1 NOR2X1_706 ( .A(u2_o_256_), .B(u2__abc_52138_new_n5697_), .Y(u2__abc_52138_new_n5698_));
NOR2X1 NOR2X1_707 ( .A(u2_remHi_256_), .B(u2__abc_52138_new_n5699_), .Y(u2__abc_52138_new_n5700_));
NOR2X1 NOR2X1_708 ( .A(u2__abc_52138_new_n5698_), .B(u2__abc_52138_new_n5700_), .Y(u2__abc_52138_new_n5701_));
NOR2X1 NOR2X1_709 ( .A(u2_o_257_), .B(u2__abc_52138_new_n5702_), .Y(u2__abc_52138_new_n5703_));
NOR2X1 NOR2X1_71 ( .A(\a[71] ), .B(\a[68] ), .Y(u1__abc_51895_new_n324_));
NOR2X1 NOR2X1_710 ( .A(u2_remHi_257_), .B(u2__abc_52138_new_n5704_), .Y(u2__abc_52138_new_n5705_));
NOR2X1 NOR2X1_711 ( .A(u2__abc_52138_new_n5703_), .B(u2__abc_52138_new_n5705_), .Y(u2__abc_52138_new_n5706_));
NOR2X1 NOR2X1_712 ( .A(u2__abc_52138_new_n5707_), .B(u2__abc_52138_new_n5696_), .Y(u2__abc_52138_new_n5708_));
NOR2X1 NOR2X1_713 ( .A(u2_o_260_), .B(u2__abc_52138_new_n5709_), .Y(u2__abc_52138_new_n5710_));
NOR2X1 NOR2X1_714 ( .A(u2_remHi_260_), .B(u2__abc_52138_new_n5711_), .Y(u2__abc_52138_new_n5712_));
NOR2X1 NOR2X1_715 ( .A(u2__abc_52138_new_n5710_), .B(u2__abc_52138_new_n5712_), .Y(u2__abc_52138_new_n5713_));
NOR2X1 NOR2X1_716 ( .A(u2_o_261_), .B(u2__abc_52138_new_n5714_), .Y(u2__abc_52138_new_n5715_));
NOR2X1 NOR2X1_717 ( .A(u2_remHi_261_), .B(u2__abc_52138_new_n5716_), .Y(u2__abc_52138_new_n5717_));
NOR2X1 NOR2X1_718 ( .A(u2__abc_52138_new_n5715_), .B(u2__abc_52138_new_n5717_), .Y(u2__abc_52138_new_n5718_));
NOR2X1 NOR2X1_719 ( .A(u2_o_258_), .B(u2__abc_52138_new_n5720_), .Y(u2__abc_52138_new_n5721_));
NOR2X1 NOR2X1_72 ( .A(u1__abc_51895_new_n322_), .B(u1__abc_51895_new_n325_), .Y(u1__abc_51895_new_n326_));
NOR2X1 NOR2X1_720 ( .A(u2_remHi_258_), .B(u2__abc_52138_new_n5722_), .Y(u2__abc_52138_new_n5723_));
NOR2X1 NOR2X1_721 ( .A(u2__abc_52138_new_n5721_), .B(u2__abc_52138_new_n5723_), .Y(u2__abc_52138_new_n5724_));
NOR2X1 NOR2X1_722 ( .A(u2_o_259_), .B(u2__abc_52138_new_n5725_), .Y(u2__abc_52138_new_n5726_));
NOR2X1 NOR2X1_723 ( .A(u2_remHi_259_), .B(u2__abc_52138_new_n5727_), .Y(u2__abc_52138_new_n5728_));
NOR2X1 NOR2X1_724 ( .A(u2__abc_52138_new_n5726_), .B(u2__abc_52138_new_n5728_), .Y(u2__abc_52138_new_n5729_));
NOR2X1 NOR2X1_725 ( .A(u2__abc_52138_new_n5719_), .B(u2__abc_52138_new_n5730_), .Y(u2__abc_52138_new_n5731_));
NOR2X1 NOR2X1_726 ( .A(u2__abc_52138_new_n5733_), .B(u2__abc_52138_new_n5639_), .Y(u2__abc_52138_new_n5734_));
NOR2X1 NOR2X1_727 ( .A(u2__abc_52138_new_n5735_), .B(u2__abc_52138_new_n5367_), .Y(u2__abc_52138_new_n5736_));
NOR2X1 NOR2X1_728 ( .A(u2__abc_52138_new_n5686_), .B(u2__abc_52138_new_n5745_), .Y(u2__abc_52138_new_n5746_));
NOR2X1 NOR2X1_729 ( .A(u2__abc_52138_new_n5594_), .B(u2__abc_52138_new_n5766_), .Y(u2__abc_52138_new_n5767_));
NOR2X1 NOR2X1_73 ( .A(u1__abc_51895_new_n312_), .B(u1__abc_51895_new_n327_), .Y(u1__abc_51895_new_n328_));
NOR2X1 NOR2X1_730 ( .A(u2__abc_52138_new_n5779_), .B(u2__abc_52138_new_n5767_), .Y(u2__abc_52138_new_n5780_));
NOR2X1 NOR2X1_731 ( .A(u2__abc_52138_new_n5501_), .B(u2__abc_52138_new_n5793_), .Y(u2__abc_52138_new_n5794_));
NOR2X1 NOR2X1_732 ( .A(u2__abc_52138_new_n5369_), .B(u2__abc_52138_new_n5381_), .Y(u2__abc_52138_new_n5814_));
NOR2X1 NOR2X1_733 ( .A(u2__abc_52138_new_n5406_), .B(u2__abc_52138_new_n5831_), .Y(u2__abc_52138_new_n5832_));
NOR2X1 NOR2X1_734 ( .A(u2__abc_52138_new_n5823_), .B(u2__abc_52138_new_n5832_), .Y(u2__abc_52138_new_n5833_));
NOR2X1 NOR2X1_735 ( .A(u2__abc_52138_new_n5869_), .B(u2__abc_52138_new_n5867_), .Y(u2__abc_52138_new_n5870_));
NOR2X1 NOR2X1_736 ( .A(u2__abc_52138_new_n5926_), .B(u2__abc_52138_new_n5133_), .Y(u2__abc_52138_new_n5927_));
NOR2X1 NOR2X1_737 ( .A(u2_o_444_), .B(u2__abc_52138_new_n5944_), .Y(u2__abc_52138_new_n5945_));
NOR2X1 NOR2X1_738 ( .A(u2_remHi_444_), .B(u2__abc_52138_new_n5946_), .Y(u2__abc_52138_new_n5947_));
NOR2X1 NOR2X1_739 ( .A(u2__abc_52138_new_n5945_), .B(u2__abc_52138_new_n5947_), .Y(u2__abc_52138_new_n5948_));
NOR2X1 NOR2X1_74 ( .A(\a[26] ), .B(\a[25] ), .Y(u1__abc_51895_new_n330_));
NOR2X1 NOR2X1_740 ( .A(u2_remHi_445_), .B(u2__abc_52138_new_n5949_), .Y(u2__abc_52138_new_n5950_));
NOR2X1 NOR2X1_741 ( .A(u2_o_445_), .B(u2__abc_52138_new_n5951_), .Y(u2__abc_52138_new_n5952_));
NOR2X1 NOR2X1_742 ( .A(u2__abc_52138_new_n5950_), .B(u2__abc_52138_new_n5952_), .Y(u2__abc_52138_new_n5953_));
NOR2X1 NOR2X1_743 ( .A(u2_remHi_443_), .B(u2__abc_52138_new_n5955_), .Y(u2__abc_52138_new_n5956_));
NOR2X1 NOR2X1_744 ( .A(u2_o_443_), .B(u2__abc_52138_new_n5957_), .Y(u2__abc_52138_new_n5958_));
NOR2X1 NOR2X1_745 ( .A(u2__abc_52138_new_n5956_), .B(u2__abc_52138_new_n5958_), .Y(u2__abc_52138_new_n5959_));
NOR2X1 NOR2X1_746 ( .A(u2_o_442_), .B(u2__abc_52138_new_n5960_), .Y(u2__abc_52138_new_n5961_));
NOR2X1 NOR2X1_747 ( .A(u2_remHi_442_), .B(u2__abc_52138_new_n5962_), .Y(u2__abc_52138_new_n5963_));
NOR2X1 NOR2X1_748 ( .A(u2__abc_52138_new_n5961_), .B(u2__abc_52138_new_n5963_), .Y(u2__abc_52138_new_n5964_));
NOR2X1 NOR2X1_749 ( .A(u2__abc_52138_new_n5954_), .B(u2__abc_52138_new_n5965_), .Y(u2__abc_52138_new_n5966_));
NOR2X1 NOR2X1_75 ( .A(\a[31] ), .B(\a[28] ), .Y(u1__abc_51895_new_n331_));
NOR2X1 NOR2X1_750 ( .A(u2_o_438_), .B(u2__abc_52138_new_n5967_), .Y(u2__abc_52138_new_n5968_));
NOR2X1 NOR2X1_751 ( .A(u2_remHi_438_), .B(u2__abc_52138_new_n5969_), .Y(u2__abc_52138_new_n5970_));
NOR2X1 NOR2X1_752 ( .A(u2__abc_52138_new_n5968_), .B(u2__abc_52138_new_n5970_), .Y(u2__abc_52138_new_n5971_));
NOR2X1 NOR2X1_753 ( .A(u2_o_440_), .B(u2__abc_52138_new_n5974_), .Y(u2__abc_52138_new_n5975_));
NOR2X1 NOR2X1_754 ( .A(u2_remHi_440_), .B(u2__abc_52138_new_n5976_), .Y(u2__abc_52138_new_n5977_));
NOR2X1 NOR2X1_755 ( .A(u2__abc_52138_new_n5975_), .B(u2__abc_52138_new_n5977_), .Y(u2__abc_52138_new_n5978_));
NOR2X1 NOR2X1_756 ( .A(u2_remHi_441_), .B(u2__abc_52138_new_n5979_), .Y(u2__abc_52138_new_n5980_));
NOR2X1 NOR2X1_757 ( .A(u2_o_441_), .B(u2__abc_52138_new_n5981_), .Y(u2__abc_52138_new_n5982_));
NOR2X1 NOR2X1_758 ( .A(u2__abc_52138_new_n5980_), .B(u2__abc_52138_new_n5982_), .Y(u2__abc_52138_new_n5983_));
NOR2X1 NOR2X1_759 ( .A(u2__abc_52138_new_n5973_), .B(u2__abc_52138_new_n5984_), .Y(u2__abc_52138_new_n5985_));
NOR2X1 NOR2X1_76 ( .A(\a[19] ), .B(\a[16] ), .Y(u1__abc_51895_new_n333_));
NOR2X1 NOR2X1_760 ( .A(u2_o_436_), .B(u2__abc_52138_new_n5987_), .Y(u2__abc_52138_new_n5988_));
NOR2X1 NOR2X1_761 ( .A(u2_remHi_436_), .B(u2__abc_52138_new_n5989_), .Y(u2__abc_52138_new_n5990_));
NOR2X1 NOR2X1_762 ( .A(u2__abc_52138_new_n5988_), .B(u2__abc_52138_new_n5990_), .Y(u2__abc_52138_new_n5991_));
NOR2X1 NOR2X1_763 ( .A(u2_o_437_), .B(u2__abc_52138_new_n5992_), .Y(u2__abc_52138_new_n5993_));
NOR2X1 NOR2X1_764 ( .A(u2_remHi_437_), .B(u2__abc_52138_new_n5994_), .Y(u2__abc_52138_new_n5995_));
NOR2X1 NOR2X1_765 ( .A(u2__abc_52138_new_n5993_), .B(u2__abc_52138_new_n5995_), .Y(u2__abc_52138_new_n5996_));
NOR2X1 NOR2X1_766 ( .A(u2_remHi_435_), .B(u2__abc_52138_new_n5998_), .Y(u2__abc_52138_new_n5999_));
NOR2X1 NOR2X1_767 ( .A(u2_o_435_), .B(u2__abc_52138_new_n6000_), .Y(u2__abc_52138_new_n6001_));
NOR2X1 NOR2X1_768 ( .A(u2__abc_52138_new_n5999_), .B(u2__abc_52138_new_n6001_), .Y(u2__abc_52138_new_n6002_));
NOR2X1 NOR2X1_769 ( .A(u2_o_434_), .B(u2__abc_52138_new_n6003_), .Y(u2__abc_52138_new_n6004_));
NOR2X1 NOR2X1_77 ( .A(\a[22] ), .B(\a[21] ), .Y(u1__abc_51895_new_n334_));
NOR2X1 NOR2X1_770 ( .A(u2_remHi_434_), .B(u2__abc_52138_new_n6005_), .Y(u2__abc_52138_new_n6006_));
NOR2X1 NOR2X1_771 ( .A(u2__abc_52138_new_n6004_), .B(u2__abc_52138_new_n6006_), .Y(u2__abc_52138_new_n6007_));
NOR2X1 NOR2X1_772 ( .A(u2__abc_52138_new_n5997_), .B(u2__abc_52138_new_n6008_), .Y(u2__abc_52138_new_n6009_));
NOR2X1 NOR2X1_773 ( .A(u2_o_430_), .B(u2__abc_52138_new_n6010_), .Y(u2__abc_52138_new_n6011_));
NOR2X1 NOR2X1_774 ( .A(u2_remHi_430_), .B(u2__abc_52138_new_n6012_), .Y(u2__abc_52138_new_n6013_));
NOR2X1 NOR2X1_775 ( .A(u2__abc_52138_new_n6011_), .B(u2__abc_52138_new_n6013_), .Y(u2__abc_52138_new_n6014_));
NOR2X1 NOR2X1_776 ( .A(u2_remHi_431_), .B(u2__abc_52138_new_n6015_), .Y(u2__abc_52138_new_n6016_));
NOR2X1 NOR2X1_777 ( .A(u2_o_431_), .B(u2__abc_52138_new_n6017_), .Y(u2__abc_52138_new_n6018_));
NOR2X1 NOR2X1_778 ( .A(u2__abc_52138_new_n6016_), .B(u2__abc_52138_new_n6018_), .Y(u2__abc_52138_new_n6019_));
NOR2X1 NOR2X1_779 ( .A(u2_o_432_), .B(u2__abc_52138_new_n6021_), .Y(u2__abc_52138_new_n6022_));
NOR2X1 NOR2X1_78 ( .A(u1__abc_51895_new_n332_), .B(u1__abc_51895_new_n335_), .Y(u1__abc_51895_new_n336_));
NOR2X1 NOR2X1_780 ( .A(u2_remHi_432_), .B(u2__abc_52138_new_n6023_), .Y(u2__abc_52138_new_n6024_));
NOR2X1 NOR2X1_781 ( .A(u2__abc_52138_new_n6022_), .B(u2__abc_52138_new_n6024_), .Y(u2__abc_52138_new_n6025_));
NOR2X1 NOR2X1_782 ( .A(u2_remHi_433_), .B(u2__abc_52138_new_n6026_), .Y(u2__abc_52138_new_n6027_));
NOR2X1 NOR2X1_783 ( .A(u2_o_433_), .B(u2__abc_52138_new_n6028_), .Y(u2__abc_52138_new_n6029_));
NOR2X1 NOR2X1_784 ( .A(u2__abc_52138_new_n6027_), .B(u2__abc_52138_new_n6029_), .Y(u2__abc_52138_new_n6030_));
NOR2X1 NOR2X1_785 ( .A(u2__abc_52138_new_n6020_), .B(u2__abc_52138_new_n6031_), .Y(u2__abc_52138_new_n6032_));
NOR2X1 NOR2X1_786 ( .A(u2__abc_52138_new_n5986_), .B(u2__abc_52138_new_n6033_), .Y(u2__abc_52138_new_n6034_));
NOR2X1 NOR2X1_787 ( .A(u2__abc_52138_new_n6040_), .B(u2__abc_52138_new_n6045_), .Y(u2__abc_52138_new_n6046_));
NOR2X1 NOR2X1_788 ( .A(u2_o_422_), .B(u2__abc_52138_new_n6047_), .Y(u2__abc_52138_new_n6048_));
NOR2X1 NOR2X1_789 ( .A(u2_remHi_422_), .B(u2__abc_52138_new_n6049_), .Y(u2__abc_52138_new_n6050_));
NOR2X1 NOR2X1_79 ( .A(\a[43] ), .B(\a[40] ), .Y(u1__abc_51895_new_n337_));
NOR2X1 NOR2X1_790 ( .A(u2__abc_52138_new_n6048_), .B(u2__abc_52138_new_n6050_), .Y(u2__abc_52138_new_n6051_));
NOR2X1 NOR2X1_791 ( .A(u2_remHi_423_), .B(u2__abc_52138_new_n6052_), .Y(u2__abc_52138_new_n6053_));
NOR2X1 NOR2X1_792 ( .A(u2_o_423_), .B(u2__abc_52138_new_n6054_), .Y(u2__abc_52138_new_n6055_));
NOR2X1 NOR2X1_793 ( .A(u2__abc_52138_new_n6053_), .B(u2__abc_52138_new_n6055_), .Y(u2__abc_52138_new_n6056_));
NOR2X1 NOR2X1_794 ( .A(u2__abc_52138_new_n6062_), .B(u2__abc_52138_new_n6067_), .Y(u2__abc_52138_new_n6068_));
NOR2X1 NOR2X1_795 ( .A(u2_remHi_427_), .B(u2__abc_52138_new_n6070_), .Y(u2__abc_52138_new_n6071_));
NOR2X1 NOR2X1_796 ( .A(u2_o_427_), .B(u2__abc_52138_new_n6072_), .Y(u2__abc_52138_new_n6073_));
NOR2X1 NOR2X1_797 ( .A(u2__abc_52138_new_n6071_), .B(u2__abc_52138_new_n6073_), .Y(u2__abc_52138_new_n6074_));
NOR2X1 NOR2X1_798 ( .A(u2_o_426_), .B(u2__abc_52138_new_n6075_), .Y(u2__abc_52138_new_n6076_));
NOR2X1 NOR2X1_799 ( .A(u2_remHi_426_), .B(u2__abc_52138_new_n6077_), .Y(u2__abc_52138_new_n6078_));
NOR2X1 NOR2X1_8 ( .A(_abc_65734_new_n1481_), .B(_abc_65734_new_n1472_), .Y(_abc_65734_new_n1482_));
NOR2X1 NOR2X1_80 ( .A(\a[46] ), .B(\a[45] ), .Y(u1__abc_51895_new_n338_));
NOR2X1 NOR2X1_800 ( .A(u2__abc_52138_new_n6076_), .B(u2__abc_52138_new_n6078_), .Y(u2__abc_52138_new_n6079_));
NOR2X1 NOR2X1_801 ( .A(u2__abc_52138_new_n6080_), .B(u2__abc_52138_new_n6069_), .Y(u2__abc_52138_new_n6081_));
NOR2X1 NOR2X1_802 ( .A(u2__abc_52138_new_n6057_), .B(u2__abc_52138_new_n6082_), .Y(u2__abc_52138_new_n6083_));
NOR2X1 NOR2X1_803 ( .A(u2__abc_52138_new_n6088_), .B(u2__abc_52138_new_n6093_), .Y(u2__abc_52138_new_n6094_));
NOR2X1 NOR2X1_804 ( .A(u2_remHi_419_), .B(u2__abc_52138_new_n6096_), .Y(u2__abc_52138_new_n6097_));
NOR2X1 NOR2X1_805 ( .A(u2_o_419_), .B(u2__abc_52138_new_n6098_), .Y(u2__abc_52138_new_n6099_));
NOR2X1 NOR2X1_806 ( .A(u2__abc_52138_new_n6097_), .B(u2__abc_52138_new_n6099_), .Y(u2__abc_52138_new_n6100_));
NOR2X1 NOR2X1_807 ( .A(u2_o_418_), .B(u2__abc_52138_new_n6101_), .Y(u2__abc_52138_new_n6102_));
NOR2X1 NOR2X1_808 ( .A(u2_remHi_418_), .B(u2__abc_52138_new_n6103_), .Y(u2__abc_52138_new_n6104_));
NOR2X1 NOR2X1_809 ( .A(u2__abc_52138_new_n6102_), .B(u2__abc_52138_new_n6104_), .Y(u2__abc_52138_new_n6105_));
NOR2X1 NOR2X1_81 ( .A(\a[34] ), .B(\a[33] ), .Y(u1__abc_51895_new_n340_));
NOR2X1 NOR2X1_810 ( .A(u2__abc_52138_new_n6106_), .B(u2__abc_52138_new_n6095_), .Y(u2__abc_52138_new_n6107_));
NOR2X1 NOR2X1_811 ( .A(u2__abc_52138_new_n6112_), .B(u2__abc_52138_new_n6117_), .Y(u2__abc_52138_new_n6118_));
NOR2X1 NOR2X1_812 ( .A(u2_remHi_415_), .B(u2__abc_52138_new_n6120_), .Y(u2__abc_52138_new_n6121_));
NOR2X1 NOR2X1_813 ( .A(u2_o_415_), .B(u2__abc_52138_new_n6122_), .Y(u2__abc_52138_new_n6123_));
NOR2X1 NOR2X1_814 ( .A(u2__abc_52138_new_n6121_), .B(u2__abc_52138_new_n6123_), .Y(u2__abc_52138_new_n6124_));
NOR2X1 NOR2X1_815 ( .A(u2_o_414_), .B(u2__abc_52138_new_n6125_), .Y(u2__abc_52138_new_n6126_));
NOR2X1 NOR2X1_816 ( .A(u2_remHi_414_), .B(u2__abc_52138_new_n6127_), .Y(u2__abc_52138_new_n6128_));
NOR2X1 NOR2X1_817 ( .A(u2__abc_52138_new_n6126_), .B(u2__abc_52138_new_n6128_), .Y(u2__abc_52138_new_n6129_));
NOR2X1 NOR2X1_818 ( .A(u2__abc_52138_new_n6130_), .B(u2__abc_52138_new_n6119_), .Y(u2__abc_52138_new_n6131_));
NOR2X1 NOR2X1_819 ( .A(u2__abc_52138_new_n6035_), .B(u2__abc_52138_new_n6134_), .Y(u2__abc_52138_new_n6135_));
NOR2X1 NOR2X1_82 ( .A(\a[39] ), .B(\a[36] ), .Y(u1__abc_51895_new_n341_));
NOR2X1 NOR2X1_820 ( .A(u2_o_388_), .B(u2__abc_52138_new_n6136_), .Y(u2__abc_52138_new_n6137_));
NOR2X1 NOR2X1_821 ( .A(u2_remHi_388_), .B(u2__abc_52138_new_n6138_), .Y(u2__abc_52138_new_n6139_));
NOR2X1 NOR2X1_822 ( .A(u2__abc_52138_new_n6137_), .B(u2__abc_52138_new_n6139_), .Y(u2__abc_52138_new_n6140_));
NOR2X1 NOR2X1_823 ( .A(u2_o_389_), .B(u2__abc_52138_new_n6141_), .Y(u2__abc_52138_new_n6142_));
NOR2X1 NOR2X1_824 ( .A(u2_remHi_389_), .B(u2__abc_52138_new_n6143_), .Y(u2__abc_52138_new_n6144_));
NOR2X1 NOR2X1_825 ( .A(u2__abc_52138_new_n6142_), .B(u2__abc_52138_new_n6144_), .Y(u2__abc_52138_new_n6145_));
NOR2X1 NOR2X1_826 ( .A(u2_remHi_387_), .B(u2__abc_52138_new_n6147_), .Y(u2__abc_52138_new_n6148_));
NOR2X1 NOR2X1_827 ( .A(u2_o_387_), .B(u2__abc_52138_new_n6149_), .Y(u2__abc_52138_new_n6150_));
NOR2X1 NOR2X1_828 ( .A(u2__abc_52138_new_n6148_), .B(u2__abc_52138_new_n6150_), .Y(u2__abc_52138_new_n6151_));
NOR2X1 NOR2X1_829 ( .A(u2_o_386_), .B(u2__abc_52138_new_n6152_), .Y(u2__abc_52138_new_n6153_));
NOR2X1 NOR2X1_83 ( .A(u1__abc_51895_new_n339_), .B(u1__abc_51895_new_n342_), .Y(u1__abc_51895_new_n343_));
NOR2X1 NOR2X1_830 ( .A(u2_remHi_386_), .B(u2__abc_52138_new_n6154_), .Y(u2__abc_52138_new_n6155_));
NOR2X1 NOR2X1_831 ( .A(u2__abc_52138_new_n6153_), .B(u2__abc_52138_new_n6155_), .Y(u2__abc_52138_new_n6156_));
NOR2X1 NOR2X1_832 ( .A(u2__abc_52138_new_n6146_), .B(u2__abc_52138_new_n6157_), .Y(u2__abc_52138_new_n6158_));
NOR2X1 NOR2X1_833 ( .A(u2_o_384_), .B(u2__abc_52138_new_n6160_), .Y(u2__abc_52138_new_n6161_));
NOR2X1 NOR2X1_834 ( .A(u2_remHi_384_), .B(u2__abc_52138_new_n6162_), .Y(u2__abc_52138_new_n6163_));
NOR2X1 NOR2X1_835 ( .A(u2__abc_52138_new_n6161_), .B(u2__abc_52138_new_n6163_), .Y(u2__abc_52138_new_n6164_));
NOR2X1 NOR2X1_836 ( .A(u2_remHi_385_), .B(u2__abc_52138_new_n6165_), .Y(u2__abc_52138_new_n6166_));
NOR2X1 NOR2X1_837 ( .A(u2_o_385_), .B(u2__abc_52138_new_n6167_), .Y(u2__abc_52138_new_n6168_));
NOR2X1 NOR2X1_838 ( .A(u2__abc_52138_new_n6166_), .B(u2__abc_52138_new_n6168_), .Y(u2__abc_52138_new_n6169_));
NOR2X1 NOR2X1_839 ( .A(u2_remHi_383_), .B(u2__abc_52138_new_n6171_), .Y(u2__abc_52138_new_n6172_));
NOR2X1 NOR2X1_84 ( .A(\a[90] ), .B(\a[89] ), .Y(u1__abc_51895_new_n345_));
NOR2X1 NOR2X1_840 ( .A(u2_o_383_), .B(u2__abc_52138_new_n6173_), .Y(u2__abc_52138_new_n6174_));
NOR2X1 NOR2X1_841 ( .A(u2__abc_52138_new_n6172_), .B(u2__abc_52138_new_n6174_), .Y(u2__abc_52138_new_n6175_));
NOR2X1 NOR2X1_842 ( .A(u2_o_382_), .B(u2__abc_52138_new_n6176_), .Y(u2__abc_52138_new_n6177_));
NOR2X1 NOR2X1_843 ( .A(u2_remHi_382_), .B(u2__abc_52138_new_n6178_), .Y(u2__abc_52138_new_n6179_));
NOR2X1 NOR2X1_844 ( .A(u2__abc_52138_new_n6177_), .B(u2__abc_52138_new_n6179_), .Y(u2__abc_52138_new_n6180_));
NOR2X1 NOR2X1_845 ( .A(u2__abc_52138_new_n6170_), .B(u2__abc_52138_new_n6181_), .Y(u2__abc_52138_new_n6182_));
NOR2X1 NOR2X1_846 ( .A(u2__abc_52138_new_n6159_), .B(u2__abc_52138_new_n6183_), .Y(u2__abc_52138_new_n6184_));
NOR2X1 NOR2X1_847 ( .A(u2_o_408_), .B(u2__abc_52138_new_n6185_), .Y(u2__abc_52138_new_n6186_));
NOR2X1 NOR2X1_848 ( .A(u2_remHi_408_), .B(u2__abc_52138_new_n6187_), .Y(u2__abc_52138_new_n6188_));
NOR2X1 NOR2X1_849 ( .A(u2__abc_52138_new_n6186_), .B(u2__abc_52138_new_n6188_), .Y(u2__abc_52138_new_n6189_));
NOR2X1 NOR2X1_85 ( .A(\a[95] ), .B(\a[92] ), .Y(u1__abc_51895_new_n346_));
NOR2X1 NOR2X1_850 ( .A(u2_remHi_409_), .B(u2__abc_52138_new_n6190_), .Y(u2__abc_52138_new_n6191_));
NOR2X1 NOR2X1_851 ( .A(u2_o_409_), .B(u2__abc_52138_new_n6192_), .Y(u2__abc_52138_new_n6193_));
NOR2X1 NOR2X1_852 ( .A(u2__abc_52138_new_n6191_), .B(u2__abc_52138_new_n6193_), .Y(u2__abc_52138_new_n6194_));
NOR2X1 NOR2X1_853 ( .A(u2_remHi_407_), .B(u2__abc_52138_new_n6196_), .Y(u2__abc_52138_new_n6197_));
NOR2X1 NOR2X1_854 ( .A(u2_o_407_), .B(u2__abc_52138_new_n6198_), .Y(u2__abc_52138_new_n6199_));
NOR2X1 NOR2X1_855 ( .A(u2__abc_52138_new_n6197_), .B(u2__abc_52138_new_n6199_), .Y(u2__abc_52138_new_n6200_));
NOR2X1 NOR2X1_856 ( .A(u2_o_406_), .B(u2__abc_52138_new_n6201_), .Y(u2__abc_52138_new_n6202_));
NOR2X1 NOR2X1_857 ( .A(u2_remHi_406_), .B(u2__abc_52138_new_n6203_), .Y(u2__abc_52138_new_n6204_));
NOR2X1 NOR2X1_858 ( .A(u2__abc_52138_new_n6202_), .B(u2__abc_52138_new_n6204_), .Y(u2__abc_52138_new_n6205_));
NOR2X1 NOR2X1_859 ( .A(u2__abc_52138_new_n6195_), .B(u2__abc_52138_new_n6206_), .Y(u2__abc_52138_new_n6207_));
NOR2X1 NOR2X1_86 ( .A(\a[83] ), .B(\a[80] ), .Y(u1__abc_51895_new_n348_));
NOR2X1 NOR2X1_860 ( .A(u2_o_412_), .B(u2__abc_52138_new_n6208_), .Y(u2__abc_52138_new_n6209_));
NOR2X1 NOR2X1_861 ( .A(u2_remHi_412_), .B(u2__abc_52138_new_n6210_), .Y(u2__abc_52138_new_n6211_));
NOR2X1 NOR2X1_862 ( .A(u2__abc_52138_new_n6209_), .B(u2__abc_52138_new_n6211_), .Y(u2__abc_52138_new_n6212_));
NOR2X1 NOR2X1_863 ( .A(u2_o_413_), .B(u2__abc_52138_new_n6213_), .Y(u2__abc_52138_new_n6214_));
NOR2X1 NOR2X1_864 ( .A(u2_remHi_413_), .B(u2__abc_52138_new_n6215_), .Y(u2__abc_52138_new_n6216_));
NOR2X1 NOR2X1_865 ( .A(u2__abc_52138_new_n6214_), .B(u2__abc_52138_new_n6216_), .Y(u2__abc_52138_new_n6217_));
NOR2X1 NOR2X1_866 ( .A(u2_remHi_411_), .B(u2__abc_52138_new_n6219_), .Y(u2__abc_52138_new_n6220_));
NOR2X1 NOR2X1_867 ( .A(u2_o_411_), .B(u2__abc_52138_new_n6221_), .Y(u2__abc_52138_new_n6222_));
NOR2X1 NOR2X1_868 ( .A(u2__abc_52138_new_n6220_), .B(u2__abc_52138_new_n6222_), .Y(u2__abc_52138_new_n6223_));
NOR2X1 NOR2X1_869 ( .A(u2_o_410_), .B(u2__abc_52138_new_n6224_), .Y(u2__abc_52138_new_n6225_));
NOR2X1 NOR2X1_87 ( .A(\a[86] ), .B(\a[85] ), .Y(u1__abc_51895_new_n349_));
NOR2X1 NOR2X1_870 ( .A(u2_remHi_410_), .B(u2__abc_52138_new_n6226_), .Y(u2__abc_52138_new_n6227_));
NOR2X1 NOR2X1_871 ( .A(u2__abc_52138_new_n6225_), .B(u2__abc_52138_new_n6227_), .Y(u2__abc_52138_new_n6228_));
NOR2X1 NOR2X1_872 ( .A(u2__abc_52138_new_n6218_), .B(u2__abc_52138_new_n6229_), .Y(u2__abc_52138_new_n6230_));
NOR2X1 NOR2X1_873 ( .A(u2_o_398_), .B(u2__abc_52138_new_n6232_), .Y(u2__abc_52138_new_n6233_));
NOR2X1 NOR2X1_874 ( .A(u2_remHi_398_), .B(u2__abc_52138_new_n6234_), .Y(u2__abc_52138_new_n6235_));
NOR2X1 NOR2X1_875 ( .A(u2__abc_52138_new_n6233_), .B(u2__abc_52138_new_n6235_), .Y(u2__abc_52138_new_n6236_));
NOR2X1 NOR2X1_876 ( .A(u2_remHi_399_), .B(u2__abc_52138_new_n6237_), .Y(u2__abc_52138_new_n6238_));
NOR2X1 NOR2X1_877 ( .A(u2_o_399_), .B(u2__abc_52138_new_n6239_), .Y(u2__abc_52138_new_n6240_));
NOR2X1 NOR2X1_878 ( .A(u2__abc_52138_new_n6238_), .B(u2__abc_52138_new_n6240_), .Y(u2__abc_52138_new_n6241_));
NOR2X1 NOR2X1_879 ( .A(u2_o_400_), .B(u2__abc_52138_new_n6243_), .Y(u2__abc_52138_new_n6244_));
NOR2X1 NOR2X1_88 ( .A(u1__abc_51895_new_n347_), .B(u1__abc_51895_new_n350_), .Y(u1__abc_51895_new_n351_));
NOR2X1 NOR2X1_880 ( .A(u2_remHi_400_), .B(u2__abc_52138_new_n6245_), .Y(u2__abc_52138_new_n6246_));
NOR2X1 NOR2X1_881 ( .A(u2__abc_52138_new_n6244_), .B(u2__abc_52138_new_n6246_), .Y(u2__abc_52138_new_n6247_));
NOR2X1 NOR2X1_882 ( .A(u2_remHi_401_), .B(u2__abc_52138_new_n6248_), .Y(u2__abc_52138_new_n6249_));
NOR2X1 NOR2X1_883 ( .A(u2_o_401_), .B(u2__abc_52138_new_n6250_), .Y(u2__abc_52138_new_n6251_));
NOR2X1 NOR2X1_884 ( .A(u2__abc_52138_new_n6249_), .B(u2__abc_52138_new_n6251_), .Y(u2__abc_52138_new_n6252_));
NOR2X1 NOR2X1_885 ( .A(u2__abc_52138_new_n6242_), .B(u2__abc_52138_new_n6253_), .Y(u2__abc_52138_new_n6254_));
NOR2X1 NOR2X1_886 ( .A(u2_o_404_), .B(u2__abc_52138_new_n6255_), .Y(u2__abc_52138_new_n6256_));
NOR2X1 NOR2X1_887 ( .A(u2_remHi_404_), .B(u2__abc_52138_new_n6257_), .Y(u2__abc_52138_new_n6258_));
NOR2X1 NOR2X1_888 ( .A(u2__abc_52138_new_n6256_), .B(u2__abc_52138_new_n6258_), .Y(u2__abc_52138_new_n6259_));
NOR2X1 NOR2X1_889 ( .A(u2_o_405_), .B(u2__abc_52138_new_n6260_), .Y(u2__abc_52138_new_n6261_));
NOR2X1 NOR2X1_89 ( .A(\a[107] ), .B(\a[104] ), .Y(u1__abc_51895_new_n352_));
NOR2X1 NOR2X1_890 ( .A(u2_remHi_405_), .B(u2__abc_52138_new_n6262_), .Y(u2__abc_52138_new_n6263_));
NOR2X1 NOR2X1_891 ( .A(u2__abc_52138_new_n6261_), .B(u2__abc_52138_new_n6263_), .Y(u2__abc_52138_new_n6264_));
NOR2X1 NOR2X1_892 ( .A(u2_remHi_403_), .B(u2__abc_52138_new_n6266_), .Y(u2__abc_52138_new_n6267_));
NOR2X1 NOR2X1_893 ( .A(u2_o_403_), .B(u2__abc_52138_new_n6268_), .Y(u2__abc_52138_new_n6269_));
NOR2X1 NOR2X1_894 ( .A(u2__abc_52138_new_n6267_), .B(u2__abc_52138_new_n6269_), .Y(u2__abc_52138_new_n6270_));
NOR2X1 NOR2X1_895 ( .A(u2_o_402_), .B(u2__abc_52138_new_n6271_), .Y(u2__abc_52138_new_n6272_));
NOR2X1 NOR2X1_896 ( .A(u2_remHi_402_), .B(u2__abc_52138_new_n6273_), .Y(u2__abc_52138_new_n6274_));
NOR2X1 NOR2X1_897 ( .A(u2__abc_52138_new_n6272_), .B(u2__abc_52138_new_n6274_), .Y(u2__abc_52138_new_n6275_));
NOR2X1 NOR2X1_898 ( .A(u2__abc_52138_new_n6265_), .B(u2__abc_52138_new_n6276_), .Y(u2__abc_52138_new_n6277_));
NOR2X1 NOR2X1_899 ( .A(u2__abc_52138_new_n6231_), .B(u2__abc_52138_new_n6278_), .Y(u2__abc_52138_new_n6279_));
NOR2X1 NOR2X1_9 ( .A(_abc_65734_new_n1475_), .B(_abc_65734_new_n1488_), .Y(_abc_65734_new_n1489_));
NOR2X1 NOR2X1_90 ( .A(\a[110] ), .B(\a[109] ), .Y(u1__abc_51895_new_n353_));
NOR2X1 NOR2X1_900 ( .A(u2_o_392_), .B(u2__abc_52138_new_n6280_), .Y(u2__abc_52138_new_n6281_));
NOR2X1 NOR2X1_901 ( .A(u2_remHi_392_), .B(u2__abc_52138_new_n6282_), .Y(u2__abc_52138_new_n6283_));
NOR2X1 NOR2X1_902 ( .A(u2__abc_52138_new_n6281_), .B(u2__abc_52138_new_n6283_), .Y(u2__abc_52138_new_n6284_));
NOR2X1 NOR2X1_903 ( .A(u2_remHi_393_), .B(u2__abc_52138_new_n6285_), .Y(u2__abc_52138_new_n6286_));
NOR2X1 NOR2X1_904 ( .A(u2_o_390_), .B(u2__abc_52138_new_n6292_), .Y(u2__abc_52138_new_n6293_));
NOR2X1 NOR2X1_905 ( .A(u2__abc_52138_new_n6293_), .B(u2__abc_52138_new_n6295_), .Y(u2__abc_52138_new_n6296_));
NOR2X1 NOR2X1_906 ( .A(u2_o_391_), .B(u2__abc_52138_new_n6297_), .Y(u2__abc_52138_new_n6300_));
NOR2X1 NOR2X1_907 ( .A(u2__abc_52138_new_n6300_), .B(u2__abc_52138_new_n6299_), .Y(u2__abc_52138_new_n6301_));
NOR2X1 NOR2X1_908 ( .A(u2__abc_52138_new_n6302_), .B(u2__abc_52138_new_n6291_), .Y(u2__abc_52138_new_n6303_));
NOR2X1 NOR2X1_909 ( .A(u2_o_396_), .B(u2__abc_52138_new_n6304_), .Y(u2__abc_52138_new_n6305_));
NOR2X1 NOR2X1_91 ( .A(\a[98] ), .B(\a[97] ), .Y(u1__abc_51895_new_n355_));
NOR2X1 NOR2X1_910 ( .A(u2_remHi_396_), .B(u2__abc_52138_new_n6306_), .Y(u2__abc_52138_new_n6307_));
NOR2X1 NOR2X1_911 ( .A(u2__abc_52138_new_n6305_), .B(u2__abc_52138_new_n6307_), .Y(u2__abc_52138_new_n6308_));
NOR2X1 NOR2X1_912 ( .A(u2_o_397_), .B(u2__abc_52138_new_n6309_), .Y(u2__abc_52138_new_n6310_));
NOR2X1 NOR2X1_913 ( .A(u2_remHi_397_), .B(u2__abc_52138_new_n6311_), .Y(u2__abc_52138_new_n6312_));
NOR2X1 NOR2X1_914 ( .A(u2__abc_52138_new_n6310_), .B(u2__abc_52138_new_n6312_), .Y(u2__abc_52138_new_n6313_));
NOR2X1 NOR2X1_915 ( .A(u2_remHi_395_), .B(u2__abc_52138_new_n6315_), .Y(u2__abc_52138_new_n6316_));
NOR2X1 NOR2X1_916 ( .A(u2_o_395_), .B(u2__abc_52138_new_n6317_), .Y(u2__abc_52138_new_n6318_));
NOR2X1 NOR2X1_917 ( .A(u2__abc_52138_new_n6316_), .B(u2__abc_52138_new_n6318_), .Y(u2__abc_52138_new_n6319_));
NOR2X1 NOR2X1_918 ( .A(u2_o_394_), .B(u2__abc_52138_new_n6320_), .Y(u2__abc_52138_new_n6321_));
NOR2X1 NOR2X1_919 ( .A(u2__abc_52138_new_n6314_), .B(u2__abc_52138_new_n6325_), .Y(u2__abc_52138_new_n6326_));
NOR2X1 NOR2X1_92 ( .A(\a[103] ), .B(\a[100] ), .Y(u1__abc_51895_new_n356_));
NOR2X1 NOR2X1_920 ( .A(u2__abc_52138_new_n6343_), .B(u2__abc_52138_new_n6327_), .Y(u2__abc_52138_new_n6344_));
NOR2X1 NOR2X1_921 ( .A(u2__abc_52138_new_n6231_), .B(u2__abc_52138_new_n6383_), .Y(u2__abc_52138_new_n6384_));
NOR2X1 NOR2X1_922 ( .A(u2__abc_52138_new_n6372_), .B(u2__abc_52138_new_n6384_), .Y(u2__abc_52138_new_n6385_));
NOR2X1 NOR2X1_923 ( .A(u2__abc_52138_new_n6402_), .B(u2__abc_52138_new_n6400_), .Y(u2__abc_52138_new_n6403_));
NOR2X1 NOR2X1_924 ( .A(u2__abc_52138_new_n5986_), .B(u2__abc_52138_new_n6436_), .Y(u2__abc_52138_new_n6437_));
NOR2X1 NOR2X1_925 ( .A(u2__abc_52138_new_n6437_), .B(u2__abc_52138_new_n6426_), .Y(u2__abc_52138_new_n6438_));
NOR2X1 NOR2X1_926 ( .A(u2__abc_52138_new_n6439_), .B(u2__abc_52138_new_n6386_), .Y(u2__abc_52138_new_n6440_));
NOR2X1 NOR2X1_927 ( .A(u2__abc_52138_new_n3006_), .B(u2__abc_52138_new_n3011_), .Y(u2__abc_52138_new_n6443_));
NOR2X1 NOR2X1_928 ( .A(u2__abc_52138_new_n6443_), .B(u2__abc_52138_new_n6444_), .Y(u2__abc_52138_new_n6445_));
NOR2X1 NOR2X1_929 ( .A(u2__abc_52138_new_n6449_), .B(u2__abc_52138_new_n6445_), .Y(u2__abc_52138_new_n6450_));
NOR2X1 NOR2X1_93 ( .A(u1__abc_51895_new_n354_), .B(u1__abc_51895_new_n357_), .Y(u1__abc_51895_new_n358_));
NOR2X1 NOR2X1_930 ( .A(u2_remHiShift_1_), .B(u2__abc_52138_new_n3069_), .Y(u2__abc_52138_new_n6454_));
NOR2X1 NOR2X1_931 ( .A(u2__abc_52138_new_n6454_), .B(u2__abc_52138_new_n3071_), .Y(u2__abc_52138_new_n6455_));
NOR2X1 NOR2X1_932 ( .A(u2__abc_52138_new_n3068_), .B(u2__abc_52138_new_n6456_), .Y(u2__abc_52138_new_n6457_));
NOR2X1 NOR2X1_933 ( .A(u2__abc_52138_new_n6460_), .B(u2__abc_52138_new_n6461_), .Y(u2__abc_52138_new_n6462_));
NOR2X1 NOR2X1_934 ( .A(u2__abc_52138_new_n6463_), .B(u2__abc_52138_new_n6464_), .Y(u2__abc_52138_new_n6465_));
NOR2X1 NOR2X1_935 ( .A(u2__abc_52138_new_n6466_), .B(u2__abc_52138_new_n6467_), .Y(u2__abc_52138_new_n6468_));
NOR2X1 NOR2X1_936 ( .A(u2__abc_52138_new_n6453_), .B(u2__abc_52138_new_n6469_), .Y(u2__abc_52138_new_n6470_));
NOR2X1 NOR2X1_937 ( .A(u2__abc_52138_new_n6471_), .B(u2__abc_52138_new_n6452_), .Y(u2__abc_52138_new_n6472_));
NOR2X1 NOR2X1_938 ( .A(u2__abc_52138_new_n5365_), .B(u2__abc_52138_new_n5639_), .Y(u2__abc_52138_new_n6473_));
NOR2X1 NOR2X1_939 ( .A(u2__abc_52138_new_n6474_), .B(u2__abc_52138_new_n6477_), .Y(u2__abc_52138_new_n6478_));
NOR2X1 NOR2X1_94 ( .A(\a[59] ), .B(\a[56] ), .Y(u1__abc_51895_new_n360_));
NOR2X1 NOR2X1_940 ( .A(u2__abc_52138_new_n5733_), .B(u2__abc_52138_new_n6480_), .Y(u2__abc_52138_new_n6481_));
NOR2X1 NOR2X1_941 ( .A(u2__abc_52138_new_n3784_), .B(u2__abc_52138_new_n4049_), .Y(u2__abc_52138_new_n6485_));
NOR2X1 NOR2X1_942 ( .A(u2__abc_52138_new_n6487_), .B(u2__abc_52138_new_n6488_), .Y(u2__abc_52138_new_n6489_));
NOR2X1 NOR2X1_943 ( .A(u2__abc_52138_new_n3052_), .B(u2__abc_52138_new_n3427_), .Y(u2__abc_52138_new_n6490_));
NOR2X1 NOR2X1_944 ( .A(u2__abc_52138_new_n6491_), .B(u2__abc_52138_new_n6486_), .Y(u2__abc_52138_new_n6492_));
NOR2X1 NOR2X1_945 ( .A(u2__abc_52138_new_n4240_), .B(u2__abc_52138_new_n4097_), .Y(u2__abc_52138_new_n6493_));
NOR2X1 NOR2X1_946 ( .A(u2__abc_52138_new_n4287_), .B(u2__abc_52138_new_n4330_), .Y(u2__abc_52138_new_n6494_));
NOR2X1 NOR2X1_947 ( .A(u2__abc_52138_new_n6496_), .B(u2__abc_52138_new_n6482_), .Y(u2__abc_52138_new_n6497_));
NOR2X1 NOR2X1_948 ( .A(u2__abc_52138_new_n2996_), .B(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6500_));
NOR2X1 NOR2X1_949 ( .A(u2__abc_52138_new_n6503_), .B(u2__abc_52138_new_n2966_), .Y(u2__abc_52138_new_n6504_));
NOR2X1 NOR2X1_95 ( .A(\a[62] ), .B(\a[61] ), .Y(u1__abc_51895_new_n361_));
NOR2X1 NOR2X1_950 ( .A(u2__abc_52138_new_n6466_), .B(u2__abc_52138_new_n6550_), .Y(u2__abc_52138_new_n6576_));
NOR2X1 NOR2X1_951 ( .A(u2__abc_52138_new_n6581_), .B(u2__abc_52138_new_n6576_), .Y(u2__abc_52138_new_n6582_));
NOR2X1 NOR2X1_952 ( .A(u2__abc_52138_new_n6592_), .B(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n6593_));
NOR2X1 NOR2X1_953 ( .A(u2__abc_52138_new_n6599_), .B(u2__abc_52138_new_n6604_), .Y(u2__abc_52138_new_n6606_));
NOR2X1 NOR2X1_954 ( .A(u2__abc_52138_new_n6636_), .B(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n6637_));
NOR2X1 NOR2X1_955 ( .A(u2__abc_52138_new_n6667_), .B(u2__abc_52138_new_n6653_), .Y(u2__abc_52138_new_n6668_));
NOR2X1 NOR2X1_956 ( .A(u2__abc_52138_new_n6684_), .B(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n6685_));
NOR2X1 NOR2X1_957 ( .A(u2__abc_52138_new_n3193_), .B(u2__abc_52138_new_n6716_), .Y(u2__abc_52138_new_n6736_));
NOR2X1 NOR2X1_958 ( .A(u2__abc_52138_new_n6737_), .B(u2__abc_52138_new_n6736_), .Y(u2__abc_52138_new_n6738_));
NOR2X1 NOR2X1_959 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6749_), .Y(u2__abc_52138_new_n6750_));
NOR2X1 NOR2X1_96 ( .A(\a[50] ), .B(\a[49] ), .Y(u1__abc_51895_new_n363_));
NOR2X1 NOR2X1_960 ( .A(u2__abc_52138_new_n3195_), .B(u2__abc_52138_new_n6674_), .Y(u2__abc_52138_new_n6756_));
NOR2X1 NOR2X1_961 ( .A(u2__abc_52138_new_n6735_), .B(u2__abc_52138_new_n6747_), .Y(u2__abc_52138_new_n6758_));
NOR2X1 NOR2X1_962 ( .A(u2__abc_52138_new_n6762_), .B(u2__abc_52138_new_n6756_), .Y(u2__abc_52138_new_n6763_));
NOR2X1 NOR2X1_963 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6794_), .Y(u2__abc_52138_new_n6795_));
NOR2X1 NOR2X1_964 ( .A(u2__abc_52138_new_n3155_), .B(u2__abc_52138_new_n6806_), .Y(u2__abc_52138_new_n6808_));
NOR2X1 NOR2X1_965 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6817_), .Y(u2__abc_52138_new_n6818_));
NOR2X1 NOR2X1_966 ( .A(u2__abc_52138_new_n3233_), .B(u2__abc_52138_new_n3229_), .Y(u2__abc_52138_new_n6841_));
NOR2X1 NOR2X1_967 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6855_), .Y(u2__abc_52138_new_n6856_));
NOR2X1 NOR2X1_968 ( .A(u2__abc_52138_new_n3387_), .B(u2__abc_52138_new_n6872_), .Y(u2__abc_52138_new_n6873_));
NOR2X1 NOR2X1_969 ( .A(u2__abc_52138_new_n3417_), .B(u2__abc_52138_new_n6885_), .Y(u2__abc_52138_new_n6886_));
NOR2X1 NOR2X1_97 ( .A(\a[55] ), .B(\a[52] ), .Y(u1__abc_51895_new_n364_));
NOR2X1 NOR2X1_970 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6916_), .Y(u2__abc_52138_new_n6917_));
NOR2X1 NOR2X1_971 ( .A(u2__abc_52138_new_n6926_), .B(u2__abc_52138_new_n6924_), .Y(u2__abc_52138_new_n6927_));
NOR2X1 NOR2X1_972 ( .A(u2__abc_52138_new_n6923_), .B(u2__abc_52138_new_n6929_), .Y(u2__abc_52138_new_n6930_));
NOR2X1 NOR2X1_973 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6940_), .Y(u2__abc_52138_new_n6941_));
NOR2X1 NOR2X1_974 ( .A(u2_remHi_41_), .B(u2__abc_52138_new_n3340_), .Y(u2__abc_52138_new_n6956_));
NOR2X1 NOR2X1_975 ( .A(u2__abc_52138_new_n3456_), .B(u2__abc_52138_new_n6956_), .Y(u2__abc_52138_new_n6957_));
NOR2X1 NOR2X1_976 ( .A(u2__abc_52138_new_n3336_), .B(u2__abc_52138_new_n6956_), .Y(u2__abc_52138_new_n6968_));
NOR2X1 NOR2X1_977 ( .A(u2__abc_52138_new_n3456_), .B(u2__abc_52138_new_n6968_), .Y(u2__abc_52138_new_n6969_));
NOR2X1 NOR2X1_978 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6981_), .Y(u2__abc_52138_new_n6982_));
NOR2X1 NOR2X1_979 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6991_), .Y(u2__abc_52138_new_n6992_));
NOR2X1 NOR2X1_98 ( .A(u1__abc_51895_new_n362_), .B(u1__abc_51895_new_n365_), .Y(u1__abc_51895_new_n366_));
NOR2X1 NOR2X1_980 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7000_), .Y(u2__abc_52138_new_n7001_));
NOR2X1 NOR2X1_981 ( .A(u2__abc_52138_new_n3308_), .B(u2__abc_52138_new_n7012_), .Y(u2__abc_52138_new_n7013_));
NOR2X1 NOR2X1_982 ( .A(u2__abc_52138_new_n3307_), .B(u2__abc_52138_new_n7014_), .Y(u2__abc_52138_new_n7015_));
NOR2X1 NOR2X1_983 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7066_), .Y(u2__abc_52138_new_n7067_));
NOR2X1 NOR2X1_984 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7077_), .Y(u2__abc_52138_new_n7078_));
NOR2X1 NOR2X1_985 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7086_), .Y(u2__abc_52138_new_n7087_));
NOR2X1 NOR2X1_986 ( .A(u2__abc_52138_new_n3423_), .B(u2__abc_52138_new_n7014_), .Y(u2__abc_52138_new_n7099_));
NOR2X1 NOR2X1_987 ( .A(u2__abc_52138_new_n7098_), .B(u2__abc_52138_new_n7099_), .Y(u2__abc_52138_new_n7100_));
NOR2X1 NOR2X1_988 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7111_), .Y(u2__abc_52138_new_n7112_));
NOR2X1 NOR2X1_989 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7119_), .Y(u2__abc_52138_new_n7120_));
NOR2X1 NOR2X1_99 ( .A(\a[74] ), .B(\a[73] ), .Y(u1__abc_51895_new_n367_));
NOR2X1 NOR2X1_990 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7128_), .Y(u2__abc_52138_new_n7129_));
NOR2X1 NOR2X1_991 ( .A(u2__abc_52138_new_n7135_), .B(u2__abc_52138_new_n7139_), .Y(u2__abc_52138_new_n7142_));
NOR2X1 NOR2X1_992 ( .A(u2__abc_52138_new_n3494_), .B(u2__abc_52138_new_n7152_), .Y(u2__abc_52138_new_n7160_));
NOR2X1 NOR2X1_993 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7170_), .Y(u2__abc_52138_new_n7171_));
NOR2X1 NOR2X1_994 ( .A(u2__abc_52138_new_n3334_), .B(u2__abc_52138_new_n7011_), .Y(u2__abc_52138_new_n7183_));
NOR2X1 NOR2X1_995 ( .A(u2__abc_52138_new_n7182_), .B(u2__abc_52138_new_n7183_), .Y(u2__abc_52138_new_n7184_));
NOR2X1 NOR2X1_996 ( .A(u2__abc_52138_new_n7212_), .B(u2__abc_52138_new_n3878_), .Y(u2__abc_52138_new_n7213_));
NOR2X1 NOR2X1_997 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7236_), .Y(u2__abc_52138_new_n7237_));
NOR2X1 NOR2X1_998 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7255_), .Y(u2__abc_52138_new_n7256_));
NOR2X1 NOR2X1_999 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n7291_), .Y(u2__abc_52138_new_n7292_));
NOR3X1 NOR3X1_1 ( .A(_abc_65734_new_n1473_), .B(_abc_65734_new_n1461_), .C(_abc_65734_new_n1462_), .Y(_abc_65734_new_n1486_));
NOR3X1 NOR3X1_10 ( .A(u2__abc_52138_new_n4712_), .B(u2__abc_52138_new_n4665_), .C(u2__abc_52138_new_n4751_), .Y(u2__abc_52138_new_n4752_));
NOR3X1 NOR3X1_100 ( .A(u2__abc_52138_new_n3575_), .B(u2__abc_52138_new_n3583_), .C(u2__abc_52138_new_n13936_), .Y(u2__abc_52138_new_n13952_));
NOR3X1 NOR3X1_101 ( .A(u2__abc_52138_new_n3578_), .B(u2__abc_52138_new_n3575_), .C(u2__abc_52138_new_n13958_), .Y(u2__abc_52138_new_n13959_));
NOR3X1 NOR3X1_102 ( .A(u2__abc_52138_new_n3511_), .B(u2__abc_52138_new_n13962_), .C(u2__abc_52138_new_n13976_), .Y(u2__abc_52138_new_n13977_));
NOR3X1 NOR3X1_103 ( .A(u2__abc_52138_new_n3516_), .B(u2__abc_52138_new_n3511_), .C(u2__abc_52138_new_n13968_), .Y(u2__abc_52138_new_n13984_));
NOR3X1 NOR3X1_104 ( .A(u2__abc_52138_new_n3521_), .B(u2__abc_52138_new_n3516_), .C(u2__abc_52138_new_n13990_), .Y(u2__abc_52138_new_n13991_));
NOR3X1 NOR3X1_105 ( .A(u2__abc_52138_new_n3538_), .B(u2__abc_52138_new_n3544_), .C(u2__abc_52138_new_n14007_), .Y(u2__abc_52138_new_n14008_));
NOR3X1 NOR3X1_106 ( .A(u2__abc_52138_new_n3527_), .B(u2__abc_52138_new_n3538_), .C(u2__abc_52138_new_n13999_), .Y(u2__abc_52138_new_n14015_));
NOR3X1 NOR3X1_107 ( .A(u2__abc_52138_new_n3534_), .B(u2__abc_52138_new_n3527_), .C(u2__abc_52138_new_n14021_), .Y(u2__abc_52138_new_n14022_));
NOR3X1 NOR3X1_108 ( .A(u2__abc_52138_new_n4719_), .B(u2__abc_52138_new_n4713_), .C(u2__abc_52138_new_n14038_), .Y(u2__abc_52138_new_n14039_));
NOR3X1 NOR3X1_109 ( .A(u2__abc_52138_new_n4770_), .B(u2__abc_52138_new_n4719_), .C(u2__abc_52138_new_n14030_), .Y(u2__abc_52138_new_n14046_));
NOR3X1 NOR3X1_11 ( .A(u2__abc_52138_new_n3809_), .B(u2__abc_52138_new_n3811_), .C(u2__abc_52138_new_n7353_), .Y(u2__abc_52138_new_n7354_));
NOR3X1 NOR3X1_110 ( .A(u2__abc_52138_new_n4727_), .B(u2__abc_52138_new_n4770_), .C(u2__abc_52138_new_n14053_), .Y(u2__abc_52138_new_n14054_));
NOR3X1 NOR3X1_111 ( .A(u2__abc_52138_new_n4744_), .B(u2__abc_52138_new_n14056_), .C(u2__abc_52138_new_n14070_), .Y(u2__abc_52138_new_n14071_));
NOR3X1 NOR3X1_112 ( .A(u2__abc_52138_new_n4733_), .B(u2__abc_52138_new_n4744_), .C(u2__abc_52138_new_n14062_), .Y(u2__abc_52138_new_n14078_));
NOR3X1 NOR3X1_113 ( .A(u2__abc_52138_new_n4738_), .B(u2__abc_52138_new_n4733_), .C(u2__abc_52138_new_n14085_), .Y(u2__abc_52138_new_n14086_));
NOR3X1 NOR3X1_114 ( .A(u2__abc_52138_new_n4682_), .B(u2__abc_52138_new_n4677_), .C(u2__abc_52138_new_n14100_), .Y(u2__abc_52138_new_n14101_));
NOR3X1 NOR3X1_115 ( .A(u2__abc_52138_new_n4666_), .B(u2__abc_52138_new_n4682_), .C(u2__abc_52138_new_n14093_), .Y(u2__abc_52138_new_n14109_));
NOR3X1 NOR3X1_116 ( .A(u2__abc_52138_new_n4671_), .B(u2__abc_52138_new_n4666_), .C(u2__abc_52138_new_n14116_), .Y(u2__abc_52138_new_n14117_));
NOR3X1 NOR3X1_117 ( .A(u2__abc_52138_new_n4700_), .B(u2__abc_52138_new_n4705_), .C(u2__abc_52138_new_n14131_), .Y(u2__abc_52138_new_n14132_));
NOR3X1 NOR3X1_118 ( .A(u2__abc_52138_new_n4689_), .B(u2__abc_52138_new_n4700_), .C(u2__abc_52138_new_n14124_), .Y(u2__abc_52138_new_n14140_));
NOR3X1 NOR3X1_119 ( .A(u2__abc_52138_new_n4694_), .B(u2__abc_52138_new_n4689_), .C(u2__abc_52138_new_n14146_), .Y(u2__abc_52138_new_n14147_));
NOR3X1 NOR3X1_12 ( .A(u2__abc_52138_new_n3607_), .B(u2__abc_52138_new_n3617_), .C(u2__abc_52138_new_n7714_), .Y(u2__abc_52138_new_n7715_));
NOR3X1 NOR3X1_120 ( .A(u2__abc_52138_new_n4655_), .B(u2__abc_52138_new_n4660_), .C(u2__abc_52138_new_n14163_), .Y(u2__abc_52138_new_n14164_));
NOR3X1 NOR3X1_121 ( .A(u2__abc_52138_new_n4642_), .B(u2__abc_52138_new_n4655_), .C(u2__abc_52138_new_n14155_), .Y(u2__abc_52138_new_n14171_));
NOR3X1 NOR3X1_122 ( .A(u2__abc_52138_new_n4647_), .B(u2__abc_52138_new_n4642_), .C(u2__abc_52138_new_n14178_), .Y(u2__abc_52138_new_n14179_));
NOR3X1 NOR3X1_123 ( .A(u2__abc_52138_new_n4630_), .B(u2__abc_52138_new_n4635_), .C(u2__abc_52138_new_n14193_), .Y(u2__abc_52138_new_n14194_));
NOR3X1 NOR3X1_124 ( .A(u2__abc_52138_new_n4619_), .B(u2__abc_52138_new_n4630_), .C(u2__abc_52138_new_n14186_), .Y(u2__abc_52138_new_n14202_));
NOR3X1 NOR3X1_125 ( .A(u2__abc_52138_new_n4624_), .B(u2__abc_52138_new_n4619_), .C(u2__abc_52138_new_n14208_), .Y(u2__abc_52138_new_n14209_));
NOR3X1 NOR3X1_126 ( .A(u2__abc_52138_new_n4584_), .B(u2__abc_52138_new_n4589_), .C(u2__abc_52138_new_n14225_), .Y(u2__abc_52138_new_n14226_));
NOR3X1 NOR3X1_127 ( .A(u2__abc_52138_new_n4573_), .B(u2__abc_52138_new_n4584_), .C(u2__abc_52138_new_n14217_), .Y(u2__abc_52138_new_n14233_));
NOR3X1 NOR3X1_128 ( .A(u2__abc_52138_new_n4578_), .B(u2__abc_52138_new_n4573_), .C(u2__abc_52138_new_n14239_), .Y(u2__abc_52138_new_n14240_));
NOR3X1 NOR3X1_129 ( .A(u2__abc_52138_new_n4609_), .B(u2__abc_52138_new_n4614_), .C(u2__abc_52138_new_n14256_), .Y(u2__abc_52138_new_n14257_));
NOR3X1 NOR3X1_13 ( .A(u2__abc_52138_new_n3072_), .B(u2__abc_52138_new_n3069_), .C(u2__abc_52138_new_n6498_), .Y(u2__abc_52138_new_n13051_));
NOR3X1 NOR3X1_130 ( .A(u2__abc_52138_new_n4596_), .B(u2__abc_52138_new_n4609_), .C(u2__abc_52138_new_n14248_), .Y(u2__abc_52138_new_n14264_));
NOR3X1 NOR3X1_131 ( .A(u2__abc_52138_new_n4601_), .B(u2__abc_52138_new_n4596_), .C(u2__abc_52138_new_n14270_), .Y(u2__abc_52138_new_n14271_));
NOR3X1 NOR3X1_132 ( .A(u2__abc_52138_new_n4536_), .B(u2__abc_52138_new_n4543_), .C(u2__abc_52138_new_n14287_), .Y(u2__abc_52138_new_n14288_));
NOR3X1 NOR3X1_133 ( .A(u2__abc_52138_new_n4525_), .B(u2__abc_52138_new_n4536_), .C(u2__abc_52138_new_n14279_), .Y(u2__abc_52138_new_n14295_));
NOR3X1 NOR3X1_134 ( .A(u2__abc_52138_new_n4530_), .B(u2__abc_52138_new_n4525_), .C(u2__abc_52138_new_n14302_), .Y(u2__abc_52138_new_n14303_));
NOR3X1 NOR3X1_135 ( .A(u2__abc_52138_new_n4559_), .B(u2__abc_52138_new_n4564_), .C(u2__abc_52138_new_n14317_), .Y(u2__abc_52138_new_n14318_));
NOR3X1 NOR3X1_136 ( .A(u2__abc_52138_new_n4548_), .B(u2__abc_52138_new_n4559_), .C(u2__abc_52138_new_n14310_), .Y(u2__abc_52138_new_n14326_));
NOR3X1 NOR3X1_137 ( .A(u2__abc_52138_new_n4553_), .B(u2__abc_52138_new_n4548_), .C(u2__abc_52138_new_n14332_), .Y(u2__abc_52138_new_n14333_));
NOR3X1 NOR3X1_138 ( .A(u2__abc_52138_new_n4512_), .B(u2__abc_52138_new_n4519_), .C(u2__abc_52138_new_n14349_), .Y(u2__abc_52138_new_n14350_));
NOR3X1 NOR3X1_139 ( .A(u2__abc_52138_new_n4501_), .B(u2__abc_52138_new_n4512_), .C(u2__abc_52138_new_n14341_), .Y(u2__abc_52138_new_n14357_));
NOR3X1 NOR3X1_14 ( .A(u2__abc_52138_new_n3074_), .B(u2__abc_52138_new_n3072_), .C(u2__abc_52138_new_n13059_), .Y(u2__abc_52138_new_n13060_));
NOR3X1 NOR3X1_140 ( .A(u2__abc_52138_new_n4506_), .B(u2__abc_52138_new_n4501_), .C(u2__abc_52138_new_n14363_), .Y(u2__abc_52138_new_n14364_));
NOR3X1 NOR3X1_141 ( .A(u2__abc_52138_new_n4489_), .B(u2__abc_52138_new_n4494_), .C(u2__abc_52138_new_n14380_), .Y(u2__abc_52138_new_n14381_));
NOR3X1 NOR3X1_142 ( .A(u2__abc_52138_new_n4478_), .B(u2__abc_52138_new_n4489_), .C(u2__abc_52138_new_n14372_), .Y(u2__abc_52138_new_n14388_));
NOR3X1 NOR3X1_143 ( .A(u2__abc_52138_new_n4483_), .B(u2__abc_52138_new_n4478_), .C(u2__abc_52138_new_n14394_), .Y(u2__abc_52138_new_n14395_));
NOR3X1 NOR3X1_144 ( .A(u2__abc_52138_new_n4469_), .B(u2__abc_52138_new_n4463_), .C(u2__abc_52138_new_n14411_), .Y(u2__abc_52138_new_n14412_));
NOR3X1 NOR3X1_145 ( .A(u2__abc_52138_new_n4452_), .B(u2__abc_52138_new_n4469_), .C(u2__abc_52138_new_n14403_), .Y(u2__abc_52138_new_n14419_));
NOR3X1 NOR3X1_146 ( .A(u2__abc_52138_new_n4457_), .B(u2__abc_52138_new_n4452_), .C(u2__abc_52138_new_n14425_), .Y(u2__abc_52138_new_n14426_));
NOR3X1 NOR3X1_147 ( .A(u2__abc_52138_new_n4440_), .B(u2__abc_52138_new_n4445_), .C(u2__abc_52138_new_n14442_), .Y(u2__abc_52138_new_n14443_));
NOR3X1 NOR3X1_148 ( .A(u2__abc_52138_new_n4429_), .B(u2__abc_52138_new_n4440_), .C(u2__abc_52138_new_n14434_), .Y(u2__abc_52138_new_n14450_));
NOR3X1 NOR3X1_149 ( .A(u2__abc_52138_new_n4434_), .B(u2__abc_52138_new_n4429_), .C(u2__abc_52138_new_n14456_), .Y(u2__abc_52138_new_n14457_));
NOR3X1 NOR3X1_15 ( .A(u2__abc_52138_new_n3079_), .B(u2__abc_52138_new_n3060_), .C(u2__abc_52138_new_n13075_), .Y(u2__abc_52138_new_n13076_));
NOR3X1 NOR3X1_150 ( .A(u2__abc_52138_new_n4387_), .B(u2__abc_52138_new_n4382_), .C(u2__abc_52138_new_n14473_), .Y(u2__abc_52138_new_n14474_));
NOR3X1 NOR3X1_151 ( .A(u2__abc_52138_new_n4393_), .B(u2__abc_52138_new_n4387_), .C(u2__abc_52138_new_n14465_), .Y(u2__abc_52138_new_n14481_));
NOR3X1 NOR3X1_152 ( .A(u2__abc_52138_new_n4398_), .B(u2__abc_52138_new_n4393_), .C(u2__abc_52138_new_n14487_), .Y(u2__abc_52138_new_n14488_));
NOR3X1 NOR3X1_153 ( .A(u2__abc_52138_new_n4416_), .B(u2__abc_52138_new_n4421_), .C(u2__abc_52138_new_n14504_), .Y(u2__abc_52138_new_n14505_));
NOR3X1 NOR3X1_154 ( .A(u2__abc_52138_new_n4405_), .B(u2__abc_52138_new_n4416_), .C(u2__abc_52138_new_n14496_), .Y(u2__abc_52138_new_n14512_));
NOR3X1 NOR3X1_155 ( .A(u2__abc_52138_new_n4410_), .B(u2__abc_52138_new_n4405_), .C(u2__abc_52138_new_n14518_), .Y(u2__abc_52138_new_n14519_));
NOR3X1 NOR3X1_156 ( .A(u2__abc_52138_new_n4372_), .B(u2__abc_52138_new_n4366_), .C(u2__abc_52138_new_n14534_), .Y(u2__abc_52138_new_n14535_));
NOR3X1 NOR3X1_157 ( .A(u2__abc_52138_new_n4356_), .B(u2__abc_52138_new_n4372_), .C(u2__abc_52138_new_n14527_), .Y(u2__abc_52138_new_n14543_));
NOR3X1 NOR3X1_158 ( .A(u2__abc_52138_new_n4358_), .B(u2__abc_52138_new_n4356_), .C(u2__abc_52138_new_n14550_), .Y(u2__abc_52138_new_n14551_));
NOR3X1 NOR3X1_159 ( .A(u2__abc_52138_new_n4342_), .B(u2__abc_52138_new_n4347_), .C(u2__abc_52138_new_n14565_), .Y(u2__abc_52138_new_n14566_));
NOR3X1 NOR3X1_16 ( .A(u2__abc_52138_new_n6458_), .B(u2__abc_52138_new_n3079_), .C(u2__abc_52138_new_n13067_), .Y(u2__abc_52138_new_n13083_));
NOR3X1 NOR3X1_160 ( .A(u2__abc_52138_new_n4331_), .B(u2__abc_52138_new_n4342_), .C(u2__abc_52138_new_n14558_), .Y(u2__abc_52138_new_n14574_));
NOR3X1 NOR3X1_161 ( .A(u2__abc_52138_new_n4336_), .B(u2__abc_52138_new_n4331_), .C(u2__abc_52138_new_n14580_), .Y(u2__abc_52138_new_n14581_));
NOR3X1 NOR3X1_162 ( .A(u2__abc_52138_new_n4300_), .B(u2__abc_52138_new_n4305_), .C(u2__abc_52138_new_n14597_), .Y(u2__abc_52138_new_n14598_));
NOR3X1 NOR3X1_163 ( .A(u2__abc_52138_new_n4289_), .B(u2__abc_52138_new_n4300_), .C(u2__abc_52138_new_n14589_), .Y(u2__abc_52138_new_n14605_));
NOR3X1 NOR3X1_164 ( .A(u2__abc_52138_new_n4294_), .B(u2__abc_52138_new_n4289_), .C(u2__abc_52138_new_n14611_), .Y(u2__abc_52138_new_n14612_));
NOR3X1 NOR3X1_165 ( .A(u2__abc_52138_new_n4325_), .B(u2__abc_52138_new_n14615_), .C(u2__abc_52138_new_n14629_), .Y(u2__abc_52138_new_n14630_));
NOR3X1 NOR3X1_166 ( .A(u2__abc_52138_new_n4312_), .B(u2__abc_52138_new_n4325_), .C(u2__abc_52138_new_n14621_), .Y(u2__abc_52138_new_n14637_));
NOR3X1 NOR3X1_167 ( .A(u2__abc_52138_new_n4317_), .B(u2__abc_52138_new_n4312_), .C(u2__abc_52138_new_n14643_), .Y(u2__abc_52138_new_n14644_));
NOR3X1 NOR3X1_168 ( .A(u2__abc_52138_new_n4257_), .B(u2__abc_52138_new_n4252_), .C(u2__abc_52138_new_n14660_), .Y(u2__abc_52138_new_n14661_));
NOR3X1 NOR3X1_169 ( .A(u2__abc_52138_new_n4241_), .B(u2__abc_52138_new_n4257_), .C(u2__abc_52138_new_n14652_), .Y(u2__abc_52138_new_n14668_));
NOR3X1 NOR3X1_17 ( .A(u2__abc_52138_new_n3056_), .B(u2__abc_52138_new_n6458_), .C(u2__abc_52138_new_n13090_), .Y(u2__abc_52138_new_n13091_));
NOR3X1 NOR3X1_170 ( .A(u2__abc_52138_new_n4246_), .B(u2__abc_52138_new_n4241_), .C(u2__abc_52138_new_n14674_), .Y(u2__abc_52138_new_n14675_));
NOR3X1 NOR3X1_171 ( .A(u2__abc_52138_new_n4277_), .B(u2__abc_52138_new_n4282_), .C(u2__abc_52138_new_n14691_), .Y(u2__abc_52138_new_n14692_));
NOR3X1 NOR3X1_172 ( .A(u2__abc_52138_new_n4266_), .B(u2__abc_52138_new_n4277_), .C(u2__abc_52138_new_n14683_), .Y(u2__abc_52138_new_n14699_));
NOR3X1 NOR3X1_173 ( .A(u2__abc_52138_new_n4271_), .B(u2__abc_52138_new_n4266_), .C(u2__abc_52138_new_n14705_), .Y(u2__abc_52138_new_n14706_));
NOR3X1 NOR3X1_174 ( .A(u2__abc_52138_new_n4210_), .B(u2__abc_52138_new_n4205_), .C(u2__abc_52138_new_n14722_), .Y(u2__abc_52138_new_n14723_));
NOR3X1 NOR3X1_175 ( .A(u2__abc_52138_new_n4194_), .B(u2__abc_52138_new_n4210_), .C(u2__abc_52138_new_n14714_), .Y(u2__abc_52138_new_n14730_));
NOR3X1 NOR3X1_176 ( .A(u2__abc_52138_new_n4199_), .B(u2__abc_52138_new_n4194_), .C(u2__abc_52138_new_n14736_), .Y(u2__abc_52138_new_n14737_));
NOR3X1 NOR3X1_177 ( .A(u2__abc_52138_new_n4230_), .B(u2__abc_52138_new_n4233_), .C(u2__abc_52138_new_n14753_), .Y(u2__abc_52138_new_n14754_));
NOR3X1 NOR3X1_178 ( .A(u2__abc_52138_new_n4217_), .B(u2__abc_52138_new_n4230_), .C(u2__abc_52138_new_n14745_), .Y(u2__abc_52138_new_n14761_));
NOR3X1 NOR3X1_179 ( .A(u2__abc_52138_new_n4222_), .B(u2__abc_52138_new_n4217_), .C(u2__abc_52138_new_n14767_), .Y(u2__abc_52138_new_n14768_));
NOR3X1 NOR3X1_18 ( .A(u2__abc_52138_new_n3040_), .B(u2__abc_52138_new_n3045_), .C(u2__abc_52138_new_n13106_), .Y(u2__abc_52138_new_n13107_));
NOR3X1 NOR3X1_180 ( .A(u2__abc_52138_new_n4157_), .B(u2__abc_52138_new_n4162_), .C(u2__abc_52138_new_n14783_), .Y(u2__abc_52138_new_n14784_));
NOR3X1 NOR3X1_181 ( .A(u2__abc_52138_new_n4146_), .B(u2__abc_52138_new_n4157_), .C(u2__abc_52138_new_n14776_), .Y(u2__abc_52138_new_n14792_));
NOR3X1 NOR3X1_182 ( .A(u2__abc_52138_new_n4151_), .B(u2__abc_52138_new_n4146_), .C(u2__abc_52138_new_n14798_), .Y(u2__abc_52138_new_n14799_));
NOR3X1 NOR3X1_183 ( .A(u2__abc_52138_new_n4182_), .B(u2__abc_52138_new_n4187_), .C(u2__abc_52138_new_n14815_), .Y(u2__abc_52138_new_n14816_));
NOR3X1 NOR3X1_184 ( .A(u2__abc_52138_new_n4169_), .B(u2__abc_52138_new_n4182_), .C(u2__abc_52138_new_n14807_), .Y(u2__abc_52138_new_n14823_));
NOR3X1 NOR3X1_185 ( .A(u2__abc_52138_new_n4174_), .B(u2__abc_52138_new_n4169_), .C(u2__abc_52138_new_n14829_), .Y(u2__abc_52138_new_n14830_));
NOR3X1 NOR3X1_186 ( .A(u2__abc_52138_new_n4960_), .B(u2__abc_52138_new_n4140_), .C(u2__abc_52138_new_n14846_), .Y(u2__abc_52138_new_n14847_));
NOR3X1 NOR3X1_187 ( .A(u2__abc_52138_new_n4123_), .B(u2__abc_52138_new_n4960_), .C(u2__abc_52138_new_n14838_), .Y(u2__abc_52138_new_n14854_));
NOR3X1 NOR3X1_188 ( .A(u2__abc_52138_new_n4128_), .B(u2__abc_52138_new_n4123_), .C(u2__abc_52138_new_n14860_), .Y(u2__abc_52138_new_n14861_));
NOR3X1 NOR3X1_189 ( .A(u2__abc_52138_new_n4110_), .B(u2__abc_52138_new_n4115_), .C(u2__abc_52138_new_n14877_), .Y(u2__abc_52138_new_n14878_));
NOR3X1 NOR3X1_19 ( .A(u2__abc_52138_new_n3096_), .B(u2__abc_52138_new_n3040_), .C(u2__abc_52138_new_n13098_), .Y(u2__abc_52138_new_n13114_));
NOR3X1 NOR3X1_190 ( .A(u2__abc_52138_new_n4099_), .B(u2__abc_52138_new_n4110_), .C(u2__abc_52138_new_n14869_), .Y(u2__abc_52138_new_n14885_));
NOR3X1 NOR3X1_191 ( .A(u2__abc_52138_new_n4104_), .B(u2__abc_52138_new_n4099_), .C(u2__abc_52138_new_n14891_), .Y(u2__abc_52138_new_n14892_));
NOR3X1 NOR3X1_192 ( .A(u2__abc_52138_new_n4055_), .B(u2__abc_52138_new_n4050_), .C(u2__abc_52138_new_n14907_), .Y(u2__abc_52138_new_n14908_));
NOR3X1 NOR3X1_193 ( .A(u2__abc_52138_new_n4061_), .B(u2__abc_52138_new_n4055_), .C(u2__abc_52138_new_n14900_), .Y(u2__abc_52138_new_n14916_));
NOR3X1 NOR3X1_194 ( .A(u2__abc_52138_new_n4066_), .B(u2__abc_52138_new_n4061_), .C(u2__abc_52138_new_n14922_), .Y(u2__abc_52138_new_n14923_));
NOR3X1 NOR3X1_195 ( .A(u2__abc_52138_new_n4087_), .B(u2__abc_52138_new_n4090_), .C(u2__abc_52138_new_n14939_), .Y(u2__abc_52138_new_n14940_));
NOR3X1 NOR3X1_196 ( .A(u2__abc_52138_new_n4074_), .B(u2__abc_52138_new_n4087_), .C(u2__abc_52138_new_n14931_), .Y(u2__abc_52138_new_n14947_));
NOR3X1 NOR3X1_197 ( .A(u2__abc_52138_new_n4079_), .B(u2__abc_52138_new_n4074_), .C(u2__abc_52138_new_n14953_), .Y(u2__abc_52138_new_n14954_));
NOR3X1 NOR3X1_198 ( .A(u2__abc_52138_new_n4008_), .B(u2__abc_52138_new_n4003_), .C(u2__abc_52138_new_n14969_), .Y(u2__abc_52138_new_n14970_));
NOR3X1 NOR3X1_199 ( .A(u2__abc_52138_new_n4014_), .B(u2__abc_52138_new_n4008_), .C(u2__abc_52138_new_n14962_), .Y(u2__abc_52138_new_n14978_));
NOR3X1 NOR3X1_2 ( .A(_abc_65734_new_n1481_), .B(_abc_65734_new_n1493_), .C(_abc_65734_new_n1472_), .Y(_abc_65734_new_n1511_));
NOR3X1 NOR3X1_20 ( .A(u2__abc_52138_new_n3035_), .B(u2__abc_52138_new_n3096_), .C(u2__abc_52138_new_n13121_), .Y(u2__abc_52138_new_n13122_));
NOR3X1 NOR3X1_200 ( .A(u2__abc_52138_new_n4019_), .B(u2__abc_52138_new_n4014_), .C(u2__abc_52138_new_n14984_), .Y(u2__abc_52138_new_n14985_));
NOR3X1 NOR3X1_201 ( .A(u2__abc_52138_new_n4037_), .B(u2__abc_52138_new_n4042_), .C(u2__abc_52138_new_n15000_), .Y(u2__abc_52138_new_n15001_));
NOR3X1 NOR3X1_202 ( .A(u2__abc_52138_new_n4026_), .B(u2__abc_52138_new_n4037_), .C(u2__abc_52138_new_n14993_), .Y(u2__abc_52138_new_n15009_));
NOR3X1 NOR3X1_203 ( .A(u2__abc_52138_new_n4033_), .B(u2__abc_52138_new_n4026_), .C(u2__abc_52138_new_n15015_), .Y(u2__abc_52138_new_n15016_));
NOR3X1 NOR3X1_204 ( .A(u2__abc_52138_new_n5692_), .B(u2__abc_52138_new_n5687_), .C(u2__abc_52138_new_n15031_), .Y(u2__abc_52138_new_n15032_));
NOR3X1 NOR3X1_205 ( .A(u2__abc_52138_new_n5699_), .B(u2__abc_52138_new_n5692_), .C(u2__abc_52138_new_n15024_), .Y(u2__abc_52138_new_n15040_));
NOR3X1 NOR3X1_206 ( .A(u2__abc_52138_new_n5704_), .B(u2__abc_52138_new_n5699_), .C(u2__abc_52138_new_n15047_), .Y(u2__abc_52138_new_n15048_));
NOR3X1 NOR3X1_207 ( .A(u2__abc_52138_new_n5727_), .B(u2__abc_52138_new_n5722_), .C(u2__abc_52138_new_n15062_), .Y(u2__abc_52138_new_n15063_));
NOR3X1 NOR3X1_208 ( .A(u2__abc_52138_new_n5711_), .B(u2__abc_52138_new_n5727_), .C(u2__abc_52138_new_n15055_), .Y(u2__abc_52138_new_n15071_));
NOR3X1 NOR3X1_209 ( .A(u2__abc_52138_new_n5716_), .B(u2__abc_52138_new_n5711_), .C(u2__abc_52138_new_n15077_), .Y(u2__abc_52138_new_n15078_));
NOR3X1 NOR3X1_21 ( .A(u2__abc_52138_new_n3022_), .B(u2__abc_52138_new_n3027_), .C(u2__abc_52138_new_n13137_), .Y(u2__abc_52138_new_n13138_));
NOR3X1 NOR3X1_210 ( .A(u2__abc_52138_new_n5679_), .B(u2__abc_52138_new_n5674_), .C(u2__abc_52138_new_n15094_), .Y(u2__abc_52138_new_n15095_));
NOR3X1 NOR3X1_211 ( .A(u2__abc_52138_new_n5665_), .B(u2__abc_52138_new_n5679_), .C(u2__abc_52138_new_n15086_), .Y(u2__abc_52138_new_n15102_));
NOR3X1 NOR3X1_212 ( .A(u2__abc_52138_new_n5670_), .B(u2__abc_52138_new_n5665_), .C(u2__abc_52138_new_n15108_), .Y(u2__abc_52138_new_n15109_));
NOR3X1 NOR3X1_213 ( .A(u2__abc_52138_new_n5658_), .B(u2__abc_52138_new_n5653_), .C(u2__abc_52138_new_n15125_), .Y(u2__abc_52138_new_n15126_));
NOR3X1 NOR3X1_214 ( .A(u2__abc_52138_new_n5640_), .B(u2__abc_52138_new_n5658_), .C(u2__abc_52138_new_n15117_), .Y(u2__abc_52138_new_n15133_));
NOR3X1 NOR3X1_215 ( .A(u2__abc_52138_new_n5645_), .B(u2__abc_52138_new_n5640_), .C(u2__abc_52138_new_n15139_), .Y(u2__abc_52138_new_n15140_));
NOR3X1 NOR3X1_216 ( .A(u2__abc_52138_new_n5613_), .B(u2__abc_52138_new_n5608_), .C(u2__abc_52138_new_n15156_), .Y(u2__abc_52138_new_n15157_));
NOR3X1 NOR3X1_217 ( .A(u2__abc_52138_new_n5597_), .B(u2__abc_52138_new_n5613_), .C(u2__abc_52138_new_n15148_), .Y(u2__abc_52138_new_n15164_));
NOR3X1 NOR3X1_218 ( .A(u2__abc_52138_new_n5602_), .B(u2__abc_52138_new_n5597_), .C(u2__abc_52138_new_n15170_), .Y(u2__abc_52138_new_n15171_));
NOR3X1 NOR3X1_219 ( .A(u2__abc_52138_new_n5632_), .B(u2__abc_52138_new_n5761_), .C(u2__abc_52138_new_n15187_), .Y(u2__abc_52138_new_n15188_));
NOR3X1 NOR3X1_22 ( .A(u2__abc_52138_new_n6654_), .B(u2__abc_52138_new_n3022_), .C(u2__abc_52138_new_n13129_), .Y(u2__abc_52138_new_n13145_));
NOR3X1 NOR3X1_220 ( .A(u2__abc_52138_new_n5620_), .B(u2__abc_52138_new_n5632_), .C(u2__abc_52138_new_n15179_), .Y(u2__abc_52138_new_n15195_));
NOR3X1 NOR3X1_221 ( .A(u2__abc_52138_new_n5625_), .B(u2__abc_52138_new_n5620_), .C(u2__abc_52138_new_n15201_), .Y(u2__abc_52138_new_n15202_));
NOR3X1 NOR3X1_222 ( .A(u2__abc_52138_new_n5566_), .B(u2__abc_52138_new_n5561_), .C(u2__abc_52138_new_n15218_), .Y(u2__abc_52138_new_n15219_));
NOR3X1 NOR3X1_223 ( .A(u2__abc_52138_new_n5550_), .B(u2__abc_52138_new_n5566_), .C(u2__abc_52138_new_n15210_), .Y(u2__abc_52138_new_n15226_));
NOR3X1 NOR3X1_224 ( .A(u2__abc_52138_new_n5555_), .B(u2__abc_52138_new_n5550_), .C(u2__abc_52138_new_n15232_), .Y(u2__abc_52138_new_n15233_));
NOR3X1 NOR3X1_225 ( .A(u2__abc_52138_new_n5589_), .B(u2__abc_52138_new_n5584_), .C(u2__abc_52138_new_n15249_), .Y(u2__abc_52138_new_n15250_));
NOR3X1 NOR3X1_226 ( .A(u2__abc_52138_new_n5573_), .B(u2__abc_52138_new_n5589_), .C(u2__abc_52138_new_n15241_), .Y(u2__abc_52138_new_n15257_));
NOR3X1 NOR3X1_227 ( .A(u2__abc_52138_new_n5578_), .B(u2__abc_52138_new_n5573_), .C(u2__abc_52138_new_n15263_), .Y(u2__abc_52138_new_n15264_));
NOR3X1 NOR3X1_228 ( .A(u2__abc_52138_new_n5520_), .B(u2__abc_52138_new_n5515_), .C(u2__abc_52138_new_n15279_), .Y(u2__abc_52138_new_n15280_));
NOR3X1 NOR3X1_229 ( .A(u2__abc_52138_new_n5504_), .B(u2__abc_52138_new_n5520_), .C(u2__abc_52138_new_n15272_), .Y(u2__abc_52138_new_n15288_));
NOR3X1 NOR3X1_23 ( .A(u2__abc_52138_new_n3019_), .B(u2__abc_52138_new_n6654_), .C(u2__abc_52138_new_n13152_), .Y(u2__abc_52138_new_n13153_));
NOR3X1 NOR3X1_230 ( .A(u2__abc_52138_new_n5509_), .B(u2__abc_52138_new_n5504_), .C(u2__abc_52138_new_n15294_), .Y(u2__abc_52138_new_n15295_));
NOR3X1 NOR3X1_231 ( .A(u2__abc_52138_new_n5539_), .B(u2__abc_52138_new_n5787_), .C(u2__abc_52138_new_n15311_), .Y(u2__abc_52138_new_n15312_));
NOR3X1 NOR3X1_232 ( .A(u2__abc_52138_new_n5527_), .B(u2__abc_52138_new_n5539_), .C(u2__abc_52138_new_n15303_), .Y(u2__abc_52138_new_n15319_));
NOR3X1 NOR3X1_233 ( .A(u2__abc_52138_new_n5532_), .B(u2__abc_52138_new_n5527_), .C(u2__abc_52138_new_n15325_), .Y(u2__abc_52138_new_n15326_));
NOR3X1 NOR3X1_234 ( .A(u2__abc_52138_new_n5462_), .B(u2__abc_52138_new_n5455_), .C(u2__abc_52138_new_n15342_), .Y(u2__abc_52138_new_n15343_));
NOR3X1 NOR3X1_235 ( .A(u2__abc_52138_new_n5468_), .B(u2__abc_52138_new_n5462_), .C(u2__abc_52138_new_n15334_), .Y(u2__abc_52138_new_n15350_));
NOR3X1 NOR3X1_236 ( .A(u2__abc_52138_new_n5473_), .B(u2__abc_52138_new_n5468_), .C(u2__abc_52138_new_n15356_), .Y(u2__abc_52138_new_n15357_));
NOR3X1 NOR3X1_237 ( .A(u2__abc_52138_new_n5496_), .B(u2__abc_52138_new_n5491_), .C(u2__abc_52138_new_n15373_), .Y(u2__abc_52138_new_n15374_));
NOR3X1 NOR3X1_238 ( .A(u2__abc_52138_new_n5480_), .B(u2__abc_52138_new_n5496_), .C(u2__abc_52138_new_n15365_), .Y(u2__abc_52138_new_n15381_));
NOR3X1 NOR3X1_239 ( .A(u2__abc_52138_new_n5485_), .B(u2__abc_52138_new_n5480_), .C(u2__abc_52138_new_n15387_), .Y(u2__abc_52138_new_n15388_));
NOR3X1 NOR3X1_24 ( .A(u2__abc_52138_new_n3175_), .B(u2__abc_52138_new_n3170_), .C(u2__abc_52138_new_n13168_), .Y(u2__abc_52138_new_n13169_));
NOR3X1 NOR3X1_240 ( .A(u2__abc_52138_new_n5412_), .B(u2__abc_52138_new_n5407_), .C(u2__abc_52138_new_n15403_), .Y(u2__abc_52138_new_n15404_));
NOR3X1 NOR3X1_241 ( .A(u2__abc_52138_new_n5420_), .B(u2__abc_52138_new_n5412_), .C(u2__abc_52138_new_n15396_), .Y(u2__abc_52138_new_n15412_));
NOR3X1 NOR3X1_242 ( .A(u2__abc_52138_new_n5425_), .B(u2__abc_52138_new_n5420_), .C(u2__abc_52138_new_n15418_), .Y(u2__abc_52138_new_n15419_));
NOR3X1 NOR3X1_243 ( .A(u2__abc_52138_new_n5443_), .B(u2__abc_52138_new_n5448_), .C(u2__abc_52138_new_n15435_), .Y(u2__abc_52138_new_n15436_));
NOR3X1 NOR3X1_244 ( .A(u2__abc_52138_new_n5432_), .B(u2__abc_52138_new_n5443_), .C(u2__abc_52138_new_n15427_), .Y(u2__abc_52138_new_n15443_));
NOR3X1 NOR3X1_245 ( .A(u2__abc_52138_new_n5437_), .B(u2__abc_52138_new_n5432_), .C(u2__abc_52138_new_n15449_), .Y(u2__abc_52138_new_n15450_));
NOR3X1 NOR3X1_246 ( .A(u2__abc_52138_new_n5382_), .B(u2__abc_52138_new_n5811_), .C(u2__abc_52138_new_n15465_), .Y(u2__abc_52138_new_n15466_));
NOR3X1 NOR3X1_247 ( .A(u2__abc_52138_new_n5370_), .B(u2__abc_52138_new_n5382_), .C(u2__abc_52138_new_n15458_), .Y(u2__abc_52138_new_n15474_));
NOR3X1 NOR3X1_248 ( .A(u2__abc_52138_new_n5375_), .B(u2__abc_52138_new_n5370_), .C(u2__abc_52138_new_n15480_), .Y(u2__abc_52138_new_n15481_));
NOR3X1 NOR3X1_249 ( .A(u2__abc_52138_new_n5401_), .B(u2__abc_52138_new_n15484_), .C(u2__abc_52138_new_n15497_), .Y(u2__abc_52138_new_n15498_));
NOR3X1 NOR3X1_25 ( .A(u2__abc_52138_new_n3159_), .B(u2__abc_52138_new_n3175_), .C(u2__abc_52138_new_n13160_), .Y(u2__abc_52138_new_n13176_));
NOR3X1 NOR3X1_250 ( .A(u2__abc_52138_new_n5389_), .B(u2__abc_52138_new_n5401_), .C(u2__abc_52138_new_n15490_), .Y(u2__abc_52138_new_n15506_));
NOR3X1 NOR3X1_251 ( .A(u2__abc_52138_new_n5394_), .B(u2__abc_52138_new_n5389_), .C(u2__abc_52138_new_n15512_), .Y(u2__abc_52138_new_n15513_));
NOR3X1 NOR3X1_252 ( .A(u2__abc_52138_new_n5348_), .B(u2__abc_52138_new_n5341_), .C(u2__abc_52138_new_n15528_), .Y(u2__abc_52138_new_n15529_));
NOR3X1 NOR3X1_253 ( .A(u2__abc_52138_new_n5354_), .B(u2__abc_52138_new_n5348_), .C(u2__abc_52138_new_n15521_), .Y(u2__abc_52138_new_n15537_));
NOR3X1 NOR3X1_254 ( .A(u2__abc_52138_new_n5359_), .B(u2__abc_52138_new_n5354_), .C(u2__abc_52138_new_n15543_), .Y(u2__abc_52138_new_n15544_));
NOR3X1 NOR3X1_255 ( .A(u2__abc_52138_new_n5333_), .B(u2__abc_52138_new_n5844_), .C(u2__abc_52138_new_n15560_), .Y(u2__abc_52138_new_n15561_));
NOR3X1 NOR3X1_256 ( .A(u2__abc_52138_new_n5321_), .B(u2__abc_52138_new_n5333_), .C(u2__abc_52138_new_n15552_), .Y(u2__abc_52138_new_n15568_));
NOR3X1 NOR3X1_257 ( .A(u2__abc_52138_new_n5326_), .B(u2__abc_52138_new_n5321_), .C(u2__abc_52138_new_n15574_), .Y(u2__abc_52138_new_n15575_));
NOR3X1 NOR3X1_258 ( .A(u2__abc_52138_new_n5281_), .B(u2__abc_52138_new_n5274_), .C(u2__abc_52138_new_n15591_), .Y(u2__abc_52138_new_n15592_));
NOR3X1 NOR3X1_259 ( .A(u2__abc_52138_new_n5287_), .B(u2__abc_52138_new_n5281_), .C(u2__abc_52138_new_n15583_), .Y(u2__abc_52138_new_n15599_));
NOR3X1 NOR3X1_26 ( .A(u2__abc_52138_new_n3164_), .B(u2__abc_52138_new_n3159_), .C(u2__abc_52138_new_n13183_), .Y(u2__abc_52138_new_n13184_));
NOR3X1 NOR3X1_260 ( .A(u2__abc_52138_new_n5292_), .B(u2__abc_52138_new_n5287_), .C(u2__abc_52138_new_n15605_), .Y(u2__abc_52138_new_n15606_));
NOR3X1 NOR3X1_261 ( .A(u2__abc_52138_new_n5315_), .B(u2__abc_52138_new_n5310_), .C(u2__abc_52138_new_n15622_), .Y(u2__abc_52138_new_n15623_));
NOR3X1 NOR3X1_262 ( .A(u2__abc_52138_new_n5299_), .B(u2__abc_52138_new_n5315_), .C(u2__abc_52138_new_n15614_), .Y(u2__abc_52138_new_n15630_));
NOR3X1 NOR3X1_263 ( .A(u2__abc_52138_new_n5304_), .B(u2__abc_52138_new_n5299_), .C(u2__abc_52138_new_n15636_), .Y(u2__abc_52138_new_n15637_));
NOR3X1 NOR3X1_264 ( .A(u2__abc_52138_new_n5242_), .B(u2__abc_52138_new_n15640_), .C(u2__abc_52138_new_n15653_), .Y(u2__abc_52138_new_n15654_));
NOR3X1 NOR3X1_265 ( .A(u2__abc_52138_new_n5231_), .B(u2__abc_52138_new_n5242_), .C(u2__abc_52138_new_n15646_), .Y(u2__abc_52138_new_n15662_));
NOR3X1 NOR3X1_266 ( .A(u2__abc_52138_new_n5236_), .B(u2__abc_52138_new_n5231_), .C(u2__abc_52138_new_n15668_), .Y(u2__abc_52138_new_n15669_));
NOR3X1 NOR3X1_267 ( .A(u2__abc_52138_new_n5268_), .B(u2__abc_52138_new_n15672_), .C(u2__abc_52138_new_n15686_), .Y(u2__abc_52138_new_n15687_));
NOR3X1 NOR3X1_268 ( .A(u2__abc_52138_new_n5249_), .B(u2__abc_52138_new_n5268_), .C(u2__abc_52138_new_n15678_), .Y(u2__abc_52138_new_n15694_));
NOR3X1 NOR3X1_269 ( .A(u2__abc_52138_new_n5256_), .B(u2__abc_52138_new_n5249_), .C(u2__abc_52138_new_n15700_), .Y(u2__abc_52138_new_n15701_));
NOR3X1 NOR3X1_27 ( .A(u2__abc_52138_new_n3206_), .B(u2__abc_52138_new_n3189_), .C(u2__abc_52138_new_n13199_), .Y(u2__abc_52138_new_n13200_));
NOR3X1 NOR3X1_270 ( .A(u2__abc_52138_new_n5202_), .B(u2__abc_52138_new_n5197_), .C(u2__abc_52138_new_n15716_), .Y(u2__abc_52138_new_n15717_));
NOR3X1 NOR3X1_271 ( .A(u2__abc_52138_new_n5183_), .B(u2__abc_52138_new_n5202_), .C(u2__abc_52138_new_n15709_), .Y(u2__abc_52138_new_n15725_));
NOR3X1 NOR3X1_272 ( .A(u2__abc_52138_new_n5190_), .B(u2__abc_52138_new_n5183_), .C(u2__abc_52138_new_n15731_), .Y(u2__abc_52138_new_n15732_));
NOR3X1 NOR3X1_273 ( .A(u2__abc_52138_new_n5223_), .B(u2__abc_52138_new_n5218_), .C(u2__abc_52138_new_n15747_), .Y(u2__abc_52138_new_n15748_));
NOR3X1 NOR3X1_274 ( .A(u2__abc_52138_new_n5206_), .B(u2__abc_52138_new_n5223_), .C(u2__abc_52138_new_n15740_), .Y(u2__abc_52138_new_n15756_));
NOR3X1 NOR3X1_275 ( .A(u2__abc_52138_new_n5212_), .B(u2__abc_52138_new_n5206_), .C(u2__abc_52138_new_n15762_), .Y(u2__abc_52138_new_n15763_));
NOR3X1 NOR3X1_276 ( .A(u2__abc_52138_new_n5152_), .B(u2__abc_52138_new_n5147_), .C(u2__abc_52138_new_n15778_), .Y(u2__abc_52138_new_n15779_));
NOR3X1 NOR3X1_277 ( .A(u2__abc_52138_new_n5136_), .B(u2__abc_52138_new_n5152_), .C(u2__abc_52138_new_n15771_), .Y(u2__abc_52138_new_n15787_));
NOR3X1 NOR3X1_278 ( .A(u2__abc_52138_new_n5141_), .B(u2__abc_52138_new_n5136_), .C(u2__abc_52138_new_n15793_), .Y(u2__abc_52138_new_n15794_));
NOR3X1 NOR3X1_279 ( .A(u2__abc_52138_new_n5175_), .B(u2__abc_52138_new_n5170_), .C(u2__abc_52138_new_n15810_), .Y(u2__abc_52138_new_n15811_));
NOR3X1 NOR3X1_28 ( .A(u2__abc_52138_new_n6733_), .B(u2__abc_52138_new_n3206_), .C(u2__abc_52138_new_n13191_), .Y(u2__abc_52138_new_n13207_));
NOR3X1 NOR3X1_280 ( .A(u2__abc_52138_new_n5159_), .B(u2__abc_52138_new_n5175_), .C(u2__abc_52138_new_n15802_), .Y(u2__abc_52138_new_n15818_));
NOR3X1 NOR3X1_281 ( .A(u2__abc_52138_new_n5164_), .B(u2__abc_52138_new_n5159_), .C(u2__abc_52138_new_n15824_), .Y(u2__abc_52138_new_n15825_));
NOR3X1 NOR3X1_282 ( .A(u2__abc_52138_new_n5098_), .B(u2__abc_52138_new_n5091_), .C(u2__abc_52138_new_n15840_), .Y(u2__abc_52138_new_n15841_));
NOR3X1 NOR3X1_283 ( .A(u2__abc_52138_new_n5104_), .B(u2__abc_52138_new_n5098_), .C(u2__abc_52138_new_n15833_), .Y(u2__abc_52138_new_n15849_));
NOR3X1 NOR3X1_284 ( .A(u2__abc_52138_new_n5107_), .B(u2__abc_52138_new_n5104_), .C(u2__abc_52138_new_n15855_), .Y(u2__abc_52138_new_n15856_));
NOR3X1 NOR3X1_285 ( .A(u2__abc_52138_new_n5128_), .B(u2__abc_52138_new_n5911_), .C(u2__abc_52138_new_n15871_), .Y(u2__abc_52138_new_n15872_));
NOR3X1 NOR3X1_286 ( .A(u2__abc_52138_new_n5116_), .B(u2__abc_52138_new_n5128_), .C(u2__abc_52138_new_n15864_), .Y(u2__abc_52138_new_n15880_));
NOR3X1 NOR3X1_287 ( .A(u2__abc_52138_new_n5121_), .B(u2__abc_52138_new_n5116_), .C(u2__abc_52138_new_n15886_), .Y(u2__abc_52138_new_n15887_));
NOR3X1 NOR3X1_288 ( .A(u2__abc_52138_new_n5057_), .B(u2__abc_52138_new_n5890_), .C(u2__abc_52138_new_n15902_), .Y(u2__abc_52138_new_n15903_));
NOR3X1 NOR3X1_289 ( .A(u2__abc_52138_new_n5047_), .B(u2__abc_52138_new_n5057_), .C(u2__abc_52138_new_n15895_), .Y(u2__abc_52138_new_n15911_));
NOR3X1 NOR3X1_29 ( .A(u2__abc_52138_new_n3183_), .B(u2__abc_52138_new_n6733_), .C(u2__abc_52138_new_n13214_), .Y(u2__abc_52138_new_n13215_));
NOR3X1 NOR3X1_290 ( .A(u2__abc_52138_new_n15913_), .B(u2__abc_52138_new_n5047_), .C(u2__abc_52138_new_n15918_), .Y(u2__abc_52138_new_n15919_));
NOR3X1 NOR3X1_291 ( .A(u2__abc_52138_new_n5076_), .B(u2__abc_52138_new_n5082_), .C(u2__abc_52138_new_n15934_), .Y(u2__abc_52138_new_n15935_));
NOR3X1 NOR3X1_292 ( .A(u2__abc_52138_new_n5067_), .B(u2__abc_52138_new_n5076_), .C(u2__abc_52138_new_n15927_), .Y(u2__abc_52138_new_n15943_));
NOR3X1 NOR3X1_293 ( .A(u2__abc_52138_new_n5072_), .B(u2__abc_52138_new_n5067_), .C(u2__abc_52138_new_n15949_), .Y(u2__abc_52138_new_n15950_));
NOR3X1 NOR3X1_294 ( .A(u2__abc_52138_new_n5025_), .B(u2__abc_52138_new_n5018_), .C(u2__abc_52138_new_n15965_), .Y(u2__abc_52138_new_n15966_));
NOR3X1 NOR3X1_295 ( .A(u2__abc_52138_new_n5032_), .B(u2__abc_52138_new_n5025_), .C(u2__abc_52138_new_n15958_), .Y(u2__abc_52138_new_n15974_));
NOR3X1 NOR3X1_296 ( .A(u2__abc_52138_new_n5038_), .B(u2__abc_52138_new_n5032_), .C(u2__abc_52138_new_n15980_), .Y(u2__abc_52138_new_n15981_));
NOR3X1 NOR3X1_297 ( .A(u2__abc_52138_new_n5013_), .B(u2__abc_52138_new_n5933_), .C(u2__abc_52138_new_n15996_), .Y(u2__abc_52138_new_n15997_));
NOR3X1 NOR3X1_298 ( .A(u2__abc_52138_new_n5001_), .B(u2__abc_52138_new_n5013_), .C(u2__abc_52138_new_n15989_), .Y(u2__abc_52138_new_n16005_));
NOR3X1 NOR3X1_299 ( .A(u2__abc_52138_new_n5004_), .B(u2__abc_52138_new_n5001_), .C(u2__abc_52138_new_n16011_), .Y(u2__abc_52138_new_n16012_));
NOR3X1 NOR3X1_3 ( .A(_abc_65734_new_n1505_), .B(_abc_65734_new_n1506_), .C(_abc_65734_new_n1514_), .Y(_abc_65734_new_n1515_));
NOR3X1 NOR3X1_30 ( .A(u2__abc_52138_new_n3123_), .B(u2__abc_52138_new_n3128_), .C(u2__abc_52138_new_n13230_), .Y(u2__abc_52138_new_n13231_));
NOR3X1 NOR3X1_300 ( .A(u2__abc_52138_new_n6171_), .B(u2__abc_52138_new_n6178_), .C(u2__abc_52138_new_n16027_), .Y(u2__abc_52138_new_n16028_));
NOR3X1 NOR3X1_301 ( .A(u2__abc_52138_new_n6162_), .B(u2__abc_52138_new_n6171_), .C(u2__abc_52138_new_n16020_), .Y(u2__abc_52138_new_n16036_));
NOR3X1 NOR3X1_302 ( .A(u2__abc_52138_new_n6165_), .B(u2__abc_52138_new_n6162_), .C(u2__abc_52138_new_n16042_), .Y(u2__abc_52138_new_n16043_));
NOR3X1 NOR3X1_303 ( .A(u2__abc_52138_new_n6147_), .B(u2__abc_52138_new_n6154_), .C(u2__abc_52138_new_n16059_), .Y(u2__abc_52138_new_n16060_));
NOR3X1 NOR3X1_304 ( .A(u2__abc_52138_new_n6138_), .B(u2__abc_52138_new_n6147_), .C(u2__abc_52138_new_n16051_), .Y(u2__abc_52138_new_n16067_));
NOR3X1 NOR3X1_305 ( .A(u2__abc_52138_new_n6143_), .B(u2__abc_52138_new_n6138_), .C(u2__abc_52138_new_n16073_), .Y(u2__abc_52138_new_n16074_));
NOR3X1 NOR3X1_306 ( .A(u2__abc_52138_new_n16086_), .B(u2__abc_52138_new_n16077_), .C(u2__abc_52138_new_n16092_), .Y(u2__abc_52138_new_n16093_));
NOR3X1 NOR3X1_307 ( .A(u2__abc_52138_new_n6282_), .B(u2__abc_52138_new_n16086_), .C(u2__abc_52138_new_n16083_), .Y(u2__abc_52138_new_n16100_));
NOR3X1 NOR3X1_308 ( .A(u2__abc_52138_new_n6285_), .B(u2__abc_52138_new_n6282_), .C(u2__abc_52138_new_n16106_), .Y(u2__abc_52138_new_n16107_));
NOR3X1 NOR3X1_309 ( .A(u2__abc_52138_new_n6315_), .B(u2__abc_52138_new_n16110_), .C(u2__abc_52138_new_n16124_), .Y(u2__abc_52138_new_n16125_));
NOR3X1 NOR3X1_31 ( .A(u2__abc_52138_new_n3112_), .B(u2__abc_52138_new_n3123_), .C(u2__abc_52138_new_n13222_), .Y(u2__abc_52138_new_n13238_));
NOR3X1 NOR3X1_310 ( .A(u2__abc_52138_new_n6306_), .B(u2__abc_52138_new_n6315_), .C(u2__abc_52138_new_n16116_), .Y(u2__abc_52138_new_n16132_));
NOR3X1 NOR3X1_311 ( .A(u2__abc_52138_new_n6311_), .B(u2__abc_52138_new_n6306_), .C(u2__abc_52138_new_n16138_), .Y(u2__abc_52138_new_n16139_));
NOR3X1 NOR3X1_312 ( .A(u2__abc_52138_new_n6237_), .B(u2__abc_52138_new_n6234_), .C(u2__abc_52138_new_n16154_), .Y(u2__abc_52138_new_n16155_));
NOR3X1 NOR3X1_313 ( .A(u2__abc_52138_new_n6245_), .B(u2__abc_52138_new_n6237_), .C(u2__abc_52138_new_n16147_), .Y(u2__abc_52138_new_n16163_));
NOR3X1 NOR3X1_314 ( .A(u2__abc_52138_new_n6248_), .B(u2__abc_52138_new_n6245_), .C(u2__abc_52138_new_n16169_), .Y(u2__abc_52138_new_n16170_));
NOR3X1 NOR3X1_315 ( .A(u2__abc_52138_new_n6266_), .B(u2__abc_52138_new_n6273_), .C(u2__abc_52138_new_n16186_), .Y(u2__abc_52138_new_n16187_));
NOR3X1 NOR3X1_316 ( .A(u2__abc_52138_new_n6257_), .B(u2__abc_52138_new_n6266_), .C(u2__abc_52138_new_n16178_), .Y(u2__abc_52138_new_n16194_));
NOR3X1 NOR3X1_317 ( .A(u2__abc_52138_new_n6262_), .B(u2__abc_52138_new_n6257_), .C(u2__abc_52138_new_n16200_), .Y(u2__abc_52138_new_n16201_));
NOR3X1 NOR3X1_318 ( .A(u2__abc_52138_new_n6196_), .B(u2__abc_52138_new_n6203_), .C(u2__abc_52138_new_n16216_), .Y(u2__abc_52138_new_n16217_));
NOR3X1 NOR3X1_319 ( .A(u2__abc_52138_new_n6187_), .B(u2__abc_52138_new_n6196_), .C(u2__abc_52138_new_n16209_), .Y(u2__abc_52138_new_n16225_));
NOR3X1 NOR3X1_32 ( .A(u2__abc_52138_new_n3117_), .B(u2__abc_52138_new_n3112_), .C(u2__abc_52138_new_n13245_), .Y(u2__abc_52138_new_n13246_));
NOR3X1 NOR3X1_320 ( .A(u2__abc_52138_new_n6190_), .B(u2__abc_52138_new_n6187_), .C(u2__abc_52138_new_n16231_), .Y(u2__abc_52138_new_n16232_));
NOR3X1 NOR3X1_321 ( .A(u2__abc_52138_new_n6219_), .B(u2__abc_52138_new_n6226_), .C(u2__abc_52138_new_n16247_), .Y(u2__abc_52138_new_n16248_));
NOR3X1 NOR3X1_322 ( .A(u2__abc_52138_new_n6210_), .B(u2__abc_52138_new_n6219_), .C(u2__abc_52138_new_n16240_), .Y(u2__abc_52138_new_n16256_));
NOR3X1 NOR3X1_323 ( .A(u2__abc_52138_new_n6215_), .B(u2__abc_52138_new_n6210_), .C(u2__abc_52138_new_n16262_), .Y(u2__abc_52138_new_n16263_));
NOR3X1 NOR3X1_324 ( .A(u2__abc_52138_new_n6120_), .B(u2__abc_52138_new_n6127_), .C(u2__abc_52138_new_n16278_), .Y(u2__abc_52138_new_n16279_));
NOR3X1 NOR3X1_325 ( .A(u2__abc_52138_new_n6108_), .B(u2__abc_52138_new_n6120_), .C(u2__abc_52138_new_n16271_), .Y(u2__abc_52138_new_n16287_));
NOR3X1 NOR3X1_326 ( .A(u2__abc_52138_new_n6115_), .B(u2__abc_52138_new_n6108_), .C(u2__abc_52138_new_n16293_), .Y(u2__abc_52138_new_n16294_));
NOR3X1 NOR3X1_327 ( .A(u2__abc_52138_new_n6096_), .B(u2__abc_52138_new_n6103_), .C(u2__abc_52138_new_n16310_), .Y(u2__abc_52138_new_n16311_));
NOR3X1 NOR3X1_328 ( .A(u2__abc_52138_new_n6084_), .B(u2__abc_52138_new_n6096_), .C(u2__abc_52138_new_n16302_), .Y(u2__abc_52138_new_n16318_));
NOR3X1 NOR3X1_329 ( .A(u2__abc_52138_new_n6089_), .B(u2__abc_52138_new_n6084_), .C(u2__abc_52138_new_n16324_), .Y(u2__abc_52138_new_n16325_));
NOR3X1 NOR3X1_33 ( .A(u2__abc_52138_new_n3146_), .B(u2__abc_52138_new_n3151_), .C(u2__abc_52138_new_n13261_), .Y(u2__abc_52138_new_n13262_));
NOR3X1 NOR3X1_330 ( .A(u2__abc_52138_new_n6052_), .B(u2__abc_52138_new_n6049_), .C(u2__abc_52138_new_n16340_), .Y(u2__abc_52138_new_n16341_));
NOR3X1 NOR3X1_331 ( .A(u2__abc_52138_new_n6036_), .B(u2__abc_52138_new_n6052_), .C(u2__abc_52138_new_n16333_), .Y(u2__abc_52138_new_n16349_));
NOR3X1 NOR3X1_332 ( .A(u2__abc_52138_new_n6043_), .B(u2__abc_52138_new_n6036_), .C(u2__abc_52138_new_n16355_), .Y(u2__abc_52138_new_n16356_));
NOR3X1 NOR3X1_333 ( .A(u2__abc_52138_new_n6070_), .B(u2__abc_52138_new_n6077_), .C(u2__abc_52138_new_n16371_), .Y(u2__abc_52138_new_n16372_));
NOR3X1 NOR3X1_334 ( .A(u2__abc_52138_new_n6058_), .B(u2__abc_52138_new_n6070_), .C(u2__abc_52138_new_n16364_), .Y(u2__abc_52138_new_n16380_));
NOR3X1 NOR3X1_335 ( .A(u2__abc_52138_new_n6063_), .B(u2__abc_52138_new_n6058_), .C(u2__abc_52138_new_n16386_), .Y(u2__abc_52138_new_n16387_));
NOR3X1 NOR3X1_336 ( .A(u2__abc_52138_new_n6015_), .B(u2__abc_52138_new_n6012_), .C(u2__abc_52138_new_n16402_), .Y(u2__abc_52138_new_n16403_));
NOR3X1 NOR3X1_337 ( .A(u2__abc_52138_new_n6023_), .B(u2__abc_52138_new_n6015_), .C(u2__abc_52138_new_n16395_), .Y(u2__abc_52138_new_n16411_));
NOR3X1 NOR3X1_338 ( .A(u2__abc_52138_new_n6026_), .B(u2__abc_52138_new_n6023_), .C(u2__abc_52138_new_n16417_), .Y(u2__abc_52138_new_n16418_));
NOR3X1 NOR3X1_339 ( .A(u2__abc_52138_new_n5998_), .B(u2__abc_52138_new_n6005_), .C(u2__abc_52138_new_n16433_), .Y(u2__abc_52138_new_n16434_));
NOR3X1 NOR3X1_34 ( .A(u2__abc_52138_new_n3135_), .B(u2__abc_52138_new_n3146_), .C(u2__abc_52138_new_n13253_), .Y(u2__abc_52138_new_n13269_));
NOR3X1 NOR3X1_340 ( .A(u2__abc_52138_new_n5989_), .B(u2__abc_52138_new_n5998_), .C(u2__abc_52138_new_n16426_), .Y(u2__abc_52138_new_n16442_));
NOR3X1 NOR3X1_341 ( .A(u2__abc_52138_new_n5994_), .B(u2__abc_52138_new_n5989_), .C(u2__abc_52138_new_n16448_), .Y(u2__abc_52138_new_n16449_));
NOR3X1 NOR3X1_342 ( .A(u2__abc_52138_new_n6414_), .B(u2__abc_52138_new_n5969_), .C(u2__abc_52138_new_n16464_), .Y(u2__abc_52138_new_n16465_));
NOR3X1 NOR3X1_343 ( .A(u2__abc_52138_new_n5976_), .B(u2__abc_52138_new_n6414_), .C(u2__abc_52138_new_n16457_), .Y(u2__abc_52138_new_n16473_));
NOR3X1 NOR3X1_344 ( .A(u2__abc_52138_new_n5979_), .B(u2__abc_52138_new_n5976_), .C(u2__abc_52138_new_n16479_), .Y(u2__abc_52138_new_n16480_));
NOR3X1 NOR3X1_345 ( .A(u2__abc_52138_new_n5955_), .B(u2__abc_52138_new_n5962_), .C(u2__abc_52138_new_n16495_), .Y(u2__abc_52138_new_n16496_));
NOR3X1 NOR3X1_346 ( .A(u2__abc_52138_new_n5946_), .B(u2__abc_52138_new_n5955_), .C(u2__abc_52138_new_n16488_), .Y(u2__abc_52138_new_n16504_));
NOR3X1 NOR3X1_347 ( .A(u2__abc_52138_new_n5949_), .B(u2__abc_52138_new_n5946_), .C(u2__abc_52138_new_n16510_), .Y(u2__abc_52138_new_n16511_));
NOR3X1 NOR3X1_348 ( .A(u2__abc_52138_new_n3005_), .B(u2__abc_52138_new_n3010_), .C(u2__abc_52138_new_n16527_), .Y(u2__abc_52138_new_n16528_));
NOR3X1 NOR3X1_349 ( .A(u2__abc_52138_new_n2997_), .B(u2__abc_52138_new_n3005_), .C(u2__abc_52138_new_n16519_), .Y(u2__abc_52138_new_n16535_));
NOR3X1 NOR3X1_35 ( .A(u2__abc_52138_new_n3142_), .B(u2__abc_52138_new_n3135_), .C(u2__abc_52138_new_n13276_), .Y(u2__abc_52138_new_n13277_));
NOR3X1 NOR3X1_36 ( .A(u2__abc_52138_new_n3394_), .B(u2__abc_52138_new_n3389_), .C(u2__abc_52138_new_n13292_), .Y(u2__abc_52138_new_n13293_));
NOR3X1 NOR3X1_37 ( .A(u2__abc_52138_new_n3437_), .B(u2__abc_52138_new_n3394_), .C(u2__abc_52138_new_n13284_), .Y(u2__abc_52138_new_n13300_));
NOR3X1 NOR3X1_38 ( .A(u2__abc_52138_new_n3383_), .B(u2__abc_52138_new_n3437_), .C(u2__abc_52138_new_n13307_), .Y(u2__abc_52138_new_n13308_));
NOR3X1 NOR3X1_39 ( .A(u2__abc_52138_new_n3412_), .B(u2__abc_52138_new_n13310_), .C(u2__abc_52138_new_n13324_), .Y(u2__abc_52138_new_n13325_));
NOR3X1 NOR3X1_4 ( .A(_abc_65734_new_n1527_), .B(_abc_65734_new_n1538_), .C(_abc_65734_new_n1522_), .Y(_abc_65734_new_n1539_));
NOR3X1 NOR3X1_40 ( .A(u2__abc_52138_new_n3401_), .B(u2__abc_52138_new_n3412_), .C(u2__abc_52138_new_n13316_), .Y(u2__abc_52138_new_n13332_));
NOR3X1 NOR3X1_41 ( .A(u2__abc_52138_new_n3406_), .B(u2__abc_52138_new_n3401_), .C(u2__abc_52138_new_n13339_), .Y(u2__abc_52138_new_n13340_));
NOR3X1 NOR3X1_42 ( .A(u2__abc_52138_new_n3351_), .B(u2__abc_52138_new_n3346_), .C(u2__abc_52138_new_n13355_), .Y(u2__abc_52138_new_n13356_));
NOR3X1 NOR3X1_43 ( .A(u2__abc_52138_new_n3335_), .B(u2__abc_52138_new_n3351_), .C(u2__abc_52138_new_n13347_), .Y(u2__abc_52138_new_n13363_));
NOR3X1 NOR3X1_44 ( .A(u2__abc_52138_new_n3340_), .B(u2__abc_52138_new_n3335_), .C(u2__abc_52138_new_n13370_), .Y(u2__abc_52138_new_n13371_));
NOR3X1 NOR3X1_45 ( .A(u2__abc_52138_new_n3369_), .B(u2__abc_52138_new_n3374_), .C(u2__abc_52138_new_n13386_), .Y(u2__abc_52138_new_n13387_));
NOR3X1 NOR3X1_46 ( .A(u2__abc_52138_new_n3358_), .B(u2__abc_52138_new_n3369_), .C(u2__abc_52138_new_n13378_), .Y(u2__abc_52138_new_n13394_));
NOR3X1 NOR3X1_47 ( .A(u2__abc_52138_new_n3363_), .B(u2__abc_52138_new_n3358_), .C(u2__abc_52138_new_n13401_), .Y(u2__abc_52138_new_n13402_));
NOR3X1 NOR3X1_48 ( .A(u2__abc_52138_new_n3300_), .B(u2__abc_52138_new_n3303_), .C(u2__abc_52138_new_n13417_), .Y(u2__abc_52138_new_n13418_));
NOR3X1 NOR3X1_49 ( .A(u2__abc_52138_new_n3289_), .B(u2__abc_52138_new_n3300_), .C(u2__abc_52138_new_n13409_), .Y(u2__abc_52138_new_n13425_));
NOR3X1 NOR3X1_5 ( .A(_abc_65734_new_n1500_), .B(_abc_65734_new_n1534_), .C(_abc_65734_new_n1492_), .Y(_abc_65734_new_n1548_));
NOR3X1 NOR3X1_50 ( .A(u2__abc_52138_new_n3294_), .B(u2__abc_52138_new_n3289_), .C(u2__abc_52138_new_n13432_), .Y(u2__abc_52138_new_n13433_));
NOR3X1 NOR3X1_51 ( .A(u2__abc_52138_new_n3322_), .B(u2__abc_52138_new_n3327_), .C(u2__abc_52138_new_n13448_), .Y(u2__abc_52138_new_n13449_));
NOR3X1 NOR3X1_52 ( .A(u2__abc_52138_new_n3311_), .B(u2__abc_52138_new_n3322_), .C(u2__abc_52138_new_n13440_), .Y(u2__abc_52138_new_n13456_));
NOR3X1 NOR3X1_53 ( .A(u2__abc_52138_new_n3316_), .B(u2__abc_52138_new_n3311_), .C(u2__abc_52138_new_n13463_), .Y(u2__abc_52138_new_n13464_));
NOR3X1 NOR3X1_54 ( .A(u2__abc_52138_new_n3256_), .B(u2__abc_52138_new_n3251_), .C(u2__abc_52138_new_n13479_), .Y(u2__abc_52138_new_n13480_));
NOR3X1 NOR3X1_55 ( .A(u2__abc_52138_new_n3240_), .B(u2__abc_52138_new_n3256_), .C(u2__abc_52138_new_n13471_), .Y(u2__abc_52138_new_n13487_));
NOR3X1 NOR3X1_56 ( .A(u2__abc_52138_new_n3245_), .B(u2__abc_52138_new_n3240_), .C(u2__abc_52138_new_n13494_), .Y(u2__abc_52138_new_n13495_));
NOR3X1 NOR3X1_57 ( .A(u2__abc_52138_new_n3274_), .B(u2__abc_52138_new_n3279_), .C(u2__abc_52138_new_n13510_), .Y(u2__abc_52138_new_n13511_));
NOR3X1 NOR3X1_58 ( .A(u2__abc_52138_new_n3263_), .B(u2__abc_52138_new_n3274_), .C(u2__abc_52138_new_n13502_), .Y(u2__abc_52138_new_n13518_));
NOR3X1 NOR3X1_59 ( .A(u2__abc_52138_new_n3270_), .B(u2__abc_52138_new_n3263_), .C(u2__abc_52138_new_n13525_), .Y(u2__abc_52138_new_n13526_));
NOR3X1 NOR3X1_6 ( .A(_abc_65734_new_n1533_), .B(_abc_65734_new_n1545_), .C(_abc_65734_new_n1546_), .Y(_abc_65734_new_n1565_));
NOR3X1 NOR3X1_60 ( .A(u2__abc_52138_new_n3837_), .B(u2__abc_52138_new_n3832_), .C(u2__abc_52138_new_n13541_), .Y(u2__abc_52138_new_n13542_));
NOR3X1 NOR3X1_61 ( .A(u2__abc_52138_new_n3843_), .B(u2__abc_52138_new_n3837_), .C(u2__abc_52138_new_n13533_), .Y(u2__abc_52138_new_n13549_));
NOR3X1 NOR3X1_62 ( .A(u2__abc_52138_new_n3848_), .B(u2__abc_52138_new_n3843_), .C(u2__abc_52138_new_n13556_), .Y(u2__abc_52138_new_n13557_));
NOR3X1 NOR3X1_63 ( .A(u2__abc_52138_new_n3881_), .B(u2__abc_52138_new_n3862_), .C(u2__abc_52138_new_n13572_), .Y(u2__abc_52138_new_n13573_));
NOR3X1 NOR3X1_64 ( .A(u2__abc_52138_new_n7264_), .B(u2__abc_52138_new_n3881_), .C(u2__abc_52138_new_n13564_), .Y(u2__abc_52138_new_n13580_));
NOR3X1 NOR3X1_65 ( .A(u2__abc_52138_new_n3856_), .B(u2__abc_52138_new_n7264_), .C(u2__abc_52138_new_n13587_), .Y(u2__abc_52138_new_n13588_));
NOR3X1 NOR3X1_66 ( .A(u2__abc_52138_new_n3793_), .B(u2__abc_52138_new_n3788_), .C(u2__abc_52138_new_n13603_), .Y(u2__abc_52138_new_n13604_));
NOR3X1 NOR3X1_67 ( .A(u2__abc_52138_new_n3797_), .B(u2__abc_52138_new_n3793_), .C(u2__abc_52138_new_n13595_), .Y(u2__abc_52138_new_n13611_));
NOR3X1 NOR3X1_68 ( .A(u2__abc_52138_new_n3802_), .B(u2__abc_52138_new_n3797_), .C(u2__abc_52138_new_n13618_), .Y(u2__abc_52138_new_n13619_));
NOR3X1 NOR3X1_69 ( .A(u2__abc_52138_new_n3821_), .B(u2__abc_52138_new_n3826_), .C(u2__abc_52138_new_n13634_), .Y(u2__abc_52138_new_n13635_));
NOR3X1 NOR3X1_7 ( .A(_abc_65734_new_n1558_), .B(_abc_65734_new_n1559_), .C(_abc_65734_new_n1544_), .Y(_abc_65734_new_n1574_));
NOR3X1 NOR3X1_70 ( .A(u2__abc_52138_new_n3810_), .B(u2__abc_52138_new_n3821_), .C(u2__abc_52138_new_n13626_), .Y(u2__abc_52138_new_n13642_));
NOR3X1 NOR3X1_71 ( .A(u2__abc_52138_new_n3815_), .B(u2__abc_52138_new_n3810_), .C(u2__abc_52138_new_n13649_), .Y(u2__abc_52138_new_n13650_));
NOR3X1 NOR3X1_72 ( .A(u2__abc_52138_new_n3743_), .B(u2__abc_52138_new_n3738_), .C(u2__abc_52138_new_n13664_), .Y(u2__abc_52138_new_n13665_));
NOR3X1 NOR3X1_73 ( .A(u2__abc_52138_new_n3749_), .B(u2__abc_52138_new_n3743_), .C(u2__abc_52138_new_n13657_), .Y(u2__abc_52138_new_n13673_));
NOR3X1 NOR3X1_74 ( .A(u2__abc_52138_new_n3754_), .B(u2__abc_52138_new_n3749_), .C(u2__abc_52138_new_n13680_), .Y(u2__abc_52138_new_n13681_));
NOR3X1 NOR3X1_75 ( .A(u2__abc_52138_new_n3772_), .B(u2__abc_52138_new_n3777_), .C(u2__abc_52138_new_n13696_), .Y(u2__abc_52138_new_n13697_));
NOR3X1 NOR3X1_76 ( .A(u2__abc_52138_new_n3761_), .B(u2__abc_52138_new_n3772_), .C(u2__abc_52138_new_n13688_), .Y(u2__abc_52138_new_n13704_));
NOR3X1 NOR3X1_77 ( .A(u2__abc_52138_new_n3766_), .B(u2__abc_52138_new_n3761_), .C(u2__abc_52138_new_n13711_), .Y(u2__abc_52138_new_n13712_));
NOR3X1 NOR3X1_78 ( .A(u2__abc_52138_new_n3727_), .B(u2__abc_52138_new_n3732_), .C(u2__abc_52138_new_n13726_), .Y(u2__abc_52138_new_n13727_));
NOR3X1 NOR3X1_79 ( .A(u2__abc_52138_new_n3713_), .B(u2__abc_52138_new_n3727_), .C(u2__abc_52138_new_n13719_), .Y(u2__abc_52138_new_n13735_));
NOR3X1 NOR3X1_8 ( .A(u1__abc_51895_new_n344_), .B(u1__abc_51895_new_n359_), .C(u1__abc_51895_new_n374_), .Y(u1__abc_51895_new_n375_));
NOR3X1 NOR3X1_80 ( .A(u2__abc_52138_new_n3718_), .B(u2__abc_52138_new_n3713_), .C(u2__abc_52138_new_n13742_), .Y(u2__abc_52138_new_n13743_));
NOR3X1 NOR3X1_81 ( .A(u2__abc_52138_new_n3702_), .B(u2__abc_52138_new_n3708_), .C(u2__abc_52138_new_n13757_), .Y(u2__abc_52138_new_n13758_));
NOR3X1 NOR3X1_82 ( .A(u2__abc_52138_new_n3691_), .B(u2__abc_52138_new_n3702_), .C(u2__abc_52138_new_n13750_), .Y(u2__abc_52138_new_n13766_));
NOR3X1 NOR3X1_83 ( .A(u2__abc_52138_new_n3696_), .B(u2__abc_52138_new_n3691_), .C(u2__abc_52138_new_n13772_), .Y(u2__abc_52138_new_n13773_));
NOR3X1 NOR3X1_84 ( .A(u2__abc_52138_new_n3653_), .B(u2__abc_52138_new_n3658_), .C(u2__abc_52138_new_n13789_), .Y(u2__abc_52138_new_n13790_));
NOR3X1 NOR3X1_85 ( .A(u2__abc_52138_new_n3644_), .B(u2__abc_52138_new_n3653_), .C(u2__abc_52138_new_n13781_), .Y(u2__abc_52138_new_n13797_));
NOR3X1 NOR3X1_86 ( .A(u2__abc_52138_new_n3649_), .B(u2__abc_52138_new_n3644_), .C(u2__abc_52138_new_n13804_), .Y(u2__abc_52138_new_n13805_));
NOR3X1 NOR3X1_87 ( .A(u2__abc_52138_new_n3676_), .B(u2__abc_52138_new_n3681_), .C(u2__abc_52138_new_n13820_), .Y(u2__abc_52138_new_n13821_));
NOR3X1 NOR3X1_88 ( .A(u2__abc_52138_new_n3665_), .B(u2__abc_52138_new_n3676_), .C(u2__abc_52138_new_n13812_), .Y(u2__abc_52138_new_n13828_));
NOR3X1 NOR3X1_89 ( .A(u2__abc_52138_new_n3670_), .B(u2__abc_52138_new_n3665_), .C(u2__abc_52138_new_n13835_), .Y(u2__abc_52138_new_n13836_));
NOR3X1 NOR3X1_9 ( .A(u2__abc_52138_new_n4355_), .B(u2__abc_52138_new_n4357_), .C(u2__abc_52138_new_n4362_), .Y(u2__abc_52138_new_n4363_));
NOR3X1 NOR3X1_90 ( .A(u2__abc_52138_new_n3608_), .B(u2__abc_52138_new_n3614_), .C(u2__abc_52138_new_n13850_), .Y(u2__abc_52138_new_n13851_));
NOR3X1 NOR3X1_91 ( .A(u2__abc_52138_new_n3597_), .B(u2__abc_52138_new_n3608_), .C(u2__abc_52138_new_n13843_), .Y(u2__abc_52138_new_n13859_));
NOR3X1 NOR3X1_92 ( .A(u2__abc_52138_new_n3602_), .B(u2__abc_52138_new_n3597_), .C(u2__abc_52138_new_n13866_), .Y(u2__abc_52138_new_n13867_));
NOR3X1 NOR3X1_93 ( .A(u2__abc_52138_new_n3630_), .B(u2__abc_52138_new_n3636_), .C(u2__abc_52138_new_n13881_), .Y(u2__abc_52138_new_n13882_));
NOR3X1 NOR3X1_94 ( .A(u2__abc_52138_new_n3619_), .B(u2__abc_52138_new_n3630_), .C(u2__abc_52138_new_n13874_), .Y(u2__abc_52138_new_n13890_));
NOR3X1 NOR3X1_95 ( .A(u2__abc_52138_new_n3624_), .B(u2__abc_52138_new_n3619_), .C(u2__abc_52138_new_n13896_), .Y(u2__abc_52138_new_n13897_));
NOR3X1 NOR3X1_96 ( .A(u2__abc_52138_new_n3555_), .B(u2__abc_52138_new_n3550_), .C(u2__abc_52138_new_n13913_), .Y(u2__abc_52138_new_n13914_));
NOR3X1 NOR3X1_97 ( .A(u2__abc_52138_new_n3561_), .B(u2__abc_52138_new_n3555_), .C(u2__abc_52138_new_n13905_), .Y(u2__abc_52138_new_n13921_));
NOR3X1 NOR3X1_98 ( .A(u2__abc_52138_new_n3566_), .B(u2__abc_52138_new_n3561_), .C(u2__abc_52138_new_n13928_), .Y(u2__abc_52138_new_n13929_));
NOR3X1 NOR3X1_99 ( .A(u2__abc_52138_new_n3583_), .B(u2__abc_52138_new_n3588_), .C(u2__abc_52138_new_n13943_), .Y(u2__abc_52138_new_n13944_));
OAI21X1 OAI21X1_1 ( .A(aNan), .B(_abc_65734_new_n830_), .C(_abc_65734_new_n831_), .Y(\o[112] ));
OAI21X1 OAI21X1_10 ( .A(aNan), .B(_abc_65734_new_n857_), .C(_abc_65734_new_n858_), .Y(\o[121] ));
OAI21X1 OAI21X1_100 ( .A(aNan), .B(_abc_65734_new_n1127_), .C(_abc_65734_new_n1128_), .Y(\o[211] ));
OAI21X1 OAI21X1_1000 ( .A(u2__abc_52138_new_n3655_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7554_));
OAI21X1 OAI21X1_1001 ( .A(u2__abc_52138_new_n7554_), .B(u2__abc_52138_new_n7553_), .C(u2__abc_52138_new_n7555_), .Y(u2__abc_52138_new_n7556_));
OAI21X1 OAI21X1_1002 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_98_), .Y(u2__abc_52138_new_n7558_));
OAI21X1 OAI21X1_1003 ( .A(sqrto_95_), .B(u2__abc_52138_new_n3655_), .C(u2__abc_52138_new_n3659_), .Y(u2__abc_52138_new_n7559_));
OAI21X1 OAI21X1_1004 ( .A(u2__abc_52138_new_n3653_), .B(u2_remHi_95_), .C(u2__abc_52138_new_n7559_), .Y(u2__abc_52138_new_n7560_));
OAI21X1 OAI21X1_1005 ( .A(u2__abc_52138_new_n3663_), .B(u2__abc_52138_new_n7541_), .C(u2__abc_52138_new_n7560_), .Y(u2__abc_52138_new_n7561_));
OAI21X1 OAI21X1_1006 ( .A(u2__abc_52138_new_n3642_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7564_));
OAI21X1 OAI21X1_1007 ( .A(u2__abc_52138_new_n7564_), .B(u2__abc_52138_new_n7563_), .C(u2__abc_52138_new_n7565_), .Y(u2__abc_52138_new_n7566_));
OAI21X1 OAI21X1_1008 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_99_), .Y(u2__abc_52138_new_n7568_));
OAI21X1 OAI21X1_1009 ( .A(u2__abc_52138_new_n3647_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7574_));
OAI21X1 OAI21X1_101 ( .A(aNan), .B(_abc_65734_new_n1130_), .C(_abc_65734_new_n1131_), .Y(\o[212] ));
OAI21X1 OAI21X1_1010 ( .A(u2__abc_52138_new_n7574_), .B(u2__abc_52138_new_n7573_), .C(u2__abc_52138_new_n7575_), .Y(u2__abc_52138_new_n7576_));
OAI21X1 OAI21X1_1011 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_100_), .Y(u2__abc_52138_new_n7578_));
OAI21X1 OAI21X1_1012 ( .A(u2__abc_52138_new_n7580_), .B(u2__abc_52138_new_n3650_), .C(u2__abc_52138_new_n7569_), .Y(u2__abc_52138_new_n7581_));
OAI21X1 OAI21X1_1013 ( .A(u2__abc_52138_new_n7560_), .B(u2__abc_52138_new_n3652_), .C(u2__abc_52138_new_n7582_), .Y(u2__abc_52138_new_n7583_));
OAI21X1 OAI21X1_1014 ( .A(u2__abc_52138_new_n7539_), .B(u2__abc_52138_new_n7540_), .C(u2__abc_52138_new_n3664_), .Y(u2__abc_52138_new_n7585_));
OAI21X1 OAI21X1_1015 ( .A(u2__abc_52138_new_n7589_), .B(u2__abc_52138_new_n7588_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7590_));
OAI21X1 OAI21X1_1016 ( .A(u2_remHi_98_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7590_), .Y(u2__abc_52138_new_n7591_));
OAI21X1 OAI21X1_1017 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_101_), .Y(u2__abc_52138_new_n7596_));
OAI21X1 OAI21X1_1018 ( .A(sqrto_98_), .B(u2__abc_52138_new_n3683_), .C(u2__abc_52138_new_n7587_), .Y(u2__abc_52138_new_n7597_));
OAI21X1 OAI21X1_1019 ( .A(u2__abc_52138_new_n3678_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7600_));
OAI21X1 OAI21X1_102 ( .A(aNan), .B(_abc_65734_new_n1133_), .C(_abc_65734_new_n1134_), .Y(\o[213] ));
OAI21X1 OAI21X1_1020 ( .A(u2__abc_52138_new_n7600_), .B(u2__abc_52138_new_n7599_), .C(u2__abc_52138_new_n7601_), .Y(u2__abc_52138_new_n7602_));
OAI21X1 OAI21X1_1021 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_102_), .Y(u2__abc_52138_new_n7604_));
OAI21X1 OAI21X1_1022 ( .A(sqrto_98_), .B(u2__abc_52138_new_n3683_), .C(u2__abc_52138_new_n3677_), .Y(u2__abc_52138_new_n7605_));
OAI21X1 OAI21X1_1023 ( .A(u2__abc_52138_new_n7605_), .B(u2__abc_52138_new_n7588_), .C(u2__abc_52138_new_n3679_), .Y(u2__abc_52138_new_n7606_));
OAI21X1 OAI21X1_1024 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7608_), .Y(u2__abc_52138_new_n7609_));
OAI21X1 OAI21X1_1025 ( .A(u2__abc_52138_new_n3667_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7611_));
OAI21X1 OAI21X1_1026 ( .A(u2__abc_52138_new_n7611_), .B(u2__abc_52138_new_n7610_), .C(u2__abc_52138_new_n7612_), .Y(u2__abc_52138_new_n7613_));
OAI21X1 OAI21X1_1027 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_103_), .Y(u2__abc_52138_new_n7615_));
OAI21X1 OAI21X1_1028 ( .A(u2__abc_52138_new_n3951_), .B(u2__abc_52138_new_n7606_), .C(u2__abc_52138_new_n3666_), .Y(u2__abc_52138_new_n7617_));
OAI21X1 OAI21X1_1029 ( .A(u2__abc_52138_new_n7616_), .B(u2__abc_52138_new_n7617_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7618_));
OAI21X1 OAI21X1_103 ( .A(aNan), .B(_abc_65734_new_n1136_), .C(_abc_65734_new_n1137_), .Y(\o[214] ));
OAI21X1 OAI21X1_1030 ( .A(u2__abc_52138_new_n3672_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7620_));
OAI21X1 OAI21X1_1031 ( .A(u2__abc_52138_new_n7620_), .B(u2__abc_52138_new_n7619_), .C(u2__abc_52138_new_n7621_), .Y(u2__abc_52138_new_n7622_));
OAI21X1 OAI21X1_1032 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_104_), .Y(u2__abc_52138_new_n7624_));
OAI21X1 OAI21X1_1033 ( .A(u2__abc_52138_new_n3666_), .B(u2__abc_52138_new_n3952_), .C(u2__abc_52138_new_n3671_), .Y(u2__abc_52138_new_n7627_));
OAI21X1 OAI21X1_1034 ( .A(u2__abc_52138_new_n7625_), .B(u2__abc_52138_new_n7584_), .C(u2__abc_52138_new_n7628_), .Y(u2__abc_52138_new_n7629_));
OAI21X1 OAI21X1_1035 ( .A(u2__abc_52138_new_n3688_), .B(u2__abc_52138_new_n7541_), .C(u2__abc_52138_new_n7630_), .Y(u2__abc_52138_new_n7631_));
OAI21X1 OAI21X1_1036 ( .A(u2__abc_52138_new_n7634_), .B(u2__abc_52138_new_n7633_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7635_));
OAI21X1 OAI21X1_1037 ( .A(u2_remHi_102_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7635_), .Y(u2__abc_52138_new_n7636_));
OAI21X1 OAI21X1_1038 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_105_), .Y(u2__abc_52138_new_n7641_));
OAI21X1 OAI21X1_1039 ( .A(sqrto_102_), .B(u2__abc_52138_new_n3612_), .C(u2__abc_52138_new_n7632_), .Y(u2__abc_52138_new_n7643_));
OAI21X1 OAI21X1_104 ( .A(aNan), .B(_abc_65734_new_n1139_), .C(_abc_65734_new_n1140_), .Y(\o[215] ));
OAI21X1 OAI21X1_1040 ( .A(u2__abc_52138_new_n3610_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7646_));
OAI21X1 OAI21X1_1041 ( .A(u2__abc_52138_new_n7646_), .B(u2__abc_52138_new_n7645_), .C(u2__abc_52138_new_n7647_), .Y(u2__abc_52138_new_n7648_));
OAI21X1 OAI21X1_1042 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_106_), .Y(u2__abc_52138_new_n7650_));
OAI21X1 OAI21X1_1043 ( .A(sqrto_102_), .B(u2__abc_52138_new_n3612_), .C(u2__abc_52138_new_n3609_), .Y(u2__abc_52138_new_n7651_));
OAI21X1 OAI21X1_1044 ( .A(u2__abc_52138_new_n7651_), .B(u2__abc_52138_new_n7633_), .C(u2__abc_52138_new_n3611_), .Y(u2__abc_52138_new_n7652_));
OAI21X1 OAI21X1_1045 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7654_), .Y(u2__abc_52138_new_n7655_));
OAI21X1 OAI21X1_1046 ( .A(u2__abc_52138_new_n3599_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7657_));
OAI21X1 OAI21X1_1047 ( .A(u2__abc_52138_new_n7657_), .B(u2__abc_52138_new_n7656_), .C(u2__abc_52138_new_n7658_), .Y(u2__abc_52138_new_n7659_));
OAI21X1 OAI21X1_1048 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_107_), .Y(u2__abc_52138_new_n7661_));
OAI21X1 OAI21X1_1049 ( .A(u2__abc_52138_new_n3601_), .B(u2__abc_52138_new_n7652_), .C(u2__abc_52138_new_n3598_), .Y(u2__abc_52138_new_n7662_));
OAI21X1 OAI21X1_105 ( .A(aNan), .B(_abc_65734_new_n1142_), .C(_abc_65734_new_n1143_), .Y(\o[216] ));
OAI21X1 OAI21X1_1050 ( .A(u2__abc_52138_new_n3604_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7665_));
OAI21X1 OAI21X1_1051 ( .A(u2__abc_52138_new_n7665_), .B(u2__abc_52138_new_n7664_), .C(u2__abc_52138_new_n7666_), .Y(u2__abc_52138_new_n7667_));
OAI21X1 OAI21X1_1052 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_108_), .Y(u2__abc_52138_new_n7669_));
OAI21X1 OAI21X1_1053 ( .A(u2__abc_52138_new_n3608_), .B(u2_remHi_103_), .C(u2__abc_52138_new_n7651_), .Y(u2__abc_52138_new_n7670_));
OAI21X1 OAI21X1_1054 ( .A(u2__abc_52138_new_n7670_), .B(u2__abc_52138_new_n3607_), .C(u2__abc_52138_new_n7672_), .Y(u2__abc_52138_new_n7673_));
OAI21X1 OAI21X1_1055 ( .A(u2__abc_52138_new_n7673_), .B(u2__abc_52138_new_n7674_), .C(u2__abc_52138_new_n3638_), .Y(u2__abc_52138_new_n7675_));
OAI21X1 OAI21X1_1056 ( .A(u2__abc_52138_new_n3635_), .B(u2__abc_52138_new_n3637_), .C(u2__abc_52138_new_n7676_), .Y(u2__abc_52138_new_n7677_));
OAI21X1 OAI21X1_1057 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7679_), .C(u2__abc_52138_new_n7680_), .Y(u2__abc_52138_new_n7681_));
OAI21X1 OAI21X1_1058 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_109_), .Y(u2__abc_52138_new_n7683_));
OAI21X1 OAI21X1_1059 ( .A(sqrto_106_), .B(u2__abc_52138_new_n3634_), .C(u2__abc_52138_new_n7675_), .Y(u2__abc_52138_new_n7685_));
OAI21X1 OAI21X1_106 ( .A(aNan), .B(_abc_65734_new_n1145_), .C(_abc_65734_new_n1146_), .Y(\o[217] ));
OAI21X1 OAI21X1_1060 ( .A(u2__abc_52138_new_n3632_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7688_));
OAI21X1 OAI21X1_1061 ( .A(u2__abc_52138_new_n7688_), .B(u2__abc_52138_new_n7687_), .C(u2__abc_52138_new_n7689_), .Y(u2__abc_52138_new_n7690_));
OAI21X1 OAI21X1_1062 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_110_), .Y(u2__abc_52138_new_n7692_));
OAI21X1 OAI21X1_1063 ( .A(sqrto_106_), .B(u2__abc_52138_new_n3634_), .C(u2__abc_52138_new_n3631_), .Y(u2__abc_52138_new_n7693_));
OAI21X1 OAI21X1_1064 ( .A(u2__abc_52138_new_n3630_), .B(u2_remHi_107_), .C(u2__abc_52138_new_n7693_), .Y(u2__abc_52138_new_n7694_));
OAI21X1 OAI21X1_1065 ( .A(u2__abc_52138_new_n3639_), .B(u2__abc_52138_new_n7676_), .C(u2__abc_52138_new_n7694_), .Y(u2__abc_52138_new_n7695_));
OAI21X1 OAI21X1_1066 ( .A(u2__abc_52138_new_n3621_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7698_));
OAI21X1 OAI21X1_1067 ( .A(u2__abc_52138_new_n7698_), .B(u2__abc_52138_new_n7697_), .C(u2__abc_52138_new_n7699_), .Y(u2__abc_52138_new_n7700_));
OAI21X1 OAI21X1_1068 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_111_), .Y(u2__abc_52138_new_n7702_));
OAI21X1 OAI21X1_1069 ( .A(u2__abc_52138_new_n3623_), .B(u2__abc_52138_new_n7705_), .C(u2__abc_52138_new_n3620_), .Y(u2__abc_52138_new_n7706_));
OAI21X1 OAI21X1_107 ( .A(aNan), .B(_abc_65734_new_n1148_), .C(_abc_65734_new_n1149_), .Y(\o[218] ));
OAI21X1 OAI21X1_1070 ( .A(u2__abc_52138_new_n7704_), .B(u2__abc_52138_new_n7706_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7707_));
OAI21X1 OAI21X1_1071 ( .A(u2__abc_52138_new_n3626_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7709_));
OAI21X1 OAI21X1_1072 ( .A(u2__abc_52138_new_n7709_), .B(u2__abc_52138_new_n7708_), .C(u2__abc_52138_new_n7710_), .Y(u2__abc_52138_new_n7711_));
OAI21X1 OAI21X1_1073 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_112_), .Y(u2__abc_52138_new_n7713_));
OAI21X1 OAI21X1_1074 ( .A(u2__abc_52138_new_n7694_), .B(u2__abc_52138_new_n3629_), .C(u2__abc_52138_new_n3625_), .Y(u2__abc_52138_new_n7716_));
OAI21X1 OAI21X1_1075 ( .A(u2__abc_52138_new_n3620_), .B(u2__abc_52138_new_n7703_), .C(u2__abc_52138_new_n7717_), .Y(u2__abc_52138_new_n7718_));
OAI21X1 OAI21X1_1076 ( .A(u2__abc_52138_new_n7539_), .B(u2__abc_52138_new_n7540_), .C(u2__abc_52138_new_n3689_), .Y(u2__abc_52138_new_n7720_));
OAI21X1 OAI21X1_1077 ( .A(u2__abc_52138_new_n3552_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7724_));
OAI21X1 OAI21X1_1078 ( .A(u2__abc_52138_new_n7724_), .B(u2__abc_52138_new_n7723_), .C(u2__abc_52138_new_n7725_), .Y(u2__abc_52138_new_n7726_));
OAI21X1 OAI21X1_1079 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_113_), .Y(u2__abc_52138_new_n7728_));
OAI21X1 OAI21X1_108 ( .A(aNan), .B(_abc_65734_new_n1151_), .C(_abc_65734_new_n1152_), .Y(\o[219] ));
OAI21X1 OAI21X1_1080 ( .A(u2__abc_52138_new_n3972_), .B(u2__abc_52138_new_n7729_), .C(u2__abc_52138_new_n3551_), .Y(u2__abc_52138_new_n7730_));
OAI21X1 OAI21X1_1081 ( .A(u2__abc_52138_new_n3557_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7733_));
OAI21X1 OAI21X1_1082 ( .A(u2__abc_52138_new_n7733_), .B(u2__abc_52138_new_n7732_), .C(u2__abc_52138_new_n7734_), .Y(u2__abc_52138_new_n7735_));
OAI21X1 OAI21X1_1083 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_114_), .Y(u2__abc_52138_new_n7737_));
OAI21X1 OAI21X1_1084 ( .A(u2__abc_52138_new_n3551_), .B(u2__abc_52138_new_n3973_), .C(u2__abc_52138_new_n3556_), .Y(u2__abc_52138_new_n7738_));
OAI21X1 OAI21X1_1085 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7741_), .Y(u2__abc_52138_new_n7742_));
OAI21X1 OAI21X1_1086 ( .A(u2__abc_52138_new_n3563_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7744_));
OAI21X1 OAI21X1_1087 ( .A(u2__abc_52138_new_n7744_), .B(u2__abc_52138_new_n7743_), .C(u2__abc_52138_new_n7745_), .Y(u2__abc_52138_new_n7746_));
OAI21X1 OAI21X1_1088 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_115_), .Y(u2__abc_52138_new_n7748_));
OAI21X1 OAI21X1_1089 ( .A(u2__abc_52138_new_n3565_), .B(u2__abc_52138_new_n7739_), .C(u2__abc_52138_new_n3562_), .Y(u2__abc_52138_new_n7749_));
OAI21X1 OAI21X1_109 ( .A(aNan), .B(_abc_65734_new_n1154_), .C(_abc_65734_new_n1155_), .Y(\o[220] ));
OAI21X1 OAI21X1_1090 ( .A(u2__abc_52138_new_n3568_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7752_));
OAI21X1 OAI21X1_1091 ( .A(u2__abc_52138_new_n7752_), .B(u2__abc_52138_new_n7751_), .C(u2__abc_52138_new_n7753_), .Y(u2__abc_52138_new_n7754_));
OAI21X1 OAI21X1_1092 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_116_), .Y(u2__abc_52138_new_n7756_));
OAI21X1 OAI21X1_1093 ( .A(u2__abc_52138_new_n7757_), .B(u2__abc_52138_new_n3971_), .C(u2__abc_52138_new_n7759_), .Y(u2__abc_52138_new_n7760_));
OAI21X1 OAI21X1_1094 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7763_), .Y(u2__abc_52138_new_n7764_));
OAI21X1 OAI21X1_1095 ( .A(u2__abc_52138_new_n3590_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7766_));
OAI21X1 OAI21X1_1096 ( .A(u2__abc_52138_new_n7766_), .B(u2__abc_52138_new_n7765_), .C(u2__abc_52138_new_n7767_), .Y(u2__abc_52138_new_n7768_));
OAI21X1 OAI21X1_1097 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_117_), .Y(u2__abc_52138_new_n7770_));
OAI21X1 OAI21X1_1098 ( .A(u2__abc_52138_new_n3592_), .B(u2__abc_52138_new_n7761_), .C(u2__abc_52138_new_n3589_), .Y(u2__abc_52138_new_n7772_));
OAI21X1 OAI21X1_1099 ( .A(u2__abc_52138_new_n7771_), .B(u2__abc_52138_new_n7772_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7773_));
OAI21X1 OAI21X1_11 ( .A(aNan), .B(_abc_65734_new_n860_), .C(_abc_65734_new_n861_), .Y(\o[122] ));
OAI21X1 OAI21X1_110 ( .A(aNan), .B(_abc_65734_new_n1157_), .C(_abc_65734_new_n1158_), .Y(\o[221] ));
OAI21X1 OAI21X1_1100 ( .A(u2__abc_52138_new_n3585_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7775_));
OAI21X1 OAI21X1_1101 ( .A(u2__abc_52138_new_n7775_), .B(u2__abc_52138_new_n7774_), .C(u2__abc_52138_new_n7776_), .Y(u2__abc_52138_new_n7777_));
OAI21X1 OAI21X1_1102 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_118_), .Y(u2__abc_52138_new_n7780_));
OAI21X1 OAI21X1_1103 ( .A(sqrto_115_), .B(u2__abc_52138_new_n3585_), .C(u2__abc_52138_new_n7781_), .Y(u2__abc_52138_new_n7782_));
OAI21X1 OAI21X1_1104 ( .A(u2__abc_52138_new_n3573_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7786_));
OAI21X1 OAI21X1_1105 ( .A(u2_remHi_118_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n7788_));
OAI21X1 OAI21X1_1106 ( .A(u2__abc_52138_new_n7788_), .B(u2__abc_52138_new_n7787_), .C(u2__abc_52138_new_n7780_), .Y(u2__abc_52138_new_n7789_));
OAI21X1 OAI21X1_1107 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_119_), .Y(u2__abc_52138_new_n7791_));
OAI21X1 OAI21X1_1108 ( .A(sqrto_116_), .B(u2__abc_52138_new_n3573_), .C(u2__abc_52138_new_n7783_), .Y(u2__abc_52138_new_n7793_));
OAI21X1 OAI21X1_1109 ( .A(u2__abc_52138_new_n3580_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7796_));
OAI21X1 OAI21X1_111 ( .A(aNan), .B(_abc_65734_new_n1160_), .C(_abc_65734_new_n1161_), .Y(\o[222] ));
OAI21X1 OAI21X1_1110 ( .A(u2__abc_52138_new_n7796_), .B(u2__abc_52138_new_n7795_), .C(u2__abc_52138_new_n7797_), .Y(u2__abc_52138_new_n7798_));
OAI21X1 OAI21X1_1111 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_120_), .Y(u2__abc_52138_new_n7800_));
OAI21X1 OAI21X1_1112 ( .A(u2__abc_52138_new_n3589_), .B(u2__abc_52138_new_n3587_), .C(u2__abc_52138_new_n3584_), .Y(u2__abc_52138_new_n7804_));
OAI21X1 OAI21X1_1113 ( .A(u2__abc_52138_new_n3578_), .B(u2_remHi_117_), .C(u2__abc_52138_new_n3574_), .Y(u2__abc_52138_new_n7806_));
OAI21X1 OAI21X1_1114 ( .A(u2__abc_52138_new_n3503_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7814_));
OAI21X1 OAI21X1_1115 ( .A(u2__abc_52138_new_n7814_), .B(u2__abc_52138_new_n7813_), .C(u2__abc_52138_new_n7815_), .Y(u2__abc_52138_new_n7816_));
OAI21X1 OAI21X1_1116 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_121_), .Y(u2__abc_52138_new_n7818_));
OAI21X1 OAI21X1_1117 ( .A(u2__abc_52138_new_n3507_), .B(u2__abc_52138_new_n7810_), .C(u2__abc_52138_new_n3505_), .Y(u2__abc_52138_new_n7820_));
OAI21X1 OAI21X1_1118 ( .A(u2__abc_52138_new_n7819_), .B(u2__abc_52138_new_n7820_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7821_));
OAI21X1 OAI21X1_1119 ( .A(u2__abc_52138_new_n3508_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7823_));
OAI21X1 OAI21X1_112 ( .A(aNan), .B(_abc_65734_new_n1163_), .C(_abc_65734_new_n1164_), .Y(\o[223] ));
OAI21X1 OAI21X1_1120 ( .A(u2__abc_52138_new_n7823_), .B(u2__abc_52138_new_n7822_), .C(u2__abc_52138_new_n7824_), .Y(u2__abc_52138_new_n7825_));
OAI21X1 OAI21X1_1121 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_122_), .Y(u2__abc_52138_new_n7827_));
OAI21X1 OAI21X1_1122 ( .A(u2__abc_52138_new_n3512_), .B(u2__abc_52138_new_n3505_), .C(u2__abc_52138_new_n3510_), .Y(u2__abc_52138_new_n7829_));
OAI21X1 OAI21X1_1123 ( .A(u2__abc_52138_new_n7808_), .B(u2__abc_52138_new_n7809_), .C(u2__abc_52138_new_n3515_), .Y(u2__abc_52138_new_n7831_));
OAI21X1 OAI21X1_1124 ( .A(u2__abc_52138_new_n7828_), .B(u2__abc_52138_new_n7832_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7833_));
OAI21X1 OAI21X1_1125 ( .A(u2__abc_52138_new_n3518_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7835_));
OAI21X1 OAI21X1_1126 ( .A(u2__abc_52138_new_n7835_), .B(u2__abc_52138_new_n7834_), .C(u2__abc_52138_new_n7836_), .Y(u2__abc_52138_new_n7837_));
OAI21X1 OAI21X1_1127 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_123_), .Y(u2__abc_52138_new_n7839_));
OAI21X1 OAI21X1_1128 ( .A(sqrto_120_), .B(u2__abc_52138_new_n3518_), .C(u2__abc_52138_new_n7840_), .Y(u2__abc_52138_new_n7841_));
OAI21X1 OAI21X1_1129 ( .A(u2__abc_52138_new_n3523_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7844_));
OAI21X1 OAI21X1_113 ( .A(\a[112] ), .B(_abc_65734_new_n1169_), .C(_abc_65734_new_n1171_), .Y(fracta1_1_));
OAI21X1 OAI21X1_1130 ( .A(u2__abc_52138_new_n7844_), .B(u2__abc_52138_new_n7843_), .C(u2__abc_52138_new_n7845_), .Y(u2__abc_52138_new_n7846_));
OAI21X1 OAI21X1_1131 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_124_), .Y(u2__abc_52138_new_n7848_));
OAI21X1 OAI21X1_1132 ( .A(u2__abc_52138_new_n3517_), .B(u2__abc_52138_new_n3525_), .C(u2__abc_52138_new_n3522_), .Y(u2__abc_52138_new_n7849_));
OAI21X1 OAI21X1_1133 ( .A(u2__abc_52138_new_n6487_), .B(u2__abc_52138_new_n7810_), .C(u2__abc_52138_new_n7850_), .Y(u2__abc_52138_new_n7851_));
OAI21X1 OAI21X1_1134 ( .A(u2__abc_52138_new_n3546_), .B(u2__abc_52138_new_n7851_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7854_));
OAI21X1 OAI21X1_1135 ( .A(u2__abc_52138_new_n3542_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7856_));
OAI21X1 OAI21X1_1136 ( .A(u2_remHi_124_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n7858_));
OAI21X1 OAI21X1_1137 ( .A(u2__abc_52138_new_n7858_), .B(u2__abc_52138_new_n7857_), .C(u2__abc_52138_new_n7848_), .Y(u2__abc_52138_new_n7859_));
OAI21X1 OAI21X1_1138 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_125_), .Y(u2__abc_52138_new_n7861_));
OAI21X1 OAI21X1_1139 ( .A(sqrto_122_), .B(u2__abc_52138_new_n3542_), .C(u2__abc_52138_new_n7852_), .Y(u2__abc_52138_new_n7863_));
OAI21X1 OAI21X1_114 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1173_), .C(_abc_65734_new_n1174_), .Y(fracta1_2_));
OAI21X1 OAI21X1_1140 ( .A(u2__abc_52138_new_n3540_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7866_));
OAI21X1 OAI21X1_1141 ( .A(u2__abc_52138_new_n7866_), .B(u2__abc_52138_new_n7865_), .C(u2__abc_52138_new_n7867_), .Y(u2__abc_52138_new_n7868_));
OAI21X1 OAI21X1_1142 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_126_), .Y(u2__abc_52138_new_n7870_));
OAI21X1 OAI21X1_1143 ( .A(sqrto_122_), .B(u2__abc_52138_new_n3542_), .C(u2__abc_52138_new_n3539_), .Y(u2__abc_52138_new_n7871_));
OAI21X1 OAI21X1_1144 ( .A(u2__abc_52138_new_n7871_), .B(u2__abc_52138_new_n7853_), .C(u2__abc_52138_new_n3541_), .Y(u2__abc_52138_new_n7872_));
OAI21X1 OAI21X1_1145 ( .A(u2__abc_52138_new_n3529_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7875_));
OAI21X1 OAI21X1_1146 ( .A(u2__abc_52138_new_n7875_), .B(u2__abc_52138_new_n7874_), .C(u2__abc_52138_new_n7876_), .Y(u2__abc_52138_new_n7877_));
OAI21X1 OAI21X1_1147 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_127_), .Y(u2__abc_52138_new_n7879_));
OAI21X1 OAI21X1_1148 ( .A(u2__abc_52138_new_n3531_), .B(u2__abc_52138_new_n7872_), .C(u2__abc_52138_new_n3528_), .Y(u2__abc_52138_new_n7880_));
OAI21X1 OAI21X1_1149 ( .A(u2__abc_52138_new_n3532_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7883_));
OAI21X1 OAI21X1_115 ( .A(\a[112] ), .B(_abc_65734_new_n1173_), .C(_abc_65734_new_n1176_), .Y(fracta1_3_));
OAI21X1 OAI21X1_1150 ( .A(u2__abc_52138_new_n7883_), .B(u2__abc_52138_new_n7882_), .C(u2__abc_52138_new_n7884_), .Y(u2__abc_52138_new_n7885_));
OAI21X1 OAI21X1_1151 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_128_), .Y(u2__abc_52138_new_n7887_));
OAI21X1 OAI21X1_1152 ( .A(u2__abc_52138_new_n7890_), .B(u2__abc_52138_new_n3992_), .C(u2__abc_52138_new_n3533_), .Y(u2__abc_52138_new_n7891_));
OAI21X1 OAI21X1_1153 ( .A(u2__abc_52138_new_n3538_), .B(u2_remHi_123_), .C(u2__abc_52138_new_n7871_), .Y(u2__abc_52138_new_n7894_));
OAI21X1 OAI21X1_1154 ( .A(u2__abc_52138_new_n7893_), .B(u2__abc_52138_new_n7719_), .C(u2__abc_52138_new_n7896_), .Y(u2__abc_52138_new_n7897_));
OAI21X1 OAI21X1_1155 ( .A(u2__abc_52138_new_n7899_), .B(u2__abc_52138_new_n7889_), .C(u2__abc_52138_new_n4718_), .Y(u2__abc_52138_new_n7900_));
OAI21X1 OAI21X1_1156 ( .A(u2__abc_52138_new_n4715_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7903_), .Y(u2__abc_52138_new_n7904_));
OAI21X1 OAI21X1_1157 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7904_), .C(u2__abc_52138_new_n7906_), .Y(u2__abc_52138_new_n7907_));
OAI21X1 OAI21X1_1158 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_129_), .Y(u2__abc_52138_new_n7909_));
OAI21X1 OAI21X1_1159 ( .A(sqrto_126_), .B(u2__abc_52138_new_n4715_), .C(u2__abc_52138_new_n7900_), .Y(u2__abc_52138_new_n7910_));
OAI21X1 OAI21X1_116 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1178_), .C(_abc_65734_new_n1179_), .Y(fracta1_4_));
OAI21X1 OAI21X1_1160 ( .A(u2__abc_52138_new_n4724_), .B(u2__abc_52138_new_n7910_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7911_));
OAI21X1 OAI21X1_1161 ( .A(u2__abc_52138_new_n4721_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7913_));
OAI21X1 OAI21X1_1162 ( .A(u2__abc_52138_new_n7913_), .B(u2__abc_52138_new_n7912_), .C(u2__abc_52138_new_n7914_), .Y(u2__abc_52138_new_n7915_));
OAI21X1 OAI21X1_1163 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_130_), .Y(u2__abc_52138_new_n7917_));
OAI21X1 OAI21X1_1164 ( .A(u2__abc_52138_new_n4714_), .B(u2__abc_52138_new_n4768_), .C(u2__abc_52138_new_n4720_), .Y(u2__abc_52138_new_n7918_));
OAI21X1 OAI21X1_1165 ( .A(u2__abc_52138_new_n4725_), .B(u2__abc_52138_new_n7901_), .C(u2__abc_52138_new_n7919_), .Y(u2__abc_52138_new_n7920_));
OAI21X1 OAI21X1_1166 ( .A(u2__abc_52138_new_n7905_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7923_));
OAI21X1 OAI21X1_1167 ( .A(u2__abc_52138_new_n7923_), .B(u2__abc_52138_new_n7922_), .C(u2__abc_52138_new_n7924_), .Y(u2__abc_52138_new_n7925_));
OAI21X1 OAI21X1_1168 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_131_), .Y(u2__abc_52138_new_n7927_));
OAI21X1 OAI21X1_1169 ( .A(sqrto_128_), .B(u2__abc_52138_new_n7905_), .C(u2__abc_52138_new_n7929_), .Y(u2__abc_52138_new_n7930_));
OAI21X1 OAI21X1_117 ( .A(\a[112] ), .B(_abc_65734_new_n1178_), .C(_abc_65734_new_n1181_), .Y(fracta1_5_));
OAI21X1 OAI21X1_1170 ( .A(u2__abc_52138_new_n4729_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7933_));
OAI21X1 OAI21X1_1171 ( .A(u2__abc_52138_new_n7933_), .B(u2__abc_52138_new_n7932_), .C(u2__abc_52138_new_n7934_), .Y(u2__abc_52138_new_n7935_));
OAI21X1 OAI21X1_1172 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_132_), .Y(u2__abc_52138_new_n7937_));
OAI21X1 OAI21X1_1173 ( .A(u2__abc_52138_new_n7940_), .B(u2__abc_52138_new_n4772_), .C(u2__abc_52138_new_n4728_), .Y(u2__abc_52138_new_n7941_));
OAI21X1 OAI21X1_1174 ( .A(u2__abc_52138_new_n4732_), .B(u2__abc_52138_new_n7901_), .C(u2__abc_52138_new_n7942_), .Y(u2__abc_52138_new_n7943_));
OAI21X1 OAI21X1_1175 ( .A(u2__abc_52138_new_n7946_), .B(u2__abc_52138_new_n7945_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7947_));
OAI21X1 OAI21X1_1176 ( .A(u2_remHi_130_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7947_), .Y(u2__abc_52138_new_n7948_));
OAI21X1 OAI21X1_1177 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_133_), .Y(u2__abc_52138_new_n7953_));
OAI21X1 OAI21X1_1178 ( .A(sqrto_130_), .B(u2__abc_52138_new_n4776_), .C(u2__abc_52138_new_n7944_), .Y(u2__abc_52138_new_n7954_));
OAI21X1 OAI21X1_1179 ( .A(u2__abc_52138_new_n4746_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7957_));
OAI21X1 OAI21X1_118 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1183_), .C(_abc_65734_new_n1184_), .Y(fracta1_6_));
OAI21X1 OAI21X1_1180 ( .A(u2__abc_52138_new_n7957_), .B(u2__abc_52138_new_n7956_), .C(u2__abc_52138_new_n7958_), .Y(u2__abc_52138_new_n7959_));
OAI21X1 OAI21X1_1181 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_134_), .Y(u2__abc_52138_new_n7961_));
OAI21X1 OAI21X1_1182 ( .A(sqrto_130_), .B(u2__abc_52138_new_n4776_), .C(u2__abc_52138_new_n4745_), .Y(u2__abc_52138_new_n7962_));
OAI21X1 OAI21X1_1183 ( .A(u2__abc_52138_new_n7962_), .B(u2__abc_52138_new_n7945_), .C(u2__abc_52138_new_n4747_), .Y(u2__abc_52138_new_n7963_));
OAI21X1 OAI21X1_1184 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7965_), .Y(u2__abc_52138_new_n7966_));
OAI21X1 OAI21X1_1185 ( .A(u2__abc_52138_new_n4735_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7968_));
OAI21X1 OAI21X1_1186 ( .A(u2__abc_52138_new_n7968_), .B(u2__abc_52138_new_n7967_), .C(u2__abc_52138_new_n7969_), .Y(u2__abc_52138_new_n7970_));
OAI21X1 OAI21X1_1187 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_135_), .Y(u2__abc_52138_new_n7972_));
OAI21X1 OAI21X1_1188 ( .A(u2__abc_52138_new_n4737_), .B(u2__abc_52138_new_n7963_), .C(u2__abc_52138_new_n4734_), .Y(u2__abc_52138_new_n7973_));
OAI21X1 OAI21X1_1189 ( .A(u2__abc_52138_new_n4740_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7976_));
OAI21X1 OAI21X1_119 ( .A(\a[112] ), .B(_abc_65734_new_n1183_), .C(_abc_65734_new_n1186_), .Y(fracta1_7_));
OAI21X1 OAI21X1_1190 ( .A(u2__abc_52138_new_n7976_), .B(u2__abc_52138_new_n7975_), .C(u2__abc_52138_new_n7977_), .Y(u2__abc_52138_new_n7978_));
OAI21X1 OAI21X1_1191 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_136_), .Y(u2__abc_52138_new_n7980_));
OAI21X1 OAI21X1_1192 ( .A(u2__abc_52138_new_n4744_), .B(u2_remHi_131_), .C(u2__abc_52138_new_n7962_), .Y(u2__abc_52138_new_n7983_));
OAI21X1 OAI21X1_1193 ( .A(u2__abc_52138_new_n4764_), .B(u2__abc_52138_new_n7983_), .C(u2__abc_52138_new_n7985_), .Y(u2__abc_52138_new_n7986_));
OAI21X1 OAI21X1_1194 ( .A(u2__abc_52138_new_n4751_), .B(u2__abc_52138_new_n7901_), .C(u2__abc_52138_new_n7987_), .Y(u2__abc_52138_new_n7988_));
OAI21X1 OAI21X1_1195 ( .A(u2__abc_52138_new_n7991_), .B(u2__abc_52138_new_n7990_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7992_));
OAI21X1 OAI21X1_1196 ( .A(u2_remHi_134_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7992_), .Y(u2__abc_52138_new_n7993_));
OAI21X1 OAI21X1_1197 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_137_), .Y(u2__abc_52138_new_n7998_));
OAI21X1 OAI21X1_1198 ( .A(sqrto_134_), .B(u2__abc_52138_new_n4679_), .C(u2__abc_52138_new_n7989_), .Y(u2__abc_52138_new_n7999_));
OAI21X1 OAI21X1_1199 ( .A(u2__abc_52138_new_n4684_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8002_));
OAI21X1 OAI21X1_12 ( .A(aNan), .B(_abc_65734_new_n863_), .C(_abc_65734_new_n864_), .Y(\o[123] ));
OAI21X1 OAI21X1_120 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1188_), .C(_abc_65734_new_n1189_), .Y(fracta1_8_));
OAI21X1 OAI21X1_1200 ( .A(u2__abc_52138_new_n8002_), .B(u2__abc_52138_new_n8001_), .C(u2__abc_52138_new_n8003_), .Y(u2__abc_52138_new_n8004_));
OAI21X1 OAI21X1_1201 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_138_), .Y(u2__abc_52138_new_n8006_));
OAI21X1 OAI21X1_1202 ( .A(u2__abc_52138_new_n8010_), .B(u2__abc_52138_new_n8011_), .C(u2__abc_52138_new_n8008_), .Y(u2__abc_52138_new_n8012_));
OAI21X1 OAI21X1_1203 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n8012_), .Y(u2__abc_52138_new_n8013_));
OAI21X1 OAI21X1_1204 ( .A(u2__abc_52138_new_n4668_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8015_));
OAI21X1 OAI21X1_1205 ( .A(u2__abc_52138_new_n8015_), .B(u2__abc_52138_new_n8014_), .C(u2__abc_52138_new_n8016_), .Y(u2__abc_52138_new_n8017_));
OAI21X1 OAI21X1_1206 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_139_), .Y(u2__abc_52138_new_n8019_));
OAI21X1 OAI21X1_1207 ( .A(u2__abc_52138_new_n8011_), .B(u2__abc_52138_new_n8008_), .C(u2__abc_52138_new_n4667_), .Y(u2__abc_52138_new_n8022_));
OAI21X1 OAI21X1_1208 ( .A(u2__abc_52138_new_n8021_), .B(u2__abc_52138_new_n8022_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8023_));
OAI21X1 OAI21X1_1209 ( .A(u2__abc_52138_new_n4673_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8025_));
OAI21X1 OAI21X1_121 ( .A(\a[112] ), .B(_abc_65734_new_n1188_), .C(_abc_65734_new_n1191_), .Y(fracta1_9_));
OAI21X1 OAI21X1_1210 ( .A(u2__abc_52138_new_n8025_), .B(u2__abc_52138_new_n8024_), .C(u2__abc_52138_new_n8026_), .Y(u2__abc_52138_new_n8027_));
OAI21X1 OAI21X1_1211 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_140_), .Y(u2__abc_52138_new_n8029_));
OAI21X1 OAI21X1_1212 ( .A(u2__abc_52138_new_n8030_), .B(u2__abc_52138_new_n8007_), .C(u2__abc_52138_new_n4685_), .Y(u2__abc_52138_new_n8031_));
OAI21X1 OAI21X1_1213 ( .A(u2__abc_52138_new_n8031_), .B(u2__abc_52138_new_n4785_), .C(u2__abc_52138_new_n8032_), .Y(u2__abc_52138_new_n8033_));
OAI21X1 OAI21X1_1214 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n8036_), .Y(u2__abc_52138_new_n8037_));
OAI21X1 OAI21X1_1215 ( .A(u2__abc_52138_new_n4707_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8039_));
OAI21X1 OAI21X1_1216 ( .A(u2__abc_52138_new_n8039_), .B(u2__abc_52138_new_n8038_), .C(u2__abc_52138_new_n8040_), .Y(u2__abc_52138_new_n8041_));
OAI21X1 OAI21X1_1217 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_141_), .Y(u2__abc_52138_new_n8043_));
OAI21X1 OAI21X1_1218 ( .A(u2__abc_52138_new_n4709_), .B(u2__abc_52138_new_n8034_), .C(u2__abc_52138_new_n4706_), .Y(u2__abc_52138_new_n8044_));
OAI21X1 OAI21X1_1219 ( .A(u2__abc_52138_new_n4702_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8047_));
OAI21X1 OAI21X1_122 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1193_), .C(_abc_65734_new_n1194_), .Y(fracta1_10_));
OAI21X1 OAI21X1_1220 ( .A(u2__abc_52138_new_n8047_), .B(u2__abc_52138_new_n8046_), .C(u2__abc_52138_new_n8048_), .Y(u2__abc_52138_new_n8049_));
OAI21X1 OAI21X1_1221 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_142_), .Y(u2__abc_52138_new_n8051_));
OAI21X1 OAI21X1_1222 ( .A(sqrto_138_), .B(u2__abc_52138_new_n4707_), .C(u2__abc_52138_new_n4701_), .Y(u2__abc_52138_new_n8052_));
OAI21X1 OAI21X1_1223 ( .A(u2__abc_52138_new_n8052_), .B(u2__abc_52138_new_n8035_), .C(u2__abc_52138_new_n4703_), .Y(u2__abc_52138_new_n8053_));
OAI21X1 OAI21X1_1224 ( .A(u2__abc_52138_new_n4691_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8056_));
OAI21X1 OAI21X1_1225 ( .A(u2__abc_52138_new_n8056_), .B(u2__abc_52138_new_n8055_), .C(u2__abc_52138_new_n8057_), .Y(u2__abc_52138_new_n8058_));
OAI21X1 OAI21X1_1226 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_143_), .Y(u2__abc_52138_new_n8060_));
OAI21X1 OAI21X1_1227 ( .A(u2__abc_52138_new_n4693_), .B(u2__abc_52138_new_n8053_), .C(u2__abc_52138_new_n4690_), .Y(u2__abc_52138_new_n8061_));
OAI21X1 OAI21X1_1228 ( .A(u2__abc_52138_new_n4696_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8064_));
OAI21X1 OAI21X1_1229 ( .A(u2__abc_52138_new_n8064_), .B(u2__abc_52138_new_n8063_), .C(u2__abc_52138_new_n8065_), .Y(u2__abc_52138_new_n8066_));
OAI21X1 OAI21X1_123 ( .A(\a[112] ), .B(_abc_65734_new_n1193_), .C(_abc_65734_new_n1196_), .Y(fracta1_11_));
OAI21X1 OAI21X1_1230 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_144_), .Y(u2__abc_52138_new_n8068_));
OAI21X1 OAI21X1_1231 ( .A(u2__abc_52138_new_n4706_), .B(u2__abc_52138_new_n4704_), .C(u2__abc_52138_new_n4701_), .Y(u2__abc_52138_new_n8074_));
OAI21X1 OAI21X1_1232 ( .A(u2__abc_52138_new_n4690_), .B(u2__abc_52138_new_n4698_), .C(u2__abc_52138_new_n4695_), .Y(u2__abc_52138_new_n8075_));
OAI21X1 OAI21X1_1233 ( .A(u2__abc_52138_new_n7899_), .B(u2__abc_52138_new_n7889_), .C(u2__abc_52138_new_n8079_), .Y(u2__abc_52138_new_n8080_));
OAI21X1 OAI21X1_1234 ( .A(u2__abc_52138_new_n8084_), .B(u2__abc_52138_new_n8083_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8085_));
OAI21X1 OAI21X1_1235 ( .A(u2_remHi_142_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n8085_), .Y(u2__abc_52138_new_n8086_));
OAI21X1 OAI21X1_1236 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_145_), .Y(u2__abc_52138_new_n8091_));
OAI21X1 OAI21X1_1237 ( .A(sqrto_142_), .B(u2__abc_52138_new_n4658_), .C(u2__abc_52138_new_n8082_), .Y(u2__abc_52138_new_n8093_));
OAI21X1 OAI21X1_1238 ( .A(u2__abc_52138_new_n4652_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8096_));
OAI21X1 OAI21X1_1239 ( .A(u2__abc_52138_new_n8096_), .B(u2__abc_52138_new_n8095_), .C(u2__abc_52138_new_n8097_), .Y(u2__abc_52138_new_n8098_));
OAI21X1 OAI21X1_124 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1198_), .C(_abc_65734_new_n1199_), .Y(fracta1_12_));
OAI21X1 OAI21X1_1240 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_146_), .Y(u2__abc_52138_new_n8100_));
OAI21X1 OAI21X1_1241 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n8104_), .Y(u2__abc_52138_new_n8105_));
OAI21X1 OAI21X1_1242 ( .A(u2__abc_52138_new_n4644_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8107_));
OAI21X1 OAI21X1_1243 ( .A(u2__abc_52138_new_n8107_), .B(u2__abc_52138_new_n8106_), .C(u2__abc_52138_new_n8108_), .Y(u2__abc_52138_new_n8109_));
OAI21X1 OAI21X1_1244 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_147_), .Y(u2__abc_52138_new_n8111_));
OAI21X1 OAI21X1_1245 ( .A(u2__abc_52138_new_n4802_), .B(u2__abc_52138_new_n8102_), .C(u2__abc_52138_new_n4643_), .Y(u2__abc_52138_new_n8113_));
OAI21X1 OAI21X1_1246 ( .A(u2__abc_52138_new_n4649_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8116_));
OAI21X1 OAI21X1_1247 ( .A(u2__abc_52138_new_n8116_), .B(u2__abc_52138_new_n8115_), .C(u2__abc_52138_new_n8117_), .Y(u2__abc_52138_new_n8118_));
OAI21X1 OAI21X1_1248 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_148_), .Y(u2__abc_52138_new_n8120_));
OAI21X1 OAI21X1_1249 ( .A(sqrto_145_), .B(u2__abc_52138_new_n4649_), .C(u2__abc_52138_new_n4643_), .Y(u2__abc_52138_new_n8121_));
OAI21X1 OAI21X1_125 ( .A(\a[112] ), .B(_abc_65734_new_n1198_), .C(_abc_65734_new_n1201_), .Y(fracta1_13_));
OAI21X1 OAI21X1_1250 ( .A(u2__abc_52138_new_n8121_), .B(u2__abc_52138_new_n8103_), .C(u2__abc_52138_new_n4650_), .Y(u2__abc_52138_new_n8122_));
OAI21X1 OAI21X1_1251 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n8124_), .Y(u2__abc_52138_new_n8125_));
OAI21X1 OAI21X1_1252 ( .A(u2__abc_52138_new_n4637_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8127_));
OAI21X1 OAI21X1_1253 ( .A(u2__abc_52138_new_n8127_), .B(u2__abc_52138_new_n8126_), .C(u2__abc_52138_new_n8128_), .Y(u2__abc_52138_new_n8129_));
OAI21X1 OAI21X1_1254 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_149_), .Y(u2__abc_52138_new_n8131_));
OAI21X1 OAI21X1_1255 ( .A(u2__abc_52138_new_n4639_), .B(u2__abc_52138_new_n8122_), .C(u2__abc_52138_new_n4636_), .Y(u2__abc_52138_new_n8133_));
OAI21X1 OAI21X1_1256 ( .A(u2__abc_52138_new_n8132_), .B(u2__abc_52138_new_n8133_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8134_));
OAI21X1 OAI21X1_1257 ( .A(u2__abc_52138_new_n4632_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8136_));
OAI21X1 OAI21X1_1258 ( .A(u2__abc_52138_new_n8136_), .B(u2__abc_52138_new_n8135_), .C(u2__abc_52138_new_n8137_), .Y(u2__abc_52138_new_n8138_));
OAI21X1 OAI21X1_1259 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_150_), .Y(u2__abc_52138_new_n8140_));
OAI21X1 OAI21X1_126 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1203_), .C(_abc_65734_new_n1204_), .Y(fracta1_14_));
OAI21X1 OAI21X1_1260 ( .A(sqrto_147_), .B(u2__abc_52138_new_n4632_), .C(u2__abc_52138_new_n8143_), .Y(u2__abc_52138_new_n8144_));
OAI21X1 OAI21X1_1261 ( .A(u2__abc_52138_new_n4621_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8148_));
OAI21X1 OAI21X1_1262 ( .A(u2_remHi_150_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8150_));
OAI21X1 OAI21X1_1263 ( .A(u2__abc_52138_new_n8150_), .B(u2__abc_52138_new_n8149_), .C(u2__abc_52138_new_n8140_), .Y(u2__abc_52138_new_n8151_));
OAI21X1 OAI21X1_1264 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_151_), .Y(u2__abc_52138_new_n8153_));
OAI21X1 OAI21X1_1265 ( .A(sqrto_148_), .B(u2__abc_52138_new_n4621_), .C(u2__abc_52138_new_n8145_), .Y(u2__abc_52138_new_n8154_));
OAI21X1 OAI21X1_1266 ( .A(u2__abc_52138_new_n4626_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8157_));
OAI21X1 OAI21X1_1267 ( .A(u2__abc_52138_new_n8157_), .B(u2__abc_52138_new_n8156_), .C(u2__abc_52138_new_n8158_), .Y(u2__abc_52138_new_n8159_));
OAI21X1 OAI21X1_1268 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_152_), .Y(u2__abc_52138_new_n8161_));
OAI21X1 OAI21X1_1269 ( .A(u2__abc_52138_new_n4807_), .B(u2__abc_52138_new_n8163_), .C(u2__abc_52138_new_n4629_), .Y(u2__abc_52138_new_n8164_));
OAI21X1 OAI21X1_127 ( .A(\a[112] ), .B(_abc_65734_new_n1203_), .C(_abc_65734_new_n1206_), .Y(fracta1_15_));
OAI21X1 OAI21X1_1270 ( .A(u2__abc_52138_new_n4653_), .B(u2__abc_52138_new_n4659_), .C(u2__abc_52138_new_n4657_), .Y(u2__abc_52138_new_n8165_));
OAI21X1 OAI21X1_1271 ( .A(u2__abc_52138_new_n4647_), .B(u2_remHi_145_), .C(u2__abc_52138_new_n8121_), .Y(u2__abc_52138_new_n8166_));
OAI21X1 OAI21X1_1272 ( .A(u2__abc_52138_new_n8165_), .B(u2__abc_52138_new_n4651_), .C(u2__abc_52138_new_n8166_), .Y(u2__abc_52138_new_n8167_));
OAI21X1 OAI21X1_1273 ( .A(u2__abc_52138_new_n4620_), .B(u2__abc_52138_new_n4811_), .C(u2__abc_52138_new_n4625_), .Y(u2__abc_52138_new_n8168_));
OAI21X1 OAI21X1_1274 ( .A(u2__abc_52138_new_n8170_), .B(u2__abc_52138_new_n8171_), .C(u2__abc_52138_new_n8162_), .Y(u2__abc_52138_new_n8172_));
OAI21X1 OAI21X1_1275 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n8176_), .C(u2__abc_52138_new_n8177_), .Y(u2__abc_52138_new_n8178_));
OAI21X1 OAI21X1_1276 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_153_), .Y(u2__abc_52138_new_n8180_));
OAI21X1 OAI21X1_1277 ( .A(sqrto_150_), .B(u2__abc_52138_new_n4591_), .C(u2__abc_52138_new_n8172_), .Y(u2__abc_52138_new_n8181_));
OAI21X1 OAI21X1_1278 ( .A(u2__abc_52138_new_n4586_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8184_));
OAI21X1 OAI21X1_1279 ( .A(u2__abc_52138_new_n8184_), .B(u2__abc_52138_new_n8183_), .C(u2__abc_52138_new_n8185_), .Y(u2__abc_52138_new_n8186_));
OAI21X1 OAI21X1_128 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1208_), .C(_abc_65734_new_n1209_), .Y(fracta1_16_));
OAI21X1 OAI21X1_1280 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_154_), .Y(u2__abc_52138_new_n8188_));
OAI21X1 OAI21X1_1281 ( .A(sqrto_150_), .B(u2__abc_52138_new_n4591_), .C(u2__abc_52138_new_n4585_), .Y(u2__abc_52138_new_n8190_));
OAI21X1 OAI21X1_1282 ( .A(u2__abc_52138_new_n8190_), .B(u2__abc_52138_new_n8189_), .C(u2__abc_52138_new_n4587_), .Y(u2__abc_52138_new_n8191_));
OAI21X1 OAI21X1_1283 ( .A(u2__abc_52138_new_n4575_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8194_));
OAI21X1 OAI21X1_1284 ( .A(u2__abc_52138_new_n8194_), .B(u2__abc_52138_new_n8193_), .C(u2__abc_52138_new_n8195_), .Y(u2__abc_52138_new_n8196_));
OAI21X1 OAI21X1_1285 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_155_), .Y(u2__abc_52138_new_n8198_));
OAI21X1 OAI21X1_1286 ( .A(u2__abc_52138_new_n4577_), .B(u2__abc_52138_new_n8191_), .C(u2__abc_52138_new_n4574_), .Y(u2__abc_52138_new_n8199_));
OAI21X1 OAI21X1_1287 ( .A(u2__abc_52138_new_n4580_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8202_));
OAI21X1 OAI21X1_1288 ( .A(u2__abc_52138_new_n8202_), .B(u2__abc_52138_new_n8201_), .C(u2__abc_52138_new_n8203_), .Y(u2__abc_52138_new_n8204_));
OAI21X1 OAI21X1_1289 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_156_), .Y(u2__abc_52138_new_n8206_));
OAI21X1 OAI21X1_129 ( .A(\a[112] ), .B(_abc_65734_new_n1208_), .C(_abc_65734_new_n1211_), .Y(fracta1_17_));
OAI21X1 OAI21X1_1290 ( .A(u2__abc_52138_new_n4590_), .B(u2__abc_52138_new_n4588_), .C(u2__abc_52138_new_n4585_), .Y(u2__abc_52138_new_n8207_));
OAI21X1 OAI21X1_1291 ( .A(u2__abc_52138_new_n4574_), .B(u2__abc_52138_new_n4582_), .C(u2__abc_52138_new_n4579_), .Y(u2__abc_52138_new_n8208_));
OAI21X1 OAI21X1_1292 ( .A(u2__abc_52138_new_n4595_), .B(u2__abc_52138_new_n8173_), .C(u2__abc_52138_new_n8209_), .Y(u2__abc_52138_new_n8210_));
OAI21X1 OAI21X1_1293 ( .A(u2__abc_52138_new_n4616_), .B(u2__abc_52138_new_n8210_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8213_));
OAI21X1 OAI21X1_1294 ( .A(u2__abc_52138_new_n4612_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8215_));
OAI21X1 OAI21X1_1295 ( .A(u2_remHi_156_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8217_));
OAI21X1 OAI21X1_1296 ( .A(u2__abc_52138_new_n8217_), .B(u2__abc_52138_new_n8216_), .C(u2__abc_52138_new_n8206_), .Y(u2__abc_52138_new_n8218_));
OAI21X1 OAI21X1_1297 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_157_), .Y(u2__abc_52138_new_n8220_));
OAI21X1 OAI21X1_1298 ( .A(sqrto_154_), .B(u2__abc_52138_new_n4612_), .C(u2__abc_52138_new_n8211_), .Y(u2__abc_52138_new_n8221_));
OAI21X1 OAI21X1_1299 ( .A(u2__abc_52138_new_n4607_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8224_));
OAI21X1 OAI21X1_13 ( .A(aNan), .B(_abc_65734_new_n866_), .C(_abc_65734_new_n867_), .Y(\o[124] ));
OAI21X1 OAI21X1_130 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1213_), .C(_abc_65734_new_n1214_), .Y(fracta1_18_));
OAI21X1 OAI21X1_1300 ( .A(u2__abc_52138_new_n8224_), .B(u2__abc_52138_new_n8223_), .C(u2__abc_52138_new_n8225_), .Y(u2__abc_52138_new_n8226_));
OAI21X1 OAI21X1_1301 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_158_), .Y(u2__abc_52138_new_n8228_));
OAI21X1 OAI21X1_1302 ( .A(u2__abc_52138_new_n8230_), .B(u2__abc_52138_new_n8212_), .C(u2__abc_52138_new_n8229_), .Y(u2__abc_52138_new_n8231_));
OAI21X1 OAI21X1_1303 ( .A(u2__abc_52138_new_n4598_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8234_));
OAI21X1 OAI21X1_1304 ( .A(u2__abc_52138_new_n8234_), .B(u2__abc_52138_new_n8233_), .C(u2__abc_52138_new_n8235_), .Y(u2__abc_52138_new_n8236_));
OAI21X1 OAI21X1_1305 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_159_), .Y(u2__abc_52138_new_n8238_));
OAI21X1 OAI21X1_1306 ( .A(u2__abc_52138_new_n4600_), .B(u2__abc_52138_new_n8231_), .C(u2__abc_52138_new_n4597_), .Y(u2__abc_52138_new_n8239_));
OAI21X1 OAI21X1_1307 ( .A(u2__abc_52138_new_n4603_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8242_));
OAI21X1 OAI21X1_1308 ( .A(u2__abc_52138_new_n8242_), .B(u2__abc_52138_new_n8241_), .C(u2__abc_52138_new_n8244_), .Y(u2__abc_52138_new_n8245_));
OAI21X1 OAI21X1_1309 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_160_), .Y(u2__abc_52138_new_n8247_));
OAI21X1 OAI21X1_131 ( .A(\a[112] ), .B(_abc_65734_new_n1213_), .C(_abc_65734_new_n1216_), .Y(fracta1_19_));
OAI21X1 OAI21X1_1310 ( .A(u2__abc_52138_new_n4597_), .B(u2__abc_52138_new_n4605_), .C(u2__abc_52138_new_n4602_), .Y(u2__abc_52138_new_n8250_));
OAI21X1 OAI21X1_1311 ( .A(u2__abc_52138_new_n4617_), .B(u2__abc_52138_new_n8209_), .C(u2__abc_52138_new_n8251_), .Y(u2__abc_52138_new_n8252_));
OAI21X1 OAI21X1_1312 ( .A(u2__abc_52138_new_n7899_), .B(u2__abc_52138_new_n7889_), .C(u2__abc_52138_new_n4752_), .Y(u2__abc_52138_new_n8255_));
OAI21X1 OAI21X1_1313 ( .A(u2__abc_52138_new_n4542_), .B(u2__abc_52138_new_n4544_), .C(u2__abc_52138_new_n8257_), .Y(u2__abc_52138_new_n8260_));
OAI21X1 OAI21X1_1314 ( .A(u2__abc_52138_new_n4541_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8263_));
OAI21X1 OAI21X1_1315 ( .A(u2__abc_52138_new_n8263_), .B(u2__abc_52138_new_n8262_), .C(u2__abc_52138_new_n8264_), .Y(u2__abc_52138_new_n8265_));
OAI21X1 OAI21X1_1316 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_161_), .Y(u2__abc_52138_new_n8267_));
OAI21X1 OAI21X1_1317 ( .A(sqrto_158_), .B(u2__abc_52138_new_n4541_), .C(u2__abc_52138_new_n8259_), .Y(u2__abc_52138_new_n8268_));
OAI21X1 OAI21X1_1318 ( .A(u2__abc_52138_new_n8243_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8271_));
OAI21X1 OAI21X1_1319 ( .A(u2__abc_52138_new_n8271_), .B(u2__abc_52138_new_n8270_), .C(u2__abc_52138_new_n8272_), .Y(u2__abc_52138_new_n8273_));
OAI21X1 OAI21X1_132 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1218_), .C(_abc_65734_new_n1219_), .Y(fracta1_20_));
OAI21X1 OAI21X1_1320 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_162_), .Y(u2__abc_52138_new_n8275_));
OAI21X1 OAI21X1_1321 ( .A(sqrto_158_), .B(u2__abc_52138_new_n4541_), .C(u2__abc_52138_new_n4537_), .Y(u2__abc_52138_new_n8276_));
OAI21X1 OAI21X1_1322 ( .A(u2__abc_52138_new_n8276_), .B(u2__abc_52138_new_n8258_), .C(u2__abc_52138_new_n4539_), .Y(u2__abc_52138_new_n8277_));
OAI21X1 OAI21X1_1323 ( .A(u2__abc_52138_new_n8279_), .B(u2__abc_52138_new_n8280_), .C(u2__abc_52138_new_n8277_), .Y(u2__abc_52138_new_n8281_));
OAI21X1 OAI21X1_1324 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n8281_), .Y(u2__abc_52138_new_n8282_));
OAI21X1 OAI21X1_1325 ( .A(u2__abc_52138_new_n4527_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8284_));
OAI21X1 OAI21X1_1326 ( .A(u2__abc_52138_new_n8284_), .B(u2__abc_52138_new_n8283_), .C(u2__abc_52138_new_n8285_), .Y(u2__abc_52138_new_n8286_));
OAI21X1 OAI21X1_1327 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_163_), .Y(u2__abc_52138_new_n8288_));
OAI21X1 OAI21X1_1328 ( .A(u2__abc_52138_new_n8280_), .B(u2__abc_52138_new_n8277_), .C(u2__abc_52138_new_n4526_), .Y(u2__abc_52138_new_n8291_));
OAI21X1 OAI21X1_1329 ( .A(u2__abc_52138_new_n8290_), .B(u2__abc_52138_new_n8291_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8292_));
OAI21X1 OAI21X1_133 ( .A(\a[112] ), .B(_abc_65734_new_n1218_), .C(_abc_65734_new_n1221_), .Y(fracta1_21_));
OAI21X1 OAI21X1_1330 ( .A(u2__abc_52138_new_n4532_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8294_));
OAI21X1 OAI21X1_1331 ( .A(u2__abc_52138_new_n8294_), .B(u2__abc_52138_new_n8293_), .C(u2__abc_52138_new_n8295_), .Y(u2__abc_52138_new_n8296_));
OAI21X1 OAI21X1_1332 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_164_), .Y(u2__abc_52138_new_n8298_));
OAI21X1 OAI21X1_1333 ( .A(u2__abc_52138_new_n4536_), .B(u2_remHi_159_), .C(u2__abc_52138_new_n8276_), .Y(u2__abc_52138_new_n8299_));
OAI21X1 OAI21X1_1334 ( .A(u2__abc_52138_new_n8299_), .B(u2__abc_52138_new_n4831_), .C(u2__abc_52138_new_n8300_), .Y(u2__abc_52138_new_n8301_));
OAI21X1 OAI21X1_1335 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n8307_), .C(u2__abc_52138_new_n8308_), .Y(u2__abc_52138_new_n8309_));
OAI21X1 OAI21X1_1336 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_165_), .Y(u2__abc_52138_new_n8311_));
OAI21X1 OAI21X1_1337 ( .A(u2__abc_52138_new_n4568_), .B(u2__abc_52138_new_n8302_), .C(u2__abc_52138_new_n4565_), .Y(u2__abc_52138_new_n8313_));
OAI21X1 OAI21X1_1338 ( .A(u2__abc_52138_new_n8312_), .B(u2__abc_52138_new_n8313_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8314_));
OAI21X1 OAI21X1_1339 ( .A(u2__abc_52138_new_n4561_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8316_));
OAI21X1 OAI21X1_134 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1223_), .C(_abc_65734_new_n1224_), .Y(fracta1_22_));
OAI21X1 OAI21X1_1340 ( .A(u2__abc_52138_new_n8316_), .B(u2__abc_52138_new_n8315_), .C(u2__abc_52138_new_n8317_), .Y(u2__abc_52138_new_n8318_));
OAI21X1 OAI21X1_1341 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_166_), .Y(u2__abc_52138_new_n8320_));
OAI21X1 OAI21X1_1342 ( .A(u2__abc_52138_new_n4565_), .B(u2__abc_52138_new_n4563_), .C(u2__abc_52138_new_n4560_), .Y(u2__abc_52138_new_n8321_));
OAI21X1 OAI21X1_1343 ( .A(u2__abc_52138_new_n4563_), .B(u2__abc_52138_new_n8304_), .C(u2__abc_52138_new_n8322_), .Y(u2__abc_52138_new_n8323_));
OAI21X1 OAI21X1_1344 ( .A(u2__abc_52138_new_n4550_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8326_));
OAI21X1 OAI21X1_1345 ( .A(u2__abc_52138_new_n8326_), .B(u2__abc_52138_new_n8325_), .C(u2__abc_52138_new_n8327_), .Y(u2__abc_52138_new_n8328_));
OAI21X1 OAI21X1_1346 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_167_), .Y(u2__abc_52138_new_n8330_));
OAI21X1 OAI21X1_1347 ( .A(u2__abc_52138_new_n4555_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8335_));
OAI21X1 OAI21X1_1348 ( .A(u2__abc_52138_new_n8335_), .B(u2__abc_52138_new_n8334_), .C(u2__abc_52138_new_n8336_), .Y(u2__abc_52138_new_n8337_));
OAI21X1 OAI21X1_1349 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_168_), .Y(u2__abc_52138_new_n8339_));
OAI21X1 OAI21X1_135 ( .A(\a[112] ), .B(_abc_65734_new_n1223_), .C(_abc_65734_new_n1226_), .Y(fracta1_23_));
OAI21X1 OAI21X1_1350 ( .A(u2__abc_52138_new_n4549_), .B(u2__abc_52138_new_n4557_), .C(u2__abc_52138_new_n4554_), .Y(u2__abc_52138_new_n8340_));
OAI21X1 OAI21X1_1351 ( .A(u2__abc_52138_new_n4837_), .B(u2__abc_52138_new_n8322_), .C(u2__abc_52138_new_n8341_), .Y(u2__abc_52138_new_n8342_));
OAI21X1 OAI21X1_1352 ( .A(u2__abc_52138_new_n4757_), .B(u2__abc_52138_new_n8257_), .C(u2__abc_52138_new_n8343_), .Y(u2__abc_52138_new_n8344_));
OAI21X1 OAI21X1_1353 ( .A(u2__abc_52138_new_n4517_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8350_));
OAI21X1 OAI21X1_1354 ( .A(u2__abc_52138_new_n8350_), .B(u2__abc_52138_new_n8349_), .C(u2__abc_52138_new_n8351_), .Y(u2__abc_52138_new_n8352_));
OAI21X1 OAI21X1_1355 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_169_), .Y(u2__abc_52138_new_n8354_));
OAI21X1 OAI21X1_1356 ( .A(sqrto_166_), .B(u2__abc_52138_new_n4517_), .C(u2__abc_52138_new_n8347_), .Y(u2__abc_52138_new_n8355_));
OAI21X1 OAI21X1_1357 ( .A(u2__abc_52138_new_n4514_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8358_));
OAI21X1 OAI21X1_1358 ( .A(u2__abc_52138_new_n8358_), .B(u2__abc_52138_new_n8357_), .C(u2__abc_52138_new_n8359_), .Y(u2__abc_52138_new_n8360_));
OAI21X1 OAI21X1_1359 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_170_), .Y(u2__abc_52138_new_n8362_));
OAI21X1 OAI21X1_136 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1228_), .C(_abc_65734_new_n1229_), .Y(fracta1_24_));
OAI21X1 OAI21X1_1360 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n8366_), .Y(u2__abc_52138_new_n8367_));
OAI21X1 OAI21X1_1361 ( .A(u2__abc_52138_new_n4503_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8369_));
OAI21X1 OAI21X1_1362 ( .A(u2__abc_52138_new_n8369_), .B(u2__abc_52138_new_n8368_), .C(u2__abc_52138_new_n8370_), .Y(u2__abc_52138_new_n8371_));
OAI21X1 OAI21X1_1363 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_171_), .Y(u2__abc_52138_new_n8373_));
OAI21X1 OAI21X1_1364 ( .A(u2__abc_52138_new_n4505_), .B(u2__abc_52138_new_n8364_), .C(u2__abc_52138_new_n4502_), .Y(u2__abc_52138_new_n8374_));
OAI21X1 OAI21X1_1365 ( .A(u2__abc_52138_new_n4508_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8377_));
OAI21X1 OAI21X1_1366 ( .A(u2__abc_52138_new_n8377_), .B(u2__abc_52138_new_n8376_), .C(u2__abc_52138_new_n8378_), .Y(u2__abc_52138_new_n8379_));
OAI21X1 OAI21X1_1367 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_172_), .Y(u2__abc_52138_new_n8381_));
OAI21X1 OAI21X1_1368 ( .A(sqrto_169_), .B(u2__abc_52138_new_n4508_), .C(u2__abc_52138_new_n4502_), .Y(u2__abc_52138_new_n8382_));
OAI21X1 OAI21X1_1369 ( .A(u2__abc_52138_new_n8382_), .B(u2__abc_52138_new_n8365_), .C(u2__abc_52138_new_n4509_), .Y(u2__abc_52138_new_n8383_));
OAI21X1 OAI21X1_137 ( .A(\a[112] ), .B(_abc_65734_new_n1228_), .C(_abc_65734_new_n1231_), .Y(fracta1_25_));
OAI21X1 OAI21X1_1370 ( .A(u2__abc_52138_new_n4496_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8387_));
OAI21X1 OAI21X1_1371 ( .A(u2_remHi_172_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8389_));
OAI21X1 OAI21X1_1372 ( .A(u2__abc_52138_new_n8389_), .B(u2__abc_52138_new_n8388_), .C(u2__abc_52138_new_n8381_), .Y(u2__abc_52138_new_n8390_));
OAI21X1 OAI21X1_1373 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_173_), .Y(u2__abc_52138_new_n8392_));
OAI21X1 OAI21X1_1374 ( .A(u2__abc_52138_new_n4498_), .B(u2__abc_52138_new_n8383_), .C(u2__abc_52138_new_n4495_), .Y(u2__abc_52138_new_n8393_));
OAI21X1 OAI21X1_1375 ( .A(u2__abc_52138_new_n4491_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8396_));
OAI21X1 OAI21X1_1376 ( .A(u2__abc_52138_new_n8396_), .B(u2__abc_52138_new_n8395_), .C(u2__abc_52138_new_n8397_), .Y(u2__abc_52138_new_n8398_));
OAI21X1 OAI21X1_1377 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_174_), .Y(u2__abc_52138_new_n8400_));
OAI21X1 OAI21X1_1378 ( .A(sqrto_170_), .B(u2__abc_52138_new_n4496_), .C(u2__abc_52138_new_n4490_), .Y(u2__abc_52138_new_n8401_));
OAI21X1 OAI21X1_1379 ( .A(u2__abc_52138_new_n8401_), .B(u2__abc_52138_new_n8384_), .C(u2__abc_52138_new_n4492_), .Y(u2__abc_52138_new_n8402_));
OAI21X1 OAI21X1_138 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1233_), .C(_abc_65734_new_n1234_), .Y(fracta1_26_));
OAI21X1 OAI21X1_1380 ( .A(u2__abc_52138_new_n4480_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8405_));
OAI21X1 OAI21X1_1381 ( .A(u2__abc_52138_new_n8405_), .B(u2__abc_52138_new_n8404_), .C(u2__abc_52138_new_n8406_), .Y(u2__abc_52138_new_n8407_));
OAI21X1 OAI21X1_1382 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_175_), .Y(u2__abc_52138_new_n8409_));
OAI21X1 OAI21X1_1383 ( .A(u2__abc_52138_new_n4853_), .B(u2__abc_52138_new_n8402_), .C(u2__abc_52138_new_n4479_), .Y(u2__abc_52138_new_n8410_));
OAI21X1 OAI21X1_1384 ( .A(u2__abc_52138_new_n4485_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8413_));
OAI21X1 OAI21X1_1385 ( .A(u2__abc_52138_new_n8413_), .B(u2__abc_52138_new_n8412_), .C(u2__abc_52138_new_n8414_), .Y(u2__abc_52138_new_n8415_));
OAI21X1 OAI21X1_1386 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_176_), .Y(u2__abc_52138_new_n8417_));
OAI21X1 OAI21X1_1387 ( .A(u2__abc_52138_new_n4518_), .B(u2__abc_52138_new_n8363_), .C(u2__abc_52138_new_n4515_), .Y(u2__abc_52138_new_n8419_));
OAI21X1 OAI21X1_1388 ( .A(u2__abc_52138_new_n4506_), .B(u2_remHi_169_), .C(u2__abc_52138_new_n8382_), .Y(u2__abc_52138_new_n8420_));
OAI21X1 OAI21X1_1389 ( .A(u2__abc_52138_new_n8419_), .B(u2__abc_52138_new_n8418_), .C(u2__abc_52138_new_n8420_), .Y(u2__abc_52138_new_n8421_));
OAI21X1 OAI21X1_139 ( .A(\a[112] ), .B(_abc_65734_new_n1233_), .C(_abc_65734_new_n1236_), .Y(fracta1_27_));
OAI21X1 OAI21X1_1390 ( .A(u2__abc_52138_new_n4489_), .B(u2_remHi_171_), .C(u2__abc_52138_new_n8401_), .Y(u2__abc_52138_new_n8423_));
OAI21X1 OAI21X1_1391 ( .A(u2__abc_52138_new_n8424_), .B(u2__abc_52138_new_n8425_), .C(u2__abc_52138_new_n4486_), .Y(u2__abc_52138_new_n8426_));
OAI21X1 OAI21X1_1392 ( .A(u2__abc_52138_new_n8423_), .B(u2__abc_52138_new_n8422_), .C(u2__abc_52138_new_n8426_), .Y(u2__abc_52138_new_n8427_));
OAI21X1 OAI21X1_1393 ( .A(u2__abc_52138_new_n4756_), .B(u2__abc_52138_new_n8343_), .C(u2__abc_52138_new_n8428_), .Y(u2__abc_52138_new_n8429_));
OAI21X1 OAI21X1_1394 ( .A(u2__abc_52138_new_n8429_), .B(u2__abc_52138_new_n8430_), .C(u2__abc_52138_new_n4468_), .Y(u2__abc_52138_new_n8431_));
OAI21X1 OAI21X1_1395 ( .A(u2__abc_52138_new_n4465_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8435_));
OAI21X1 OAI21X1_1396 ( .A(u2__abc_52138_new_n8435_), .B(u2__abc_52138_new_n8434_), .C(u2__abc_52138_new_n8436_), .Y(u2__abc_52138_new_n8437_));
OAI21X1 OAI21X1_1397 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_177_), .Y(u2__abc_52138_new_n8439_));
OAI21X1 OAI21X1_1398 ( .A(sqrto_174_), .B(u2__abc_52138_new_n4465_), .C(u2__abc_52138_new_n8431_), .Y(u2__abc_52138_new_n8440_));
OAI21X1 OAI21X1_1399 ( .A(u2__abc_52138_new_n4474_), .B(u2__abc_52138_new_n8440_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8441_));
OAI21X1 OAI21X1_14 ( .A(aNan), .B(_abc_65734_new_n869_), .C(_abc_65734_new_n870_), .Y(\o[125] ));
OAI21X1 OAI21X1_140 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1238_), .C(_abc_65734_new_n1239_), .Y(fracta1_28_));
OAI21X1 OAI21X1_1400 ( .A(u2__abc_52138_new_n4471_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8443_));
OAI21X1 OAI21X1_1401 ( .A(u2__abc_52138_new_n8443_), .B(u2__abc_52138_new_n8442_), .C(u2__abc_52138_new_n8444_), .Y(u2__abc_52138_new_n8445_));
OAI21X1 OAI21X1_1402 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_178_), .Y(u2__abc_52138_new_n8447_));
OAI21X1 OAI21X1_1403 ( .A(u2__abc_52138_new_n4464_), .B(u2__abc_52138_new_n8450_), .C(u2__abc_52138_new_n4470_), .Y(u2__abc_52138_new_n8451_));
OAI21X1 OAI21X1_1404 ( .A(u2__abc_52138_new_n8449_), .B(u2__abc_52138_new_n8432_), .C(u2__abc_52138_new_n8452_), .Y(u2__abc_52138_new_n8453_));
OAI21X1 OAI21X1_1405 ( .A(u2__abc_52138_new_n4454_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8457_));
OAI21X1 OAI21X1_1406 ( .A(u2_remHi_178_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8459_));
OAI21X1 OAI21X1_1407 ( .A(u2__abc_52138_new_n8459_), .B(u2__abc_52138_new_n8458_), .C(u2__abc_52138_new_n8447_), .Y(u2__abc_52138_new_n8460_));
OAI21X1 OAI21X1_1408 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_179_), .Y(u2__abc_52138_new_n8462_));
OAI21X1 OAI21X1_1409 ( .A(sqrto_176_), .B(u2__abc_52138_new_n4454_), .C(u2__abc_52138_new_n8454_), .Y(u2__abc_52138_new_n8463_));
OAI21X1 OAI21X1_141 ( .A(\a[112] ), .B(_abc_65734_new_n1238_), .C(_abc_65734_new_n1241_), .Y(fracta1_29_));
OAI21X1 OAI21X1_1410 ( .A(u2__abc_52138_new_n4459_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8466_));
OAI21X1 OAI21X1_1411 ( .A(u2__abc_52138_new_n8466_), .B(u2__abc_52138_new_n8465_), .C(u2__abc_52138_new_n8467_), .Y(u2__abc_52138_new_n8468_));
OAI21X1 OAI21X1_1412 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_180_), .Y(u2__abc_52138_new_n8470_));
OAI21X1 OAI21X1_1413 ( .A(u2__abc_52138_new_n4453_), .B(u2__abc_52138_new_n4461_), .C(u2__abc_52138_new_n4458_), .Y(u2__abc_52138_new_n8471_));
OAI21X1 OAI21X1_1414 ( .A(u2__abc_52138_new_n4475_), .B(u2__abc_52138_new_n8432_), .C(u2__abc_52138_new_n8472_), .Y(u2__abc_52138_new_n8473_));
OAI21X1 OAI21X1_1415 ( .A(u2__abc_52138_new_n4447_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8478_));
OAI21X1 OAI21X1_1416 ( .A(u2_remHi_180_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8480_));
OAI21X1 OAI21X1_1417 ( .A(u2__abc_52138_new_n8480_), .B(u2__abc_52138_new_n8479_), .C(u2__abc_52138_new_n8470_), .Y(u2__abc_52138_new_n8481_));
OAI21X1 OAI21X1_1418 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_181_), .Y(u2__abc_52138_new_n8483_));
OAI21X1 OAI21X1_1419 ( .A(u2__abc_52138_new_n4449_), .B(u2__abc_52138_new_n8474_), .C(u2__abc_52138_new_n4446_), .Y(u2__abc_52138_new_n8484_));
OAI21X1 OAI21X1_142 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1243_), .C(_abc_65734_new_n1244_), .Y(fracta1_30_));
OAI21X1 OAI21X1_1420 ( .A(u2__abc_52138_new_n4442_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8487_));
OAI21X1 OAI21X1_1421 ( .A(u2__abc_52138_new_n8487_), .B(u2__abc_52138_new_n8486_), .C(u2__abc_52138_new_n8488_), .Y(u2__abc_52138_new_n8489_));
OAI21X1 OAI21X1_1422 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_182_), .Y(u2__abc_52138_new_n8491_));
OAI21X1 OAI21X1_1423 ( .A(sqrto_178_), .B(u2__abc_52138_new_n4447_), .C(u2__abc_52138_new_n4441_), .Y(u2__abc_52138_new_n8492_));
OAI21X1 OAI21X1_1424 ( .A(u2__abc_52138_new_n8492_), .B(u2__abc_52138_new_n8475_), .C(u2__abc_52138_new_n4443_), .Y(u2__abc_52138_new_n8493_));
OAI21X1 OAI21X1_1425 ( .A(u2__abc_52138_new_n4431_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8496_));
OAI21X1 OAI21X1_1426 ( .A(u2__abc_52138_new_n8496_), .B(u2__abc_52138_new_n8495_), .C(u2__abc_52138_new_n8497_), .Y(u2__abc_52138_new_n8498_));
OAI21X1 OAI21X1_1427 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_183_), .Y(u2__abc_52138_new_n8500_));
OAI21X1 OAI21X1_1428 ( .A(u2__abc_52138_new_n4433_), .B(u2__abc_52138_new_n8493_), .C(u2__abc_52138_new_n4430_), .Y(u2__abc_52138_new_n8501_));
OAI21X1 OAI21X1_1429 ( .A(u2__abc_52138_new_n4436_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8504_));
OAI21X1 OAI21X1_143 ( .A(\a[112] ), .B(_abc_65734_new_n1243_), .C(_abc_65734_new_n1246_), .Y(fracta1_31_));
OAI21X1 OAI21X1_1430 ( .A(u2__abc_52138_new_n8504_), .B(u2__abc_52138_new_n8503_), .C(u2__abc_52138_new_n8505_), .Y(u2__abc_52138_new_n8506_));
OAI21X1 OAI21X1_1431 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_184_), .Y(u2__abc_52138_new_n8508_));
OAI21X1 OAI21X1_1432 ( .A(u2__abc_52138_new_n4446_), .B(u2__abc_52138_new_n4444_), .C(u2__abc_52138_new_n4441_), .Y(u2__abc_52138_new_n8509_));
OAI21X1 OAI21X1_1433 ( .A(u2__abc_52138_new_n4451_), .B(u2__abc_52138_new_n8472_), .C(u2__abc_52138_new_n8511_), .Y(u2__abc_52138_new_n8512_));
OAI21X1 OAI21X1_1434 ( .A(u2__abc_52138_new_n8429_), .B(u2__abc_52138_new_n8430_), .C(u2__abc_52138_new_n4476_), .Y(u2__abc_52138_new_n8514_));
OAI21X1 OAI21X1_1435 ( .A(u2__abc_52138_new_n4384_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8517_));
OAI21X1 OAI21X1_1436 ( .A(u2_remHi_184_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8519_));
OAI21X1 OAI21X1_1437 ( .A(u2__abc_52138_new_n8519_), .B(u2__abc_52138_new_n8518_), .C(u2__abc_52138_new_n8508_), .Y(u2__abc_52138_new_n8520_));
OAI21X1 OAI21X1_1438 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_185_), .Y(u2__abc_52138_new_n8522_));
OAI21X1 OAI21X1_1439 ( .A(u2__abc_52138_new_n4386_), .B(u2__abc_52138_new_n8523_), .C(u2__abc_52138_new_n4383_), .Y(u2__abc_52138_new_n8524_));
OAI21X1 OAI21X1_144 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1248_), .C(_abc_65734_new_n1249_), .Y(fracta1_32_));
OAI21X1 OAI21X1_1440 ( .A(u2__abc_52138_new_n4389_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8527_));
OAI21X1 OAI21X1_1441 ( .A(u2__abc_52138_new_n8527_), .B(u2__abc_52138_new_n8526_), .C(u2__abc_52138_new_n8528_), .Y(u2__abc_52138_new_n8529_));
OAI21X1 OAI21X1_1442 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_186_), .Y(u2__abc_52138_new_n8531_));
OAI21X1 OAI21X1_1443 ( .A(u2__abc_52138_new_n4383_), .B(u2__abc_52138_new_n4391_), .C(u2__abc_52138_new_n4388_), .Y(u2__abc_52138_new_n8532_));
OAI21X1 OAI21X1_1444 ( .A(u2__abc_52138_new_n4395_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8538_));
OAI21X1 OAI21X1_1445 ( .A(u2__abc_52138_new_n8538_), .B(u2__abc_52138_new_n8537_), .C(u2__abc_52138_new_n8539_), .Y(u2__abc_52138_new_n8540_));
OAI21X1 OAI21X1_1446 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_187_), .Y(u2__abc_52138_new_n8542_));
OAI21X1 OAI21X1_1447 ( .A(u2__abc_52138_new_n4397_), .B(u2__abc_52138_new_n8543_), .C(u2__abc_52138_new_n4394_), .Y(u2__abc_52138_new_n8544_));
OAI21X1 OAI21X1_1448 ( .A(u2__abc_52138_new_n4400_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8547_));
OAI21X1 OAI21X1_1449 ( .A(u2__abc_52138_new_n8547_), .B(u2__abc_52138_new_n8546_), .C(u2__abc_52138_new_n8548_), .Y(u2__abc_52138_new_n8549_));
OAI21X1 OAI21X1_145 ( .A(\a[112] ), .B(_abc_65734_new_n1248_), .C(_abc_65734_new_n1251_), .Y(fracta1_33_));
OAI21X1 OAI21X1_1450 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_188_), .Y(u2__abc_52138_new_n8551_));
OAI21X1 OAI21X1_1451 ( .A(u2__abc_52138_new_n4394_), .B(u2__abc_52138_new_n4402_), .C(u2__abc_52138_new_n4399_), .Y(u2__abc_52138_new_n8552_));
OAI21X1 OAI21X1_1452 ( .A(u2__abc_52138_new_n4404_), .B(u2__abc_52138_new_n8523_), .C(u2__abc_52138_new_n8553_), .Y(u2__abc_52138_new_n8554_));
OAI21X1 OAI21X1_1453 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n8557_), .Y(u2__abc_52138_new_n8558_));
OAI21X1 OAI21X1_1454 ( .A(u2__abc_52138_new_n4423_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8560_));
OAI21X1 OAI21X1_1455 ( .A(u2__abc_52138_new_n8560_), .B(u2__abc_52138_new_n8559_), .C(u2__abc_52138_new_n8561_), .Y(u2__abc_52138_new_n8562_));
OAI21X1 OAI21X1_1456 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_189_), .Y(u2__abc_52138_new_n8564_));
OAI21X1 OAI21X1_1457 ( .A(u2__abc_52138_new_n4425_), .B(u2__abc_52138_new_n8555_), .C(u2__abc_52138_new_n4422_), .Y(u2__abc_52138_new_n8565_));
OAI21X1 OAI21X1_1458 ( .A(u2__abc_52138_new_n4418_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8568_));
OAI21X1 OAI21X1_1459 ( .A(u2__abc_52138_new_n8568_), .B(u2__abc_52138_new_n8567_), .C(u2__abc_52138_new_n8569_), .Y(u2__abc_52138_new_n8570_));
OAI21X1 OAI21X1_146 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1253_), .C(_abc_65734_new_n1254_), .Y(fracta1_34_));
OAI21X1 OAI21X1_1460 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_190_), .Y(u2__abc_52138_new_n8572_));
OAI21X1 OAI21X1_1461 ( .A(sqrto_187_), .B(u2__abc_52138_new_n4418_), .C(u2__abc_52138_new_n4422_), .Y(u2__abc_52138_new_n8573_));
OAI21X1 OAI21X1_1462 ( .A(u2__abc_52138_new_n8573_), .B(u2__abc_52138_new_n8556_), .C(u2__abc_52138_new_n4419_), .Y(u2__abc_52138_new_n8574_));
OAI21X1 OAI21X1_1463 ( .A(u2__abc_52138_new_n4407_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8577_));
OAI21X1 OAI21X1_1464 ( .A(u2__abc_52138_new_n8577_), .B(u2__abc_52138_new_n8576_), .C(u2__abc_52138_new_n8578_), .Y(u2__abc_52138_new_n8579_));
OAI21X1 OAI21X1_1465 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_191_), .Y(u2__abc_52138_new_n8581_));
OAI21X1 OAI21X1_1466 ( .A(u2__abc_52138_new_n4409_), .B(u2__abc_52138_new_n8574_), .C(u2__abc_52138_new_n4406_), .Y(u2__abc_52138_new_n8582_));
OAI21X1 OAI21X1_1467 ( .A(u2__abc_52138_new_n4412_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8585_));
OAI21X1 OAI21X1_1468 ( .A(u2__abc_52138_new_n8585_), .B(u2__abc_52138_new_n8584_), .C(u2__abc_52138_new_n8586_), .Y(u2__abc_52138_new_n8587_));
OAI21X1 OAI21X1_1469 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_192_), .Y(u2__abc_52138_new_n8589_));
OAI21X1 OAI21X1_147 ( .A(\a[112] ), .B(_abc_65734_new_n1253_), .C(_abc_65734_new_n1256_), .Y(fracta1_35_));
OAI21X1 OAI21X1_1470 ( .A(u2__abc_52138_new_n4416_), .B(u2_remHi_187_), .C(u2__abc_52138_new_n4415_), .Y(u2__abc_52138_new_n8595_));
OAI21X1 OAI21X1_1471 ( .A(u2__abc_52138_new_n8594_), .B(u2__abc_52138_new_n8595_), .C(u2__abc_52138_new_n8597_), .Y(u2__abc_52138_new_n8598_));
OAI21X1 OAI21X1_1472 ( .A(u2__abc_52138_new_n4759_), .B(u2__abc_52138_new_n8254_), .C(u2__abc_52138_new_n8600_), .Y(u2__abc_52138_new_n8601_));
OAI21X1 OAI21X1_1473 ( .A(u2__abc_52138_new_n8590_), .B(u2__abc_52138_new_n7901_), .C(u2__abc_52138_new_n8602_), .Y(u2__abc_52138_new_n8603_));
OAI21X1 OAI21X1_1474 ( .A(u2__abc_52138_new_n4365_), .B(u2__abc_52138_new_n4367_), .C(u2__abc_52138_new_n8604_), .Y(u2__abc_52138_new_n8607_));
OAI21X1 OAI21X1_1475 ( .A(u2__abc_52138_new_n4364_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8610_));
OAI21X1 OAI21X1_1476 ( .A(u2__abc_52138_new_n8610_), .B(u2__abc_52138_new_n8609_), .C(u2__abc_52138_new_n8611_), .Y(u2__abc_52138_new_n8612_));
OAI21X1 OAI21X1_1477 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_193_), .Y(u2__abc_52138_new_n8614_));
OAI21X1 OAI21X1_1478 ( .A(sqrto_190_), .B(u2__abc_52138_new_n4364_), .C(u2__abc_52138_new_n8606_), .Y(u2__abc_52138_new_n8615_));
OAI21X1 OAI21X1_1479 ( .A(u2__abc_52138_new_n4369_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8618_));
OAI21X1 OAI21X1_148 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1258_), .C(_abc_65734_new_n1259_), .Y(fracta1_36_));
OAI21X1 OAI21X1_1480 ( .A(u2__abc_52138_new_n8618_), .B(u2__abc_52138_new_n8617_), .C(u2__abc_52138_new_n8619_), .Y(u2__abc_52138_new_n8620_));
OAI21X1 OAI21X1_1481 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_194_), .Y(u2__abc_52138_new_n8622_));
OAI21X1 OAI21X1_1482 ( .A(u2__abc_52138_new_n4355_), .B(u2__abc_52138_new_n4357_), .C(u2__abc_52138_new_n8623_), .Y(u2__abc_52138_new_n8626_));
OAI21X1 OAI21X1_1483 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n8628_), .C(u2__abc_52138_new_n8629_), .Y(u2__abc_52138_new_n8630_));
OAI21X1 OAI21X1_1484 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_195_), .Y(u2__abc_52138_new_n8632_));
OAI21X1 OAI21X1_1485 ( .A(sqrto_192_), .B(u2__abc_52138_new_n4354_), .C(u2__abc_52138_new_n8625_), .Y(u2__abc_52138_new_n8633_));
OAI21X1 OAI21X1_1486 ( .A(u2__abc_52138_new_n4883_), .B(u2__abc_52138_new_n8633_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8634_));
OAI21X1 OAI21X1_1487 ( .A(u2__abc_52138_new_n4360_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8636_));
OAI21X1 OAI21X1_1488 ( .A(u2__abc_52138_new_n8636_), .B(u2__abc_52138_new_n8635_), .C(u2__abc_52138_new_n8637_), .Y(u2__abc_52138_new_n8638_));
OAI21X1 OAI21X1_1489 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_196_), .Y(u2__abc_52138_new_n8640_));
OAI21X1 OAI21X1_149 ( .A(\a[112] ), .B(_abc_65734_new_n1258_), .C(_abc_65734_new_n1261_), .Y(fracta1_37_));
OAI21X1 OAI21X1_1490 ( .A(u2__abc_52138_new_n4365_), .B(u2__abc_52138_new_n4370_), .C(u2__abc_52138_new_n4374_), .Y(u2__abc_52138_new_n8641_));
OAI21X1 OAI21X1_1491 ( .A(u2__abc_52138_new_n8641_), .B(u2__abc_52138_new_n4884_), .C(u2__abc_52138_new_n8642_), .Y(u2__abc_52138_new_n8643_));
OAI21X1 OAI21X1_1492 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n8646_), .Y(u2__abc_52138_new_n8647_));
OAI21X1 OAI21X1_1493 ( .A(u2__abc_52138_new_n4349_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8649_));
OAI21X1 OAI21X1_1494 ( .A(u2__abc_52138_new_n8649_), .B(u2__abc_52138_new_n8648_), .C(u2__abc_52138_new_n8650_), .Y(u2__abc_52138_new_n8651_));
OAI21X1 OAI21X1_1495 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_197_), .Y(u2__abc_52138_new_n8653_));
OAI21X1 OAI21X1_1496 ( .A(u2__abc_52138_new_n4351_), .B(u2__abc_52138_new_n8644_), .C(u2__abc_52138_new_n4348_), .Y(u2__abc_52138_new_n8655_));
OAI21X1 OAI21X1_1497 ( .A(u2__abc_52138_new_n8654_), .B(u2__abc_52138_new_n8655_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8656_));
OAI21X1 OAI21X1_1498 ( .A(u2__abc_52138_new_n4344_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8658_));
OAI21X1 OAI21X1_1499 ( .A(u2__abc_52138_new_n8658_), .B(u2__abc_52138_new_n8657_), .C(u2__abc_52138_new_n8659_), .Y(u2__abc_52138_new_n8660_));
OAI21X1 OAI21X1_15 ( .A(aNan), .B(_abc_65734_new_n872_), .C(_abc_65734_new_n873_), .Y(\o[126] ));
OAI21X1 OAI21X1_150 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1263_), .C(_abc_65734_new_n1264_), .Y(fracta1_38_));
OAI21X1 OAI21X1_1500 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_198_), .Y(u2__abc_52138_new_n8662_));
OAI21X1 OAI21X1_1501 ( .A(sqrto_195_), .B(u2__abc_52138_new_n4344_), .C(u2__abc_52138_new_n8666_), .Y(u2__abc_52138_new_n8667_));
OAI21X1 OAI21X1_1502 ( .A(u2__abc_52138_new_n4333_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8671_));
OAI21X1 OAI21X1_1503 ( .A(u2_remHi_198_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8673_));
OAI21X1 OAI21X1_1504 ( .A(u2__abc_52138_new_n8673_), .B(u2__abc_52138_new_n8672_), .C(u2__abc_52138_new_n8662_), .Y(u2__abc_52138_new_n8674_));
OAI21X1 OAI21X1_1505 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_199_), .Y(u2__abc_52138_new_n8676_));
OAI21X1 OAI21X1_1506 ( .A(sqrto_196_), .B(u2__abc_52138_new_n4333_), .C(u2__abc_52138_new_n8668_), .Y(u2__abc_52138_new_n8677_));
OAI21X1 OAI21X1_1507 ( .A(u2__abc_52138_new_n4338_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8680_));
OAI21X1 OAI21X1_1508 ( .A(u2__abc_52138_new_n8680_), .B(u2__abc_52138_new_n8679_), .C(u2__abc_52138_new_n8681_), .Y(u2__abc_52138_new_n8682_));
OAI21X1 OAI21X1_1509 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_200_), .Y(u2__abc_52138_new_n8684_));
OAI21X1 OAI21X1_151 ( .A(\a[112] ), .B(_abc_65734_new_n1263_), .C(_abc_65734_new_n1266_), .Y(fracta1_39_));
OAI21X1 OAI21X1_1510 ( .A(u2__abc_52138_new_n4348_), .B(u2__abc_52138_new_n4346_), .C(u2__abc_52138_new_n4343_), .Y(u2__abc_52138_new_n8687_));
OAI21X1 OAI21X1_1511 ( .A(u2__abc_52138_new_n8690_), .B(u2__abc_52138_new_n8691_), .C(u2__abc_52138_new_n8685_), .Y(u2__abc_52138_new_n8692_));
OAI21X1 OAI21X1_1512 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n8696_), .C(u2__abc_52138_new_n8697_), .Y(u2__abc_52138_new_n8698_));
OAI21X1 OAI21X1_1513 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_201_), .Y(u2__abc_52138_new_n8700_));
OAI21X1 OAI21X1_1514 ( .A(sqrto_198_), .B(u2__abc_52138_new_n4307_), .C(u2__abc_52138_new_n8692_), .Y(u2__abc_52138_new_n8701_));
OAI21X1 OAI21X1_1515 ( .A(u2__abc_52138_new_n4302_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8704_));
OAI21X1 OAI21X1_1516 ( .A(u2__abc_52138_new_n8704_), .B(u2__abc_52138_new_n8703_), .C(u2__abc_52138_new_n8705_), .Y(u2__abc_52138_new_n8706_));
OAI21X1 OAI21X1_1517 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_202_), .Y(u2__abc_52138_new_n8708_));
OAI21X1 OAI21X1_1518 ( .A(sqrto_198_), .B(u2__abc_52138_new_n4307_), .C(u2__abc_52138_new_n4301_), .Y(u2__abc_52138_new_n8710_));
OAI21X1 OAI21X1_1519 ( .A(u2__abc_52138_new_n8710_), .B(u2__abc_52138_new_n8709_), .C(u2__abc_52138_new_n4303_), .Y(u2__abc_52138_new_n8711_));
OAI21X1 OAI21X1_152 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1268_), .C(_abc_65734_new_n1269_), .Y(fracta1_40_));
OAI21X1 OAI21X1_1520 ( .A(u2__abc_52138_new_n4291_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8714_));
OAI21X1 OAI21X1_1521 ( .A(u2__abc_52138_new_n8714_), .B(u2__abc_52138_new_n8713_), .C(u2__abc_52138_new_n8715_), .Y(u2__abc_52138_new_n8716_));
OAI21X1 OAI21X1_1522 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_203_), .Y(u2__abc_52138_new_n8718_));
OAI21X1 OAI21X1_1523 ( .A(u2__abc_52138_new_n4293_), .B(u2__abc_52138_new_n8711_), .C(u2__abc_52138_new_n4290_), .Y(u2__abc_52138_new_n8719_));
OAI21X1 OAI21X1_1524 ( .A(u2__abc_52138_new_n4296_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8722_));
OAI21X1 OAI21X1_1525 ( .A(u2__abc_52138_new_n8722_), .B(u2__abc_52138_new_n8721_), .C(u2__abc_52138_new_n8723_), .Y(u2__abc_52138_new_n8724_));
OAI21X1 OAI21X1_1526 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_204_), .Y(u2__abc_52138_new_n8726_));
OAI21X1 OAI21X1_1527 ( .A(u2__abc_52138_new_n4306_), .B(u2__abc_52138_new_n4304_), .C(u2__abc_52138_new_n4301_), .Y(u2__abc_52138_new_n8727_));
OAI21X1 OAI21X1_1528 ( .A(u2__abc_52138_new_n4290_), .B(u2__abc_52138_new_n4298_), .C(u2__abc_52138_new_n4295_), .Y(u2__abc_52138_new_n8728_));
OAI21X1 OAI21X1_1529 ( .A(u2__abc_52138_new_n4311_), .B(u2__abc_52138_new_n8693_), .C(u2__abc_52138_new_n8729_), .Y(u2__abc_52138_new_n8730_));
OAI21X1 OAI21X1_153 ( .A(\a[112] ), .B(_abc_65734_new_n1268_), .C(_abc_65734_new_n1271_), .Y(fracta1_41_));
OAI21X1 OAI21X1_1530 ( .A(u2__abc_52138_new_n4328_), .B(u2__abc_52138_new_n8730_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8733_));
OAI21X1 OAI21X1_1531 ( .A(u2__abc_52138_new_n4905_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8735_));
OAI21X1 OAI21X1_1532 ( .A(u2_remHi_204_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8737_));
OAI21X1 OAI21X1_1533 ( .A(u2__abc_52138_new_n8737_), .B(u2__abc_52138_new_n8736_), .C(u2__abc_52138_new_n8726_), .Y(u2__abc_52138_new_n8738_));
OAI21X1 OAI21X1_1534 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_205_), .Y(u2__abc_52138_new_n8740_));
OAI21X1 OAI21X1_1535 ( .A(sqrto_202_), .B(u2__abc_52138_new_n4905_), .C(u2__abc_52138_new_n8731_), .Y(u2__abc_52138_new_n8741_));
OAI21X1 OAI21X1_1536 ( .A(u2__abc_52138_new_n4323_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8744_));
OAI21X1 OAI21X1_1537 ( .A(u2__abc_52138_new_n8744_), .B(u2__abc_52138_new_n8743_), .C(u2__abc_52138_new_n8745_), .Y(u2__abc_52138_new_n8746_));
OAI21X1 OAI21X1_1538 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_206_), .Y(u2__abc_52138_new_n8748_));
OAI21X1 OAI21X1_1539 ( .A(sqrto_202_), .B(u2__abc_52138_new_n4905_), .C(u2__abc_52138_new_n8749_), .Y(u2__abc_52138_new_n8750_));
OAI21X1 OAI21X1_154 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1273_), .C(_abc_65734_new_n1274_), .Y(fracta1_42_));
OAI21X1 OAI21X1_1540 ( .A(u2__abc_52138_new_n8750_), .B(u2__abc_52138_new_n8732_), .C(u2__abc_52138_new_n4904_), .Y(u2__abc_52138_new_n8751_));
OAI21X1 OAI21X1_1541 ( .A(u2__abc_52138_new_n4314_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8754_));
OAI21X1 OAI21X1_1542 ( .A(u2__abc_52138_new_n8754_), .B(u2__abc_52138_new_n8753_), .C(u2__abc_52138_new_n8755_), .Y(u2__abc_52138_new_n8756_));
OAI21X1 OAI21X1_1543 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_207_), .Y(u2__abc_52138_new_n8758_));
OAI21X1 OAI21X1_1544 ( .A(u2__abc_52138_new_n4316_), .B(u2__abc_52138_new_n8751_), .C(u2__abc_52138_new_n4313_), .Y(u2__abc_52138_new_n8759_));
OAI21X1 OAI21X1_1545 ( .A(u2__abc_52138_new_n4319_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8762_));
OAI21X1 OAI21X1_1546 ( .A(u2__abc_52138_new_n8762_), .B(u2__abc_52138_new_n8761_), .C(u2__abc_52138_new_n8763_), .Y(u2__abc_52138_new_n8764_));
OAI21X1 OAI21X1_1547 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_208_), .Y(u2__abc_52138_new_n8766_));
OAI21X1 OAI21X1_1548 ( .A(u2__abc_52138_new_n4313_), .B(u2__abc_52138_new_n4321_), .C(u2__abc_52138_new_n4318_), .Y(u2__abc_52138_new_n8771_));
OAI21X1 OAI21X1_1549 ( .A(u2__abc_52138_new_n4329_), .B(u2__abc_52138_new_n8729_), .C(u2__abc_52138_new_n8773_), .Y(u2__abc_52138_new_n8774_));
OAI21X1 OAI21X1_155 ( .A(\a[112] ), .B(_abc_65734_new_n1273_), .C(_abc_65734_new_n1276_), .Y(fracta1_43_));
OAI21X1 OAI21X1_1550 ( .A(u2__abc_52138_new_n8774_), .B(u2__abc_52138_new_n8775_), .C(u2__abc_52138_new_n8767_), .Y(u2__abc_52138_new_n8776_));
OAI21X1 OAI21X1_1551 ( .A(u2__abc_52138_new_n4254_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8779_));
OAI21X1 OAI21X1_1552 ( .A(u2_remHi_208_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8781_));
OAI21X1 OAI21X1_1553 ( .A(u2__abc_52138_new_n8781_), .B(u2__abc_52138_new_n8780_), .C(u2__abc_52138_new_n8766_), .Y(u2__abc_52138_new_n8782_));
OAI21X1 OAI21X1_1554 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_209_), .Y(u2__abc_52138_new_n8784_));
OAI21X1 OAI21X1_1555 ( .A(sqrto_206_), .B(u2__abc_52138_new_n4254_), .C(u2__abc_52138_new_n8776_), .Y(u2__abc_52138_new_n8785_));
OAI21X1 OAI21X1_1556 ( .A(u2__abc_52138_new_n4259_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8788_));
OAI21X1 OAI21X1_1557 ( .A(u2__abc_52138_new_n8788_), .B(u2__abc_52138_new_n8787_), .C(u2__abc_52138_new_n8789_), .Y(u2__abc_52138_new_n8790_));
OAI21X1 OAI21X1_1558 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_210_), .Y(u2__abc_52138_new_n8792_));
OAI21X1 OAI21X1_1559 ( .A(u2__abc_52138_new_n4915_), .B(u2__abc_52138_new_n8793_), .C(u2__abc_52138_new_n4258_), .Y(u2__abc_52138_new_n8794_));
OAI21X1 OAI21X1_156 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1278_), .C(_abc_65734_new_n1279_), .Y(fracta1_44_));
OAI21X1 OAI21X1_1560 ( .A(u2__abc_52138_new_n4243_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8797_));
OAI21X1 OAI21X1_1561 ( .A(u2__abc_52138_new_n8797_), .B(u2__abc_52138_new_n8796_), .C(u2__abc_52138_new_n8798_), .Y(u2__abc_52138_new_n8799_));
OAI21X1 OAI21X1_1562 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_211_), .Y(u2__abc_52138_new_n8801_));
OAI21X1 OAI21X1_1563 ( .A(sqrto_208_), .B(u2__abc_52138_new_n4243_), .C(u2__abc_52138_new_n8802_), .Y(u2__abc_52138_new_n8803_));
OAI21X1 OAI21X1_1564 ( .A(u2__abc_52138_new_n4248_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8806_));
OAI21X1 OAI21X1_1565 ( .A(u2__abc_52138_new_n8806_), .B(u2__abc_52138_new_n8805_), .C(u2__abc_52138_new_n8807_), .Y(u2__abc_52138_new_n8808_));
OAI21X1 OAI21X1_1566 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_212_), .Y(u2__abc_52138_new_n8810_));
OAI21X1 OAI21X1_1567 ( .A(u2__abc_52138_new_n4253_), .B(u2__abc_52138_new_n4261_), .C(u2__abc_52138_new_n4258_), .Y(u2__abc_52138_new_n8812_));
OAI21X1 OAI21X1_1568 ( .A(u2__abc_52138_new_n4242_), .B(u2__abc_52138_new_n4918_), .C(u2__abc_52138_new_n4247_), .Y(u2__abc_52138_new_n8813_));
OAI21X1 OAI21X1_1569 ( .A(u2__abc_52138_new_n8774_), .B(u2__abc_52138_new_n8775_), .C(u2__abc_52138_new_n4263_), .Y(u2__abc_52138_new_n8815_));
OAI21X1 OAI21X1_157 ( .A(\a[112] ), .B(_abc_65734_new_n1278_), .C(_abc_65734_new_n1281_), .Y(fracta1_45_));
OAI21X1 OAI21X1_1570 ( .A(u2__abc_52138_new_n4280_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8820_));
OAI21X1 OAI21X1_1571 ( .A(u2_remHi_212_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8822_));
OAI21X1 OAI21X1_1572 ( .A(u2__abc_52138_new_n8822_), .B(u2__abc_52138_new_n8821_), .C(u2__abc_52138_new_n8810_), .Y(u2__abc_52138_new_n8823_));
OAI21X1 OAI21X1_1573 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_213_), .Y(u2__abc_52138_new_n8825_));
OAI21X1 OAI21X1_1574 ( .A(sqrto_210_), .B(u2__abc_52138_new_n4280_), .C(u2__abc_52138_new_n8817_), .Y(u2__abc_52138_new_n8826_));
OAI21X1 OAI21X1_1575 ( .A(u2__abc_52138_new_n4279_), .B(u2__abc_52138_new_n8826_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8827_));
OAI21X1 OAI21X1_1576 ( .A(u2__abc_52138_new_n4275_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8829_));
OAI21X1 OAI21X1_1577 ( .A(u2__abc_52138_new_n8829_), .B(u2__abc_52138_new_n8828_), .C(u2__abc_52138_new_n8830_), .Y(u2__abc_52138_new_n8831_));
OAI21X1 OAI21X1_1578 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_214_), .Y(u2__abc_52138_new_n8833_));
OAI21X1 OAI21X1_1579 ( .A(sqrto_211_), .B(u2__abc_52138_new_n4275_), .C(u2__abc_52138_new_n8834_), .Y(u2__abc_52138_new_n8835_));
OAI21X1 OAI21X1_158 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1283_), .C(_abc_65734_new_n1284_), .Y(fracta1_46_));
OAI21X1 OAI21X1_1580 ( .A(u2__abc_52138_new_n4268_), .B(u2__abc_52138_new_n8835_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8836_));
OAI21X1 OAI21X1_1581 ( .A(u2__abc_52138_new_n4264_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8838_));
OAI21X1 OAI21X1_1582 ( .A(u2__abc_52138_new_n8838_), .B(u2__abc_52138_new_n8837_), .C(u2__abc_52138_new_n8839_), .Y(u2__abc_52138_new_n8840_));
OAI21X1 OAI21X1_1583 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_215_), .Y(u2__abc_52138_new_n8842_));
OAI21X1 OAI21X1_1584 ( .A(u2__abc_52138_new_n4269_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8846_));
OAI21X1 OAI21X1_1585 ( .A(u2__abc_52138_new_n8846_), .B(u2__abc_52138_new_n8845_), .C(u2__abc_52138_new_n8847_), .Y(u2__abc_52138_new_n8848_));
OAI21X1 OAI21X1_1586 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_216_), .Y(u2__abc_52138_new_n8850_));
OAI21X1 OAI21X1_1587 ( .A(u2__abc_52138_new_n4278_), .B(u2__abc_52138_new_n8852_), .C(u2__abc_52138_new_n4921_), .Y(u2__abc_52138_new_n8853_));
OAI21X1 OAI21X1_1588 ( .A(u2__abc_52138_new_n8814_), .B(u2__abc_52138_new_n8854_), .C(u2__abc_52138_new_n8855_), .Y(u2__abc_52138_new_n8856_));
OAI21X1 OAI21X1_1589 ( .A(u2__abc_52138_new_n4287_), .B(u2__abc_52138_new_n8777_), .C(u2__abc_52138_new_n8857_), .Y(u2__abc_52138_new_n8858_));
OAI21X1 OAI21X1_159 ( .A(\a[112] ), .B(_abc_65734_new_n1283_), .C(_abc_65734_new_n1286_), .Y(fracta1_47_));
OAI21X1 OAI21X1_1590 ( .A(u2__abc_52138_new_n4207_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8860_));
OAI21X1 OAI21X1_1591 ( .A(u2_remHi_216_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8862_));
OAI21X1 OAI21X1_1592 ( .A(u2__abc_52138_new_n8862_), .B(u2__abc_52138_new_n8861_), .C(u2__abc_52138_new_n8850_), .Y(u2__abc_52138_new_n8863_));
OAI21X1 OAI21X1_1593 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_217_), .Y(u2__abc_52138_new_n8865_));
OAI21X1 OAI21X1_1594 ( .A(u2__abc_52138_new_n4209_), .B(u2__abc_52138_new_n8866_), .C(u2__abc_52138_new_n4206_), .Y(u2__abc_52138_new_n8867_));
OAI21X1 OAI21X1_1595 ( .A(u2__abc_52138_new_n4212_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8870_));
OAI21X1 OAI21X1_1596 ( .A(u2__abc_52138_new_n8870_), .B(u2__abc_52138_new_n8869_), .C(u2__abc_52138_new_n8871_), .Y(u2__abc_52138_new_n8872_));
OAI21X1 OAI21X1_1597 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_218_), .Y(u2__abc_52138_new_n8874_));
OAI21X1 OAI21X1_1598 ( .A(u2__abc_52138_new_n4206_), .B(u2__abc_52138_new_n4214_), .C(u2__abc_52138_new_n4211_), .Y(u2__abc_52138_new_n8875_));
OAI21X1 OAI21X1_1599 ( .A(u2__abc_52138_new_n4215_), .B(u2__abc_52138_new_n8866_), .C(u2__abc_52138_new_n8876_), .Y(u2__abc_52138_new_n8877_));
OAI21X1 OAI21X1_16 ( .A(aNan), .B(_abc_65734_new_n875_), .C(_abc_65734_new_n876_), .Y(\o[127] ));
OAI21X1 OAI21X1_160 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1288_), .C(_abc_65734_new_n1289_), .Y(fracta1_48_));
OAI21X1 OAI21X1_1600 ( .A(u2__abc_52138_new_n4196_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8880_));
OAI21X1 OAI21X1_1601 ( .A(u2__abc_52138_new_n8880_), .B(u2__abc_52138_new_n8879_), .C(u2__abc_52138_new_n8881_), .Y(u2__abc_52138_new_n8882_));
OAI21X1 OAI21X1_1602 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_219_), .Y(u2__abc_52138_new_n8884_));
OAI21X1 OAI21X1_1603 ( .A(u2__abc_52138_new_n4198_), .B(u2__abc_52138_new_n8885_), .C(u2__abc_52138_new_n4195_), .Y(u2__abc_52138_new_n8886_));
OAI21X1 OAI21X1_1604 ( .A(u2__abc_52138_new_n4201_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8889_));
OAI21X1 OAI21X1_1605 ( .A(u2__abc_52138_new_n8889_), .B(u2__abc_52138_new_n8888_), .C(u2__abc_52138_new_n8890_), .Y(u2__abc_52138_new_n8891_));
OAI21X1 OAI21X1_1606 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_220_), .Y(u2__abc_52138_new_n8893_));
OAI21X1 OAI21X1_1607 ( .A(u2__abc_52138_new_n4195_), .B(u2__abc_52138_new_n4203_), .C(u2__abc_52138_new_n4200_), .Y(u2__abc_52138_new_n8896_));
OAI21X1 OAI21X1_1608 ( .A(u2__abc_52138_new_n8895_), .B(u2__abc_52138_new_n8866_), .C(u2__abc_52138_new_n8897_), .Y(u2__abc_52138_new_n8898_));
OAI21X1 OAI21X1_1609 ( .A(u2__abc_52138_new_n4237_), .B(u2__abc_52138_new_n8898_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8901_));
OAI21X1 OAI21X1_161 ( .A(\a[112] ), .B(_abc_65734_new_n1288_), .C(_abc_65734_new_n1291_), .Y(fracta1_49_));
OAI21X1 OAI21X1_1610 ( .A(u2__abc_52138_new_n4235_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8903_));
OAI21X1 OAI21X1_1611 ( .A(u2__abc_52138_new_n8903_), .B(u2__abc_52138_new_n8902_), .C(u2__abc_52138_new_n8904_), .Y(u2__abc_52138_new_n8905_));
OAI21X1 OAI21X1_1612 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_221_), .Y(u2__abc_52138_new_n8907_));
OAI21X1 OAI21X1_1613 ( .A(u2__abc_52138_new_n8894_), .B(u2__abc_52138_new_n8899_), .C(u2__abc_52138_new_n4234_), .Y(u2__abc_52138_new_n8908_));
OAI21X1 OAI21X1_1614 ( .A(u2__abc_52138_new_n4228_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8911_));
OAI21X1 OAI21X1_1615 ( .A(u2__abc_52138_new_n8911_), .B(u2__abc_52138_new_n8910_), .C(u2__abc_52138_new_n8912_), .Y(u2__abc_52138_new_n8913_));
OAI21X1 OAI21X1_1616 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_222_), .Y(u2__abc_52138_new_n8915_));
OAI21X1 OAI21X1_1617 ( .A(sqrto_219_), .B(u2__abc_52138_new_n4228_), .C(u2__abc_52138_new_n4234_), .Y(u2__abc_52138_new_n8916_));
OAI21X1 OAI21X1_1618 ( .A(u2__abc_52138_new_n4230_), .B(u2_remHi_219_), .C(u2__abc_52138_new_n8916_), .Y(u2__abc_52138_new_n8917_));
OAI21X1 OAI21X1_1619 ( .A(u2__abc_52138_new_n4238_), .B(u2__abc_52138_new_n8899_), .C(u2__abc_52138_new_n8917_), .Y(u2__abc_52138_new_n8918_));
OAI21X1 OAI21X1_162 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1293_), .C(_abc_65734_new_n1294_), .Y(fracta1_50_));
OAI21X1 OAI21X1_1620 ( .A(u2__abc_52138_new_n4219_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8921_));
OAI21X1 OAI21X1_1621 ( .A(u2__abc_52138_new_n8921_), .B(u2__abc_52138_new_n8920_), .C(u2__abc_52138_new_n8922_), .Y(u2__abc_52138_new_n8923_));
OAI21X1 OAI21X1_1622 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_223_), .Y(u2__abc_52138_new_n8925_));
OAI21X1 OAI21X1_1623 ( .A(u2__abc_52138_new_n4224_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8930_));
OAI21X1 OAI21X1_1624 ( .A(u2__abc_52138_new_n8930_), .B(u2__abc_52138_new_n8929_), .C(u2__abc_52138_new_n8931_), .Y(u2__abc_52138_new_n8932_));
OAI21X1 OAI21X1_1625 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_224_), .Y(u2__abc_52138_new_n8934_));
OAI21X1 OAI21X1_1626 ( .A(u2__abc_52138_new_n8926_), .B(u2__abc_52138_new_n4935_), .C(u2__abc_52138_new_n4225_), .Y(u2__abc_52138_new_n8937_));
OAI21X1 OAI21X1_1627 ( .A(u2__abc_52138_new_n8942_), .B(u2__abc_52138_new_n8943_), .C(u2__abc_52138_new_n8935_), .Y(u2__abc_52138_new_n8944_));
OAI21X1 OAI21X1_1628 ( .A(u2__abc_52138_new_n8935_), .B(u2__abc_52138_new_n8947_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8948_));
OAI21X1 OAI21X1_1629 ( .A(u2__abc_52138_new_n4164_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8950_));
OAI21X1 OAI21X1_163 ( .A(\a[112] ), .B(_abc_65734_new_n1293_), .C(_abc_65734_new_n1296_), .Y(fracta1_51_));
OAI21X1 OAI21X1_1630 ( .A(u2__abc_52138_new_n8950_), .B(u2__abc_52138_new_n8949_), .C(u2__abc_52138_new_n8951_), .Y(u2__abc_52138_new_n8952_));
OAI21X1 OAI21X1_1631 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_225_), .Y(u2__abc_52138_new_n8954_));
OAI21X1 OAI21X1_1632 ( .A(sqrto_222_), .B(u2__abc_52138_new_n4164_), .C(u2__abc_52138_new_n8944_), .Y(u2__abc_52138_new_n8955_));
OAI21X1 OAI21X1_1633 ( .A(u2__abc_52138_new_n4159_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8958_));
OAI21X1 OAI21X1_1634 ( .A(u2__abc_52138_new_n8958_), .B(u2__abc_52138_new_n8957_), .C(u2__abc_52138_new_n8959_), .Y(u2__abc_52138_new_n8960_));
OAI21X1 OAI21X1_1635 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_226_), .Y(u2__abc_52138_new_n8962_));
OAI21X1 OAI21X1_1636 ( .A(u2__abc_52138_new_n4163_), .B(u2__abc_52138_new_n4161_), .C(u2__abc_52138_new_n4158_), .Y(u2__abc_52138_new_n8963_));
OAI21X1 OAI21X1_1637 ( .A(u2__abc_52138_new_n4148_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8967_));
OAI21X1 OAI21X1_1638 ( .A(u2__abc_52138_new_n8967_), .B(u2__abc_52138_new_n8966_), .C(u2__abc_52138_new_n8968_), .Y(u2__abc_52138_new_n8969_));
OAI21X1 OAI21X1_1639 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_227_), .Y(u2__abc_52138_new_n8971_));
OAI21X1 OAI21X1_164 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1298_), .C(_abc_65734_new_n1299_), .Y(fracta1_52_));
OAI21X1 OAI21X1_1640 ( .A(u2__abc_52138_new_n4150_), .B(u2__abc_52138_new_n8964_), .C(u2__abc_52138_new_n4147_), .Y(u2__abc_52138_new_n8972_));
OAI21X1 OAI21X1_1641 ( .A(u2__abc_52138_new_n4153_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8975_));
OAI21X1 OAI21X1_1642 ( .A(u2__abc_52138_new_n8975_), .B(u2__abc_52138_new_n8974_), .C(u2__abc_52138_new_n8976_), .Y(u2__abc_52138_new_n8977_));
OAI21X1 OAI21X1_1643 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_228_), .Y(u2__abc_52138_new_n8979_));
OAI21X1 OAI21X1_1644 ( .A(u2__abc_52138_new_n4147_), .B(u2__abc_52138_new_n4155_), .C(u2__abc_52138_new_n4152_), .Y(u2__abc_52138_new_n8980_));
OAI21X1 OAI21X1_1645 ( .A(u2__abc_52138_new_n4168_), .B(u2__abc_52138_new_n8946_), .C(u2__abc_52138_new_n8981_), .Y(u2__abc_52138_new_n8982_));
OAI21X1 OAI21X1_1646 ( .A(u2__abc_52138_new_n4189_), .B(u2__abc_52138_new_n8982_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n8985_));
OAI21X1 OAI21X1_1647 ( .A(u2__abc_52138_new_n4185_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8987_));
OAI21X1 OAI21X1_1648 ( .A(u2_remHi_228_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n8989_));
OAI21X1 OAI21X1_1649 ( .A(u2__abc_52138_new_n8989_), .B(u2__abc_52138_new_n8988_), .C(u2__abc_52138_new_n8979_), .Y(u2__abc_52138_new_n8990_));
OAI21X1 OAI21X1_165 ( .A(\a[112] ), .B(_abc_65734_new_n1298_), .C(_abc_65734_new_n1301_), .Y(fracta1_53_));
OAI21X1 OAI21X1_1650 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_229_), .Y(u2__abc_52138_new_n8992_));
OAI21X1 OAI21X1_1651 ( .A(u2_o_226_), .B(u2__abc_52138_new_n4185_), .C(u2__abc_52138_new_n8983_), .Y(u2__abc_52138_new_n8993_));
OAI21X1 OAI21X1_1652 ( .A(u2__abc_52138_new_n4180_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n8996_));
OAI21X1 OAI21X1_1653 ( .A(u2__abc_52138_new_n8996_), .B(u2__abc_52138_new_n8995_), .C(u2__abc_52138_new_n8997_), .Y(u2__abc_52138_new_n8998_));
OAI21X1 OAI21X1_1654 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_230_), .Y(u2__abc_52138_new_n9000_));
OAI21X1 OAI21X1_1655 ( .A(u2__abc_52138_new_n9002_), .B(u2__abc_52138_new_n8984_), .C(u2__abc_52138_new_n9001_), .Y(u2__abc_52138_new_n9003_));
OAI21X1 OAI21X1_1656 ( .A(u2__abc_52138_new_n4171_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9006_));
OAI21X1 OAI21X1_1657 ( .A(u2__abc_52138_new_n9006_), .B(u2__abc_52138_new_n9005_), .C(u2__abc_52138_new_n9007_), .Y(u2__abc_52138_new_n9008_));
OAI21X1 OAI21X1_1658 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_231_), .Y(u2__abc_52138_new_n9010_));
OAI21X1 OAI21X1_1659 ( .A(u2__abc_52138_new_n4173_), .B(u2__abc_52138_new_n9003_), .C(u2__abc_52138_new_n4170_), .Y(u2__abc_52138_new_n9011_));
OAI21X1 OAI21X1_166 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1303_), .C(_abc_65734_new_n1304_), .Y(fracta1_54_));
OAI21X1 OAI21X1_1660 ( .A(u2__abc_52138_new_n4176_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9014_));
OAI21X1 OAI21X1_1661 ( .A(u2__abc_52138_new_n9014_), .B(u2__abc_52138_new_n9013_), .C(u2__abc_52138_new_n9015_), .Y(u2__abc_52138_new_n9016_));
OAI21X1 OAI21X1_1662 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_232_), .Y(u2__abc_52138_new_n9018_));
OAI21X1 OAI21X1_1663 ( .A(u2__abc_52138_new_n4190_), .B(u2__abc_52138_new_n8981_), .C(u2__abc_52138_new_n9021_), .Y(u2__abc_52138_new_n9022_));
OAI21X1 OAI21X1_1664 ( .A(u2__abc_52138_new_n4191_), .B(u2__abc_52138_new_n8946_), .C(u2__abc_52138_new_n9023_), .Y(u2__abc_52138_new_n9024_));
OAI21X1 OAI21X1_1665 ( .A(u2__abc_52138_new_n4138_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9028_));
OAI21X1 OAI21X1_1666 ( .A(u2_remHi_232_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n9030_));
OAI21X1 OAI21X1_1667 ( .A(u2__abc_52138_new_n9030_), .B(u2__abc_52138_new_n9029_), .C(u2__abc_52138_new_n9018_), .Y(u2__abc_52138_new_n9031_));
OAI21X1 OAI21X1_1668 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_233_), .Y(u2__abc_52138_new_n9033_));
OAI21X1 OAI21X1_1669 ( .A(u2_o_230_), .B(u2__abc_52138_new_n4138_), .C(u2__abc_52138_new_n9025_), .Y(u2__abc_52138_new_n9035_));
OAI21X1 OAI21X1_167 ( .A(\a[112] ), .B(_abc_65734_new_n1303_), .C(_abc_65734_new_n1306_), .Y(fracta1_55_));
OAI21X1 OAI21X1_1670 ( .A(u2__abc_52138_new_n4134_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9038_));
OAI21X1 OAI21X1_1671 ( .A(u2__abc_52138_new_n9038_), .B(u2__abc_52138_new_n9037_), .C(u2__abc_52138_new_n9039_), .Y(u2__abc_52138_new_n9040_));
OAI21X1 OAI21X1_1672 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_234_), .Y(u2__abc_52138_new_n9042_));
OAI21X1 OAI21X1_1673 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n9045_), .Y(u2__abc_52138_new_n9046_));
OAI21X1 OAI21X1_1674 ( .A(u2__abc_52138_new_n4125_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9048_));
OAI21X1 OAI21X1_1675 ( .A(u2__abc_52138_new_n9048_), .B(u2__abc_52138_new_n9047_), .C(u2__abc_52138_new_n9049_), .Y(u2__abc_52138_new_n9050_));
OAI21X1 OAI21X1_1676 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_235_), .Y(u2__abc_52138_new_n9052_));
OAI21X1 OAI21X1_1677 ( .A(u2__abc_52138_new_n4127_), .B(u2__abc_52138_new_n9043_), .C(u2__abc_52138_new_n4124_), .Y(u2__abc_52138_new_n9053_));
OAI21X1 OAI21X1_1678 ( .A(u2__abc_52138_new_n4130_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9056_));
OAI21X1 OAI21X1_1679 ( .A(u2__abc_52138_new_n9056_), .B(u2__abc_52138_new_n9055_), .C(u2__abc_52138_new_n9057_), .Y(u2__abc_52138_new_n9058_));
OAI21X1 OAI21X1_168 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1308_), .C(_abc_65734_new_n1309_), .Y(fracta1_56_));
OAI21X1 OAI21X1_1680 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_236_), .Y(u2__abc_52138_new_n9060_));
OAI21X1 OAI21X1_1681 ( .A(u2_o_233_), .B(u2__abc_52138_new_n4130_), .C(u2__abc_52138_new_n4124_), .Y(u2__abc_52138_new_n9061_));
OAI21X1 OAI21X1_1682 ( .A(u2__abc_52138_new_n9061_), .B(u2__abc_52138_new_n9044_), .C(u2__abc_52138_new_n4131_), .Y(u2__abc_52138_new_n9062_));
OAI21X1 OAI21X1_1683 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n9064_), .Y(u2__abc_52138_new_n9065_));
OAI21X1 OAI21X1_1684 ( .A(u2__abc_52138_new_n4117_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9067_));
OAI21X1 OAI21X1_1685 ( .A(u2__abc_52138_new_n9067_), .B(u2__abc_52138_new_n9066_), .C(u2__abc_52138_new_n9068_), .Y(u2__abc_52138_new_n9069_));
OAI21X1 OAI21X1_1686 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_237_), .Y(u2__abc_52138_new_n9071_));
OAI21X1 OAI21X1_1687 ( .A(u2__abc_52138_new_n4119_), .B(u2__abc_52138_new_n9062_), .C(u2__abc_52138_new_n4116_), .Y(u2__abc_52138_new_n9072_));
OAI21X1 OAI21X1_1688 ( .A(u2__abc_52138_new_n4112_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9075_));
OAI21X1 OAI21X1_1689 ( .A(u2__abc_52138_new_n9075_), .B(u2__abc_52138_new_n9074_), .C(u2__abc_52138_new_n9076_), .Y(u2__abc_52138_new_n9077_));
OAI21X1 OAI21X1_169 ( .A(\a[112] ), .B(_abc_65734_new_n1308_), .C(_abc_65734_new_n1311_), .Y(fracta1_57_));
OAI21X1 OAI21X1_1690 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_238_), .Y(u2__abc_52138_new_n9079_));
OAI21X1 OAI21X1_1691 ( .A(u2_o_235_), .B(u2__abc_52138_new_n4112_), .C(u2__abc_52138_new_n4116_), .Y(u2__abc_52138_new_n9080_));
OAI21X1 OAI21X1_1692 ( .A(u2__abc_52138_new_n9080_), .B(u2__abc_52138_new_n9063_), .C(u2__abc_52138_new_n4113_), .Y(u2__abc_52138_new_n9081_));
OAI21X1 OAI21X1_1693 ( .A(u2__abc_52138_new_n4101_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9084_));
OAI21X1 OAI21X1_1694 ( .A(u2__abc_52138_new_n9084_), .B(u2__abc_52138_new_n9083_), .C(u2__abc_52138_new_n9085_), .Y(u2__abc_52138_new_n9086_));
OAI21X1 OAI21X1_1695 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_239_), .Y(u2__abc_52138_new_n9088_));
OAI21X1 OAI21X1_1696 ( .A(u2__abc_52138_new_n4103_), .B(u2__abc_52138_new_n9081_), .C(u2__abc_52138_new_n4100_), .Y(u2__abc_52138_new_n9089_));
OAI21X1 OAI21X1_1697 ( .A(u2__abc_52138_new_n4106_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9092_));
OAI21X1 OAI21X1_1698 ( .A(u2__abc_52138_new_n9092_), .B(u2__abc_52138_new_n9091_), .C(u2__abc_52138_new_n9093_), .Y(u2__abc_52138_new_n9094_));
OAI21X1 OAI21X1_1699 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_240_), .Y(u2__abc_52138_new_n9096_));
OAI21X1 OAI21X1_17 ( .A(aNan), .B(_abc_65734_new_n878_), .C(_abc_65734_new_n879_), .Y(\o[128] ));
OAI21X1 OAI21X1_170 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1313_), .C(_abc_65734_new_n1314_), .Y(fracta1_58_));
OAI21X1 OAI21X1_1700 ( .A(u2__abc_52138_new_n4100_), .B(u2__abc_52138_new_n4108_), .C(u2__abc_52138_new_n4105_), .Y(u2__abc_52138_new_n9097_));
OAI21X1 OAI21X1_1701 ( .A(u2__abc_52138_new_n4135_), .B(u2__abc_52138_new_n4139_), .C(u2__abc_52138_new_n4137_), .Y(u2__abc_52138_new_n9098_));
OAI21X1 OAI21X1_1702 ( .A(u2__abc_52138_new_n4128_), .B(u2_remHi_233_), .C(u2__abc_52138_new_n9061_), .Y(u2__abc_52138_new_n9099_));
OAI21X1 OAI21X1_1703 ( .A(u2__abc_52138_new_n9098_), .B(u2__abc_52138_new_n4133_), .C(u2__abc_52138_new_n9099_), .Y(u2__abc_52138_new_n9100_));
OAI21X1 OAI21X1_1704 ( .A(u2__abc_52138_new_n4110_), .B(u2_remHi_235_), .C(u2__abc_52138_new_n9080_), .Y(u2__abc_52138_new_n9101_));
OAI21X1 OAI21X1_1705 ( .A(u2__abc_52138_new_n4145_), .B(u2__abc_52138_new_n9023_), .C(u2__abc_52138_new_n9103_), .Y(u2__abc_52138_new_n9104_));
OAI21X1 OAI21X1_1706 ( .A(u2__abc_52138_new_n8942_), .B(u2__abc_52138_new_n8943_), .C(u2__abc_52138_new_n4192_), .Y(u2__abc_52138_new_n9106_));
OAI21X1 OAI21X1_1707 ( .A(u2__abc_52138_new_n4052_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9110_));
OAI21X1 OAI21X1_1708 ( .A(u2__abc_52138_new_n9110_), .B(u2__abc_52138_new_n9109_), .C(u2__abc_52138_new_n9111_), .Y(u2__abc_52138_new_n9112_));
OAI21X1 OAI21X1_1709 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_241_), .Y(u2__abc_52138_new_n9114_));
OAI21X1 OAI21X1_171 ( .A(\a[112] ), .B(_abc_65734_new_n1313_), .C(_abc_65734_new_n1316_), .Y(fracta1_59_));
OAI21X1 OAI21X1_1710 ( .A(u2__abc_52138_new_n4054_), .B(u2__abc_52138_new_n9115_), .C(u2__abc_52138_new_n4051_), .Y(u2__abc_52138_new_n9116_));
OAI21X1 OAI21X1_1711 ( .A(u2__abc_52138_new_n4057_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9119_));
OAI21X1 OAI21X1_1712 ( .A(u2__abc_52138_new_n9119_), .B(u2__abc_52138_new_n9118_), .C(u2__abc_52138_new_n9120_), .Y(u2__abc_52138_new_n9121_));
OAI21X1 OAI21X1_1713 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_242_), .Y(u2__abc_52138_new_n9123_));
OAI21X1 OAI21X1_1714 ( .A(u2__abc_52138_new_n4051_), .B(u2__abc_52138_new_n4059_), .C(u2__abc_52138_new_n4056_), .Y(u2__abc_52138_new_n9124_));
OAI21X1 OAI21X1_1715 ( .A(u2__abc_52138_new_n4060_), .B(u2__abc_52138_new_n9115_), .C(u2__abc_52138_new_n9125_), .Y(u2__abc_52138_new_n9126_));
OAI21X1 OAI21X1_1716 ( .A(u2__abc_52138_new_n4063_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9129_));
OAI21X1 OAI21X1_1717 ( .A(u2__abc_52138_new_n9129_), .B(u2__abc_52138_new_n9128_), .C(u2__abc_52138_new_n9130_), .Y(u2__abc_52138_new_n9131_));
OAI21X1 OAI21X1_1718 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_243_), .Y(u2__abc_52138_new_n9133_));
OAI21X1 OAI21X1_1719 ( .A(u2__abc_52138_new_n4065_), .B(u2__abc_52138_new_n9134_), .C(u2__abc_52138_new_n4062_), .Y(u2__abc_52138_new_n9135_));
OAI21X1 OAI21X1_172 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1318_), .C(_abc_65734_new_n1319_), .Y(fracta1_60_));
OAI21X1 OAI21X1_1720 ( .A(u2__abc_52138_new_n4068_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9138_));
OAI21X1 OAI21X1_1721 ( .A(u2__abc_52138_new_n9138_), .B(u2__abc_52138_new_n9137_), .C(u2__abc_52138_new_n9139_), .Y(u2__abc_52138_new_n9140_));
OAI21X1 OAI21X1_1722 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_244_), .Y(u2__abc_52138_new_n9142_));
OAI21X1 OAI21X1_1723 ( .A(u2__abc_52138_new_n4062_), .B(u2__abc_52138_new_n4070_), .C(u2__abc_52138_new_n4067_), .Y(u2__abc_52138_new_n9144_));
OAI21X1 OAI21X1_1724 ( .A(u2__abc_52138_new_n4092_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9150_));
OAI21X1 OAI21X1_1725 ( .A(u2__abc_52138_new_n9150_), .B(u2__abc_52138_new_n9149_), .C(u2__abc_52138_new_n9151_), .Y(u2__abc_52138_new_n9152_));
OAI21X1 OAI21X1_1726 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_245_), .Y(u2__abc_52138_new_n9154_));
OAI21X1 OAI21X1_1727 ( .A(u2__abc_52138_new_n9143_), .B(u2__abc_52138_new_n9147_), .C(u2__abc_52138_new_n4091_), .Y(u2__abc_52138_new_n9155_));
OAI21X1 OAI21X1_1728 ( .A(u2__abc_52138_new_n4089_), .B(u2__abc_52138_new_n9155_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9156_));
OAI21X1 OAI21X1_1729 ( .A(u2__abc_52138_new_n4085_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9158_));
OAI21X1 OAI21X1_173 ( .A(\a[112] ), .B(_abc_65734_new_n1318_), .C(_abc_65734_new_n1321_), .Y(fracta1_61_));
OAI21X1 OAI21X1_1730 ( .A(u2__abc_52138_new_n9158_), .B(u2__abc_52138_new_n9157_), .C(u2__abc_52138_new_n9159_), .Y(u2__abc_52138_new_n9160_));
OAI21X1 OAI21X1_1731 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_246_), .Y(u2__abc_52138_new_n9162_));
OAI21X1 OAI21X1_1732 ( .A(u2_o_243_), .B(u2__abc_52138_new_n4085_), .C(u2__abc_52138_new_n9164_), .Y(u2__abc_52138_new_n9165_));
OAI21X1 OAI21X1_1733 ( .A(u2__abc_52138_new_n9163_), .B(u2__abc_52138_new_n9165_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9166_));
OAI21X1 OAI21X1_1734 ( .A(u2__abc_52138_new_n4076_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9168_));
OAI21X1 OAI21X1_1735 ( .A(u2__abc_52138_new_n9168_), .B(u2__abc_52138_new_n9167_), .C(u2__abc_52138_new_n9169_), .Y(u2__abc_52138_new_n9170_));
OAI21X1 OAI21X1_1736 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_247_), .Y(u2__abc_52138_new_n9172_));
OAI21X1 OAI21X1_1737 ( .A(u2__abc_52138_new_n4081_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9177_));
OAI21X1 OAI21X1_1738 ( .A(u2__abc_52138_new_n9177_), .B(u2__abc_52138_new_n9176_), .C(u2__abc_52138_new_n9178_), .Y(u2__abc_52138_new_n9179_));
OAI21X1 OAI21X1_1739 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_248_), .Y(u2__abc_52138_new_n9181_));
OAI21X1 OAI21X1_174 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1323_), .C(_abc_65734_new_n1324_), .Y(fracta1_62_));
OAI21X1 OAI21X1_1740 ( .A(u2__abc_52138_new_n4091_), .B(u2__abc_52138_new_n4088_), .C(u2__abc_52138_new_n9182_), .Y(u2__abc_52138_new_n9183_));
OAI21X1 OAI21X1_1741 ( .A(u2__abc_52138_new_n4075_), .B(u2__abc_52138_new_n4083_), .C(u2__abc_52138_new_n4080_), .Y(u2__abc_52138_new_n9184_));
OAI21X1 OAI21X1_1742 ( .A(u2__abc_52138_new_n9145_), .B(u2__abc_52138_new_n4983_), .C(u2__abc_52138_new_n9185_), .Y(u2__abc_52138_new_n9186_));
OAI21X1 OAI21X1_1743 ( .A(u2__abc_52138_new_n4005_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9192_));
OAI21X1 OAI21X1_1744 ( .A(u2__abc_52138_new_n9192_), .B(u2__abc_52138_new_n9191_), .C(u2__abc_52138_new_n9193_), .Y(u2__abc_52138_new_n9194_));
OAI21X1 OAI21X1_1745 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_249_), .Y(u2__abc_52138_new_n9196_));
OAI21X1 OAI21X1_1746 ( .A(u2__abc_52138_new_n4007_), .B(u2__abc_52138_new_n9188_), .C(u2__abc_52138_new_n4004_), .Y(u2__abc_52138_new_n9197_));
OAI21X1 OAI21X1_1747 ( .A(u2__abc_52138_new_n4010_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9200_));
OAI21X1 OAI21X1_1748 ( .A(u2__abc_52138_new_n9200_), .B(u2__abc_52138_new_n9199_), .C(u2__abc_52138_new_n9201_), .Y(u2__abc_52138_new_n9202_));
OAI21X1 OAI21X1_1749 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_250_), .Y(u2__abc_52138_new_n9204_));
OAI21X1 OAI21X1_175 ( .A(\a[112] ), .B(_abc_65734_new_n1323_), .C(_abc_65734_new_n1326_), .Y(fracta1_63_));
OAI21X1 OAI21X1_1750 ( .A(u2__abc_52138_new_n4004_), .B(u2__abc_52138_new_n4012_), .C(u2__abc_52138_new_n4009_), .Y(u2__abc_52138_new_n9206_));
OAI21X1 OAI21X1_1751 ( .A(u2__abc_52138_new_n9186_), .B(u2__abc_52138_new_n9187_), .C(u2__abc_52138_new_n4013_), .Y(u2__abc_52138_new_n9208_));
OAI21X1 OAI21X1_1752 ( .A(u2__abc_52138_new_n9205_), .B(u2__abc_52138_new_n9209_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9210_));
OAI21X1 OAI21X1_1753 ( .A(u2__abc_52138_new_n4016_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9212_));
OAI21X1 OAI21X1_1754 ( .A(u2__abc_52138_new_n9212_), .B(u2__abc_52138_new_n9211_), .C(u2__abc_52138_new_n9213_), .Y(u2__abc_52138_new_n9214_));
OAI21X1 OAI21X1_1755 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_251_), .Y(u2__abc_52138_new_n9216_));
OAI21X1 OAI21X1_1756 ( .A(u2_o_248_), .B(u2__abc_52138_new_n4016_), .C(u2__abc_52138_new_n9217_), .Y(u2__abc_52138_new_n9218_));
OAI21X1 OAI21X1_1757 ( .A(u2__abc_52138_new_n4021_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9221_));
OAI21X1 OAI21X1_1758 ( .A(u2__abc_52138_new_n9221_), .B(u2__abc_52138_new_n9220_), .C(u2__abc_52138_new_n9222_), .Y(u2__abc_52138_new_n9223_));
OAI21X1 OAI21X1_1759 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_252_), .Y(u2__abc_52138_new_n9225_));
OAI21X1 OAI21X1_176 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1328_), .C(_abc_65734_new_n1329_), .Y(fracta1_64_));
OAI21X1 OAI21X1_1760 ( .A(u2__abc_52138_new_n4015_), .B(u2__abc_52138_new_n4023_), .C(u2__abc_52138_new_n4020_), .Y(u2__abc_52138_new_n9227_));
OAI21X1 OAI21X1_1761 ( .A(u2__abc_52138_new_n4025_), .B(u2__abc_52138_new_n9188_), .C(u2__abc_52138_new_n9228_), .Y(u2__abc_52138_new_n9229_));
OAI21X1 OAI21X1_1762 ( .A(u2__abc_52138_new_n9226_), .B(u2__abc_52138_new_n9229_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9232_));
OAI21X1 OAI21X1_1763 ( .A(u2__abc_52138_new_n4044_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9234_));
OAI21X1 OAI21X1_1764 ( .A(u2__abc_52138_new_n9234_), .B(u2__abc_52138_new_n9233_), .C(u2__abc_52138_new_n9235_), .Y(u2__abc_52138_new_n9236_));
OAI21X1 OAI21X1_1765 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_253_), .Y(u2__abc_52138_new_n9238_));
OAI21X1 OAI21X1_1766 ( .A(u2_o_250_), .B(u2__abc_52138_new_n4044_), .C(u2__abc_52138_new_n9230_), .Y(u2__abc_52138_new_n9239_));
OAI21X1 OAI21X1_1767 ( .A(u2__abc_52138_new_n4039_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9242_));
OAI21X1 OAI21X1_1768 ( .A(u2__abc_52138_new_n9242_), .B(u2__abc_52138_new_n9241_), .C(u2__abc_52138_new_n9243_), .Y(u2__abc_52138_new_n9244_));
OAI21X1 OAI21X1_1769 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_254_), .Y(u2__abc_52138_new_n9246_));
OAI21X1 OAI21X1_177 ( .A(\a[112] ), .B(_abc_65734_new_n1328_), .C(_abc_65734_new_n1331_), .Y(fracta1_65_));
OAI21X1 OAI21X1_1770 ( .A(u2__abc_52138_new_n4043_), .B(u2__abc_52138_new_n4041_), .C(u2__abc_52138_new_n4038_), .Y(u2__abc_52138_new_n9247_));
OAI21X1 OAI21X1_1771 ( .A(u2__abc_52138_new_n4028_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9250_));
OAI21X1 OAI21X1_1772 ( .A(u2_remHi_254_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6504_), .Y(u2__abc_52138_new_n9252_));
OAI21X1 OAI21X1_1773 ( .A(u2__abc_52138_new_n9252_), .B(u2__abc_52138_new_n9251_), .C(u2__abc_52138_new_n9246_), .Y(u2__abc_52138_new_n9253_));
OAI21X1 OAI21X1_1774 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_255_), .Y(u2__abc_52138_new_n9255_));
OAI21X1 OAI21X1_1775 ( .A(u2__abc_52138_new_n4030_), .B(u2__abc_52138_new_n9248_), .C(u2__abc_52138_new_n4027_), .Y(u2__abc_52138_new_n9256_));
OAI21X1 OAI21X1_1776 ( .A(u2__abc_52138_new_n4031_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9259_));
OAI21X1 OAI21X1_1777 ( .A(u2__abc_52138_new_n9259_), .B(u2__abc_52138_new_n9258_), .C(u2__abc_52138_new_n9260_), .Y(u2__abc_52138_new_n9261_));
OAI21X1 OAI21X1_1778 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_256_), .Y(u2__abc_52138_new_n9263_));
OAI21X1 OAI21X1_1779 ( .A(u2__abc_52138_new_n4027_), .B(u2__abc_52138_new_n4035_), .C(u2__abc_52138_new_n4034_), .Y(u2__abc_52138_new_n9271_));
OAI21X1 OAI21X1_178 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1333_), .C(_abc_65734_new_n1334_), .Y(fracta1_66_));
OAI21X1 OAI21X1_1780 ( .A(u2__abc_52138_new_n9269_), .B(u2__abc_52138_new_n9105_), .C(u2__abc_52138_new_n9273_), .Y(u2__abc_52138_new_n9274_));
OAI21X1 OAI21X1_1781 ( .A(u2__abc_52138_new_n9268_), .B(u2__abc_52138_new_n8602_), .C(u2__abc_52138_new_n9275_), .Y(u2__abc_52138_new_n9276_));
OAI21X1 OAI21X1_1782 ( .A(u2__abc_52138_new_n4753_), .B(u2__abc_52138_new_n7901_), .C(u2__abc_52138_new_n9277_), .Y(u2__abc_52138_new_n9278_));
OAI21X1 OAI21X1_1783 ( .A(u2__abc_52138_new_n9266_), .B(u2__abc_52138_new_n9278_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9279_));
OAI21X1 OAI21X1_1784 ( .A(u2__abc_52138_new_n5691_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9281_));
OAI21X1 OAI21X1_1785 ( .A(u2__abc_52138_new_n9281_), .B(u2__abc_52138_new_n9280_), .C(u2__abc_52138_new_n9282_), .Y(u2__abc_52138_new_n9283_));
OAI21X1 OAI21X1_1786 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_257_), .Y(u2__abc_52138_new_n9285_));
OAI21X1 OAI21X1_1787 ( .A(u2__abc_52138_new_n9264_), .B(u2__abc_52138_new_n9288_), .C(u2__abc_52138_new_n9287_), .Y(u2__abc_52138_new_n9289_));
OAI21X1 OAI21X1_1788 ( .A(u2__abc_52138_new_n9286_), .B(u2__abc_52138_new_n9289_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9290_));
OAI21X1 OAI21X1_1789 ( .A(u2__abc_52138_new_n5688_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9292_));
OAI21X1 OAI21X1_179 ( .A(\a[112] ), .B(_abc_65734_new_n1333_), .C(_abc_65734_new_n1336_), .Y(fracta1_67_));
OAI21X1 OAI21X1_1790 ( .A(u2__abc_52138_new_n9292_), .B(u2__abc_52138_new_n9291_), .C(u2__abc_52138_new_n9293_), .Y(u2__abc_52138_new_n9294_));
OAI21X1 OAI21X1_1791 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_258_), .Y(u2__abc_52138_new_n9296_));
OAI21X1 OAI21X1_1792 ( .A(u2_remHi_255_), .B(u2__abc_52138_new_n5692_), .C(u2__abc_52138_new_n5694_), .Y(u2__abc_52138_new_n9297_));
OAI21X1 OAI21X1_1793 ( .A(u2__abc_52138_new_n5696_), .B(u2__abc_52138_new_n9288_), .C(u2__abc_52138_new_n9297_), .Y(u2__abc_52138_new_n9298_));
OAI21X1 OAI21X1_1794 ( .A(u2__abc_52138_new_n5701_), .B(u2__abc_52138_new_n9298_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9299_));
OAI21X1 OAI21X1_1795 ( .A(u2__abc_52138_new_n5697_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9301_));
OAI21X1 OAI21X1_1796 ( .A(u2__abc_52138_new_n9301_), .B(u2__abc_52138_new_n9300_), .C(u2__abc_52138_new_n9302_), .Y(u2__abc_52138_new_n9303_));
OAI21X1 OAI21X1_1797 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_259_), .Y(u2__abc_52138_new_n9305_));
OAI21X1 OAI21X1_1798 ( .A(u2__abc_52138_new_n5700_), .B(u2__abc_52138_new_n9307_), .C(u2__abc_52138_new_n9306_), .Y(u2__abc_52138_new_n9308_));
OAI21X1 OAI21X1_1799 ( .A(u2__abc_52138_new_n5706_), .B(u2__abc_52138_new_n9308_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9309_));
OAI21X1 OAI21X1_18 ( .A(aNan), .B(_abc_65734_new_n881_), .C(_abc_65734_new_n882_), .Y(\o[129] ));
OAI21X1 OAI21X1_180 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1338_), .C(_abc_65734_new_n1339_), .Y(fracta1_68_));
OAI21X1 OAI21X1_1800 ( .A(u2__abc_52138_new_n5702_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9311_));
OAI21X1 OAI21X1_1801 ( .A(u2__abc_52138_new_n9311_), .B(u2__abc_52138_new_n9310_), .C(u2__abc_52138_new_n9312_), .Y(u2__abc_52138_new_n9313_));
OAI21X1 OAI21X1_1802 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_260_), .Y(u2__abc_52138_new_n9315_));
OAI21X1 OAI21X1_1803 ( .A(u2__abc_52138_new_n5705_), .B(u2__abc_52138_new_n9306_), .C(u2__abc_52138_new_n5738_), .Y(u2__abc_52138_new_n9317_));
OAI21X1 OAI21X1_1804 ( .A(u2__abc_52138_new_n9297_), .B(u2__abc_52138_new_n5707_), .C(u2__abc_52138_new_n9318_), .Y(u2__abc_52138_new_n9319_));
OAI21X1 OAI21X1_1805 ( .A(u2__abc_52138_new_n9316_), .B(u2__abc_52138_new_n9288_), .C(u2__abc_52138_new_n9320_), .Y(u2__abc_52138_new_n9321_));
OAI21X1 OAI21X1_1806 ( .A(u2__abc_52138_new_n5724_), .B(u2__abc_52138_new_n9321_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9324_));
OAI21X1 OAI21X1_1807 ( .A(u2__abc_52138_new_n5720_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9326_));
OAI21X1 OAI21X1_1808 ( .A(u2__abc_52138_new_n9326_), .B(u2__abc_52138_new_n9325_), .C(u2__abc_52138_new_n9327_), .Y(u2__abc_52138_new_n9328_));
OAI21X1 OAI21X1_1809 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_261_), .Y(u2__abc_52138_new_n9330_));
OAI21X1 OAI21X1_181 ( .A(\a[112] ), .B(_abc_65734_new_n1338_), .C(_abc_65734_new_n1341_), .Y(fracta1_69_));
OAI21X1 OAI21X1_1810 ( .A(u2__abc_52138_new_n5720_), .B(u2_o_258_), .C(u2__abc_52138_new_n9322_), .Y(u2__abc_52138_new_n9331_));
OAI21X1 OAI21X1_1811 ( .A(u2__abc_52138_new_n5725_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9334_));
OAI21X1 OAI21X1_1812 ( .A(u2__abc_52138_new_n9334_), .B(u2__abc_52138_new_n9333_), .C(u2__abc_52138_new_n9335_), .Y(u2__abc_52138_new_n9336_));
OAI21X1 OAI21X1_1813 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_262_), .Y(u2__abc_52138_new_n9338_));
OAI21X1 OAI21X1_1814 ( .A(u2__abc_52138_new_n5720_), .B(u2_o_258_), .C(u2__abc_52138_new_n5741_), .Y(u2__abc_52138_new_n9339_));
OAI21X1 OAI21X1_1815 ( .A(u2__abc_52138_new_n9339_), .B(u2__abc_52138_new_n9323_), .C(u2__abc_52138_new_n9340_), .Y(u2__abc_52138_new_n9341_));
OAI21X1 OAI21X1_1816 ( .A(u2__abc_52138_new_n5713_), .B(u2__abc_52138_new_n9342_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9344_));
OAI21X1 OAI21X1_1817 ( .A(u2__abc_52138_new_n5709_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9346_));
OAI21X1 OAI21X1_1818 ( .A(u2__abc_52138_new_n9346_), .B(u2__abc_52138_new_n9345_), .C(u2__abc_52138_new_n9347_), .Y(u2__abc_52138_new_n9348_));
OAI21X1 OAI21X1_1819 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_263_), .Y(u2__abc_52138_new_n9350_));
OAI21X1 OAI21X1_182 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1343_), .C(_abc_65734_new_n1344_), .Y(fracta1_70_));
OAI21X1 OAI21X1_1820 ( .A(u2__abc_52138_new_n5718_), .B(u2__abc_52138_new_n9352_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9353_));
OAI21X1 OAI21X1_1821 ( .A(u2__abc_52138_new_n5714_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9355_));
OAI21X1 OAI21X1_1822 ( .A(u2__abc_52138_new_n9355_), .B(u2__abc_52138_new_n9354_), .C(u2__abc_52138_new_n9356_), .Y(u2__abc_52138_new_n9357_));
OAI21X1 OAI21X1_1823 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_264_), .Y(u2__abc_52138_new_n9359_));
OAI21X1 OAI21X1_1824 ( .A(u2_remHi_259_), .B(u2__abc_52138_new_n5727_), .C(u2__abc_52138_new_n9339_), .Y(u2__abc_52138_new_n9360_));
OAI21X1 OAI21X1_1825 ( .A(u2__abc_52138_new_n5719_), .B(u2__abc_52138_new_n9360_), .C(u2__abc_52138_new_n9361_), .Y(u2__abc_52138_new_n9362_));
OAI21X1 OAI21X1_1826 ( .A(u2__abc_52138_new_n5732_), .B(u2__abc_52138_new_n9288_), .C(u2__abc_52138_new_n9363_), .Y(u2__abc_52138_new_n9364_));
OAI21X1 OAI21X1_1827 ( .A(u2__abc_52138_new_n5678_), .B(u2__abc_52138_new_n9364_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9365_));
OAI21X1 OAI21X1_1828 ( .A(u2__abc_52138_new_n5676_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9367_));
OAI21X1 OAI21X1_1829 ( .A(u2__abc_52138_new_n9367_), .B(u2__abc_52138_new_n9366_), .C(u2__abc_52138_new_n9368_), .Y(u2__abc_52138_new_n9369_));
OAI21X1 OAI21X1_183 ( .A(\a[112] ), .B(_abc_65734_new_n1343_), .C(_abc_65734_new_n1346_), .Y(fracta1_71_));
OAI21X1 OAI21X1_1830 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_265_), .Y(u2__abc_52138_new_n9371_));
OAI21X1 OAI21X1_1831 ( .A(u2__abc_52138_new_n5675_), .B(u2__abc_52138_new_n9373_), .C(u2__abc_52138_new_n9372_), .Y(u2__abc_52138_new_n9374_));
OAI21X1 OAI21X1_1832 ( .A(u2__abc_52138_new_n5683_), .B(u2__abc_52138_new_n9374_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9375_));
OAI21X1 OAI21X1_1833 ( .A(u2__abc_52138_new_n5681_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9377_));
OAI21X1 OAI21X1_1834 ( .A(u2__abc_52138_new_n9377_), .B(u2__abc_52138_new_n9376_), .C(u2__abc_52138_new_n9378_), .Y(u2__abc_52138_new_n9379_));
OAI21X1 OAI21X1_1835 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_266_), .Y(u2__abc_52138_new_n9381_));
OAI21X1 OAI21X1_1836 ( .A(u2__abc_52138_new_n5684_), .B(u2__abc_52138_new_n9373_), .C(u2__abc_52138_new_n9382_), .Y(u2__abc_52138_new_n9383_));
OAI21X1 OAI21X1_1837 ( .A(u2__abc_52138_new_n5667_), .B(u2__abc_52138_new_n9383_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9384_));
OAI21X1 OAI21X1_1838 ( .A(u2__abc_52138_new_n5663_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9386_));
OAI21X1 OAI21X1_1839 ( .A(u2__abc_52138_new_n9386_), .B(u2__abc_52138_new_n9385_), .C(u2__abc_52138_new_n9387_), .Y(u2__abc_52138_new_n9388_));
OAI21X1 OAI21X1_184 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1348_), .C(_abc_65734_new_n1349_), .Y(fracta1_72_));
OAI21X1 OAI21X1_1840 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_267_), .Y(u2__abc_52138_new_n9390_));
OAI21X1 OAI21X1_1841 ( .A(u2__abc_52138_new_n5663_), .B(u2_o_264_), .C(u2__abc_52138_new_n9391_), .Y(u2__abc_52138_new_n9392_));
OAI21X1 OAI21X1_1842 ( .A(u2__abc_52138_new_n5672_), .B(u2__abc_52138_new_n9392_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9393_));
OAI21X1 OAI21X1_1843 ( .A(u2__abc_52138_new_n5668_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9395_));
OAI21X1 OAI21X1_1844 ( .A(u2__abc_52138_new_n9395_), .B(u2__abc_52138_new_n9394_), .C(u2__abc_52138_new_n9396_), .Y(u2__abc_52138_new_n9397_));
OAI21X1 OAI21X1_1845 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_268_), .Y(u2__abc_52138_new_n9399_));
OAI21X1 OAI21X1_1846 ( .A(u2__abc_52138_new_n5655_), .B(u2__abc_52138_new_n9401_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9403_));
OAI21X1 OAI21X1_1847 ( .A(u2__abc_52138_new_n5651_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9405_));
OAI21X1 OAI21X1_1848 ( .A(u2__abc_52138_new_n9405_), .B(u2__abc_52138_new_n9404_), .C(u2__abc_52138_new_n9406_), .Y(u2__abc_52138_new_n9407_));
OAI21X1 OAI21X1_1849 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_269_), .Y(u2__abc_52138_new_n9409_));
OAI21X1 OAI21X1_185 ( .A(\a[112] ), .B(_abc_65734_new_n1348_), .C(_abc_65734_new_n1351_), .Y(fracta1_73_));
OAI21X1 OAI21X1_1850 ( .A(u2__abc_52138_new_n5656_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9413_));
OAI21X1 OAI21X1_1851 ( .A(u2__abc_52138_new_n9413_), .B(u2__abc_52138_new_n9412_), .C(u2__abc_52138_new_n9414_), .Y(u2__abc_52138_new_n9415_));
OAI21X1 OAI21X1_1852 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_270_), .Y(u2__abc_52138_new_n9417_));
OAI21X1 OAI21X1_1853 ( .A(u2__abc_52138_new_n5656_), .B(u2_o_267_), .C(u2__abc_52138_new_n9418_), .Y(u2__abc_52138_new_n9419_));
OAI21X1 OAI21X1_1854 ( .A(u2__abc_52138_new_n9419_), .B(u2__abc_52138_new_n9402_), .C(u2__abc_52138_new_n9420_), .Y(u2__abc_52138_new_n9421_));
OAI21X1 OAI21X1_1855 ( .A(u2__abc_52138_new_n5644_), .B(u2__abc_52138_new_n9422_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9423_));
OAI21X1 OAI21X1_1856 ( .A(u2__abc_52138_new_n5642_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9425_));
OAI21X1 OAI21X1_1857 ( .A(u2__abc_52138_new_n9425_), .B(u2__abc_52138_new_n9424_), .C(u2__abc_52138_new_n9426_), .Y(u2__abc_52138_new_n9427_));
OAI21X1 OAI21X1_1858 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_271_), .Y(u2__abc_52138_new_n9429_));
OAI21X1 OAI21X1_1859 ( .A(u2__abc_52138_new_n5641_), .B(u2__abc_52138_new_n9421_), .C(u2__abc_52138_new_n9430_), .Y(u2__abc_52138_new_n9431_));
OAI21X1 OAI21X1_186 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1353_), .C(_abc_65734_new_n1354_), .Y(fracta1_74_));
OAI21X1 OAI21X1_1860 ( .A(u2__abc_52138_new_n5649_), .B(u2__abc_52138_new_n9431_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9432_));
OAI21X1 OAI21X1_1861 ( .A(u2__abc_52138_new_n5647_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9434_));
OAI21X1 OAI21X1_1862 ( .A(u2__abc_52138_new_n9434_), .B(u2__abc_52138_new_n9433_), .C(u2__abc_52138_new_n9435_), .Y(u2__abc_52138_new_n9436_));
OAI21X1 OAI21X1_1863 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_272_), .Y(u2__abc_52138_new_n9438_));
OAI21X1 OAI21X1_1864 ( .A(u2_remHi_267_), .B(u2__abc_52138_new_n5658_), .C(u2__abc_52138_new_n9419_), .Y(u2__abc_52138_new_n9441_));
OAI21X1 OAI21X1_1865 ( .A(u2__abc_52138_new_n5650_), .B(u2__abc_52138_new_n9441_), .C(u2__abc_52138_new_n9440_), .Y(u2__abc_52138_new_n9442_));
OAI21X1 OAI21X1_1866 ( .A(u2__abc_52138_new_n5686_), .B(u2__abc_52138_new_n9363_), .C(u2__abc_52138_new_n9443_), .Y(u2__abc_52138_new_n9444_));
OAI21X1 OAI21X1_1867 ( .A(u2__abc_52138_new_n9444_), .B(u2__abc_52138_new_n9445_), .C(u2__abc_52138_new_n5610_), .Y(u2__abc_52138_new_n9446_));
OAI21X1 OAI21X1_1868 ( .A(u2__abc_52138_new_n5610_), .B(u2__abc_52138_new_n9449_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9450_));
OAI21X1 OAI21X1_1869 ( .A(u2__abc_52138_new_n5606_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9452_));
OAI21X1 OAI21X1_187 ( .A(\a[112] ), .B(_abc_65734_new_n1353_), .C(_abc_65734_new_n1356_), .Y(fracta1_75_));
OAI21X1 OAI21X1_1870 ( .A(u2__abc_52138_new_n9452_), .B(u2__abc_52138_new_n9451_), .C(u2__abc_52138_new_n9453_), .Y(u2__abc_52138_new_n9454_));
OAI21X1 OAI21X1_1871 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_273_), .Y(u2__abc_52138_new_n9456_));
OAI21X1 OAI21X1_1872 ( .A(u2__abc_52138_new_n5606_), .B(u2_o_270_), .C(u2__abc_52138_new_n9446_), .Y(u2__abc_52138_new_n9457_));
OAI21X1 OAI21X1_1873 ( .A(u2__abc_52138_new_n5611_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9460_));
OAI21X1 OAI21X1_1874 ( .A(u2__abc_52138_new_n9460_), .B(u2__abc_52138_new_n9459_), .C(u2__abc_52138_new_n9461_), .Y(u2__abc_52138_new_n9462_));
OAI21X1 OAI21X1_1875 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_274_), .Y(u2__abc_52138_new_n9464_));
OAI21X1 OAI21X1_1876 ( .A(u2__abc_52138_new_n5606_), .B(u2_o_270_), .C(u2__abc_52138_new_n5756_), .Y(u2__abc_52138_new_n9465_));
OAI21X1 OAI21X1_1877 ( .A(u2__abc_52138_new_n5599_), .B(u2__abc_52138_new_n9467_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9468_));
OAI21X1 OAI21X1_1878 ( .A(u2__abc_52138_new_n5595_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9470_));
OAI21X1 OAI21X1_1879 ( .A(u2__abc_52138_new_n9470_), .B(u2__abc_52138_new_n9469_), .C(u2__abc_52138_new_n9472_), .Y(u2__abc_52138_new_n9473_));
OAI21X1 OAI21X1_188 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1358_), .C(_abc_65734_new_n1359_), .Y(fracta1_76_));
OAI21X1 OAI21X1_1880 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_275_), .Y(u2__abc_52138_new_n9475_));
OAI21X1 OAI21X1_1881 ( .A(u2__abc_52138_new_n5598_), .B(u2__abc_52138_new_n9466_), .C(u2__abc_52138_new_n9476_), .Y(u2__abc_52138_new_n9477_));
OAI21X1 OAI21X1_1882 ( .A(u2__abc_52138_new_n5604_), .B(u2__abc_52138_new_n9477_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9478_));
OAI21X1 OAI21X1_1883 ( .A(u2__abc_52138_new_n5600_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9480_));
OAI21X1 OAI21X1_1884 ( .A(u2__abc_52138_new_n9480_), .B(u2__abc_52138_new_n9479_), .C(u2__abc_52138_new_n9481_), .Y(u2__abc_52138_new_n9482_));
OAI21X1 OAI21X1_1885 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_276_), .Y(u2__abc_52138_new_n9484_));
OAI21X1 OAI21X1_1886 ( .A(u2_remHi_271_), .B(u2__abc_52138_new_n5613_), .C(u2__abc_52138_new_n9465_), .Y(u2__abc_52138_new_n9487_));
OAI21X1 OAI21X1_1887 ( .A(u2__abc_52138_new_n5605_), .B(u2__abc_52138_new_n9487_), .C(u2__abc_52138_new_n9486_), .Y(u2__abc_52138_new_n9488_));
OAI21X1 OAI21X1_1888 ( .A(u2__abc_52138_new_n9485_), .B(u2__abc_52138_new_n9448_), .C(u2__abc_52138_new_n9489_), .Y(u2__abc_52138_new_n9490_));
OAI21X1 OAI21X1_1889 ( .A(u2__abc_52138_new_n5629_), .B(u2__abc_52138_new_n9490_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9493_));
OAI21X1 OAI21X1_189 ( .A(\a[112] ), .B(_abc_65734_new_n1358_), .C(_abc_65734_new_n1361_), .Y(fracta1_77_));
OAI21X1 OAI21X1_1890 ( .A(u2__abc_52138_new_n9471_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9495_));
OAI21X1 OAI21X1_1891 ( .A(u2__abc_52138_new_n9495_), .B(u2__abc_52138_new_n9494_), .C(u2__abc_52138_new_n9496_), .Y(u2__abc_52138_new_n9497_));
OAI21X1 OAI21X1_1892 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_277_), .Y(u2__abc_52138_new_n9499_));
OAI21X1 OAI21X1_1893 ( .A(u2__abc_52138_new_n9471_), .B(u2_o_274_), .C(u2__abc_52138_new_n9491_), .Y(u2__abc_52138_new_n9500_));
OAI21X1 OAI21X1_1894 ( .A(u2__abc_52138_new_n5630_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9503_));
OAI21X1 OAI21X1_1895 ( .A(u2__abc_52138_new_n9503_), .B(u2__abc_52138_new_n9502_), .C(u2__abc_52138_new_n9504_), .Y(u2__abc_52138_new_n9505_));
OAI21X1 OAI21X1_1896 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_278_), .Y(u2__abc_52138_new_n9507_));
OAI21X1 OAI21X1_1897 ( .A(u2__abc_52138_new_n9471_), .B(u2_o_274_), .C(u2__abc_52138_new_n9508_), .Y(u2__abc_52138_new_n9509_));
OAI21X1 OAI21X1_1898 ( .A(u2__abc_52138_new_n9509_), .B(u2__abc_52138_new_n9492_), .C(u2__abc_52138_new_n5762_), .Y(u2__abc_52138_new_n9510_));
OAI21X1 OAI21X1_1899 ( .A(u2__abc_52138_new_n5622_), .B(u2__abc_52138_new_n9511_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9512_));
OAI21X1 OAI21X1_19 ( .A(aNan), .B(_abc_65734_new_n884_), .C(_abc_65734_new_n885_), .Y(\o[130] ));
OAI21X1 OAI21X1_190 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1363_), .C(_abc_65734_new_n1364_), .Y(fracta1_78_));
OAI21X1 OAI21X1_1900 ( .A(u2__abc_52138_new_n5618_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9514_));
OAI21X1 OAI21X1_1901 ( .A(u2__abc_52138_new_n9514_), .B(u2__abc_52138_new_n9513_), .C(u2__abc_52138_new_n9515_), .Y(u2__abc_52138_new_n9516_));
OAI21X1 OAI21X1_1902 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_279_), .Y(u2__abc_52138_new_n9518_));
OAI21X1 OAI21X1_1903 ( .A(u2__abc_52138_new_n5621_), .B(u2__abc_52138_new_n9510_), .C(u2__abc_52138_new_n9519_), .Y(u2__abc_52138_new_n9520_));
OAI21X1 OAI21X1_1904 ( .A(u2__abc_52138_new_n5627_), .B(u2__abc_52138_new_n9520_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9521_));
OAI21X1 OAI21X1_1905 ( .A(u2__abc_52138_new_n5623_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9523_));
OAI21X1 OAI21X1_1906 ( .A(u2__abc_52138_new_n9523_), .B(u2__abc_52138_new_n9522_), .C(u2__abc_52138_new_n9524_), .Y(u2__abc_52138_new_n9525_));
OAI21X1 OAI21X1_1907 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_280_), .Y(u2__abc_52138_new_n9527_));
OAI21X1 OAI21X1_1908 ( .A(u2_remHi_275_), .B(u2__abc_52138_new_n5632_), .C(u2__abc_52138_new_n9509_), .Y(u2__abc_52138_new_n9528_));
OAI21X1 OAI21X1_1909 ( .A(u2__abc_52138_new_n5628_), .B(u2__abc_52138_new_n9528_), .C(u2__abc_52138_new_n9529_), .Y(u2__abc_52138_new_n9530_));
OAI21X1 OAI21X1_191 ( .A(\a[112] ), .B(_abc_65734_new_n1363_), .C(_abc_65734_new_n1366_), .Y(fracta1_79_));
OAI21X1 OAI21X1_1910 ( .A(u2__abc_52138_new_n5637_), .B(u2__abc_52138_new_n9448_), .C(u2__abc_52138_new_n9531_), .Y(u2__abc_52138_new_n9532_));
OAI21X1 OAI21X1_1911 ( .A(u2__abc_52138_new_n5563_), .B(u2__abc_52138_new_n9532_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9535_));
OAI21X1 OAI21X1_1912 ( .A(u2__abc_52138_new_n5559_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9537_));
OAI21X1 OAI21X1_1913 ( .A(u2__abc_52138_new_n9537_), .B(u2__abc_52138_new_n9536_), .C(u2__abc_52138_new_n9538_), .Y(u2__abc_52138_new_n9539_));
OAI21X1 OAI21X1_1914 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_281_), .Y(u2__abc_52138_new_n9541_));
OAI21X1 OAI21X1_1915 ( .A(u2__abc_52138_new_n5559_), .B(u2_o_278_), .C(u2__abc_52138_new_n9533_), .Y(u2__abc_52138_new_n9542_));
OAI21X1 OAI21X1_1916 ( .A(u2__abc_52138_new_n5564_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9545_));
OAI21X1 OAI21X1_1917 ( .A(u2__abc_52138_new_n9545_), .B(u2__abc_52138_new_n9544_), .C(u2__abc_52138_new_n9546_), .Y(u2__abc_52138_new_n9547_));
OAI21X1 OAI21X1_1918 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_282_), .Y(u2__abc_52138_new_n9549_));
OAI21X1 OAI21X1_1919 ( .A(u2__abc_52138_new_n5559_), .B(u2_o_278_), .C(u2__abc_52138_new_n5768_), .Y(u2__abc_52138_new_n9550_));
OAI21X1 OAI21X1_192 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1368_), .C(_abc_65734_new_n1369_), .Y(fracta1_80_));
OAI21X1 OAI21X1_1920 ( .A(u2__abc_52138_new_n5552_), .B(u2__abc_52138_new_n9552_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9553_));
OAI21X1 OAI21X1_1921 ( .A(u2__abc_52138_new_n5548_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9555_));
OAI21X1 OAI21X1_1922 ( .A(u2__abc_52138_new_n9555_), .B(u2__abc_52138_new_n9554_), .C(u2__abc_52138_new_n9556_), .Y(u2__abc_52138_new_n9557_));
OAI21X1 OAI21X1_1923 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_283_), .Y(u2__abc_52138_new_n9559_));
OAI21X1 OAI21X1_1924 ( .A(u2__abc_52138_new_n5551_), .B(u2__abc_52138_new_n9551_), .C(u2__abc_52138_new_n9560_), .Y(u2__abc_52138_new_n9561_));
OAI21X1 OAI21X1_1925 ( .A(u2__abc_52138_new_n5557_), .B(u2__abc_52138_new_n9561_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9562_));
OAI21X1 OAI21X1_1926 ( .A(u2__abc_52138_new_n5553_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9564_));
OAI21X1 OAI21X1_1927 ( .A(u2__abc_52138_new_n9564_), .B(u2__abc_52138_new_n9563_), .C(u2__abc_52138_new_n9565_), .Y(u2__abc_52138_new_n9566_));
OAI21X1 OAI21X1_1928 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_284_), .Y(u2__abc_52138_new_n9568_));
OAI21X1 OAI21X1_1929 ( .A(u2_remHi_279_), .B(u2__abc_52138_new_n5566_), .C(u2__abc_52138_new_n9550_), .Y(u2__abc_52138_new_n9569_));
OAI21X1 OAI21X1_193 ( .A(\a[112] ), .B(_abc_65734_new_n1368_), .C(_abc_65734_new_n1371_), .Y(fracta1_81_));
OAI21X1 OAI21X1_1930 ( .A(u2__abc_52138_new_n5556_), .B(u2__abc_52138_new_n9560_), .C(u2__abc_52138_new_n5770_), .Y(u2__abc_52138_new_n9570_));
OAI21X1 OAI21X1_1931 ( .A(u2__abc_52138_new_n5558_), .B(u2__abc_52138_new_n9569_), .C(u2__abc_52138_new_n9571_), .Y(u2__abc_52138_new_n9572_));
OAI21X1 OAI21X1_1932 ( .A(u2__abc_52138_new_n5586_), .B(u2__abc_52138_new_n9574_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9577_));
OAI21X1 OAI21X1_1933 ( .A(u2__abc_52138_new_n5582_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9579_));
OAI21X1 OAI21X1_1934 ( .A(u2__abc_52138_new_n9579_), .B(u2__abc_52138_new_n9578_), .C(u2__abc_52138_new_n9580_), .Y(u2__abc_52138_new_n9581_));
OAI21X1 OAI21X1_1935 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_285_), .Y(u2__abc_52138_new_n9583_));
OAI21X1 OAI21X1_1936 ( .A(u2__abc_52138_new_n5585_), .B(u2__abc_52138_new_n9573_), .C(u2__abc_52138_new_n9584_), .Y(u2__abc_52138_new_n9585_));
OAI21X1 OAI21X1_1937 ( .A(u2__abc_52138_new_n5587_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9588_));
OAI21X1 OAI21X1_1938 ( .A(u2__abc_52138_new_n9588_), .B(u2__abc_52138_new_n9587_), .C(u2__abc_52138_new_n9589_), .Y(u2__abc_52138_new_n9590_));
OAI21X1 OAI21X1_1939 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_286_), .Y(u2__abc_52138_new_n9592_));
OAI21X1 OAI21X1_194 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1373_), .C(_abc_65734_new_n1374_), .Y(fracta1_82_));
OAI21X1 OAI21X1_1940 ( .A(u2__abc_52138_new_n5587_), .B(u2_o_283_), .C(u2__abc_52138_new_n9584_), .Y(u2__abc_52138_new_n9593_));
OAI21X1 OAI21X1_1941 ( .A(u2__abc_52138_new_n9593_), .B(u2__abc_52138_new_n9576_), .C(u2__abc_52138_new_n9594_), .Y(u2__abc_52138_new_n9595_));
OAI21X1 OAI21X1_1942 ( .A(u2__abc_52138_new_n5575_), .B(u2__abc_52138_new_n9596_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9597_));
OAI21X1 OAI21X1_1943 ( .A(u2__abc_52138_new_n5571_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9599_));
OAI21X1 OAI21X1_1944 ( .A(u2__abc_52138_new_n9599_), .B(u2__abc_52138_new_n9598_), .C(u2__abc_52138_new_n9600_), .Y(u2__abc_52138_new_n9601_));
OAI21X1 OAI21X1_1945 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_287_), .Y(u2__abc_52138_new_n9603_));
OAI21X1 OAI21X1_1946 ( .A(u2__abc_52138_new_n5574_), .B(u2__abc_52138_new_n9595_), .C(u2__abc_52138_new_n9604_), .Y(u2__abc_52138_new_n9605_));
OAI21X1 OAI21X1_1947 ( .A(u2__abc_52138_new_n5580_), .B(u2__abc_52138_new_n9605_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9606_));
OAI21X1 OAI21X1_1948 ( .A(u2__abc_52138_new_n5576_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9608_));
OAI21X1 OAI21X1_1949 ( .A(u2__abc_52138_new_n9608_), .B(u2__abc_52138_new_n9607_), .C(u2__abc_52138_new_n9609_), .Y(u2__abc_52138_new_n9610_));
OAI21X1 OAI21X1_195 ( .A(\a[112] ), .B(_abc_65734_new_n1373_), .C(_abc_65734_new_n1376_), .Y(fracta1_83_));
OAI21X1 OAI21X1_1950 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_288_), .Y(u2__abc_52138_new_n9612_));
OAI21X1 OAI21X1_1951 ( .A(u2__abc_52138_new_n9604_), .B(u2__abc_52138_new_n5579_), .C(u2__abc_52138_new_n9614_), .Y(u2__abc_52138_new_n9615_));
OAI21X1 OAI21X1_1952 ( .A(u2__abc_52138_new_n5594_), .B(u2__abc_52138_new_n9531_), .C(u2__abc_52138_new_n9617_), .Y(u2__abc_52138_new_n9618_));
OAI21X1 OAI21X1_1953 ( .A(u2__abc_52138_new_n9619_), .B(u2__abc_52138_new_n9620_), .C(u2__abc_52138_new_n5517_), .Y(u2__abc_52138_new_n9621_));
OAI21X1 OAI21X1_1954 ( .A(u2__abc_52138_new_n5517_), .B(u2__abc_52138_new_n9624_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9625_));
OAI21X1 OAI21X1_1955 ( .A(u2__abc_52138_new_n5513_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9627_));
OAI21X1 OAI21X1_1956 ( .A(u2__abc_52138_new_n9627_), .B(u2__abc_52138_new_n9626_), .C(u2__abc_52138_new_n9628_), .Y(u2__abc_52138_new_n9629_));
OAI21X1 OAI21X1_1957 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_289_), .Y(u2__abc_52138_new_n9631_));
OAI21X1 OAI21X1_1958 ( .A(u2__abc_52138_new_n5513_), .B(u2_o_286_), .C(u2__abc_52138_new_n9621_), .Y(u2__abc_52138_new_n9632_));
OAI21X1 OAI21X1_1959 ( .A(u2__abc_52138_new_n5518_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9635_));
OAI21X1 OAI21X1_196 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1378_), .C(_abc_65734_new_n1379_), .Y(fracta1_84_));
OAI21X1 OAI21X1_1960 ( .A(u2__abc_52138_new_n9635_), .B(u2__abc_52138_new_n9634_), .C(u2__abc_52138_new_n9636_), .Y(u2__abc_52138_new_n9637_));
OAI21X1 OAI21X1_1961 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_290_), .Y(u2__abc_52138_new_n9639_));
OAI21X1 OAI21X1_1962 ( .A(u2__abc_52138_new_n5513_), .B(u2_o_286_), .C(u2__abc_52138_new_n5784_), .Y(u2__abc_52138_new_n9640_));
OAI21X1 OAI21X1_1963 ( .A(u2__abc_52138_new_n5506_), .B(u2__abc_52138_new_n9642_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9643_));
OAI21X1 OAI21X1_1964 ( .A(u2__abc_52138_new_n5502_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9645_));
OAI21X1 OAI21X1_1965 ( .A(u2__abc_52138_new_n9645_), .B(u2__abc_52138_new_n9644_), .C(u2__abc_52138_new_n9647_), .Y(u2__abc_52138_new_n9648_));
OAI21X1 OAI21X1_1966 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_291_), .Y(u2__abc_52138_new_n9650_));
OAI21X1 OAI21X1_1967 ( .A(u2__abc_52138_new_n5505_), .B(u2__abc_52138_new_n9641_), .C(u2__abc_52138_new_n9651_), .Y(u2__abc_52138_new_n9652_));
OAI21X1 OAI21X1_1968 ( .A(u2__abc_52138_new_n5511_), .B(u2__abc_52138_new_n9652_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9653_));
OAI21X1 OAI21X1_1969 ( .A(u2__abc_52138_new_n5507_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9655_));
OAI21X1 OAI21X1_197 ( .A(\a[112] ), .B(_abc_65734_new_n1378_), .C(_abc_65734_new_n1381_), .Y(fracta1_85_));
OAI21X1 OAI21X1_1970 ( .A(u2__abc_52138_new_n9655_), .B(u2__abc_52138_new_n9654_), .C(u2__abc_52138_new_n9656_), .Y(u2__abc_52138_new_n9657_));
OAI21X1 OAI21X1_1971 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_292_), .Y(u2__abc_52138_new_n9659_));
OAI21X1 OAI21X1_1972 ( .A(u2_remHi_287_), .B(u2__abc_52138_new_n5520_), .C(u2__abc_52138_new_n9640_), .Y(u2__abc_52138_new_n9661_));
OAI21X1 OAI21X1_1973 ( .A(u2__abc_52138_new_n5510_), .B(u2__abc_52138_new_n9651_), .C(u2__abc_52138_new_n5782_), .Y(u2__abc_52138_new_n9662_));
OAI21X1 OAI21X1_1974 ( .A(u2__abc_52138_new_n5512_), .B(u2__abc_52138_new_n9661_), .C(u2__abc_52138_new_n9663_), .Y(u2__abc_52138_new_n9664_));
OAI21X1 OAI21X1_1975 ( .A(u2__abc_52138_new_n9660_), .B(u2__abc_52138_new_n9623_), .C(u2__abc_52138_new_n9665_), .Y(u2__abc_52138_new_n9666_));
OAI21X1 OAI21X1_1976 ( .A(u2__abc_52138_new_n5536_), .B(u2__abc_52138_new_n9666_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9669_));
OAI21X1 OAI21X1_1977 ( .A(u2__abc_52138_new_n9646_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9671_));
OAI21X1 OAI21X1_1978 ( .A(u2__abc_52138_new_n9671_), .B(u2__abc_52138_new_n9670_), .C(u2__abc_52138_new_n9672_), .Y(u2__abc_52138_new_n9673_));
OAI21X1 OAI21X1_1979 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_293_), .Y(u2__abc_52138_new_n9675_));
OAI21X1 OAI21X1_198 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1383_), .C(_abc_65734_new_n1384_), .Y(fracta1_86_));
OAI21X1 OAI21X1_1980 ( .A(u2__abc_52138_new_n9646_), .B(u2_o_290_), .C(u2__abc_52138_new_n9667_), .Y(u2__abc_52138_new_n9676_));
OAI21X1 OAI21X1_1981 ( .A(u2__abc_52138_new_n5537_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9679_));
OAI21X1 OAI21X1_1982 ( .A(u2__abc_52138_new_n9679_), .B(u2__abc_52138_new_n9678_), .C(u2__abc_52138_new_n9680_), .Y(u2__abc_52138_new_n9681_));
OAI21X1 OAI21X1_1983 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_294_), .Y(u2__abc_52138_new_n9683_));
OAI21X1 OAI21X1_1984 ( .A(u2__abc_52138_new_n9646_), .B(u2_o_290_), .C(u2__abc_52138_new_n9684_), .Y(u2__abc_52138_new_n9685_));
OAI21X1 OAI21X1_1985 ( .A(u2__abc_52138_new_n9685_), .B(u2__abc_52138_new_n9668_), .C(u2__abc_52138_new_n5788_), .Y(u2__abc_52138_new_n9686_));
OAI21X1 OAI21X1_1986 ( .A(u2__abc_52138_new_n5529_), .B(u2__abc_52138_new_n9687_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9688_));
OAI21X1 OAI21X1_1987 ( .A(u2__abc_52138_new_n5525_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9690_));
OAI21X1 OAI21X1_1988 ( .A(u2__abc_52138_new_n9690_), .B(u2__abc_52138_new_n9689_), .C(u2__abc_52138_new_n9691_), .Y(u2__abc_52138_new_n9692_));
OAI21X1 OAI21X1_1989 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_295_), .Y(u2__abc_52138_new_n9694_));
OAI21X1 OAI21X1_199 ( .A(\a[112] ), .B(_abc_65734_new_n1383_), .C(_abc_65734_new_n1386_), .Y(fracta1_87_));
OAI21X1 OAI21X1_1990 ( .A(u2__abc_52138_new_n5528_), .B(u2__abc_52138_new_n9686_), .C(u2__abc_52138_new_n9695_), .Y(u2__abc_52138_new_n9696_));
OAI21X1 OAI21X1_1991 ( .A(u2__abc_52138_new_n5534_), .B(u2__abc_52138_new_n9696_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9697_));
OAI21X1 OAI21X1_1992 ( .A(u2__abc_52138_new_n5530_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9699_));
OAI21X1 OAI21X1_1993 ( .A(u2__abc_52138_new_n9699_), .B(u2__abc_52138_new_n9698_), .C(u2__abc_52138_new_n9700_), .Y(u2__abc_52138_new_n9701_));
OAI21X1 OAI21X1_1994 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_296_), .Y(u2__abc_52138_new_n9703_));
OAI21X1 OAI21X1_1995 ( .A(u2_remHi_291_), .B(u2__abc_52138_new_n5539_), .C(u2__abc_52138_new_n9685_), .Y(u2__abc_52138_new_n9704_));
OAI21X1 OAI21X1_1996 ( .A(u2__abc_52138_new_n5535_), .B(u2__abc_52138_new_n9704_), .C(u2__abc_52138_new_n9705_), .Y(u2__abc_52138_new_n9706_));
OAI21X1 OAI21X1_1997 ( .A(u2__abc_52138_new_n5544_), .B(u2__abc_52138_new_n9623_), .C(u2__abc_52138_new_n9707_), .Y(u2__abc_52138_new_n9708_));
OAI21X1 OAI21X1_1998 ( .A(u2__abc_52138_new_n5459_), .B(u2__abc_52138_new_n9708_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9709_));
OAI21X1 OAI21X1_1999 ( .A(u2__abc_52138_new_n5457_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9711_));
OAI21X1 OAI21X1_2 ( .A(aNan), .B(_abc_65734_new_n833_), .C(_abc_65734_new_n834_), .Y(\o[113] ));
OAI21X1 OAI21X1_20 ( .A(aNan), .B(_abc_65734_new_n887_), .C(_abc_65734_new_n888_), .Y(\o[131] ));
OAI21X1 OAI21X1_200 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1388_), .C(_abc_65734_new_n1389_), .Y(fracta1_88_));
OAI21X1 OAI21X1_2000 ( .A(u2__abc_52138_new_n9711_), .B(u2__abc_52138_new_n9710_), .C(u2__abc_52138_new_n9712_), .Y(u2__abc_52138_new_n9713_));
OAI21X1 OAI21X1_2001 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_297_), .Y(u2__abc_52138_new_n9715_));
OAI21X1 OAI21X1_2002 ( .A(u2__abc_52138_new_n5456_), .B(u2__abc_52138_new_n9717_), .C(u2__abc_52138_new_n9716_), .Y(u2__abc_52138_new_n9718_));
OAI21X1 OAI21X1_2003 ( .A(u2__abc_52138_new_n5464_), .B(u2__abc_52138_new_n9718_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9719_));
OAI21X1 OAI21X1_2004 ( .A(u2__abc_52138_new_n5460_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9721_));
OAI21X1 OAI21X1_2005 ( .A(u2__abc_52138_new_n9721_), .B(u2__abc_52138_new_n9720_), .C(u2__abc_52138_new_n9722_), .Y(u2__abc_52138_new_n9723_));
OAI21X1 OAI21X1_2006 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_298_), .Y(u2__abc_52138_new_n9725_));
OAI21X1 OAI21X1_2007 ( .A(u2__abc_52138_new_n5457_), .B(u2_o_294_), .C(u2__abc_52138_new_n5463_), .Y(u2__abc_52138_new_n9726_));
OAI21X1 OAI21X1_2008 ( .A(u2_remHi_295_), .B(u2__abc_52138_new_n5462_), .C(u2__abc_52138_new_n9726_), .Y(u2__abc_52138_new_n9727_));
OAI21X1 OAI21X1_2009 ( .A(u2__abc_52138_new_n5465_), .B(u2__abc_52138_new_n9717_), .C(u2__abc_52138_new_n9727_), .Y(u2__abc_52138_new_n9728_));
OAI21X1 OAI21X1_201 ( .A(\a[112] ), .B(_abc_65734_new_n1388_), .C(_abc_65734_new_n1391_), .Y(fracta1_89_));
OAI21X1 OAI21X1_2010 ( .A(u2__abc_52138_new_n5470_), .B(u2__abc_52138_new_n9728_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9729_));
OAI21X1 OAI21X1_2011 ( .A(u2__abc_52138_new_n5466_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9731_));
OAI21X1 OAI21X1_2012 ( .A(u2__abc_52138_new_n9731_), .B(u2__abc_52138_new_n9730_), .C(u2__abc_52138_new_n9732_), .Y(u2__abc_52138_new_n9733_));
OAI21X1 OAI21X1_2013 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_299_), .Y(u2__abc_52138_new_n9735_));
OAI21X1 OAI21X1_2014 ( .A(u2__abc_52138_new_n5466_), .B(u2_o_296_), .C(u2__abc_52138_new_n9736_), .Y(u2__abc_52138_new_n9737_));
OAI21X1 OAI21X1_2015 ( .A(u2__abc_52138_new_n5475_), .B(u2__abc_52138_new_n9737_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9738_));
OAI21X1 OAI21X1_2016 ( .A(u2__abc_52138_new_n5471_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9740_));
OAI21X1 OAI21X1_2017 ( .A(u2__abc_52138_new_n9740_), .B(u2__abc_52138_new_n9739_), .C(u2__abc_52138_new_n9741_), .Y(u2__abc_52138_new_n9742_));
OAI21X1 OAI21X1_2018 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_300_), .Y(u2__abc_52138_new_n9744_));
OAI21X1 OAI21X1_2019 ( .A(u2__abc_52138_new_n9727_), .B(u2__abc_52138_new_n5476_), .C(u2__abc_52138_new_n9745_), .Y(u2__abc_52138_new_n9746_));
OAI21X1 OAI21X1_202 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1393_), .C(_abc_65734_new_n1394_), .Y(fracta1_90_));
OAI21X1 OAI21X1_2020 ( .A(u2__abc_52138_new_n5493_), .B(u2__abc_52138_new_n9748_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9751_));
OAI21X1 OAI21X1_2021 ( .A(u2__abc_52138_new_n5489_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9753_));
OAI21X1 OAI21X1_2022 ( .A(u2__abc_52138_new_n9753_), .B(u2__abc_52138_new_n9752_), .C(u2__abc_52138_new_n9754_), .Y(u2__abc_52138_new_n9755_));
OAI21X1 OAI21X1_2023 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_301_), .Y(u2__abc_52138_new_n9757_));
OAI21X1 OAI21X1_2024 ( .A(u2__abc_52138_new_n5489_), .B(u2_o_298_), .C(u2__abc_52138_new_n9749_), .Y(u2__abc_52138_new_n9758_));
OAI21X1 OAI21X1_2025 ( .A(u2__abc_52138_new_n5494_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9761_));
OAI21X1 OAI21X1_2026 ( .A(u2__abc_52138_new_n9761_), .B(u2__abc_52138_new_n9760_), .C(u2__abc_52138_new_n9762_), .Y(u2__abc_52138_new_n9763_));
OAI21X1 OAI21X1_2027 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_302_), .Y(u2__abc_52138_new_n9765_));
OAI21X1 OAI21X1_2028 ( .A(u2__abc_52138_new_n5489_), .B(u2_o_298_), .C(u2__abc_52138_new_n9766_), .Y(u2__abc_52138_new_n9767_));
OAI21X1 OAI21X1_2029 ( .A(u2__abc_52138_new_n9767_), .B(u2__abc_52138_new_n9750_), .C(u2__abc_52138_new_n9768_), .Y(u2__abc_52138_new_n9769_));
OAI21X1 OAI21X1_203 ( .A(\a[112] ), .B(_abc_65734_new_n1393_), .C(_abc_65734_new_n1396_), .Y(fracta1_91_));
OAI21X1 OAI21X1_2030 ( .A(u2__abc_52138_new_n5482_), .B(u2__abc_52138_new_n9770_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9771_));
OAI21X1 OAI21X1_2031 ( .A(u2__abc_52138_new_n5478_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9773_));
OAI21X1 OAI21X1_2032 ( .A(u2__abc_52138_new_n9773_), .B(u2__abc_52138_new_n9772_), .C(u2__abc_52138_new_n9774_), .Y(u2__abc_52138_new_n9775_));
OAI21X1 OAI21X1_2033 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_303_), .Y(u2__abc_52138_new_n9777_));
OAI21X1 OAI21X1_2034 ( .A(u2__abc_52138_new_n5481_), .B(u2__abc_52138_new_n9769_), .C(u2__abc_52138_new_n9778_), .Y(u2__abc_52138_new_n9779_));
OAI21X1 OAI21X1_2035 ( .A(u2__abc_52138_new_n5487_), .B(u2__abc_52138_new_n9779_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9780_));
OAI21X1 OAI21X1_2036 ( .A(u2__abc_52138_new_n5483_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9782_));
OAI21X1 OAI21X1_2037 ( .A(u2__abc_52138_new_n9782_), .B(u2__abc_52138_new_n9781_), .C(u2__abc_52138_new_n9783_), .Y(u2__abc_52138_new_n9784_));
OAI21X1 OAI21X1_2038 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_304_), .Y(u2__abc_52138_new_n9786_));
OAI21X1 OAI21X1_2039 ( .A(u2__abc_52138_new_n9619_), .B(u2__abc_52138_new_n9620_), .C(u2__abc_52138_new_n5545_), .Y(u2__abc_52138_new_n9793_));
OAI21X1 OAI21X1_204 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1398_), .C(_abc_65734_new_n1399_), .Y(fracta1_92_));
OAI21X1 OAI21X1_2040 ( .A(u2__abc_52138_new_n5411_), .B(u2__abc_52138_new_n9794_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9795_));
OAI21X1 OAI21X1_2041 ( .A(u2__abc_52138_new_n5409_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9797_));
OAI21X1 OAI21X1_2042 ( .A(u2__abc_52138_new_n9797_), .B(u2__abc_52138_new_n9796_), .C(u2__abc_52138_new_n9798_), .Y(u2__abc_52138_new_n9799_));
OAI21X1 OAI21X1_2043 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_305_), .Y(u2__abc_52138_new_n9801_));
OAI21X1 OAI21X1_2044 ( .A(u2__abc_52138_new_n5408_), .B(u2__abc_52138_new_n9803_), .C(u2__abc_52138_new_n9802_), .Y(u2__abc_52138_new_n9804_));
OAI21X1 OAI21X1_2045 ( .A(u2__abc_52138_new_n5416_), .B(u2__abc_52138_new_n9804_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9805_));
OAI21X1 OAI21X1_2046 ( .A(u2__abc_52138_new_n5414_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9807_));
OAI21X1 OAI21X1_2047 ( .A(u2__abc_52138_new_n9807_), .B(u2__abc_52138_new_n9806_), .C(u2__abc_52138_new_n9808_), .Y(u2__abc_52138_new_n9809_));
OAI21X1 OAI21X1_2048 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_306_), .Y(u2__abc_52138_new_n9811_));
OAI21X1 OAI21X1_2049 ( .A(u2__abc_52138_new_n5417_), .B(u2__abc_52138_new_n9803_), .C(u2__abc_52138_new_n9812_), .Y(u2__abc_52138_new_n9813_));
OAI21X1 OAI21X1_205 ( .A(\a[112] ), .B(_abc_65734_new_n1398_), .C(_abc_65734_new_n1401_), .Y(fracta1_93_));
OAI21X1 OAI21X1_2050 ( .A(u2__abc_52138_new_n5422_), .B(u2__abc_52138_new_n9813_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9814_));
OAI21X1 OAI21X1_2051 ( .A(u2__abc_52138_new_n5418_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9816_));
OAI21X1 OAI21X1_2052 ( .A(u2__abc_52138_new_n9816_), .B(u2__abc_52138_new_n9815_), .C(u2__abc_52138_new_n9817_), .Y(u2__abc_52138_new_n9818_));
OAI21X1 OAI21X1_2053 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_307_), .Y(u2__abc_52138_new_n9820_));
OAI21X1 OAI21X1_2054 ( .A(u2__abc_52138_new_n5418_), .B(u2_o_304_), .C(u2__abc_52138_new_n9821_), .Y(u2__abc_52138_new_n9822_));
OAI21X1 OAI21X1_2055 ( .A(u2__abc_52138_new_n5427_), .B(u2__abc_52138_new_n9822_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9823_));
OAI21X1 OAI21X1_2056 ( .A(u2__abc_52138_new_n5423_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9825_));
OAI21X1 OAI21X1_2057 ( .A(u2__abc_52138_new_n9825_), .B(u2__abc_52138_new_n9824_), .C(u2__abc_52138_new_n9826_), .Y(u2__abc_52138_new_n9827_));
OAI21X1 OAI21X1_2058 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_308_), .Y(u2__abc_52138_new_n9829_));
OAI21X1 OAI21X1_2059 ( .A(u2__abc_52138_new_n5428_), .B(u2__abc_52138_new_n9812_), .C(u2__abc_52138_new_n9831_), .Y(u2__abc_52138_new_n9832_));
OAI21X1 OAI21X1_206 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1403_), .C(_abc_65734_new_n1404_), .Y(fracta1_94_));
OAI21X1 OAI21X1_2060 ( .A(u2__abc_52138_new_n9830_), .B(u2__abc_52138_new_n9803_), .C(u2__abc_52138_new_n9833_), .Y(u2__abc_52138_new_n9834_));
OAI21X1 OAI21X1_2061 ( .A(u2__abc_52138_new_n5450_), .B(u2__abc_52138_new_n9834_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9837_));
OAI21X1 OAI21X1_2062 ( .A(u2__abc_52138_new_n5446_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9839_));
OAI21X1 OAI21X1_2063 ( .A(u2__abc_52138_new_n9839_), .B(u2__abc_52138_new_n9838_), .C(u2__abc_52138_new_n9840_), .Y(u2__abc_52138_new_n9841_));
OAI21X1 OAI21X1_2064 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_309_), .Y(u2__abc_52138_new_n9843_));
OAI21X1 OAI21X1_2065 ( .A(u2__abc_52138_new_n5447_), .B(u2__abc_52138_new_n9836_), .C(u2__abc_52138_new_n5445_), .Y(u2__abc_52138_new_n9844_));
OAI21X1 OAI21X1_2066 ( .A(u2__abc_52138_new_n5446_), .B(u2_o_306_), .C(u2__abc_52138_new_n9835_), .Y(u2__abc_52138_new_n9846_));
OAI21X1 OAI21X1_2067 ( .A(u2__abc_52138_new_n5445_), .B(u2__abc_52138_new_n9846_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9847_));
OAI21X1 OAI21X1_2068 ( .A(u2__abc_52138_new_n5441_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9849_));
OAI21X1 OAI21X1_2069 ( .A(u2__abc_52138_new_n9849_), .B(u2__abc_52138_new_n9848_), .C(u2__abc_52138_new_n9850_), .Y(u2__abc_52138_new_n9851_));
OAI21X1 OAI21X1_207 ( .A(\a[112] ), .B(_abc_65734_new_n1403_), .C(_abc_65734_new_n1406_), .Y(fracta1_95_));
OAI21X1 OAI21X1_2070 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_310_), .Y(u2__abc_52138_new_n9853_));
OAI21X1 OAI21X1_2071 ( .A(u2__abc_52138_new_n5441_), .B(u2_o_307_), .C(u2__abc_52138_new_n9844_), .Y(u2__abc_52138_new_n9854_));
OAI21X1 OAI21X1_2072 ( .A(u2__abc_52138_new_n5434_), .B(u2__abc_52138_new_n9854_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9855_));
OAI21X1 OAI21X1_2073 ( .A(u2__abc_52138_new_n5430_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9857_));
OAI21X1 OAI21X1_2074 ( .A(u2__abc_52138_new_n9857_), .B(u2__abc_52138_new_n9856_), .C(u2__abc_52138_new_n9859_), .Y(u2__abc_52138_new_n9860_));
OAI21X1 OAI21X1_2075 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_311_), .Y(u2__abc_52138_new_n9862_));
OAI21X1 OAI21X1_2076 ( .A(u2__abc_52138_new_n5442_), .B(u2__abc_52138_new_n9845_), .C(u2__abc_52138_new_n5434_), .Y(u2__abc_52138_new_n9863_));
OAI21X1 OAI21X1_2077 ( .A(u2__abc_52138_new_n5430_), .B(u2_o_308_), .C(u2__abc_52138_new_n9863_), .Y(u2__abc_52138_new_n9864_));
OAI21X1 OAI21X1_2078 ( .A(u2__abc_52138_new_n5439_), .B(u2__abc_52138_new_n9864_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9865_));
OAI21X1 OAI21X1_2079 ( .A(u2__abc_52138_new_n5435_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9867_));
OAI21X1 OAI21X1_208 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1408_), .C(_abc_65734_new_n1409_), .Y(fracta1_96_));
OAI21X1 OAI21X1_2080 ( .A(u2__abc_52138_new_n9867_), .B(u2__abc_52138_new_n9866_), .C(u2__abc_52138_new_n9868_), .Y(u2__abc_52138_new_n9869_));
OAI21X1 OAI21X1_2081 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_312_), .Y(u2__abc_52138_new_n9871_));
OAI21X1 OAI21X1_2082 ( .A(u2__abc_52138_new_n5440_), .B(u2__abc_52138_new_n9872_), .C(u2__abc_52138_new_n9873_), .Y(u2__abc_52138_new_n9874_));
OAI21X1 OAI21X1_2083 ( .A(u2__abc_52138_new_n5453_), .B(u2__abc_52138_new_n9803_), .C(u2__abc_52138_new_n9875_), .Y(u2__abc_52138_new_n9876_));
OAI21X1 OAI21X1_2084 ( .A(u2__abc_52138_new_n5379_), .B(u2__abc_52138_new_n9876_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9879_));
OAI21X1 OAI21X1_2085 ( .A(u2__abc_52138_new_n9858_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9881_));
OAI21X1 OAI21X1_2086 ( .A(u2__abc_52138_new_n9881_), .B(u2__abc_52138_new_n9880_), .C(u2__abc_52138_new_n9882_), .Y(u2__abc_52138_new_n9883_));
OAI21X1 OAI21X1_2087 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_313_), .Y(u2__abc_52138_new_n9885_));
OAI21X1 OAI21X1_2088 ( .A(u2__abc_52138_new_n9858_), .B(u2_o_310_), .C(u2__abc_52138_new_n9877_), .Y(u2__abc_52138_new_n9886_));
OAI21X1 OAI21X1_2089 ( .A(u2__abc_52138_new_n5380_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9889_));
OAI21X1 OAI21X1_209 ( .A(\a[112] ), .B(_abc_65734_new_n1408_), .C(_abc_65734_new_n1411_), .Y(fracta1_97_));
OAI21X1 OAI21X1_2090 ( .A(u2__abc_52138_new_n9889_), .B(u2__abc_52138_new_n9888_), .C(u2__abc_52138_new_n9890_), .Y(u2__abc_52138_new_n9891_));
OAI21X1 OAI21X1_2091 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_314_), .Y(u2__abc_52138_new_n9893_));
OAI21X1 OAI21X1_2092 ( .A(u2__abc_52138_new_n9858_), .B(u2_o_310_), .C(u2__abc_52138_new_n9894_), .Y(u2__abc_52138_new_n9895_));
OAI21X1 OAI21X1_2093 ( .A(u2__abc_52138_new_n9895_), .B(u2__abc_52138_new_n9878_), .C(u2__abc_52138_new_n5812_), .Y(u2__abc_52138_new_n9896_));
OAI21X1 OAI21X1_2094 ( .A(u2__abc_52138_new_n5372_), .B(u2__abc_52138_new_n9897_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9898_));
OAI21X1 OAI21X1_2095 ( .A(u2__abc_52138_new_n5368_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9900_));
OAI21X1 OAI21X1_2096 ( .A(u2__abc_52138_new_n9900_), .B(u2__abc_52138_new_n9899_), .C(u2__abc_52138_new_n9901_), .Y(u2__abc_52138_new_n9902_));
OAI21X1 OAI21X1_2097 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_315_), .Y(u2__abc_52138_new_n9904_));
OAI21X1 OAI21X1_2098 ( .A(u2__abc_52138_new_n5371_), .B(u2__abc_52138_new_n9896_), .C(u2__abc_52138_new_n9905_), .Y(u2__abc_52138_new_n9906_));
OAI21X1 OAI21X1_2099 ( .A(u2__abc_52138_new_n5377_), .B(u2__abc_52138_new_n9906_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9907_));
OAI21X1 OAI21X1_21 ( .A(aNan), .B(_abc_65734_new_n890_), .C(_abc_65734_new_n891_), .Y(\o[132] ));
OAI21X1 OAI21X1_210 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1413_), .C(_abc_65734_new_n1414_), .Y(fracta1_98_));
OAI21X1 OAI21X1_2100 ( .A(u2__abc_52138_new_n5373_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9909_));
OAI21X1 OAI21X1_2101 ( .A(u2__abc_52138_new_n9909_), .B(u2__abc_52138_new_n9908_), .C(u2__abc_52138_new_n9910_), .Y(u2__abc_52138_new_n9911_));
OAI21X1 OAI21X1_2102 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_316_), .Y(u2__abc_52138_new_n9913_));
OAI21X1 OAI21X1_2103 ( .A(u2_remHi_311_), .B(u2__abc_52138_new_n5382_), .C(u2__abc_52138_new_n9895_), .Y(u2__abc_52138_new_n9914_));
OAI21X1 OAI21X1_2104 ( .A(u2__abc_52138_new_n5378_), .B(u2__abc_52138_new_n9914_), .C(u2__abc_52138_new_n9915_), .Y(u2__abc_52138_new_n9916_));
OAI21X1 OAI21X1_2105 ( .A(u2__abc_52138_new_n5398_), .B(u2__abc_52138_new_n9919_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9922_));
OAI21X1 OAI21X1_2106 ( .A(u2__abc_52138_new_n5818_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9924_));
OAI21X1 OAI21X1_2107 ( .A(u2__abc_52138_new_n9924_), .B(u2__abc_52138_new_n9923_), .C(u2__abc_52138_new_n9925_), .Y(u2__abc_52138_new_n9926_));
OAI21X1 OAI21X1_2108 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_317_), .Y(u2__abc_52138_new_n9928_));
OAI21X1 OAI21X1_2109 ( .A(u2__abc_52138_new_n5818_), .B(u2_o_314_), .C(u2__abc_52138_new_n9920_), .Y(u2__abc_52138_new_n9929_));
OAI21X1 OAI21X1_211 ( .A(\a[112] ), .B(_abc_65734_new_n1413_), .C(_abc_65734_new_n1416_), .Y(fracta1_99_));
OAI21X1 OAI21X1_2110 ( .A(u2__abc_52138_new_n5399_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9932_));
OAI21X1 OAI21X1_2111 ( .A(u2__abc_52138_new_n9932_), .B(u2__abc_52138_new_n9931_), .C(u2__abc_52138_new_n9933_), .Y(u2__abc_52138_new_n9934_));
OAI21X1 OAI21X1_2112 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_318_), .Y(u2__abc_52138_new_n9936_));
OAI21X1 OAI21X1_2113 ( .A(u2__abc_52138_new_n5818_), .B(u2_o_314_), .C(u2__abc_52138_new_n9937_), .Y(u2__abc_52138_new_n9938_));
OAI21X1 OAI21X1_2114 ( .A(u2__abc_52138_new_n9938_), .B(u2__abc_52138_new_n9921_), .C(u2__abc_52138_new_n5820_), .Y(u2__abc_52138_new_n9939_));
OAI21X1 OAI21X1_2115 ( .A(u2__abc_52138_new_n5391_), .B(u2__abc_52138_new_n9940_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9941_));
OAI21X1 OAI21X1_2116 ( .A(u2__abc_52138_new_n5387_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9943_));
OAI21X1 OAI21X1_2117 ( .A(u2__abc_52138_new_n9943_), .B(u2__abc_52138_new_n9942_), .C(u2__abc_52138_new_n9944_), .Y(u2__abc_52138_new_n9945_));
OAI21X1 OAI21X1_2118 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_319_), .Y(u2__abc_52138_new_n9947_));
OAI21X1 OAI21X1_2119 ( .A(u2__abc_52138_new_n5390_), .B(u2__abc_52138_new_n9939_), .C(u2__abc_52138_new_n9948_), .Y(u2__abc_52138_new_n9949_));
OAI21X1 OAI21X1_212 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1418_), .C(_abc_65734_new_n1419_), .Y(fracta1_100_));
OAI21X1 OAI21X1_2120 ( .A(u2__abc_52138_new_n5396_), .B(u2__abc_52138_new_n9949_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9950_));
OAI21X1 OAI21X1_2121 ( .A(u2__abc_52138_new_n5392_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9952_));
OAI21X1 OAI21X1_2122 ( .A(u2__abc_52138_new_n9952_), .B(u2__abc_52138_new_n9951_), .C(u2__abc_52138_new_n9953_), .Y(u2__abc_52138_new_n9954_));
OAI21X1 OAI21X1_2123 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_320_), .Y(u2__abc_52138_new_n9956_));
OAI21X1 OAI21X1_2124 ( .A(u2__abc_52138_new_n9613_), .B(u2__abc_52138_new_n9618_), .C(u2__abc_52138_new_n5547_), .Y(u2__abc_52138_new_n9957_));
OAI21X1 OAI21X1_2125 ( .A(u2__abc_52138_new_n5395_), .B(u2__abc_52138_new_n9948_), .C(u2__abc_52138_new_n5808_), .Y(u2__abc_52138_new_n9961_));
OAI21X1 OAI21X1_2126 ( .A(u2__abc_52138_new_n5406_), .B(u2__abc_52138_new_n9875_), .C(u2__abc_52138_new_n9962_), .Y(u2__abc_52138_new_n9963_));
OAI21X1 OAI21X1_2127 ( .A(u2__abc_52138_new_n5345_), .B(u2__abc_52138_new_n9968_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9969_));
OAI21X1 OAI21X1_2128 ( .A(u2__abc_52138_new_n5343_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9971_));
OAI21X1 OAI21X1_2129 ( .A(u2__abc_52138_new_n9971_), .B(u2__abc_52138_new_n9970_), .C(u2__abc_52138_new_n9972_), .Y(u2__abc_52138_new_n9973_));
OAI21X1 OAI21X1_213 ( .A(\a[112] ), .B(_abc_65734_new_n1418_), .C(_abc_65734_new_n1421_), .Y(fracta1_101_));
OAI21X1 OAI21X1_2130 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_321_), .Y(u2__abc_52138_new_n9975_));
OAI21X1 OAI21X1_2131 ( .A(u2__abc_52138_new_n5342_), .B(u2__abc_52138_new_n9967_), .C(u2__abc_52138_new_n9976_), .Y(u2__abc_52138_new_n9977_));
OAI21X1 OAI21X1_2132 ( .A(u2__abc_52138_new_n5350_), .B(u2__abc_52138_new_n9977_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9978_));
OAI21X1 OAI21X1_2133 ( .A(u2__abc_52138_new_n5346_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9980_));
OAI21X1 OAI21X1_2134 ( .A(u2__abc_52138_new_n9980_), .B(u2__abc_52138_new_n9979_), .C(u2__abc_52138_new_n9981_), .Y(u2__abc_52138_new_n9982_));
OAI21X1 OAI21X1_2135 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_322_), .Y(u2__abc_52138_new_n9984_));
OAI21X1 OAI21X1_2136 ( .A(u2__abc_52138_new_n9976_), .B(u2__abc_52138_new_n9985_), .C(u2__abc_52138_new_n5349_), .Y(u2__abc_52138_new_n9986_));
OAI21X1 OAI21X1_2137 ( .A(u2__abc_52138_new_n5351_), .B(u2__abc_52138_new_n9967_), .C(u2__abc_52138_new_n9987_), .Y(u2__abc_52138_new_n9988_));
OAI21X1 OAI21X1_2138 ( .A(u2__abc_52138_new_n5356_), .B(u2__abc_52138_new_n9988_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9989_));
OAI21X1 OAI21X1_2139 ( .A(u2__abc_52138_new_n5352_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n9991_));
OAI21X1 OAI21X1_214 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1423_), .C(_abc_65734_new_n1424_), .Y(fracta1_102_));
OAI21X1 OAI21X1_2140 ( .A(u2__abc_52138_new_n9991_), .B(u2__abc_52138_new_n9990_), .C(u2__abc_52138_new_n9993_), .Y(u2__abc_52138_new_n9994_));
OAI21X1 OAI21X1_2141 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_323_), .Y(u2__abc_52138_new_n9996_));
OAI21X1 OAI21X1_2142 ( .A(u2__abc_52138_new_n5352_), .B(u2_o_320_), .C(u2__abc_52138_new_n9997_), .Y(u2__abc_52138_new_n9998_));
OAI21X1 OAI21X1_2143 ( .A(u2__abc_52138_new_n5361_), .B(u2__abc_52138_new_n9998_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n9999_));
OAI21X1 OAI21X1_2144 ( .A(u2__abc_52138_new_n5357_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10001_));
OAI21X1 OAI21X1_2145 ( .A(u2__abc_52138_new_n10001_), .B(u2__abc_52138_new_n10000_), .C(u2__abc_52138_new_n10002_), .Y(u2__abc_52138_new_n10003_));
OAI21X1 OAI21X1_2146 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_324_), .Y(u2__abc_52138_new_n10005_));
OAI21X1 OAI21X1_2147 ( .A(u2__abc_52138_new_n5362_), .B(u2__abc_52138_new_n9987_), .C(u2__abc_52138_new_n10006_), .Y(u2__abc_52138_new_n10007_));
OAI21X1 OAI21X1_2148 ( .A(u2__abc_52138_new_n5363_), .B(u2__abc_52138_new_n9967_), .C(u2__abc_52138_new_n10008_), .Y(u2__abc_52138_new_n10009_));
OAI21X1 OAI21X1_2149 ( .A(u2__abc_52138_new_n5332_), .B(u2__abc_52138_new_n10009_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10012_));
OAI21X1 OAI21X1_215 ( .A(\a[112] ), .B(_abc_65734_new_n1423_), .C(_abc_65734_new_n1426_), .Y(fracta1_103_));
OAI21X1 OAI21X1_2150 ( .A(u2__abc_52138_new_n9992_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10014_));
OAI21X1 OAI21X1_2151 ( .A(u2__abc_52138_new_n10014_), .B(u2__abc_52138_new_n10013_), .C(u2__abc_52138_new_n10015_), .Y(u2__abc_52138_new_n10016_));
OAI21X1 OAI21X1_2152 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_325_), .Y(u2__abc_52138_new_n10018_));
OAI21X1 OAI21X1_2153 ( .A(u2__abc_52138_new_n9992_), .B(u2_o_322_), .C(u2__abc_52138_new_n10010_), .Y(u2__abc_52138_new_n10019_));
OAI21X1 OAI21X1_2154 ( .A(u2__abc_52138_new_n5335_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10022_));
OAI21X1 OAI21X1_2155 ( .A(u2__abc_52138_new_n10022_), .B(u2__abc_52138_new_n10021_), .C(u2__abc_52138_new_n10023_), .Y(u2__abc_52138_new_n10024_));
OAI21X1 OAI21X1_2156 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_326_), .Y(u2__abc_52138_new_n10026_));
OAI21X1 OAI21X1_2157 ( .A(u2__abc_52138_new_n9992_), .B(u2_o_322_), .C(u2__abc_52138_new_n5334_), .Y(u2__abc_52138_new_n10027_));
OAI21X1 OAI21X1_2158 ( .A(u2__abc_52138_new_n10027_), .B(u2__abc_52138_new_n10011_), .C(u2__abc_52138_new_n5336_), .Y(u2__abc_52138_new_n10028_));
OAI21X1 OAI21X1_2159 ( .A(u2__abc_52138_new_n5325_), .B(u2__abc_52138_new_n10029_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10030_));
OAI21X1 OAI21X1_216 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1428_), .C(_abc_65734_new_n1429_), .Y(fracta1_104_));
OAI21X1 OAI21X1_2160 ( .A(u2__abc_52138_new_n5323_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10032_));
OAI21X1 OAI21X1_2161 ( .A(u2__abc_52138_new_n10032_), .B(u2__abc_52138_new_n10031_), .C(u2__abc_52138_new_n10033_), .Y(u2__abc_52138_new_n10034_));
OAI21X1 OAI21X1_2162 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_327_), .Y(u2__abc_52138_new_n10036_));
OAI21X1 OAI21X1_2163 ( .A(u2__abc_52138_new_n5322_), .B(u2__abc_52138_new_n10028_), .C(u2__abc_52138_new_n10037_), .Y(u2__abc_52138_new_n10038_));
OAI21X1 OAI21X1_2164 ( .A(u2__abc_52138_new_n5330_), .B(u2__abc_52138_new_n10038_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10039_));
OAI21X1 OAI21X1_2165 ( .A(u2__abc_52138_new_n5328_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10041_));
OAI21X1 OAI21X1_2166 ( .A(u2__abc_52138_new_n10041_), .B(u2__abc_52138_new_n10040_), .C(u2__abc_52138_new_n10042_), .Y(u2__abc_52138_new_n10043_));
OAI21X1 OAI21X1_2167 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_328_), .Y(u2__abc_52138_new_n10045_));
OAI21X1 OAI21X1_2168 ( .A(u2_remHi_323_), .B(u2__abc_52138_new_n5333_), .C(u2__abc_52138_new_n10027_), .Y(u2__abc_52138_new_n10047_));
OAI21X1 OAI21X1_2169 ( .A(u2__abc_52138_new_n10047_), .B(u2__abc_52138_new_n5331_), .C(u2__abc_52138_new_n10048_), .Y(u2__abc_52138_new_n10049_));
OAI21X1 OAI21X1_217 ( .A(\a[112] ), .B(_abc_65734_new_n1428_), .C(_abc_65734_new_n1431_), .Y(fracta1_105_));
OAI21X1 OAI21X1_2170 ( .A(u2__abc_52138_new_n9965_), .B(u2__abc_52138_new_n9966_), .C(u2__abc_52138_new_n5364_), .Y(u2__abc_52138_new_n10051_));
OAI21X1 OAI21X1_2171 ( .A(u2__abc_52138_new_n5278_), .B(u2__abc_52138_new_n10052_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10053_));
OAI21X1 OAI21X1_2172 ( .A(u2__abc_52138_new_n5276_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10055_));
OAI21X1 OAI21X1_2173 ( .A(u2__abc_52138_new_n10055_), .B(u2__abc_52138_new_n10054_), .C(u2__abc_52138_new_n10056_), .Y(u2__abc_52138_new_n10057_));
OAI21X1 OAI21X1_2174 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_329_), .Y(u2__abc_52138_new_n10059_));
OAI21X1 OAI21X1_2175 ( .A(u2__abc_52138_new_n5275_), .B(u2__abc_52138_new_n10061_), .C(u2__abc_52138_new_n10060_), .Y(u2__abc_52138_new_n10062_));
OAI21X1 OAI21X1_2176 ( .A(u2__abc_52138_new_n5283_), .B(u2__abc_52138_new_n10062_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10063_));
OAI21X1 OAI21X1_2177 ( .A(u2__abc_52138_new_n5279_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10065_));
OAI21X1 OAI21X1_2178 ( .A(u2__abc_52138_new_n10065_), .B(u2__abc_52138_new_n10064_), .C(u2__abc_52138_new_n10066_), .Y(u2__abc_52138_new_n10067_));
OAI21X1 OAI21X1_2179 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_330_), .Y(u2__abc_52138_new_n10069_));
OAI21X1 OAI21X1_218 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1433_), .C(_abc_65734_new_n1434_), .Y(fracta1_106_));
OAI21X1 OAI21X1_2180 ( .A(u2__abc_52138_new_n5276_), .B(u2_o_326_), .C(u2__abc_52138_new_n5282_), .Y(u2__abc_52138_new_n10070_));
OAI21X1 OAI21X1_2181 ( .A(u2_remHi_327_), .B(u2__abc_52138_new_n5281_), .C(u2__abc_52138_new_n10070_), .Y(u2__abc_52138_new_n10071_));
OAI21X1 OAI21X1_2182 ( .A(u2__abc_52138_new_n5284_), .B(u2__abc_52138_new_n10061_), .C(u2__abc_52138_new_n10071_), .Y(u2__abc_52138_new_n10072_));
OAI21X1 OAI21X1_2183 ( .A(u2__abc_52138_new_n5289_), .B(u2__abc_52138_new_n10072_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10073_));
OAI21X1 OAI21X1_2184 ( .A(u2__abc_52138_new_n5285_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10075_));
OAI21X1 OAI21X1_2185 ( .A(u2__abc_52138_new_n10075_), .B(u2__abc_52138_new_n10074_), .C(u2__abc_52138_new_n10076_), .Y(u2__abc_52138_new_n10077_));
OAI21X1 OAI21X1_2186 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_331_), .Y(u2__abc_52138_new_n10079_));
OAI21X1 OAI21X1_2187 ( .A(u2__abc_52138_new_n5285_), .B(u2_o_328_), .C(u2__abc_52138_new_n10080_), .Y(u2__abc_52138_new_n10081_));
OAI21X1 OAI21X1_2188 ( .A(u2__abc_52138_new_n5294_), .B(u2__abc_52138_new_n10081_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10082_));
OAI21X1 OAI21X1_2189 ( .A(u2__abc_52138_new_n5290_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10084_));
OAI21X1 OAI21X1_219 ( .A(\a[112] ), .B(_abc_65734_new_n1433_), .C(_abc_65734_new_n1436_), .Y(fracta1_107_));
OAI21X1 OAI21X1_2190 ( .A(u2__abc_52138_new_n10084_), .B(u2__abc_52138_new_n10083_), .C(u2__abc_52138_new_n10085_), .Y(u2__abc_52138_new_n10086_));
OAI21X1 OAI21X1_2191 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_332_), .Y(u2__abc_52138_new_n10088_));
OAI21X1 OAI21X1_2192 ( .A(u2__abc_52138_new_n10071_), .B(u2__abc_52138_new_n5295_), .C(u2__abc_52138_new_n10089_), .Y(u2__abc_52138_new_n10090_));
OAI21X1 OAI21X1_2193 ( .A(u2__abc_52138_new_n5312_), .B(u2__abc_52138_new_n10092_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10095_));
OAI21X1 OAI21X1_2194 ( .A(u2__abc_52138_new_n5308_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10097_));
OAI21X1 OAI21X1_2195 ( .A(u2__abc_52138_new_n10097_), .B(u2__abc_52138_new_n10096_), .C(u2__abc_52138_new_n10098_), .Y(u2__abc_52138_new_n10099_));
OAI21X1 OAI21X1_2196 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_333_), .Y(u2__abc_52138_new_n10101_));
OAI21X1 OAI21X1_2197 ( .A(u2__abc_52138_new_n5311_), .B(u2__abc_52138_new_n10091_), .C(u2__abc_52138_new_n10102_), .Y(u2__abc_52138_new_n10103_));
OAI21X1 OAI21X1_2198 ( .A(u2__abc_52138_new_n5313_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10106_));
OAI21X1 OAI21X1_2199 ( .A(u2__abc_52138_new_n10106_), .B(u2__abc_52138_new_n10105_), .C(u2__abc_52138_new_n10107_), .Y(u2__abc_52138_new_n10108_));
OAI21X1 OAI21X1_22 ( .A(aNan), .B(_abc_65734_new_n893_), .C(_abc_65734_new_n894_), .Y(\o[133] ));
OAI21X1 OAI21X1_220 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1438_), .C(_abc_65734_new_n1439_), .Y(fracta1_108_));
OAI21X1 OAI21X1_2200 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_334_), .Y(u2__abc_52138_new_n10110_));
OAI21X1 OAI21X1_2201 ( .A(u2__abc_52138_new_n5313_), .B(u2_o_331_), .C(u2__abc_52138_new_n10102_), .Y(u2__abc_52138_new_n10111_));
OAI21X1 OAI21X1_2202 ( .A(u2__abc_52138_new_n10111_), .B(u2__abc_52138_new_n10094_), .C(u2__abc_52138_new_n10112_), .Y(u2__abc_52138_new_n10113_));
OAI21X1 OAI21X1_2203 ( .A(u2__abc_52138_new_n5301_), .B(u2__abc_52138_new_n10114_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10115_));
OAI21X1 OAI21X1_2204 ( .A(u2__abc_52138_new_n5297_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10117_));
OAI21X1 OAI21X1_2205 ( .A(u2__abc_52138_new_n10117_), .B(u2__abc_52138_new_n10116_), .C(u2__abc_52138_new_n10118_), .Y(u2__abc_52138_new_n10119_));
OAI21X1 OAI21X1_2206 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_335_), .Y(u2__abc_52138_new_n10121_));
OAI21X1 OAI21X1_2207 ( .A(u2__abc_52138_new_n5300_), .B(u2__abc_52138_new_n10113_), .C(u2__abc_52138_new_n10122_), .Y(u2__abc_52138_new_n10123_));
OAI21X1 OAI21X1_2208 ( .A(u2__abc_52138_new_n5306_), .B(u2__abc_52138_new_n10123_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10124_));
OAI21X1 OAI21X1_2209 ( .A(u2__abc_52138_new_n5302_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10126_));
OAI21X1 OAI21X1_221 ( .A(\a[112] ), .B(_abc_65734_new_n1438_), .C(_abc_65734_new_n1441_), .Y(fracta1_109_));
OAI21X1 OAI21X1_2210 ( .A(u2__abc_52138_new_n10126_), .B(u2__abc_52138_new_n10125_), .C(u2__abc_52138_new_n10127_), .Y(u2__abc_52138_new_n10128_));
OAI21X1 OAI21X1_2211 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_336_), .Y(u2__abc_52138_new_n10130_));
OAI21X1 OAI21X1_2212 ( .A(u2_remHi_333_), .B(u2__abc_52138_new_n5304_), .C(u2__abc_52138_new_n5298_), .Y(u2__abc_52138_new_n10133_));
OAI21X1 OAI21X1_2213 ( .A(u2__abc_52138_new_n5365_), .B(u2__abc_52138_new_n9967_), .C(u2__abc_52138_new_n10136_), .Y(u2__abc_52138_new_n10137_));
OAI21X1 OAI21X1_2214 ( .A(u2__abc_52138_new_n5241_), .B(u2__abc_52138_new_n10137_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10140_));
OAI21X1 OAI21X1_2215 ( .A(u2__abc_52138_new_n5874_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10142_));
OAI21X1 OAI21X1_2216 ( .A(u2__abc_52138_new_n10142_), .B(u2__abc_52138_new_n10141_), .C(u2__abc_52138_new_n10143_), .Y(u2__abc_52138_new_n10144_));
OAI21X1 OAI21X1_2217 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_337_), .Y(u2__abc_52138_new_n10146_));
OAI21X1 OAI21X1_2218 ( .A(u2__abc_52138_new_n5874_), .B(u2_o_334_), .C(u2__abc_52138_new_n10138_), .Y(u2__abc_52138_new_n10147_));
OAI21X1 OAI21X1_2219 ( .A(u2__abc_52138_new_n5244_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10150_));
OAI21X1 OAI21X1_222 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1443_), .C(_abc_65734_new_n1444_), .Y(fracta1_110_));
OAI21X1 OAI21X1_2220 ( .A(u2__abc_52138_new_n10150_), .B(u2__abc_52138_new_n10149_), .C(u2__abc_52138_new_n10151_), .Y(u2__abc_52138_new_n10152_));
OAI21X1 OAI21X1_2221 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_338_), .Y(u2__abc_52138_new_n10154_));
OAI21X1 OAI21X1_2222 ( .A(u2__abc_52138_new_n5874_), .B(u2_o_334_), .C(u2__abc_52138_new_n5243_), .Y(u2__abc_52138_new_n10155_));
OAI21X1 OAI21X1_2223 ( .A(u2__abc_52138_new_n10155_), .B(u2__abc_52138_new_n10139_), .C(u2__abc_52138_new_n5245_), .Y(u2__abc_52138_new_n10156_));
OAI21X1 OAI21X1_2224 ( .A(u2__abc_52138_new_n5233_), .B(u2__abc_52138_new_n10157_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10158_));
OAI21X1 OAI21X1_2225 ( .A(u2__abc_52138_new_n5229_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10160_));
OAI21X1 OAI21X1_2226 ( .A(u2__abc_52138_new_n10160_), .B(u2__abc_52138_new_n10159_), .C(u2__abc_52138_new_n10161_), .Y(u2__abc_52138_new_n10162_));
OAI21X1 OAI21X1_2227 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_339_), .Y(u2__abc_52138_new_n10164_));
OAI21X1 OAI21X1_2228 ( .A(u2__abc_52138_new_n5232_), .B(u2__abc_52138_new_n10156_), .C(u2__abc_52138_new_n10165_), .Y(u2__abc_52138_new_n10166_));
OAI21X1 OAI21X1_2229 ( .A(u2__abc_52138_new_n5238_), .B(u2__abc_52138_new_n10166_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10167_));
OAI21X1 OAI21X1_223 ( .A(\a[112] ), .B(_abc_65734_new_n1443_), .C(_abc_65734_new_n1446_), .Y(fracta1_111_));
OAI21X1 OAI21X1_2230 ( .A(u2__abc_52138_new_n5234_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10169_));
OAI21X1 OAI21X1_2231 ( .A(u2__abc_52138_new_n10169_), .B(u2__abc_52138_new_n10168_), .C(u2__abc_52138_new_n10170_), .Y(u2__abc_52138_new_n10171_));
OAI21X1 OAI21X1_2232 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_340_), .Y(u2__abc_52138_new_n10173_));
OAI21X1 OAI21X1_2233 ( .A(u2_remHi_335_), .B(u2__abc_52138_new_n5242_), .C(u2__abc_52138_new_n10155_), .Y(u2__abc_52138_new_n10175_));
OAI21X1 OAI21X1_2234 ( .A(u2__abc_52138_new_n5237_), .B(u2__abc_52138_new_n10165_), .C(u2__abc_52138_new_n5872_), .Y(u2__abc_52138_new_n10176_));
OAI21X1 OAI21X1_2235 ( .A(u2__abc_52138_new_n10175_), .B(u2__abc_52138_new_n5239_), .C(u2__abc_52138_new_n10177_), .Y(u2__abc_52138_new_n10178_));
OAI21X1 OAI21X1_2236 ( .A(u2__abc_52138_new_n5248_), .B(u2__abc_52138_new_n10174_), .C(u2__abc_52138_new_n10179_), .Y(u2__abc_52138_new_n10180_));
OAI21X1 OAI21X1_2237 ( .A(u2__abc_52138_new_n5265_), .B(u2__abc_52138_new_n10180_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10183_));
OAI21X1 OAI21X1_2238 ( .A(u2__abc_52138_new_n5261_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10185_));
OAI21X1 OAI21X1_2239 ( .A(u2__abc_52138_new_n10185_), .B(u2__abc_52138_new_n10184_), .C(u2__abc_52138_new_n10186_), .Y(u2__abc_52138_new_n10187_));
OAI21X1 OAI21X1_224 ( .A(_abc_65734_new_n1168_), .B(_abc_65734_new_n1448_), .C(_abc_65734_new_n1449_), .Y(fracta1_112_));
OAI21X1 OAI21X1_2240 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_341_), .Y(u2__abc_52138_new_n10189_));
OAI21X1 OAI21X1_2241 ( .A(u2__abc_52138_new_n5261_), .B(u2_o_338_), .C(u2__abc_52138_new_n10181_), .Y(u2__abc_52138_new_n10190_));
OAI21X1 OAI21X1_2242 ( .A(u2__abc_52138_new_n5266_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10193_));
OAI21X1 OAI21X1_2243 ( .A(u2__abc_52138_new_n10193_), .B(u2__abc_52138_new_n10192_), .C(u2__abc_52138_new_n10194_), .Y(u2__abc_52138_new_n10195_));
OAI21X1 OAI21X1_2244 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_342_), .Y(u2__abc_52138_new_n10197_));
OAI21X1 OAI21X1_2245 ( .A(u2__abc_52138_new_n5266_), .B(u2_o_339_), .C(u2__abc_52138_new_n5263_), .Y(u2__abc_52138_new_n10198_));
OAI21X1 OAI21X1_2246 ( .A(u2__abc_52138_new_n10198_), .B(u2__abc_52138_new_n10182_), .C(u2__abc_52138_new_n5880_), .Y(u2__abc_52138_new_n10199_));
OAI21X1 OAI21X1_2247 ( .A(u2__abc_52138_new_n5253_), .B(u2__abc_52138_new_n10200_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10201_));
OAI21X1 OAI21X1_2248 ( .A(u2__abc_52138_new_n5251_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10203_));
OAI21X1 OAI21X1_2249 ( .A(u2__abc_52138_new_n10203_), .B(u2__abc_52138_new_n10202_), .C(u2__abc_52138_new_n10204_), .Y(u2__abc_52138_new_n10205_));
OAI21X1 OAI21X1_225 ( .A(_abc_65734_new_n1453_), .B(_abc_65734_new_n1452_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1454_));
OAI21X1 OAI21X1_2250 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_343_), .Y(u2__abc_52138_new_n10207_));
OAI21X1 OAI21X1_2251 ( .A(u2__abc_52138_new_n10208_), .B(u2__abc_52138_new_n10199_), .C(u2__abc_52138_new_n5250_), .Y(u2__abc_52138_new_n10209_));
OAI21X1 OAI21X1_2252 ( .A(u2__abc_52138_new_n5258_), .B(u2__abc_52138_new_n10209_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10210_));
OAI21X1 OAI21X1_2253 ( .A(u2__abc_52138_new_n5254_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10212_));
OAI21X1 OAI21X1_2254 ( .A(u2__abc_52138_new_n10212_), .B(u2__abc_52138_new_n10211_), .C(u2__abc_52138_new_n10213_), .Y(u2__abc_52138_new_n10214_));
OAI21X1 OAI21X1_2255 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_344_), .Y(u2__abc_52138_new_n10216_));
OAI21X1 OAI21X1_2256 ( .A(u2__abc_52138_new_n5250_), .B(u2__abc_52138_new_n5257_), .C(u2__abc_52138_new_n10218_), .Y(u2__abc_52138_new_n10219_));
OAI21X1 OAI21X1_2257 ( .A(u2__abc_52138_new_n5271_), .B(u2__abc_52138_new_n10179_), .C(u2__abc_52138_new_n10220_), .Y(u2__abc_52138_new_n10221_));
OAI21X1 OAI21X1_2258 ( .A(u2__abc_52138_new_n5199_), .B(u2__abc_52138_new_n10223_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10226_));
OAI21X1 OAI21X1_2259 ( .A(u2__abc_52138_new_n5195_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10228_));
OAI21X1 OAI21X1_226 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1168_), .C(_abc_65734_new_n1454_), .Y(\o[226] ));
OAI21X1 OAI21X1_2260 ( .A(u2__abc_52138_new_n10228_), .B(u2__abc_52138_new_n10227_), .C(u2__abc_52138_new_n10229_), .Y(u2__abc_52138_new_n10230_));
OAI21X1 OAI21X1_2261 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_345_), .Y(u2__abc_52138_new_n10232_));
OAI21X1 OAI21X1_2262 ( .A(u2__abc_52138_new_n5198_), .B(u2__abc_52138_new_n10222_), .C(u2__abc_52138_new_n10233_), .Y(u2__abc_52138_new_n10234_));
OAI21X1 OAI21X1_2263 ( .A(u2__abc_52138_new_n5200_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10237_));
OAI21X1 OAI21X1_2264 ( .A(u2__abc_52138_new_n10237_), .B(u2__abc_52138_new_n10236_), .C(u2__abc_52138_new_n10238_), .Y(u2__abc_52138_new_n10239_));
OAI21X1 OAI21X1_2265 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_346_), .Y(u2__abc_52138_new_n10241_));
OAI21X1 OAI21X1_2266 ( .A(u2__abc_52138_new_n5200_), .B(u2_o_343_), .C(u2__abc_52138_new_n10233_), .Y(u2__abc_52138_new_n10242_));
OAI21X1 OAI21X1_2267 ( .A(u2__abc_52138_new_n10242_), .B(u2__abc_52138_new_n10225_), .C(u2__abc_52138_new_n10243_), .Y(u2__abc_52138_new_n10244_));
OAI21X1 OAI21X1_2268 ( .A(u2__abc_52138_new_n5187_), .B(u2__abc_52138_new_n10245_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10246_));
OAI21X1 OAI21X1_2269 ( .A(u2__abc_52138_new_n5185_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10248_));
OAI21X1 OAI21X1_227 ( .A(\a[112] ), .B(_abc_65734_new_n1458_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1459_));
OAI21X1 OAI21X1_2270 ( .A(u2__abc_52138_new_n10248_), .B(u2__abc_52138_new_n10247_), .C(u2__abc_52138_new_n10249_), .Y(u2__abc_52138_new_n10250_));
OAI21X1 OAI21X1_2271 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_347_), .Y(u2__abc_52138_new_n10252_));
OAI21X1 OAI21X1_2272 ( .A(u2__abc_52138_new_n10253_), .B(u2__abc_52138_new_n10244_), .C(u2__abc_52138_new_n5184_), .Y(u2__abc_52138_new_n10254_));
OAI21X1 OAI21X1_2273 ( .A(u2__abc_52138_new_n5192_), .B(u2__abc_52138_new_n10254_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10255_));
OAI21X1 OAI21X1_2274 ( .A(u2__abc_52138_new_n5188_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10257_));
OAI21X1 OAI21X1_2275 ( .A(u2__abc_52138_new_n10257_), .B(u2__abc_52138_new_n10256_), .C(u2__abc_52138_new_n10258_), .Y(u2__abc_52138_new_n10259_));
OAI21X1 OAI21X1_2276 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_348_), .Y(u2__abc_52138_new_n10261_));
OAI21X1 OAI21X1_2277 ( .A(u2_remHi_343_), .B(u2__abc_52138_new_n5202_), .C(u2__abc_52138_new_n10242_), .Y(u2__abc_52138_new_n10262_));
OAI21X1 OAI21X1_2278 ( .A(u2__abc_52138_new_n5193_), .B(u2__abc_52138_new_n10262_), .C(u2__abc_52138_new_n10264_), .Y(u2__abc_52138_new_n10265_));
OAI21X1 OAI21X1_2279 ( .A(u2__abc_52138_new_n5205_), .B(u2__abc_52138_new_n10222_), .C(u2__abc_52138_new_n10266_), .Y(u2__abc_52138_new_n10267_));
OAI21X1 OAI21X1_228 ( .A(_abc_65734_new_n1461_), .B(_abc_65734_new_n1462_), .C(_abc_65734_new_n1464_), .Y(_abc_65734_new_n1465_));
OAI21X1 OAI21X1_2280 ( .A(u2__abc_52138_new_n5220_), .B(u2__abc_52138_new_n10267_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10270_));
OAI21X1 OAI21X1_2281 ( .A(u2__abc_52138_new_n5216_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10272_));
OAI21X1 OAI21X1_2282 ( .A(u2__abc_52138_new_n10272_), .B(u2__abc_52138_new_n10271_), .C(u2__abc_52138_new_n10273_), .Y(u2__abc_52138_new_n10274_));
OAI21X1 OAI21X1_2283 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_349_), .Y(u2__abc_52138_new_n10276_));
OAI21X1 OAI21X1_2284 ( .A(u2__abc_52138_new_n5216_), .B(u2_o_346_), .C(u2__abc_52138_new_n10268_), .Y(u2__abc_52138_new_n10277_));
OAI21X1 OAI21X1_2285 ( .A(u2__abc_52138_new_n5221_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10280_));
OAI21X1 OAI21X1_2286 ( .A(u2__abc_52138_new_n10280_), .B(u2__abc_52138_new_n10279_), .C(u2__abc_52138_new_n10281_), .Y(u2__abc_52138_new_n10282_));
OAI21X1 OAI21X1_2287 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_350_), .Y(u2__abc_52138_new_n10284_));
OAI21X1 OAI21X1_2288 ( .A(u2__abc_52138_new_n10286_), .B(u2__abc_52138_new_n10269_), .C(u2__abc_52138_new_n5865_), .Y(u2__abc_52138_new_n10287_));
OAI21X1 OAI21X1_2289 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n10289_), .Y(u2__abc_52138_new_n10290_));
OAI21X1 OAI21X1_229 ( .A(_abc_65734_new_n1465_), .B(_abc_65734_new_n1467_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1468_));
OAI21X1 OAI21X1_2290 ( .A(u2__abc_52138_new_n5208_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10292_));
OAI21X1 OAI21X1_2291 ( .A(u2__abc_52138_new_n10292_), .B(u2__abc_52138_new_n10291_), .C(u2__abc_52138_new_n10293_), .Y(u2__abc_52138_new_n10294_));
OAI21X1 OAI21X1_2292 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_351_), .Y(u2__abc_52138_new_n10296_));
OAI21X1 OAI21X1_2293 ( .A(u2__abc_52138_new_n10285_), .B(u2__abc_52138_new_n10287_), .C(u2__abc_52138_new_n5207_), .Y(u2__abc_52138_new_n10297_));
OAI21X1 OAI21X1_2294 ( .A(u2__abc_52138_new_n5214_), .B(u2__abc_52138_new_n10297_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10298_));
OAI21X1 OAI21X1_2295 ( .A(u2__abc_52138_new_n5210_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10300_));
OAI21X1 OAI21X1_2296 ( .A(u2__abc_52138_new_n10300_), .B(u2__abc_52138_new_n10299_), .C(u2__abc_52138_new_n10301_), .Y(u2__abc_52138_new_n10302_));
OAI21X1 OAI21X1_2297 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_352_), .Y(u2__abc_52138_new_n10304_));
OAI21X1 OAI21X1_2298 ( .A(u2_remHi_347_), .B(u2__abc_52138_new_n5223_), .C(u2__abc_52138_new_n10286_), .Y(u2__abc_52138_new_n10306_));
OAI21X1 OAI21X1_2299 ( .A(u2__abc_52138_new_n5273_), .B(u2__abc_52138_new_n10136_), .C(u2__abc_52138_new_n10309_), .Y(u2__abc_52138_new_n10310_));
OAI21X1 OAI21X1_23 ( .A(aNan), .B(_abc_65734_new_n896_), .C(_abc_65734_new_n897_), .Y(\o[134] ));
OAI21X1 OAI21X1_230 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1458_), .C(_abc_65734_new_n1468_), .Y(\o[228] ));
OAI21X1 OAI21X1_2300 ( .A(u2__abc_52138_new_n9965_), .B(u2__abc_52138_new_n9966_), .C(u2__abc_52138_new_n5366_), .Y(u2__abc_52138_new_n10312_));
OAI21X1 OAI21X1_2301 ( .A(u2__abc_52138_new_n5149_), .B(u2__abc_52138_new_n10313_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10316_));
OAI21X1 OAI21X1_2302 ( .A(u2__abc_52138_new_n5145_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10318_));
OAI21X1 OAI21X1_2303 ( .A(u2__abc_52138_new_n10318_), .B(u2__abc_52138_new_n10317_), .C(u2__abc_52138_new_n10319_), .Y(u2__abc_52138_new_n10320_));
OAI21X1 OAI21X1_2304 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_353_), .Y(u2__abc_52138_new_n10322_));
OAI21X1 OAI21X1_2305 ( .A(u2__abc_52138_new_n5145_), .B(u2_o_350_), .C(u2__abc_52138_new_n10314_), .Y(u2__abc_52138_new_n10323_));
OAI21X1 OAI21X1_2306 ( .A(u2__abc_52138_new_n5150_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10326_));
OAI21X1 OAI21X1_2307 ( .A(u2__abc_52138_new_n10326_), .B(u2__abc_52138_new_n10325_), .C(u2__abc_52138_new_n10327_), .Y(u2__abc_52138_new_n10328_));
OAI21X1 OAI21X1_2308 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_354_), .Y(u2__abc_52138_new_n10330_));
OAI21X1 OAI21X1_2309 ( .A(u2__abc_52138_new_n5145_), .B(u2_o_350_), .C(u2__abc_52138_new_n5920_), .Y(u2__abc_52138_new_n10331_));
OAI21X1 OAI21X1_231 ( .A(_abc_65734_new_n1461_), .B(_abc_65734_new_n1462_), .C(_abc_65734_new_n1473_), .Y(_abc_65734_new_n1474_));
OAI21X1 OAI21X1_2310 ( .A(u2__abc_52138_new_n5138_), .B(u2__abc_52138_new_n10333_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10334_));
OAI21X1 OAI21X1_2311 ( .A(u2__abc_52138_new_n5134_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10336_));
OAI21X1 OAI21X1_2312 ( .A(u2__abc_52138_new_n10336_), .B(u2__abc_52138_new_n10335_), .C(u2__abc_52138_new_n10337_), .Y(u2__abc_52138_new_n10338_));
OAI21X1 OAI21X1_2313 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_355_), .Y(u2__abc_52138_new_n10340_));
OAI21X1 OAI21X1_2314 ( .A(u2__abc_52138_new_n5137_), .B(u2__abc_52138_new_n10332_), .C(u2__abc_52138_new_n10341_), .Y(u2__abc_52138_new_n10342_));
OAI21X1 OAI21X1_2315 ( .A(u2__abc_52138_new_n5143_), .B(u2__abc_52138_new_n10342_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10343_));
OAI21X1 OAI21X1_2316 ( .A(u2__abc_52138_new_n5139_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10345_));
OAI21X1 OAI21X1_2317 ( .A(u2__abc_52138_new_n10345_), .B(u2__abc_52138_new_n10344_), .C(u2__abc_52138_new_n10346_), .Y(u2__abc_52138_new_n10347_));
OAI21X1 OAI21X1_2318 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_356_), .Y(u2__abc_52138_new_n10349_));
OAI21X1 OAI21X1_2319 ( .A(u2_remHi_351_), .B(u2__abc_52138_new_n5152_), .C(u2__abc_52138_new_n10331_), .Y(u2__abc_52138_new_n10350_));
OAI21X1 OAI21X1_232 ( .A(_abc_65734_new_n1475_), .B(_abc_65734_new_n1476_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1477_));
OAI21X1 OAI21X1_2320 ( .A(u2__abc_52138_new_n5142_), .B(u2__abc_52138_new_n10341_), .C(u2__abc_52138_new_n5918_), .Y(u2__abc_52138_new_n10351_));
OAI21X1 OAI21X1_2321 ( .A(u2__abc_52138_new_n5144_), .B(u2__abc_52138_new_n10350_), .C(u2__abc_52138_new_n10352_), .Y(u2__abc_52138_new_n10353_));
OAI21X1 OAI21X1_2322 ( .A(u2__abc_52138_new_n5172_), .B(u2__abc_52138_new_n10355_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10358_));
OAI21X1 OAI21X1_2323 ( .A(u2__abc_52138_new_n5168_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10360_));
OAI21X1 OAI21X1_2324 ( .A(u2__abc_52138_new_n10360_), .B(u2__abc_52138_new_n10359_), .C(u2__abc_52138_new_n10361_), .Y(u2__abc_52138_new_n10362_));
OAI21X1 OAI21X1_2325 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_357_), .Y(u2__abc_52138_new_n10364_));
OAI21X1 OAI21X1_2326 ( .A(u2__abc_52138_new_n5171_), .B(u2__abc_52138_new_n10354_), .C(u2__abc_52138_new_n10365_), .Y(u2__abc_52138_new_n10366_));
OAI21X1 OAI21X1_2327 ( .A(u2__abc_52138_new_n5173_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10369_));
OAI21X1 OAI21X1_2328 ( .A(u2__abc_52138_new_n10369_), .B(u2__abc_52138_new_n10368_), .C(u2__abc_52138_new_n10370_), .Y(u2__abc_52138_new_n10371_));
OAI21X1 OAI21X1_2329 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_358_), .Y(u2__abc_52138_new_n10373_));
OAI21X1 OAI21X1_233 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1463_), .C(_abc_65734_new_n1477_), .Y(\o[229] ));
OAI21X1 OAI21X1_2330 ( .A(u2__abc_52138_new_n5173_), .B(u2_o_355_), .C(u2__abc_52138_new_n10365_), .Y(u2__abc_52138_new_n10374_));
OAI21X1 OAI21X1_2331 ( .A(u2__abc_52138_new_n10374_), .B(u2__abc_52138_new_n10357_), .C(u2__abc_52138_new_n10375_), .Y(u2__abc_52138_new_n10376_));
OAI21X1 OAI21X1_2332 ( .A(u2__abc_52138_new_n5161_), .B(u2__abc_52138_new_n10377_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10378_));
OAI21X1 OAI21X1_2333 ( .A(u2__abc_52138_new_n5157_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10380_));
OAI21X1 OAI21X1_2334 ( .A(u2__abc_52138_new_n10380_), .B(u2__abc_52138_new_n10379_), .C(u2__abc_52138_new_n10381_), .Y(u2__abc_52138_new_n10382_));
OAI21X1 OAI21X1_2335 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_359_), .Y(u2__abc_52138_new_n10384_));
OAI21X1 OAI21X1_2336 ( .A(u2__abc_52138_new_n5160_), .B(u2__abc_52138_new_n10376_), .C(u2__abc_52138_new_n10385_), .Y(u2__abc_52138_new_n10386_));
OAI21X1 OAI21X1_2337 ( .A(u2__abc_52138_new_n5166_), .B(u2__abc_52138_new_n10386_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10387_));
OAI21X1 OAI21X1_2338 ( .A(u2__abc_52138_new_n5162_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10389_));
OAI21X1 OAI21X1_2339 ( .A(u2__abc_52138_new_n10389_), .B(u2__abc_52138_new_n10388_), .C(u2__abc_52138_new_n10390_), .Y(u2__abc_52138_new_n10391_));
OAI21X1 OAI21X1_234 ( .A(_abc_65734_new_n1480_), .B(_abc_65734_new_n1482_), .C(_abc_65734_new_n1475_), .Y(_abc_65734_new_n1483_));
OAI21X1 OAI21X1_2340 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_360_), .Y(u2__abc_52138_new_n10393_));
OAI21X1 OAI21X1_2341 ( .A(u2_remHi_355_), .B(u2__abc_52138_new_n5175_), .C(u2__abc_52138_new_n10374_), .Y(u2__abc_52138_new_n10394_));
OAI21X1 OAI21X1_2342 ( .A(u2__abc_52138_new_n5167_), .B(u2__abc_52138_new_n10394_), .C(u2__abc_52138_new_n10395_), .Y(u2__abc_52138_new_n10396_));
OAI21X1 OAI21X1_2343 ( .A(u2__abc_52138_new_n5095_), .B(u2__abc_52138_new_n10401_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10402_));
OAI21X1 OAI21X1_2344 ( .A(u2__abc_52138_new_n5093_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10404_));
OAI21X1 OAI21X1_2345 ( .A(u2__abc_52138_new_n10404_), .B(u2__abc_52138_new_n10403_), .C(u2__abc_52138_new_n10405_), .Y(u2__abc_52138_new_n10406_));
OAI21X1 OAI21X1_2346 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_361_), .Y(u2__abc_52138_new_n10408_));
OAI21X1 OAI21X1_2347 ( .A(u2__abc_52138_new_n10398_), .B(u2__abc_52138_new_n10399_), .C(u2__abc_52138_new_n5095_), .Y(u2__abc_52138_new_n10409_));
OAI21X1 OAI21X1_2348 ( .A(u2__abc_52138_new_n5093_), .B(u2_o_358_), .C(u2__abc_52138_new_n10409_), .Y(u2__abc_52138_new_n10410_));
OAI21X1 OAI21X1_2349 ( .A(u2__abc_52138_new_n5100_), .B(u2__abc_52138_new_n10410_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10411_));
OAI21X1 OAI21X1_235 ( .A(_abc_65734_new_n1473_), .B(_abc_65734_new_n1471_), .C(_abc_65734_new_n1481_), .Y(_abc_65734_new_n1485_));
OAI21X1 OAI21X1_2350 ( .A(u2__abc_52138_new_n5096_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10413_));
OAI21X1 OAI21X1_2351 ( .A(u2__abc_52138_new_n10413_), .B(u2__abc_52138_new_n10412_), .C(u2__abc_52138_new_n10414_), .Y(u2__abc_52138_new_n10415_));
OAI21X1 OAI21X1_2352 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_362_), .Y(u2__abc_52138_new_n10417_));
OAI21X1 OAI21X1_2353 ( .A(u2__abc_52138_new_n5096_), .B(u2_o_359_), .C(u2__abc_52138_new_n10418_), .Y(u2__abc_52138_new_n10419_));
OAI21X1 OAI21X1_2354 ( .A(u2__abc_52138_new_n5101_), .B(u2__abc_52138_new_n10400_), .C(u2__abc_52138_new_n10420_), .Y(u2__abc_52138_new_n10421_));
OAI21X1 OAI21X1_2355 ( .A(u2__abc_52138_new_n5106_), .B(u2__abc_52138_new_n10421_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10422_));
OAI21X1 OAI21X1_2356 ( .A(u2__abc_52138_new_n5102_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10424_));
OAI21X1 OAI21X1_2357 ( .A(u2__abc_52138_new_n10424_), .B(u2__abc_52138_new_n10423_), .C(u2__abc_52138_new_n10426_), .Y(u2__abc_52138_new_n10427_));
OAI21X1 OAI21X1_2358 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_363_), .Y(u2__abc_52138_new_n10429_));
OAI21X1 OAI21X1_2359 ( .A(u2__abc_52138_new_n5102_), .B(u2_o_360_), .C(u2__abc_52138_new_n10430_), .Y(u2__abc_52138_new_n10431_));
OAI21X1 OAI21X1_236 ( .A(_abc_65734_new_n1489_), .B(_abc_65734_new_n1484_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1490_));
OAI21X1 OAI21X1_2360 ( .A(u2__abc_52138_new_n5111_), .B(u2__abc_52138_new_n10431_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10432_));
OAI21X1 OAI21X1_2361 ( .A(u2__abc_52138_new_n5109_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10434_));
OAI21X1 OAI21X1_2362 ( .A(u2__abc_52138_new_n10434_), .B(u2__abc_52138_new_n10433_), .C(u2__abc_52138_new_n10435_), .Y(u2__abc_52138_new_n10436_));
OAI21X1 OAI21X1_2363 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_364_), .Y(u2__abc_52138_new_n10438_));
OAI21X1 OAI21X1_2364 ( .A(u2_remHi_361_), .B(u2__abc_52138_new_n5107_), .C(u2__abc_52138_new_n5103_), .Y(u2__abc_52138_new_n10440_));
OAI21X1 OAI21X1_2365 ( .A(u2__abc_52138_new_n5109_), .B(u2_o_361_), .C(u2__abc_52138_new_n10440_), .Y(u2__abc_52138_new_n10441_));
OAI21X1 OAI21X1_2366 ( .A(u2__abc_52138_new_n5113_), .B(u2__abc_52138_new_n10400_), .C(u2__abc_52138_new_n10442_), .Y(u2__abc_52138_new_n10443_));
OAI21X1 OAI21X1_2367 ( .A(u2__abc_52138_new_n5125_), .B(u2__abc_52138_new_n10443_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10446_));
OAI21X1 OAI21X1_2368 ( .A(u2__abc_52138_new_n10425_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10448_));
OAI21X1 OAI21X1_2369 ( .A(u2__abc_52138_new_n10448_), .B(u2__abc_52138_new_n10447_), .C(u2__abc_52138_new_n10449_), .Y(u2__abc_52138_new_n10450_));
OAI21X1 OAI21X1_237 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1473_), .C(_abc_65734_new_n1490_), .Y(\o[230] ));
OAI21X1 OAI21X1_2370 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_365_), .Y(u2__abc_52138_new_n10452_));
OAI21X1 OAI21X1_2371 ( .A(u2__abc_52138_new_n10425_), .B(u2_o_362_), .C(u2__abc_52138_new_n10444_), .Y(u2__abc_52138_new_n10453_));
OAI21X1 OAI21X1_2372 ( .A(u2__abc_52138_new_n5126_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10456_));
OAI21X1 OAI21X1_2373 ( .A(u2__abc_52138_new_n10456_), .B(u2__abc_52138_new_n10455_), .C(u2__abc_52138_new_n10457_), .Y(u2__abc_52138_new_n10458_));
OAI21X1 OAI21X1_2374 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_366_), .Y(u2__abc_52138_new_n10460_));
OAI21X1 OAI21X1_2375 ( .A(u2__abc_52138_new_n10425_), .B(u2_o_362_), .C(u2__abc_52138_new_n5910_), .Y(u2__abc_52138_new_n10461_));
OAI21X1 OAI21X1_2376 ( .A(u2__abc_52138_new_n10461_), .B(u2__abc_52138_new_n10445_), .C(u2__abc_52138_new_n5912_), .Y(u2__abc_52138_new_n10462_));
OAI21X1 OAI21X1_2377 ( .A(u2__abc_52138_new_n5118_), .B(u2__abc_52138_new_n10463_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10464_));
OAI21X1 OAI21X1_2378 ( .A(u2__abc_52138_new_n5114_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10466_));
OAI21X1 OAI21X1_2379 ( .A(u2__abc_52138_new_n10466_), .B(u2__abc_52138_new_n10465_), .C(u2__abc_52138_new_n10467_), .Y(u2__abc_52138_new_n10468_));
OAI21X1 OAI21X1_238 ( .A(_abc_65734_new_n1481_), .B(_abc_65734_new_n1472_), .C(_abc_65734_new_n1493_), .Y(_abc_65734_new_n1494_));
OAI21X1 OAI21X1_2380 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_367_), .Y(u2__abc_52138_new_n10470_));
OAI21X1 OAI21X1_2381 ( .A(u2__abc_52138_new_n5117_), .B(u2__abc_52138_new_n10462_), .C(u2__abc_52138_new_n10471_), .Y(u2__abc_52138_new_n10472_));
OAI21X1 OAI21X1_2382 ( .A(u2__abc_52138_new_n5123_), .B(u2__abc_52138_new_n10472_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10473_));
OAI21X1 OAI21X1_2383 ( .A(u2__abc_52138_new_n5119_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10475_));
OAI21X1 OAI21X1_2384 ( .A(u2__abc_52138_new_n10475_), .B(u2__abc_52138_new_n10474_), .C(u2__abc_52138_new_n10476_), .Y(u2__abc_52138_new_n10477_));
OAI21X1 OAI21X1_2385 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_368_), .Y(u2__abc_52138_new_n10479_));
OAI21X1 OAI21X1_2386 ( .A(u2__abc_52138_new_n10471_), .B(u2__abc_52138_new_n5122_), .C(u2__abc_52138_new_n10480_), .Y(u2__abc_52138_new_n10481_));
OAI21X1 OAI21X1_2387 ( .A(u2__abc_52138_new_n5132_), .B(u2__abc_52138_new_n10442_), .C(u2__abc_52138_new_n5915_), .Y(u2__abc_52138_new_n10482_));
OAI21X1 OAI21X1_2388 ( .A(u2__abc_52138_new_n5133_), .B(u2__abc_52138_new_n10397_), .C(u2__abc_52138_new_n10483_), .Y(u2__abc_52138_new_n10484_));
OAI21X1 OAI21X1_2389 ( .A(u2__abc_52138_new_n10484_), .B(u2__abc_52138_new_n10485_), .C(u2__abc_52138_new_n5056_), .Y(u2__abc_52138_new_n10486_));
OAI21X1 OAI21X1_239 ( .A(_abc_65734_new_n1495_), .B(_abc_65734_new_n1497_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1498_));
OAI21X1 OAI21X1_2390 ( .A(u2__abc_52138_new_n5056_), .B(u2__abc_52138_new_n10489_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10490_));
OAI21X1 OAI21X1_2391 ( .A(u2__abc_52138_new_n5052_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10492_));
OAI21X1 OAI21X1_2392 ( .A(u2__abc_52138_new_n10492_), .B(u2__abc_52138_new_n10491_), .C(u2__abc_52138_new_n10493_), .Y(u2__abc_52138_new_n10494_));
OAI21X1 OAI21X1_2393 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_369_), .Y(u2__abc_52138_new_n10496_));
OAI21X1 OAI21X1_2394 ( .A(u2__abc_52138_new_n5052_), .B(u2_o_366_), .C(u2__abc_52138_new_n10486_), .Y(u2__abc_52138_new_n10497_));
OAI21X1 OAI21X1_2395 ( .A(u2__abc_52138_new_n5059_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10500_));
OAI21X1 OAI21X1_2396 ( .A(u2__abc_52138_new_n10500_), .B(u2__abc_52138_new_n10499_), .C(u2__abc_52138_new_n10501_), .Y(u2__abc_52138_new_n10502_));
OAI21X1 OAI21X1_2397 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_370_), .Y(u2__abc_52138_new_n10504_));
OAI21X1 OAI21X1_2398 ( .A(u2__abc_52138_new_n5052_), .B(u2_o_366_), .C(u2__abc_52138_new_n5058_), .Y(u2__abc_52138_new_n10505_));
OAI21X1 OAI21X1_2399 ( .A(u2__abc_52138_new_n10505_), .B(u2__abc_52138_new_n10487_), .C(u2__abc_52138_new_n5060_), .Y(u2__abc_52138_new_n10506_));
OAI21X1 OAI21X1_24 ( .A(aNan), .B(_abc_65734_new_n899_), .C(_abc_65734_new_n900_), .Y(\o[135] ));
OAI21X1 OAI21X1_240 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1481_), .C(_abc_65734_new_n1498_), .Y(\o[231] ));
OAI21X1 OAI21X1_2400 ( .A(u2__abc_52138_new_n5049_), .B(u2__abc_52138_new_n10507_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10508_));
OAI21X1 OAI21X1_2401 ( .A(u2__abc_52138_new_n5045_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10510_));
OAI21X1 OAI21X1_2402 ( .A(u2__abc_52138_new_n10510_), .B(u2__abc_52138_new_n10509_), .C(u2__abc_52138_new_n10511_), .Y(u2__abc_52138_new_n10512_));
OAI21X1 OAI21X1_2403 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_371_), .Y(u2__abc_52138_new_n10514_));
OAI21X1 OAI21X1_2404 ( .A(u2__abc_52138_new_n5048_), .B(u2__abc_52138_new_n10506_), .C(u2__abc_52138_new_n10515_), .Y(u2__abc_52138_new_n10516_));
OAI21X1 OAI21X1_2405 ( .A(u2__abc_52138_new_n5050_), .B(u2__abc_52138_new_n10516_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10517_));
OAI21X1 OAI21X1_2406 ( .A(u2__abc_52138_new_n5886_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10519_));
OAI21X1 OAI21X1_2407 ( .A(u2__abc_52138_new_n10519_), .B(u2__abc_52138_new_n10518_), .C(u2__abc_52138_new_n10520_), .Y(u2__abc_52138_new_n10521_));
OAI21X1 OAI21X1_2408 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_372_), .Y(u2__abc_52138_new_n10523_));
OAI21X1 OAI21X1_2409 ( .A(u2__abc_52138_new_n5886_), .B(u2_o_369_), .C(u2__abc_52138_new_n10515_), .Y(u2__abc_52138_new_n10524_));
OAI21X1 OAI21X1_241 ( .A(_abc_65734_new_n1493_), .B(_abc_65734_new_n1487_), .C(_abc_65734_new_n1500_), .Y(_abc_65734_new_n1501_));
OAI21X1 OAI21X1_2410 ( .A(u2__abc_52138_new_n10484_), .B(u2__abc_52138_new_n10485_), .C(u2__abc_52138_new_n5064_), .Y(u2__abc_52138_new_n10527_));
OAI21X1 OAI21X1_2411 ( .A(u2__abc_52138_new_n5086_), .B(u2__abc_52138_new_n10528_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10529_));
OAI21X1 OAI21X1_2412 ( .A(u2__abc_52138_new_n5084_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10531_));
OAI21X1 OAI21X1_2413 ( .A(u2__abc_52138_new_n10531_), .B(u2__abc_52138_new_n10530_), .C(u2__abc_52138_new_n10532_), .Y(u2__abc_52138_new_n10533_));
OAI21X1 OAI21X1_2414 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_373_), .Y(u2__abc_52138_new_n10535_));
OAI21X1 OAI21X1_2415 ( .A(u2__abc_52138_new_n5084_), .B(u2_o_370_), .C(u2__abc_52138_new_n10536_), .Y(u2__abc_52138_new_n10537_));
OAI21X1 OAI21X1_2416 ( .A(u2__abc_52138_new_n5081_), .B(u2__abc_52138_new_n10537_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10538_));
OAI21X1 OAI21X1_2417 ( .A(u2__abc_52138_new_n5078_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10540_));
OAI21X1 OAI21X1_2418 ( .A(u2__abc_52138_new_n10540_), .B(u2__abc_52138_new_n10539_), .C(u2__abc_52138_new_n10541_), .Y(u2__abc_52138_new_n10542_));
OAI21X1 OAI21X1_2419 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_374_), .Y(u2__abc_52138_new_n10544_));
OAI21X1 OAI21X1_242 ( .A(_abc_65734_new_n1507_), .B(_abc_65734_new_n1504_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1508_));
OAI21X1 OAI21X1_2420 ( .A(u2__abc_52138_new_n5080_), .B(u2__abc_52138_new_n10545_), .C(u2__abc_52138_new_n5077_), .Y(u2__abc_52138_new_n10546_));
OAI21X1 OAI21X1_2421 ( .A(u2__abc_52138_new_n5069_), .B(u2__abc_52138_new_n10546_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10547_));
OAI21X1 OAI21X1_2422 ( .A(u2__abc_52138_new_n5065_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10549_));
OAI21X1 OAI21X1_2423 ( .A(u2__abc_52138_new_n10549_), .B(u2__abc_52138_new_n10548_), .C(u2__abc_52138_new_n10550_), .Y(u2__abc_52138_new_n10551_));
OAI21X1 OAI21X1_2424 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_375_), .Y(u2__abc_52138_new_n10553_));
OAI21X1 OAI21X1_2425 ( .A(u2__abc_52138_new_n5065_), .B(u2_o_372_), .C(u2__abc_52138_new_n10554_), .Y(u2__abc_52138_new_n10555_));
OAI21X1 OAI21X1_2426 ( .A(u2__abc_52138_new_n5074_), .B(u2__abc_52138_new_n10555_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10556_));
OAI21X1 OAI21X1_2427 ( .A(u2__abc_52138_new_n5070_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10558_));
OAI21X1 OAI21X1_2428 ( .A(u2__abc_52138_new_n10558_), .B(u2__abc_52138_new_n10557_), .C(u2__abc_52138_new_n10559_), .Y(u2__abc_52138_new_n10560_));
OAI21X1 OAI21X1_2429 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_376_), .Y(u2__abc_52138_new_n10562_));
OAI21X1 OAI21X1_243 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1493_), .C(_abc_65734_new_n1508_), .Y(\o[232] ));
OAI21X1 OAI21X1_2430 ( .A(u2__abc_52138_new_n5083_), .B(u2__abc_52138_new_n5080_), .C(u2__abc_52138_new_n5077_), .Y(u2__abc_52138_new_n10563_));
OAI21X1 OAI21X1_2431 ( .A(u2__abc_52138_new_n10564_), .B(u2__abc_52138_new_n10526_), .C(u2__abc_52138_new_n10565_), .Y(u2__abc_52138_new_n10566_));
OAI21X1 OAI21X1_2432 ( .A(u2__abc_52138_new_n5089_), .B(u2__abc_52138_new_n10488_), .C(u2__abc_52138_new_n10567_), .Y(u2__abc_52138_new_n10568_));
OAI21X1 OAI21X1_2433 ( .A(u2__abc_52138_new_n5022_), .B(u2__abc_52138_new_n10568_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10569_));
OAI21X1 OAI21X1_2434 ( .A(u2__abc_52138_new_n5020_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10571_));
OAI21X1 OAI21X1_2435 ( .A(u2__abc_52138_new_n10571_), .B(u2__abc_52138_new_n10570_), .C(u2__abc_52138_new_n10572_), .Y(u2__abc_52138_new_n10573_));
OAI21X1 OAI21X1_2436 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_377_), .Y(u2__abc_52138_new_n10575_));
OAI21X1 OAI21X1_2437 ( .A(u2__abc_52138_new_n5020_), .B(u2_o_374_), .C(u2__abc_52138_new_n10576_), .Y(u2__abc_52138_new_n10577_));
OAI21X1 OAI21X1_2438 ( .A(u2__abc_52138_new_n5028_), .B(u2__abc_52138_new_n10577_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10578_));
OAI21X1 OAI21X1_2439 ( .A(u2__abc_52138_new_n5023_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10580_));
OAI21X1 OAI21X1_244 ( .A(_abc_65734_new_n1500_), .B(_abc_65734_new_n1492_), .C(\a[120] ), .Y(_abc_65734_new_n1513_));
OAI21X1 OAI21X1_2440 ( .A(u2__abc_52138_new_n10580_), .B(u2__abc_52138_new_n10579_), .C(u2__abc_52138_new_n10581_), .Y(u2__abc_52138_new_n10582_));
OAI21X1 OAI21X1_2441 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_378_), .Y(u2__abc_52138_new_n10584_));
OAI21X1 OAI21X1_2442 ( .A(u2__abc_52138_new_n5027_), .B(u2__abc_52138_new_n10586_), .C(u2__abc_52138_new_n5026_), .Y(u2__abc_52138_new_n10587_));
OAI21X1 OAI21X1_2443 ( .A(u2__abc_52138_new_n5030_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10592_));
OAI21X1 OAI21X1_2444 ( .A(u2__abc_52138_new_n10592_), .B(u2__abc_52138_new_n10591_), .C(u2__abc_52138_new_n10594_), .Y(u2__abc_52138_new_n10595_));
OAI21X1 OAI21X1_2445 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_379_), .Y(u2__abc_52138_new_n10597_));
OAI21X1 OAI21X1_2446 ( .A(u2__abc_52138_new_n5030_), .B(u2_o_376_), .C(u2__abc_52138_new_n10589_), .Y(u2__abc_52138_new_n10599_));
OAI21X1 OAI21X1_2447 ( .A(u2__abc_52138_new_n10598_), .B(u2__abc_52138_new_n10599_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10600_));
OAI21X1 OAI21X1_2448 ( .A(u2__abc_52138_new_n5035_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10602_));
OAI21X1 OAI21X1_2449 ( .A(u2__abc_52138_new_n10602_), .B(u2__abc_52138_new_n10601_), .C(u2__abc_52138_new_n10603_), .Y(u2__abc_52138_new_n10604_));
OAI21X1 OAI21X1_245 ( .A(_abc_65734_new_n1500_), .B(_abc_65734_new_n1492_), .C(_abc_65734_new_n1510_), .Y(_abc_65734_new_n1517_));
OAI21X1 OAI21X1_2450 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_380_), .Y(u2__abc_52138_new_n10606_));
OAI21X1 OAI21X1_2451 ( .A(u2__abc_52138_new_n5042_), .B(u2__abc_52138_new_n10588_), .C(u2__abc_52138_new_n10607_), .Y(u2__abc_52138_new_n10608_));
OAI21X1 OAI21X1_2452 ( .A(u2__abc_52138_new_n5010_), .B(u2__abc_52138_new_n10608_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10611_));
OAI21X1 OAI21X1_2453 ( .A(u2__abc_52138_new_n10593_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10613_));
OAI21X1 OAI21X1_2454 ( .A(u2__abc_52138_new_n10613_), .B(u2__abc_52138_new_n10612_), .C(u2__abc_52138_new_n10614_), .Y(u2__abc_52138_new_n10615_));
OAI21X1 OAI21X1_2455 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_381_), .Y(u2__abc_52138_new_n10617_));
OAI21X1 OAI21X1_2456 ( .A(u2__abc_52138_new_n10593_), .B(u2_o_378_), .C(u2__abc_52138_new_n10609_), .Y(u2__abc_52138_new_n10618_));
OAI21X1 OAI21X1_2457 ( .A(u2__abc_52138_new_n5011_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10621_));
OAI21X1 OAI21X1_2458 ( .A(u2__abc_52138_new_n10621_), .B(u2__abc_52138_new_n10620_), .C(u2__abc_52138_new_n10622_), .Y(u2__abc_52138_new_n10623_));
OAI21X1 OAI21X1_2459 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_382_), .Y(u2__abc_52138_new_n10625_));
OAI21X1 OAI21X1_246 ( .A(_abc_65734_new_n1515_), .B(_abc_65734_new_n1519_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1520_));
OAI21X1 OAI21X1_2460 ( .A(u2__abc_52138_new_n10593_), .B(u2_o_378_), .C(u2__abc_52138_new_n10626_), .Y(u2__abc_52138_new_n10627_));
OAI21X1 OAI21X1_2461 ( .A(u2__abc_52138_new_n10627_), .B(u2__abc_52138_new_n10610_), .C(u2__abc_52138_new_n5934_), .Y(u2__abc_52138_new_n10628_));
OAI21X1 OAI21X1_2462 ( .A(u2__abc_52138_new_n5003_), .B(u2__abc_52138_new_n10629_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10630_));
OAI21X1 OAI21X1_2463 ( .A(u2__abc_52138_new_n4999_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10632_));
OAI21X1 OAI21X1_2464 ( .A(u2__abc_52138_new_n10632_), .B(u2__abc_52138_new_n10631_), .C(u2__abc_52138_new_n10633_), .Y(u2__abc_52138_new_n10634_));
OAI21X1 OAI21X1_2465 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_383_), .Y(u2__abc_52138_new_n10636_));
OAI21X1 OAI21X1_2466 ( .A(u2__abc_52138_new_n5002_), .B(u2__abc_52138_new_n10628_), .C(u2__abc_52138_new_n10637_), .Y(u2__abc_52138_new_n10638_));
OAI21X1 OAI21X1_2467 ( .A(u2__abc_52138_new_n5008_), .B(u2__abc_52138_new_n10638_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10639_));
OAI21X1 OAI21X1_2468 ( .A(u2__abc_52138_new_n5006_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10641_));
OAI21X1 OAI21X1_2469 ( .A(u2__abc_52138_new_n10641_), .B(u2__abc_52138_new_n10640_), .C(u2__abc_52138_new_n10642_), .Y(u2__abc_52138_new_n10643_));
OAI21X1 OAI21X1_247 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1500_), .C(_abc_65734_new_n1520_), .Y(\o[233] ));
OAI21X1 OAI21X1_2470 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_384_), .Y(u2__abc_52138_new_n10645_));
OAI21X1 OAI21X1_2471 ( .A(u2__abc_52138_new_n10305_), .B(u2__abc_52138_new_n10310_), .C(u2__abc_52138_new_n5182_), .Y(u2__abc_52138_new_n10650_));
OAI21X1 OAI21X1_2472 ( .A(u2__abc_52138_new_n10651_), .B(u2__abc_52138_new_n5042_), .C(u2__abc_52138_new_n10607_), .Y(u2__abc_52138_new_n10652_));
OAI21X1 OAI21X1_2473 ( .A(u2_remHi_379_), .B(u2__abc_52138_new_n5013_), .C(u2__abc_52138_new_n10627_), .Y(u2__abc_52138_new_n10653_));
OAI21X1 OAI21X1_2474 ( .A(u2__abc_52138_new_n5009_), .B(u2__abc_52138_new_n10653_), .C(u2__abc_52138_new_n10654_), .Y(u2__abc_52138_new_n10655_));
OAI21X1 OAI21X1_2475 ( .A(u2__abc_52138_new_n5044_), .B(u2__abc_52138_new_n10567_), .C(u2__abc_52138_new_n10656_), .Y(u2__abc_52138_new_n10657_));
OAI21X1 OAI21X1_2476 ( .A(u2__abc_52138_new_n10659_), .B(u2__abc_52138_new_n10647_), .C(u2__abc_52138_new_n6180_), .Y(u2__abc_52138_new_n10660_));
OAI21X1 OAI21X1_2477 ( .A(u2__abc_52138_new_n6180_), .B(u2__abc_52138_new_n10663_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10664_));
OAI21X1 OAI21X1_2478 ( .A(u2__abc_52138_new_n6176_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10666_));
OAI21X1 OAI21X1_2479 ( .A(u2__abc_52138_new_n10666_), .B(u2__abc_52138_new_n10665_), .C(u2__abc_52138_new_n10667_), .Y(u2__abc_52138_new_n10668_));
OAI21X1 OAI21X1_248 ( .A(_abc_65734_new_n1510_), .B(_abc_65734_new_n1502_), .C(\a[121] ), .Y(_abc_65734_new_n1526_));
OAI21X1 OAI21X1_2480 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_385_), .Y(u2__abc_52138_new_n10670_));
OAI21X1 OAI21X1_2481 ( .A(u2_o_382_), .B(u2__abc_52138_new_n6176_), .C(u2__abc_52138_new_n10660_), .Y(u2__abc_52138_new_n10671_));
OAI21X1 OAI21X1_2482 ( .A(u2__abc_52138_new_n6175_), .B(u2__abc_52138_new_n10671_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10672_));
OAI21X1 OAI21X1_2483 ( .A(u2__abc_52138_new_n6173_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10674_));
OAI21X1 OAI21X1_2484 ( .A(u2__abc_52138_new_n10674_), .B(u2__abc_52138_new_n10673_), .C(u2__abc_52138_new_n10675_), .Y(u2__abc_52138_new_n10676_));
OAI21X1 OAI21X1_2485 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_386_), .Y(u2__abc_52138_new_n10678_));
OAI21X1 OAI21X1_2486 ( .A(u2_o_382_), .B(u2__abc_52138_new_n6176_), .C(u2__abc_52138_new_n6334_), .Y(u2__abc_52138_new_n10680_));
OAI21X1 OAI21X1_2487 ( .A(u2__abc_52138_new_n10680_), .B(u2__abc_52138_new_n10661_), .C(u2__abc_52138_new_n10679_), .Y(u2__abc_52138_new_n10681_));
OAI21X1 OAI21X1_2488 ( .A(u2__abc_52138_new_n6164_), .B(u2__abc_52138_new_n10682_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10683_));
OAI21X1 OAI21X1_2489 ( .A(u2__abc_52138_new_n6160_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10685_));
OAI21X1 OAI21X1_249 ( .A(_abc_65734_new_n1528_), .B(_abc_65734_new_n1530_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1531_));
OAI21X1 OAI21X1_2490 ( .A(u2__abc_52138_new_n10685_), .B(u2__abc_52138_new_n10684_), .C(u2__abc_52138_new_n10686_), .Y(u2__abc_52138_new_n10687_));
OAI21X1 OAI21X1_2491 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_387_), .Y(u2__abc_52138_new_n10689_));
OAI21X1 OAI21X1_2492 ( .A(u2__abc_52138_new_n6163_), .B(u2__abc_52138_new_n10681_), .C(u2__abc_52138_new_n10690_), .Y(u2__abc_52138_new_n10691_));
OAI21X1 OAI21X1_2493 ( .A(u2__abc_52138_new_n6169_), .B(u2__abc_52138_new_n10691_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10692_));
OAI21X1 OAI21X1_2494 ( .A(u2__abc_52138_new_n6167_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10694_));
OAI21X1 OAI21X1_2495 ( .A(u2__abc_52138_new_n10694_), .B(u2__abc_52138_new_n10693_), .C(u2__abc_52138_new_n10695_), .Y(u2__abc_52138_new_n10696_));
OAI21X1 OAI21X1_2496 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_388_), .Y(u2__abc_52138_new_n10698_));
OAI21X1 OAI21X1_2497 ( .A(u2__abc_52138_new_n6171_), .B(u2_remHi_383_), .C(u2__abc_52138_new_n10680_), .Y(u2__abc_52138_new_n10699_));
OAI21X1 OAI21X1_2498 ( .A(u2__abc_52138_new_n6166_), .B(u2__abc_52138_new_n10690_), .C(u2__abc_52138_new_n6336_), .Y(u2__abc_52138_new_n10700_));
OAI21X1 OAI21X1_2499 ( .A(u2__abc_52138_new_n6170_), .B(u2__abc_52138_new_n10699_), .C(u2__abc_52138_new_n10701_), .Y(u2__abc_52138_new_n10702_));
OAI21X1 OAI21X1_25 ( .A(aNan), .B(_abc_65734_new_n902_), .C(_abc_65734_new_n903_), .Y(\o[136] ));
OAI21X1 OAI21X1_250 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1510_), .C(_abc_65734_new_n1531_), .Y(\o[234] ));
OAI21X1 OAI21X1_2500 ( .A(u2__abc_52138_new_n6183_), .B(u2__abc_52138_new_n10662_), .C(u2__abc_52138_new_n10703_), .Y(u2__abc_52138_new_n10704_));
OAI21X1 OAI21X1_2501 ( .A(u2__abc_52138_new_n6156_), .B(u2__abc_52138_new_n10704_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10707_));
OAI21X1 OAI21X1_2502 ( .A(u2__abc_52138_new_n6152_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10709_));
OAI21X1 OAI21X1_2503 ( .A(u2__abc_52138_new_n10709_), .B(u2__abc_52138_new_n10708_), .C(u2__abc_52138_new_n10710_), .Y(u2__abc_52138_new_n10711_));
OAI21X1 OAI21X1_2504 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_389_), .Y(u2__abc_52138_new_n10713_));
OAI21X1 OAI21X1_2505 ( .A(u2_o_386_), .B(u2__abc_52138_new_n6152_), .C(u2__abc_52138_new_n10705_), .Y(u2__abc_52138_new_n10714_));
OAI21X1 OAI21X1_2506 ( .A(u2__abc_52138_new_n6149_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10717_));
OAI21X1 OAI21X1_2507 ( .A(u2__abc_52138_new_n10717_), .B(u2__abc_52138_new_n10716_), .C(u2__abc_52138_new_n10718_), .Y(u2__abc_52138_new_n10719_));
OAI21X1 OAI21X1_2508 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_390_), .Y(u2__abc_52138_new_n10721_));
OAI21X1 OAI21X1_2509 ( .A(u2_o_386_), .B(u2__abc_52138_new_n6152_), .C(u2__abc_52138_new_n6339_), .Y(u2__abc_52138_new_n10724_));
OAI21X1 OAI21X1_251 ( .A(_abc_65734_new_n1534_), .B(_abc_65734_new_n1502_), .C(\a[122] ), .Y(_abc_65734_new_n1537_));
OAI21X1 OAI21X1_2510 ( .A(u2__abc_52138_new_n10724_), .B(u2__abc_52138_new_n10706_), .C(u2__abc_52138_new_n10723_), .Y(u2__abc_52138_new_n10725_));
OAI21X1 OAI21X1_2511 ( .A(u2__abc_52138_new_n6137_), .B(u2__abc_52138_new_n6139_), .C(u2__abc_52138_new_n10725_), .Y(u2__abc_52138_new_n10727_));
OAI21X1 OAI21X1_2512 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n10727_), .Y(u2__abc_52138_new_n10728_));
OAI21X1 OAI21X1_2513 ( .A(u2__abc_52138_new_n6136_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10730_));
OAI21X1 OAI21X1_2514 ( .A(u2__abc_52138_new_n10730_), .B(u2__abc_52138_new_n10729_), .C(u2__abc_52138_new_n10731_), .Y(u2__abc_52138_new_n10732_));
OAI21X1 OAI21X1_2515 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_391_), .Y(u2__abc_52138_new_n10734_));
OAI21X1 OAI21X1_2516 ( .A(u2__abc_52138_new_n6139_), .B(u2__abc_52138_new_n10725_), .C(u2__abc_52138_new_n10735_), .Y(u2__abc_52138_new_n10736_));
OAI21X1 OAI21X1_2517 ( .A(u2__abc_52138_new_n6145_), .B(u2__abc_52138_new_n10736_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10737_));
OAI21X1 OAI21X1_2518 ( .A(u2__abc_52138_new_n6141_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10739_));
OAI21X1 OAI21X1_2519 ( .A(u2__abc_52138_new_n10739_), .B(u2__abc_52138_new_n10738_), .C(u2__abc_52138_new_n10740_), .Y(u2__abc_52138_new_n10741_));
OAI21X1 OAI21X1_252 ( .A(_abc_65734_new_n1539_), .B(_abc_65734_new_n1541_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1542_));
OAI21X1 OAI21X1_2520 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_392_), .Y(u2__abc_52138_new_n10743_));
OAI21X1 OAI21X1_2521 ( .A(u2__abc_52138_new_n6144_), .B(u2__abc_52138_new_n10735_), .C(u2__abc_52138_new_n10745_), .Y(u2__abc_52138_new_n10746_));
OAI21X1 OAI21X1_2522 ( .A(u2__abc_52138_new_n6159_), .B(u2__abc_52138_new_n10703_), .C(u2__abc_52138_new_n10747_), .Y(u2__abc_52138_new_n10748_));
OAI21X1 OAI21X1_2523 ( .A(u2__abc_52138_new_n10659_), .B(u2__abc_52138_new_n10647_), .C(u2__abc_52138_new_n6184_), .Y(u2__abc_52138_new_n10750_));
OAI21X1 OAI21X1_2524 ( .A(u2__abc_52138_new_n6296_), .B(u2__abc_52138_new_n10751_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10752_));
OAI21X1 OAI21X1_2525 ( .A(u2__abc_52138_new_n6292_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10754_));
OAI21X1 OAI21X1_2526 ( .A(u2__abc_52138_new_n10754_), .B(u2__abc_52138_new_n10753_), .C(u2__abc_52138_new_n10755_), .Y(u2__abc_52138_new_n10756_));
OAI21X1 OAI21X1_2527 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_393_), .Y(u2__abc_52138_new_n10758_));
OAI21X1 OAI21X1_2528 ( .A(u2_o_390_), .B(u2__abc_52138_new_n6292_), .C(u2__abc_52138_new_n10759_), .Y(u2__abc_52138_new_n10760_));
OAI21X1 OAI21X1_2529 ( .A(u2__abc_52138_new_n6299_), .B(u2__abc_52138_new_n6300_), .C(u2__abc_52138_new_n10760_), .Y(u2__abc_52138_new_n10761_));
OAI21X1 OAI21X1_253 ( .A(_abc_65734_new_n753_), .B(_abc_65734_new_n1523_), .C(_abc_65734_new_n1542_), .Y(\o[235] ));
OAI21X1 OAI21X1_2530 ( .A(u2__abc_52138_new_n6297_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10765_));
OAI21X1 OAI21X1_2531 ( .A(u2__abc_52138_new_n10765_), .B(u2__abc_52138_new_n10764_), .C(u2__abc_52138_new_n10766_), .Y(u2__abc_52138_new_n10767_));
OAI21X1 OAI21X1_2532 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_394_), .Y(u2__abc_52138_new_n10769_));
OAI21X1 OAI21X1_2533 ( .A(u2__abc_52138_new_n6299_), .B(u2__abc_52138_new_n10762_), .C(u2__abc_52138_new_n6350_), .Y(u2__abc_52138_new_n10770_));
OAI21X1 OAI21X1_2534 ( .A(u2__abc_52138_new_n6284_), .B(u2__abc_52138_new_n10770_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10771_));
OAI21X1 OAI21X1_2535 ( .A(u2__abc_52138_new_n6280_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10773_));
OAI21X1 OAI21X1_2536 ( .A(u2__abc_52138_new_n10773_), .B(u2__abc_52138_new_n10772_), .C(u2__abc_52138_new_n10774_), .Y(u2__abc_52138_new_n10775_));
OAI21X1 OAI21X1_2537 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_395_), .Y(u2__abc_52138_new_n10777_));
OAI21X1 OAI21X1_2538 ( .A(u2__abc_52138_new_n6280_), .B(u2_o_392_), .C(u2__abc_52138_new_n10778_), .Y(u2__abc_52138_new_n10779_));
OAI21X1 OAI21X1_2539 ( .A(u2__abc_52138_new_n6290_), .B(u2__abc_52138_new_n10779_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10780_));
OAI21X1 OAI21X1_254 ( .A(_abc_65734_new_n1533_), .B(_abc_65734_new_n1546_), .C(_abc_65734_new_n1545_), .Y(_abc_65734_new_n1547_));
OAI21X1 OAI21X1_2540 ( .A(u2__abc_52138_new_n6352_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10782_));
OAI21X1 OAI21X1_2541 ( .A(u2__abc_52138_new_n10782_), .B(u2__abc_52138_new_n10781_), .C(u2__abc_52138_new_n10783_), .Y(u2__abc_52138_new_n10784_));
OAI21X1 OAI21X1_2542 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_396_), .Y(u2__abc_52138_new_n10786_));
OAI21X1 OAI21X1_2543 ( .A(u2__abc_52138_new_n6293_), .B(u2__abc_52138_new_n6300_), .C(u2__abc_52138_new_n6298_), .Y(u2__abc_52138_new_n10787_));
OAI21X1 OAI21X1_2544 ( .A(u2__abc_52138_new_n6286_), .B(u2__abc_52138_new_n10788_), .C(u2__abc_52138_new_n6288_), .Y(u2__abc_52138_new_n10789_));
OAI21X1 OAI21X1_2545 ( .A(u2__abc_52138_new_n10787_), .B(u2__abc_52138_new_n6291_), .C(u2__abc_52138_new_n10790_), .Y(u2__abc_52138_new_n10791_));
OAI21X1 OAI21X1_2546 ( .A(u2__abc_52138_new_n6324_), .B(u2__abc_52138_new_n10793_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10796_));
OAI21X1 OAI21X1_2547 ( .A(u2__abc_52138_new_n6320_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10798_));
OAI21X1 OAI21X1_2548 ( .A(u2__abc_52138_new_n10798_), .B(u2__abc_52138_new_n10797_), .C(u2__abc_52138_new_n10799_), .Y(u2__abc_52138_new_n10800_));
OAI21X1 OAI21X1_2549 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_397_), .Y(u2__abc_52138_new_n10802_));
OAI21X1 OAI21X1_255 ( .A(aNan), .B(_abc_65734_new_n1551_), .C(_abc_65734_new_n1552_), .Y(\o[236] ));
OAI21X1 OAI21X1_2550 ( .A(u2_o_394_), .B(u2__abc_52138_new_n6320_), .C(u2__abc_52138_new_n10794_), .Y(u2__abc_52138_new_n10803_));
OAI21X1 OAI21X1_2551 ( .A(u2__abc_52138_new_n6317_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10806_));
OAI21X1 OAI21X1_2552 ( .A(u2__abc_52138_new_n10806_), .B(u2__abc_52138_new_n10805_), .C(u2__abc_52138_new_n10807_), .Y(u2__abc_52138_new_n10808_));
OAI21X1 OAI21X1_2553 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_398_), .Y(u2__abc_52138_new_n10810_));
OAI21X1 OAI21X1_2554 ( .A(u2_o_395_), .B(u2__abc_52138_new_n6317_), .C(u2__abc_52138_new_n6322_), .Y(u2__abc_52138_new_n10811_));
OAI21X1 OAI21X1_2555 ( .A(u2__abc_52138_new_n10811_), .B(u2__abc_52138_new_n10795_), .C(u2__abc_52138_new_n6346_), .Y(u2__abc_52138_new_n10812_));
OAI21X1 OAI21X1_2556 ( .A(u2__abc_52138_new_n6308_), .B(u2__abc_52138_new_n10813_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10814_));
OAI21X1 OAI21X1_2557 ( .A(u2__abc_52138_new_n6304_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10816_));
OAI21X1 OAI21X1_2558 ( .A(u2__abc_52138_new_n10816_), .B(u2__abc_52138_new_n10815_), .C(u2__abc_52138_new_n10817_), .Y(u2__abc_52138_new_n10818_));
OAI21X1 OAI21X1_2559 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_399_), .Y(u2__abc_52138_new_n10820_));
OAI21X1 OAI21X1_256 ( .A(_abc_65734_new_n1558_), .B(_abc_65734_new_n1544_), .C(_abc_65734_new_n1559_), .Y(_abc_65734_new_n1560_));
OAI21X1 OAI21X1_2560 ( .A(u2__abc_52138_new_n6307_), .B(u2__abc_52138_new_n10812_), .C(u2__abc_52138_new_n10821_), .Y(u2__abc_52138_new_n10822_));
OAI21X1 OAI21X1_2561 ( .A(u2__abc_52138_new_n6313_), .B(u2__abc_52138_new_n10822_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10823_));
OAI21X1 OAI21X1_2562 ( .A(u2__abc_52138_new_n6309_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10825_));
OAI21X1 OAI21X1_2563 ( .A(u2__abc_52138_new_n10825_), .B(u2__abc_52138_new_n10824_), .C(u2__abc_52138_new_n10826_), .Y(u2__abc_52138_new_n10827_));
OAI21X1 OAI21X1_2564 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_400_), .Y(u2__abc_52138_new_n10829_));
OAI21X1 OAI21X1_2565 ( .A(u2_remHi_397_), .B(u2__abc_52138_new_n6311_), .C(u2__abc_52138_new_n6305_), .Y(u2__abc_52138_new_n10831_));
OAI21X1 OAI21X1_2566 ( .A(u2__abc_52138_new_n6236_), .B(u2__abc_52138_new_n10836_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10837_));
OAI21X1 OAI21X1_2567 ( .A(u2__abc_52138_new_n6232_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10839_));
OAI21X1 OAI21X1_2568 ( .A(u2__abc_52138_new_n10839_), .B(u2__abc_52138_new_n10838_), .C(u2__abc_52138_new_n10840_), .Y(u2__abc_52138_new_n10841_));
OAI21X1 OAI21X1_2569 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_401_), .Y(u2__abc_52138_new_n10843_));
OAI21X1 OAI21X1_257 ( .A(aNan), .B(_abc_65734_new_n1561_), .C(_abc_65734_new_n1554_), .Y(\o[237] ));
OAI21X1 OAI21X1_2570 ( .A(u2__abc_52138_new_n6235_), .B(u2__abc_52138_new_n10835_), .C(u2__abc_52138_new_n10844_), .Y(u2__abc_52138_new_n10845_));
OAI21X1 OAI21X1_2571 ( .A(u2__abc_52138_new_n6241_), .B(u2__abc_52138_new_n10845_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10846_));
OAI21X1 OAI21X1_2572 ( .A(u2__abc_52138_new_n6239_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10848_));
OAI21X1 OAI21X1_2573 ( .A(u2__abc_52138_new_n10848_), .B(u2__abc_52138_new_n10847_), .C(u2__abc_52138_new_n10849_), .Y(u2__abc_52138_new_n10850_));
OAI21X1 OAI21X1_2574 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_402_), .Y(u2__abc_52138_new_n10852_));
OAI21X1 OAI21X1_2575 ( .A(u2__abc_52138_new_n6238_), .B(u2__abc_52138_new_n10844_), .C(u2__abc_52138_new_n6373_), .Y(u2__abc_52138_new_n10853_));
OAI21X1 OAI21X1_2576 ( .A(u2__abc_52138_new_n6242_), .B(u2__abc_52138_new_n10835_), .C(u2__abc_52138_new_n10854_), .Y(u2__abc_52138_new_n10855_));
OAI21X1 OAI21X1_2577 ( .A(u2__abc_52138_new_n6247_), .B(u2__abc_52138_new_n10855_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10856_));
OAI21X1 OAI21X1_2578 ( .A(u2__abc_52138_new_n6243_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10858_));
OAI21X1 OAI21X1_2579 ( .A(u2__abc_52138_new_n10858_), .B(u2__abc_52138_new_n10857_), .C(u2__abc_52138_new_n10859_), .Y(u2__abc_52138_new_n10860_));
OAI21X1 OAI21X1_258 ( .A(_abc_65734_new_n1555_), .B(_abc_65734_new_n1549_), .C(_abc_65734_new_n1563_), .Y(_abc_65734_new_n1564_));
OAI21X1 OAI21X1_2580 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_403_), .Y(u2__abc_52138_new_n10862_));
OAI21X1 OAI21X1_2581 ( .A(u2__abc_52138_new_n6243_), .B(u2_o_400_), .C(u2__abc_52138_new_n10863_), .Y(u2__abc_52138_new_n10864_));
OAI21X1 OAI21X1_2582 ( .A(u2__abc_52138_new_n6252_), .B(u2__abc_52138_new_n10864_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10865_));
OAI21X1 OAI21X1_2583 ( .A(u2__abc_52138_new_n6250_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10867_));
OAI21X1 OAI21X1_2584 ( .A(u2__abc_52138_new_n10867_), .B(u2__abc_52138_new_n10866_), .C(u2__abc_52138_new_n10868_), .Y(u2__abc_52138_new_n10869_));
OAI21X1 OAI21X1_2585 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_404_), .Y(u2__abc_52138_new_n10871_));
OAI21X1 OAI21X1_2586 ( .A(u2__abc_52138_new_n6249_), .B(u2__abc_52138_new_n10874_), .C(u2__abc_52138_new_n6375_), .Y(u2__abc_52138_new_n10875_));
OAI21X1 OAI21X1_2587 ( .A(u2__abc_52138_new_n10872_), .B(u2__abc_52138_new_n10835_), .C(u2__abc_52138_new_n10876_), .Y(u2__abc_52138_new_n10877_));
OAI21X1 OAI21X1_2588 ( .A(u2__abc_52138_new_n6275_), .B(u2__abc_52138_new_n10877_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10880_));
OAI21X1 OAI21X1_2589 ( .A(u2__abc_52138_new_n6271_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10882_));
OAI21X1 OAI21X1_259 ( .A(aNan), .B(_abc_65734_new_n1568_), .C(_abc_65734_new_n1569_), .Y(\o[238] ));
OAI21X1 OAI21X1_2590 ( .A(u2__abc_52138_new_n10882_), .B(u2__abc_52138_new_n10881_), .C(u2__abc_52138_new_n10883_), .Y(u2__abc_52138_new_n10884_));
OAI21X1 OAI21X1_2591 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_405_), .Y(u2__abc_52138_new_n10886_));
OAI21X1 OAI21X1_2592 ( .A(u2_o_402_), .B(u2__abc_52138_new_n6271_), .C(u2__abc_52138_new_n10878_), .Y(u2__abc_52138_new_n10887_));
OAI21X1 OAI21X1_2593 ( .A(u2__abc_52138_new_n6268_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10890_));
OAI21X1 OAI21X1_2594 ( .A(u2__abc_52138_new_n10890_), .B(u2__abc_52138_new_n10889_), .C(u2__abc_52138_new_n10891_), .Y(u2__abc_52138_new_n10892_));
OAI21X1 OAI21X1_2595 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_406_), .Y(u2__abc_52138_new_n10894_));
OAI21X1 OAI21X1_2596 ( .A(u2_o_402_), .B(u2__abc_52138_new_n6271_), .C(u2__abc_52138_new_n6378_), .Y(u2__abc_52138_new_n10896_));
OAI21X1 OAI21X1_2597 ( .A(u2__abc_52138_new_n10896_), .B(u2__abc_52138_new_n10879_), .C(u2__abc_52138_new_n10895_), .Y(u2__abc_52138_new_n10897_));
OAI21X1 OAI21X1_2598 ( .A(u2__abc_52138_new_n6259_), .B(u2__abc_52138_new_n10898_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10899_));
OAI21X1 OAI21X1_2599 ( .A(u2__abc_52138_new_n6255_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10901_));
OAI21X1 OAI21X1_26 ( .A(aNan), .B(_abc_65734_new_n905_), .C(_abc_65734_new_n906_), .Y(\o[137] ));
OAI21X1 OAI21X1_260 ( .A(_abc_65734_new_n1571_), .B(_abc_65734_new_n1557_), .C(_abc_65734_new_n1572_), .Y(_abc_65734_new_n1573_));
OAI21X1 OAI21X1_2600 ( .A(u2__abc_52138_new_n10901_), .B(u2__abc_52138_new_n10900_), .C(u2__abc_52138_new_n10902_), .Y(u2__abc_52138_new_n10903_));
OAI21X1 OAI21X1_2601 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_407_), .Y(u2__abc_52138_new_n10905_));
OAI21X1 OAI21X1_2602 ( .A(u2__abc_52138_new_n6258_), .B(u2__abc_52138_new_n10897_), .C(u2__abc_52138_new_n10906_), .Y(u2__abc_52138_new_n10907_));
OAI21X1 OAI21X1_2603 ( .A(u2__abc_52138_new_n6264_), .B(u2__abc_52138_new_n10907_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10908_));
OAI21X1 OAI21X1_2604 ( .A(u2__abc_52138_new_n6260_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10910_));
OAI21X1 OAI21X1_2605 ( .A(u2__abc_52138_new_n10910_), .B(u2__abc_52138_new_n10909_), .C(u2__abc_52138_new_n10911_), .Y(u2__abc_52138_new_n10912_));
OAI21X1 OAI21X1_2606 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_408_), .Y(u2__abc_52138_new_n10914_));
OAI21X1 OAI21X1_2607 ( .A(u2__abc_52138_new_n6266_), .B(u2_remHi_403_), .C(u2__abc_52138_new_n10896_), .Y(u2__abc_52138_new_n10917_));
OAI21X1 OAI21X1_2608 ( .A(u2__abc_52138_new_n6265_), .B(u2__abc_52138_new_n10917_), .C(u2__abc_52138_new_n10918_), .Y(u2__abc_52138_new_n10919_));
OAI21X1 OAI21X1_2609 ( .A(u2__abc_52138_new_n6278_), .B(u2__abc_52138_new_n10835_), .C(u2__abc_52138_new_n10920_), .Y(u2__abc_52138_new_n10921_));
OAI21X1 OAI21X1_261 ( .A(_abc_65734_new_n1563_), .B(_abc_65734_new_n1582_), .C(_abc_65734_new_n753_), .Y(_abc_65734_new_n1583_));
OAI21X1 OAI21X1_2610 ( .A(u2__abc_52138_new_n6205_), .B(u2__abc_52138_new_n10921_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10924_));
OAI21X1 OAI21X1_2611 ( .A(u2__abc_52138_new_n6201_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10926_));
OAI21X1 OAI21X1_2612 ( .A(u2__abc_52138_new_n10926_), .B(u2__abc_52138_new_n10925_), .C(u2__abc_52138_new_n10927_), .Y(u2__abc_52138_new_n10928_));
OAI21X1 OAI21X1_2613 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_409_), .Y(u2__abc_52138_new_n10930_));
OAI21X1 OAI21X1_2614 ( .A(u2_o_406_), .B(u2__abc_52138_new_n6201_), .C(u2__abc_52138_new_n10922_), .Y(u2__abc_52138_new_n10931_));
OAI21X1 OAI21X1_2615 ( .A(u2__abc_52138_new_n6198_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10934_));
OAI21X1 OAI21X1_2616 ( .A(u2__abc_52138_new_n10934_), .B(u2__abc_52138_new_n10933_), .C(u2__abc_52138_new_n10935_), .Y(u2__abc_52138_new_n10936_));
OAI21X1 OAI21X1_2617 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_410_), .Y(u2__abc_52138_new_n10938_));
OAI21X1 OAI21X1_2618 ( .A(u2_o_406_), .B(u2__abc_52138_new_n6201_), .C(u2__abc_52138_new_n6358_), .Y(u2__abc_52138_new_n10940_));
OAI21X1 OAI21X1_2619 ( .A(u2__abc_52138_new_n10940_), .B(u2__abc_52138_new_n10923_), .C(u2__abc_52138_new_n10939_), .Y(u2__abc_52138_new_n10941_));
OAI21X1 OAI21X1_262 ( .A(aNan), .B(_abc_65734_new_n1573_), .C(_abc_65734_new_n1584_), .Y(\o[240] ));
OAI21X1 OAI21X1_2620 ( .A(u2__abc_52138_new_n6189_), .B(u2__abc_52138_new_n10942_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10943_));
OAI21X1 OAI21X1_2621 ( .A(u2__abc_52138_new_n6185_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10945_));
OAI21X1 OAI21X1_2622 ( .A(u2__abc_52138_new_n10945_), .B(u2__abc_52138_new_n10944_), .C(u2__abc_52138_new_n10946_), .Y(u2__abc_52138_new_n10947_));
OAI21X1 OAI21X1_2623 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_411_), .Y(u2__abc_52138_new_n10949_));
OAI21X1 OAI21X1_2624 ( .A(u2__abc_52138_new_n6188_), .B(u2__abc_52138_new_n10941_), .C(u2__abc_52138_new_n10950_), .Y(u2__abc_52138_new_n10951_));
OAI21X1 OAI21X1_2625 ( .A(u2__abc_52138_new_n6194_), .B(u2__abc_52138_new_n10951_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10952_));
OAI21X1 OAI21X1_2626 ( .A(u2__abc_52138_new_n6192_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10954_));
OAI21X1 OAI21X1_2627 ( .A(u2__abc_52138_new_n10954_), .B(u2__abc_52138_new_n10953_), .C(u2__abc_52138_new_n10955_), .Y(u2__abc_52138_new_n10956_));
OAI21X1 OAI21X1_2628 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_412_), .Y(u2__abc_52138_new_n10958_));
OAI21X1 OAI21X1_2629 ( .A(u2__abc_52138_new_n6196_), .B(u2_remHi_407_), .C(u2__abc_52138_new_n10940_), .Y(u2__abc_52138_new_n10959_));
OAI21X1 OAI21X1_263 ( .A(u2__abc_52138_new_n2966_), .B(u2__abc_52138_new_n2978_), .C(u2_state_2_), .Y(u2__abc_52138_new_n2979_));
OAI21X1 OAI21X1_2630 ( .A(u2__abc_52138_new_n6191_), .B(u2__abc_52138_new_n10950_), .C(u2__abc_52138_new_n6360_), .Y(u2__abc_52138_new_n10960_));
OAI21X1 OAI21X1_2631 ( .A(u2__abc_52138_new_n6195_), .B(u2__abc_52138_new_n10959_), .C(u2__abc_52138_new_n10961_), .Y(u2__abc_52138_new_n10962_));
OAI21X1 OAI21X1_2632 ( .A(u2__abc_52138_new_n6228_), .B(u2__abc_52138_new_n10964_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10967_));
OAI21X1 OAI21X1_2633 ( .A(u2__abc_52138_new_n6224_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10969_));
OAI21X1 OAI21X1_2634 ( .A(u2__abc_52138_new_n10969_), .B(u2__abc_52138_new_n10968_), .C(u2__abc_52138_new_n10970_), .Y(u2__abc_52138_new_n10971_));
OAI21X1 OAI21X1_2635 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_413_), .Y(u2__abc_52138_new_n10973_));
OAI21X1 OAI21X1_2636 ( .A(u2__abc_52138_new_n6227_), .B(u2__abc_52138_new_n10963_), .C(u2__abc_52138_new_n10974_), .Y(u2__abc_52138_new_n10975_));
OAI21X1 OAI21X1_2637 ( .A(u2__abc_52138_new_n6221_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10978_));
OAI21X1 OAI21X1_2638 ( .A(u2__abc_52138_new_n10978_), .B(u2__abc_52138_new_n10977_), .C(u2__abc_52138_new_n10979_), .Y(u2__abc_52138_new_n10980_));
OAI21X1 OAI21X1_2639 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_414_), .Y(u2__abc_52138_new_n10982_));
OAI21X1 OAI21X1_264 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n2992_), .C(u2__abc_52138_new_n2987_), .Y(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_1_));
OAI21X1 OAI21X1_2640 ( .A(u2_o_411_), .B(u2__abc_52138_new_n6221_), .C(u2__abc_52138_new_n10974_), .Y(u2__abc_52138_new_n10983_));
OAI21X1 OAI21X1_2641 ( .A(u2__abc_52138_new_n10983_), .B(u2__abc_52138_new_n10966_), .C(u2__abc_52138_new_n6365_), .Y(u2__abc_52138_new_n10984_));
OAI21X1 OAI21X1_2642 ( .A(u2__abc_52138_new_n6212_), .B(u2__abc_52138_new_n10985_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10986_));
OAI21X1 OAI21X1_2643 ( .A(u2__abc_52138_new_n6208_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10988_));
OAI21X1 OAI21X1_2644 ( .A(u2__abc_52138_new_n10988_), .B(u2__abc_52138_new_n10987_), .C(u2__abc_52138_new_n10989_), .Y(u2__abc_52138_new_n10990_));
OAI21X1 OAI21X1_2645 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_415_), .Y(u2__abc_52138_new_n10992_));
OAI21X1 OAI21X1_2646 ( .A(u2__abc_52138_new_n6211_), .B(u2__abc_52138_new_n10984_), .C(u2__abc_52138_new_n10993_), .Y(u2__abc_52138_new_n10994_));
OAI21X1 OAI21X1_2647 ( .A(u2__abc_52138_new_n6217_), .B(u2__abc_52138_new_n10994_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n10995_));
OAI21X1 OAI21X1_2648 ( .A(u2__abc_52138_new_n6213_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n10997_));
OAI21X1 OAI21X1_2649 ( .A(u2__abc_52138_new_n10997_), .B(u2__abc_52138_new_n10996_), .C(u2__abc_52138_new_n10998_), .Y(u2__abc_52138_new_n10999_));
OAI21X1 OAI21X1_265 ( .A(u2_state_2_), .B(u2_state_0_), .C(ce), .Y(u2__abc_52138_new_n2994_));
OAI21X1 OAI21X1_2650 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_416_), .Y(u2__abc_52138_new_n11001_));
OAI21X1 OAI21X1_2651 ( .A(u2__abc_52138_new_n10659_), .B(u2__abc_52138_new_n10647_), .C(u2__abc_52138_new_n6331_), .Y(u2__abc_52138_new_n11002_));
OAI21X1 OAI21X1_2652 ( .A(u2__abc_52138_new_n10993_), .B(u2__abc_52138_new_n6216_), .C(u2__abc_52138_new_n11003_), .Y(u2__abc_52138_new_n11004_));
OAI21X1 OAI21X1_2653 ( .A(u2__abc_52138_new_n6329_), .B(u2__abc_52138_new_n10749_), .C(u2__abc_52138_new_n11006_), .Y(u2__abc_52138_new_n11007_));
OAI21X1 OAI21X1_2654 ( .A(u2__abc_52138_new_n6231_), .B(u2__abc_52138_new_n10920_), .C(u2__abc_52138_new_n11008_), .Y(u2__abc_52138_new_n11009_));
OAI21X1 OAI21X1_2655 ( .A(u2__abc_52138_new_n6129_), .B(u2__abc_52138_new_n11011_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11014_));
OAI21X1 OAI21X1_2656 ( .A(u2__abc_52138_new_n6125_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11016_));
OAI21X1 OAI21X1_2657 ( .A(u2__abc_52138_new_n11016_), .B(u2__abc_52138_new_n11015_), .C(u2__abc_52138_new_n11017_), .Y(u2__abc_52138_new_n11018_));
OAI21X1 OAI21X1_2658 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_417_), .Y(u2__abc_52138_new_n11020_));
OAI21X1 OAI21X1_2659 ( .A(u2_o_414_), .B(u2__abc_52138_new_n6125_), .C(u2__abc_52138_new_n11012_), .Y(u2__abc_52138_new_n11021_));
OAI21X1 OAI21X1_266 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_0_), .Y(u2__abc_52138_new_n2995_));
OAI21X1 OAI21X1_2660 ( .A(u2__abc_52138_new_n6122_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11024_));
OAI21X1 OAI21X1_2661 ( .A(u2__abc_52138_new_n11024_), .B(u2__abc_52138_new_n11023_), .C(u2__abc_52138_new_n11025_), .Y(u2__abc_52138_new_n11026_));
OAI21X1 OAI21X1_2662 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_418_), .Y(u2__abc_52138_new_n11028_));
OAI21X1 OAI21X1_2663 ( .A(u2_o_414_), .B(u2__abc_52138_new_n6125_), .C(u2__abc_52138_new_n11029_), .Y(u2__abc_52138_new_n11030_));
OAI21X1 OAI21X1_2664 ( .A(u2__abc_52138_new_n11030_), .B(u2__abc_52138_new_n11013_), .C(u2__abc_52138_new_n6388_), .Y(u2__abc_52138_new_n11031_));
OAI21X1 OAI21X1_2665 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n11033_), .Y(u2__abc_52138_new_n11034_));
OAI21X1 OAI21X1_2666 ( .A(u2__abc_52138_new_n6110_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11036_));
OAI21X1 OAI21X1_2667 ( .A(u2__abc_52138_new_n11036_), .B(u2__abc_52138_new_n11035_), .C(u2__abc_52138_new_n11037_), .Y(u2__abc_52138_new_n11038_));
OAI21X1 OAI21X1_2668 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_419_), .Y(u2__abc_52138_new_n11040_));
OAI21X1 OAI21X1_2669 ( .A(u2__abc_52138_new_n6112_), .B(u2__abc_52138_new_n11031_), .C(u2__abc_52138_new_n6109_), .Y(u2__abc_52138_new_n11042_));
OAI21X1 OAI21X1_267 ( .A(u2_o_448_), .B(u2__abc_52138_new_n2999_), .C(u2__abc_52138_new_n3000_), .Y(u2__abc_52138_new_n3001_));
OAI21X1 OAI21X1_2670 ( .A(u2__abc_52138_new_n11041_), .B(u2__abc_52138_new_n11042_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11043_));
OAI21X1 OAI21X1_2671 ( .A(u2__abc_52138_new_n6113_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11045_));
OAI21X1 OAI21X1_2672 ( .A(u2__abc_52138_new_n11045_), .B(u2__abc_52138_new_n11044_), .C(u2__abc_52138_new_n11046_), .Y(u2__abc_52138_new_n11047_));
OAI21X1 OAI21X1_2673 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_420_), .Y(u2__abc_52138_new_n11049_));
OAI21X1 OAI21X1_2674 ( .A(u2__abc_52138_new_n6120_), .B(u2_remHi_415_), .C(u2__abc_52138_new_n11030_), .Y(u2__abc_52138_new_n11050_));
OAI21X1 OAI21X1_2675 ( .A(u2__abc_52138_new_n6109_), .B(u2__abc_52138_new_n6117_), .C(u2__abc_52138_new_n6116_), .Y(u2__abc_52138_new_n11051_));
OAI21X1 OAI21X1_2676 ( .A(u2__abc_52138_new_n6119_), .B(u2__abc_52138_new_n11050_), .C(u2__abc_52138_new_n11052_), .Y(u2__abc_52138_new_n11053_));
OAI21X1 OAI21X1_2677 ( .A(u2__abc_52138_new_n6105_), .B(u2__abc_52138_new_n11055_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11058_));
OAI21X1 OAI21X1_2678 ( .A(u2__abc_52138_new_n6101_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11060_));
OAI21X1 OAI21X1_2679 ( .A(u2__abc_52138_new_n11060_), .B(u2__abc_52138_new_n11059_), .C(u2__abc_52138_new_n11061_), .Y(u2__abc_52138_new_n11062_));
OAI21X1 OAI21X1_268 ( .A(u2__abc_52138_new_n3071_), .B(u2__abc_52138_new_n3068_), .C(u2__abc_52138_new_n3077_), .Y(u2__abc_52138_new_n3078_));
OAI21X1 OAI21X1_2680 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_421_), .Y(u2__abc_52138_new_n11064_));
OAI21X1 OAI21X1_2681 ( .A(u2__abc_52138_new_n6104_), .B(u2__abc_52138_new_n11054_), .C(u2__abc_52138_new_n11065_), .Y(u2__abc_52138_new_n11066_));
OAI21X1 OAI21X1_2682 ( .A(u2__abc_52138_new_n6098_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11069_));
OAI21X1 OAI21X1_2683 ( .A(u2__abc_52138_new_n11069_), .B(u2__abc_52138_new_n11068_), .C(u2__abc_52138_new_n11070_), .Y(u2__abc_52138_new_n11071_));
OAI21X1 OAI21X1_2684 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_422_), .Y(u2__abc_52138_new_n11073_));
OAI21X1 OAI21X1_2685 ( .A(u2_o_419_), .B(u2__abc_52138_new_n6098_), .C(u2__abc_52138_new_n11065_), .Y(u2__abc_52138_new_n11074_));
OAI21X1 OAI21X1_2686 ( .A(u2__abc_52138_new_n11074_), .B(u2__abc_52138_new_n11057_), .C(u2__abc_52138_new_n6393_), .Y(u2__abc_52138_new_n11075_));
OAI21X1 OAI21X1_2687 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n11077_), .Y(u2__abc_52138_new_n11078_));
OAI21X1 OAI21X1_2688 ( .A(u2__abc_52138_new_n6086_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11080_));
OAI21X1 OAI21X1_2689 ( .A(u2__abc_52138_new_n11080_), .B(u2__abc_52138_new_n11079_), .C(u2__abc_52138_new_n11081_), .Y(u2__abc_52138_new_n11082_));
OAI21X1 OAI21X1_269 ( .A(u2__abc_52138_new_n3058_), .B(u2__abc_52138_new_n3085_), .C(u2__abc_52138_new_n3090_), .Y(u2__abc_52138_new_n3091_));
OAI21X1 OAI21X1_2690 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_423_), .Y(u2__abc_52138_new_n11084_));
OAI21X1 OAI21X1_2691 ( .A(u2__abc_52138_new_n6088_), .B(u2__abc_52138_new_n11075_), .C(u2__abc_52138_new_n6085_), .Y(u2__abc_52138_new_n11086_));
OAI21X1 OAI21X1_2692 ( .A(u2__abc_52138_new_n11085_), .B(u2__abc_52138_new_n11086_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11087_));
OAI21X1 OAI21X1_2693 ( .A(u2__abc_52138_new_n6091_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11089_));
OAI21X1 OAI21X1_2694 ( .A(u2__abc_52138_new_n11089_), .B(u2__abc_52138_new_n11088_), .C(u2__abc_52138_new_n11090_), .Y(u2__abc_52138_new_n11091_));
OAI21X1 OAI21X1_2695 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_424_), .Y(u2__abc_52138_new_n11093_));
OAI21X1 OAI21X1_2696 ( .A(u2__abc_52138_new_n6085_), .B(u2__abc_52138_new_n6093_), .C(u2__abc_52138_new_n6090_), .Y(u2__abc_52138_new_n11096_));
OAI21X1 OAI21X1_2697 ( .A(u2__abc_52138_new_n6387_), .B(u2__abc_52138_new_n11094_), .C(u2__abc_52138_new_n11097_), .Y(u2__abc_52138_new_n11098_));
OAI21X1 OAI21X1_2698 ( .A(u2__abc_52138_new_n6051_), .B(u2__abc_52138_new_n11100_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11101_));
OAI21X1 OAI21X1_2699 ( .A(u2__abc_52138_new_n6047_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11103_));
OAI21X1 OAI21X1_27 ( .A(aNan), .B(_abc_65734_new_n908_), .C(_abc_65734_new_n909_), .Y(\o[138] ));
OAI21X1 OAI21X1_270 ( .A(sqrto_9_), .B(u2__abc_52138_new_n3037_), .C(u2__abc_52138_new_n3097_), .Y(u2__abc_52138_new_n3098_));
OAI21X1 OAI21X1_2700 ( .A(u2__abc_52138_new_n11103_), .B(u2__abc_52138_new_n11102_), .C(u2__abc_52138_new_n11104_), .Y(u2__abc_52138_new_n11105_));
OAI21X1 OAI21X1_2701 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_425_), .Y(u2__abc_52138_new_n11107_));
OAI21X1 OAI21X1_2702 ( .A(u2__abc_52138_new_n6050_), .B(u2__abc_52138_new_n11099_), .C(u2__abc_52138_new_n11108_), .Y(u2__abc_52138_new_n11109_));
OAI21X1 OAI21X1_2703 ( .A(u2__abc_52138_new_n6054_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11112_));
OAI21X1 OAI21X1_2704 ( .A(u2__abc_52138_new_n11112_), .B(u2__abc_52138_new_n11111_), .C(u2__abc_52138_new_n11113_), .Y(u2__abc_52138_new_n11114_));
OAI21X1 OAI21X1_2705 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_426_), .Y(u2__abc_52138_new_n11116_));
OAI21X1 OAI21X1_2706 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n11120_), .Y(u2__abc_52138_new_n11121_));
OAI21X1 OAI21X1_2707 ( .A(u2__abc_52138_new_n6038_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11123_));
OAI21X1 OAI21X1_2708 ( .A(u2__abc_52138_new_n11123_), .B(u2__abc_52138_new_n11122_), .C(u2__abc_52138_new_n11124_), .Y(u2__abc_52138_new_n11125_));
OAI21X1 OAI21X1_2709 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_427_), .Y(u2__abc_52138_new_n11127_));
OAI21X1 OAI21X1_271 ( .A(u2__abc_52138_new_n3095_), .B(u2__abc_52138_new_n3039_), .C(u2__abc_52138_new_n3099_), .Y(u2__abc_52138_new_n3100_));
OAI21X1 OAI21X1_2710 ( .A(u2__abc_52138_new_n6040_), .B(u2__abc_52138_new_n11118_), .C(u2__abc_52138_new_n6037_), .Y(u2__abc_52138_new_n11129_));
OAI21X1 OAI21X1_2711 ( .A(u2__abc_52138_new_n11128_), .B(u2__abc_52138_new_n11129_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11130_));
OAI21X1 OAI21X1_2712 ( .A(u2__abc_52138_new_n6041_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11132_));
OAI21X1 OAI21X1_2713 ( .A(u2__abc_52138_new_n11132_), .B(u2__abc_52138_new_n11131_), .C(u2__abc_52138_new_n11133_), .Y(u2__abc_52138_new_n11134_));
OAI21X1 OAI21X1_2714 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_428_), .Y(u2__abc_52138_new_n11136_));
OAI21X1 OAI21X1_2715 ( .A(u2__abc_52138_new_n6037_), .B(u2__abc_52138_new_n6045_), .C(u2__abc_52138_new_n6044_), .Y(u2__abc_52138_new_n11138_));
OAI21X1 OAI21X1_2716 ( .A(u2__abc_52138_new_n6057_), .B(u2__abc_52138_new_n11099_), .C(u2__abc_52138_new_n11139_), .Y(u2__abc_52138_new_n11140_));
OAI21X1 OAI21X1_2717 ( .A(u2__abc_52138_new_n6079_), .B(u2__abc_52138_new_n11140_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11143_));
OAI21X1 OAI21X1_2718 ( .A(u2__abc_52138_new_n6075_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11145_));
OAI21X1 OAI21X1_2719 ( .A(u2__abc_52138_new_n11145_), .B(u2__abc_52138_new_n11144_), .C(u2__abc_52138_new_n11146_), .Y(u2__abc_52138_new_n11147_));
OAI21X1 OAI21X1_272 ( .A(u2__abc_52138_new_n3021_), .B(u2__abc_52138_new_n3108_), .C(u2__abc_52138_new_n3105_), .Y(u2__abc_52138_new_n3109_));
OAI21X1 OAI21X1_2720 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_429_), .Y(u2__abc_52138_new_n11149_));
OAI21X1 OAI21X1_2721 ( .A(u2_o_426_), .B(u2__abc_52138_new_n6075_), .C(u2__abc_52138_new_n11141_), .Y(u2__abc_52138_new_n11150_));
OAI21X1 OAI21X1_2722 ( .A(u2__abc_52138_new_n6072_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11153_));
OAI21X1 OAI21X1_2723 ( .A(u2__abc_52138_new_n11153_), .B(u2__abc_52138_new_n11152_), .C(u2__abc_52138_new_n11154_), .Y(u2__abc_52138_new_n11155_));
OAI21X1 OAI21X1_2724 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_430_), .Y(u2__abc_52138_new_n11157_));
OAI21X1 OAI21X1_2725 ( .A(u2__abc_52138_new_n11159_), .B(u2__abc_52138_new_n11142_), .C(u2__abc_52138_new_n6406_), .Y(u2__abc_52138_new_n11160_));
OAI21X1 OAI21X1_2726 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n11162_), .Y(u2__abc_52138_new_n11163_));
OAI21X1 OAI21X1_2727 ( .A(u2__abc_52138_new_n6060_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11165_));
OAI21X1 OAI21X1_2728 ( .A(u2__abc_52138_new_n11165_), .B(u2__abc_52138_new_n11164_), .C(u2__abc_52138_new_n11166_), .Y(u2__abc_52138_new_n11167_));
OAI21X1 OAI21X1_2729 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_431_), .Y(u2__abc_52138_new_n11169_));
OAI21X1 OAI21X1_273 ( .A(u2__abc_52138_new_n3052_), .B(u2__abc_52138_new_n3092_), .C(u2__abc_52138_new_n3110_), .Y(u2__abc_52138_new_n3111_));
OAI21X1 OAI21X1_2730 ( .A(u2__abc_52138_new_n6062_), .B(u2__abc_52138_new_n11160_), .C(u2__abc_52138_new_n6059_), .Y(u2__abc_52138_new_n11171_));
OAI21X1 OAI21X1_2731 ( .A(u2__abc_52138_new_n11170_), .B(u2__abc_52138_new_n11171_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11172_));
OAI21X1 OAI21X1_2732 ( .A(u2__abc_52138_new_n6065_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11174_));
OAI21X1 OAI21X1_2733 ( .A(u2__abc_52138_new_n11174_), .B(u2__abc_52138_new_n11173_), .C(u2__abc_52138_new_n11175_), .Y(u2__abc_52138_new_n11176_));
OAI21X1 OAI21X1_2734 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_432_), .Y(u2__abc_52138_new_n11178_));
OAI21X1 OAI21X1_2735 ( .A(u2__abc_52138_new_n6059_), .B(u2__abc_52138_new_n6067_), .C(u2__abc_52138_new_n6064_), .Y(u2__abc_52138_new_n11181_));
OAI21X1 OAI21X1_2736 ( .A(u2__abc_52138_new_n11139_), .B(u2__abc_52138_new_n6082_), .C(u2__abc_52138_new_n11182_), .Y(u2__abc_52138_new_n11183_));
OAI21X1 OAI21X1_2737 ( .A(u2__abc_52138_new_n6134_), .B(u2__abc_52138_new_n11179_), .C(u2__abc_52138_new_n11184_), .Y(u2__abc_52138_new_n11185_));
OAI21X1 OAI21X1_2738 ( .A(u2__abc_52138_new_n6014_), .B(u2__abc_52138_new_n11185_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11186_));
OAI21X1 OAI21X1_2739 ( .A(u2__abc_52138_new_n6010_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11188_));
OAI21X1 OAI21X1_274 ( .A(u2__abc_52138_new_n3198_), .B(u2__abc_52138_new_n3201_), .C(u2__abc_52138_new_n3204_), .Y(u2__abc_52138_new_n3205_));
OAI21X1 OAI21X1_2740 ( .A(u2__abc_52138_new_n11188_), .B(u2__abc_52138_new_n11187_), .C(u2__abc_52138_new_n11189_), .Y(u2__abc_52138_new_n11190_));
OAI21X1 OAI21X1_2741 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_433_), .Y(u2__abc_52138_new_n11192_));
OAI21X1 OAI21X1_2742 ( .A(u2__abc_52138_new_n6013_), .B(u2__abc_52138_new_n11194_), .C(u2__abc_52138_new_n11193_), .Y(u2__abc_52138_new_n11195_));
OAI21X1 OAI21X1_2743 ( .A(u2__abc_52138_new_n6019_), .B(u2__abc_52138_new_n11195_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11196_));
OAI21X1 OAI21X1_2744 ( .A(u2__abc_52138_new_n6017_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11198_));
OAI21X1 OAI21X1_2745 ( .A(u2__abc_52138_new_n11198_), .B(u2__abc_52138_new_n11197_), .C(u2__abc_52138_new_n11199_), .Y(u2__abc_52138_new_n11200_));
OAI21X1 OAI21X1_2746 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_434_), .Y(u2__abc_52138_new_n11202_));
OAI21X1 OAI21X1_2747 ( .A(u2__abc_52138_new_n6016_), .B(u2__abc_52138_new_n11193_), .C(u2__abc_52138_new_n6427_), .Y(u2__abc_52138_new_n11203_));
OAI21X1 OAI21X1_2748 ( .A(u2__abc_52138_new_n6020_), .B(u2__abc_52138_new_n11194_), .C(u2__abc_52138_new_n11204_), .Y(u2__abc_52138_new_n11205_));
OAI21X1 OAI21X1_2749 ( .A(u2__abc_52138_new_n6025_), .B(u2__abc_52138_new_n11205_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11208_));
OAI21X1 OAI21X1_275 ( .A(u2__abc_52138_new_n3212_), .B(u2__abc_52138_new_n3213_), .C(u2__abc_52138_new_n3186_), .Y(u2__abc_52138_new_n3214_));
OAI21X1 OAI21X1_2750 ( .A(u2__abc_52138_new_n6021_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11210_));
OAI21X1 OAI21X1_2751 ( .A(u2__abc_52138_new_n11210_), .B(u2__abc_52138_new_n11209_), .C(u2__abc_52138_new_n11211_), .Y(u2__abc_52138_new_n11212_));
OAI21X1 OAI21X1_2752 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_435_), .Y(u2__abc_52138_new_n11214_));
OAI21X1 OAI21X1_2753 ( .A(u2__abc_52138_new_n6021_), .B(u2_o_432_), .C(u2__abc_52138_new_n11206_), .Y(u2__abc_52138_new_n11215_));
OAI21X1 OAI21X1_2754 ( .A(u2__abc_52138_new_n6030_), .B(u2__abc_52138_new_n11215_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11216_));
OAI21X1 OAI21X1_2755 ( .A(u2__abc_52138_new_n6028_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11218_));
OAI21X1 OAI21X1_2756 ( .A(u2__abc_52138_new_n11218_), .B(u2__abc_52138_new_n11217_), .C(u2__abc_52138_new_n11219_), .Y(u2__abc_52138_new_n11220_));
OAI21X1 OAI21X1_2757 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_436_), .Y(u2__abc_52138_new_n11222_));
OAI21X1 OAI21X1_2758 ( .A(u2__abc_52138_new_n11224_), .B(u2__abc_52138_new_n11207_), .C(u2__abc_52138_new_n11223_), .Y(u2__abc_52138_new_n11225_));
OAI21X1 OAI21X1_2759 ( .A(u2__abc_52138_new_n6007_), .B(u2__abc_52138_new_n11226_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11227_));
OAI21X1 OAI21X1_276 ( .A(u2__abc_52138_new_n3187_), .B(u2__abc_52138_new_n3210_), .C(u2__abc_52138_new_n3215_), .Y(u2__abc_52138_new_n3216_));
OAI21X1 OAI21X1_2760 ( .A(u2__abc_52138_new_n6003_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11229_));
OAI21X1 OAI21X1_2761 ( .A(u2__abc_52138_new_n11229_), .B(u2__abc_52138_new_n11228_), .C(u2__abc_52138_new_n11230_), .Y(u2__abc_52138_new_n11231_));
OAI21X1 OAI21X1_2762 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_437_), .Y(u2__abc_52138_new_n11233_));
OAI21X1 OAI21X1_2763 ( .A(u2__abc_52138_new_n6006_), .B(u2__abc_52138_new_n11225_), .C(u2__abc_52138_new_n11234_), .Y(u2__abc_52138_new_n11235_));
OAI21X1 OAI21X1_2764 ( .A(u2__abc_52138_new_n6002_), .B(u2__abc_52138_new_n11235_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11238_));
OAI21X1 OAI21X1_2765 ( .A(u2__abc_52138_new_n6000_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11240_));
OAI21X1 OAI21X1_2766 ( .A(u2__abc_52138_new_n11240_), .B(u2__abc_52138_new_n11239_), .C(u2__abc_52138_new_n11241_), .Y(u2__abc_52138_new_n11242_));
OAI21X1 OAI21X1_2767 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_438_), .Y(u2__abc_52138_new_n11244_));
OAI21X1 OAI21X1_2768 ( .A(u2__abc_52138_new_n6001_), .B(u2__abc_52138_new_n11237_), .C(u2__abc_52138_new_n5991_), .Y(u2__abc_52138_new_n11245_));
OAI21X1 OAI21X1_2769 ( .A(u2_o_435_), .B(u2__abc_52138_new_n6000_), .C(u2__abc_52138_new_n11236_), .Y(u2__abc_52138_new_n11246_));
OAI21X1 OAI21X1_277 ( .A(u2__abc_52138_new_n3115_), .B(u2__abc_52138_new_n3225_), .C(u2__abc_52138_new_n3120_), .Y(u2__abc_52138_new_n3226_));
OAI21X1 OAI21X1_2770 ( .A(u2__abc_52138_new_n5987_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11250_));
OAI21X1 OAI21X1_2771 ( .A(u2__abc_52138_new_n11250_), .B(u2__abc_52138_new_n11249_), .C(u2__abc_52138_new_n11251_), .Y(u2__abc_52138_new_n11252_));
OAI21X1 OAI21X1_2772 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_439_), .Y(u2__abc_52138_new_n11254_));
OAI21X1 OAI21X1_2773 ( .A(u2__abc_52138_new_n5987_), .B(u2_o_436_), .C(u2__abc_52138_new_n11245_), .Y(u2__abc_52138_new_n11255_));
OAI21X1 OAI21X1_2774 ( .A(u2__abc_52138_new_n5996_), .B(u2__abc_52138_new_n11255_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11256_));
OAI21X1 OAI21X1_2775 ( .A(u2__abc_52138_new_n5992_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11258_));
OAI21X1 OAI21X1_2776 ( .A(u2__abc_52138_new_n11258_), .B(u2__abc_52138_new_n11257_), .C(u2__abc_52138_new_n11259_), .Y(u2__abc_52138_new_n11260_));
OAI21X1 OAI21X1_2777 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_440_), .Y(u2__abc_52138_new_n11262_));
OAI21X1 OAI21X1_2778 ( .A(u2_remHi_433_), .B(u2__abc_52138_new_n6026_), .C(u2__abc_52138_new_n11224_), .Y(u2__abc_52138_new_n11263_));
OAI21X1 OAI21X1_2779 ( .A(u2__abc_52138_new_n6031_), .B(u2__abc_52138_new_n11204_), .C(u2__abc_52138_new_n11263_), .Y(u2__abc_52138_new_n11264_));
OAI21X1 OAI21X1_278 ( .A(u2__abc_52138_new_n3224_), .B(u2__abc_52138_new_n3221_), .C(u2__abc_52138_new_n3227_), .Y(u2__abc_52138_new_n3228_));
OAI21X1 OAI21X1_2780 ( .A(u2__abc_52138_new_n5997_), .B(u2__abc_52138_new_n11265_), .C(u2__abc_52138_new_n11266_), .Y(u2__abc_52138_new_n11267_));
OAI21X1 OAI21X1_2781 ( .A(u2__abc_52138_new_n6033_), .B(u2__abc_52138_new_n11194_), .C(u2__abc_52138_new_n11268_), .Y(u2__abc_52138_new_n11269_));
OAI21X1 OAI21X1_2782 ( .A(u2__abc_52138_new_n5971_), .B(u2__abc_52138_new_n11269_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11270_));
OAI21X1 OAI21X1_2783 ( .A(u2__abc_52138_new_n5967_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11272_));
OAI21X1 OAI21X1_2784 ( .A(u2__abc_52138_new_n11272_), .B(u2__abc_52138_new_n11271_), .C(u2__abc_52138_new_n11273_), .Y(u2__abc_52138_new_n11274_));
OAI21X1 OAI21X1_2785 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_441_), .Y(u2__abc_52138_new_n11276_));
OAI21X1 OAI21X1_2786 ( .A(u2_o_438_), .B(u2__abc_52138_new_n5967_), .C(u2__abc_52138_new_n11277_), .Y(u2__abc_52138_new_n11278_));
OAI21X1 OAI21X1_2787 ( .A(u2__abc_52138_new_n5972_), .B(u2__abc_52138_new_n11278_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11279_));
OAI21X1 OAI21X1_2788 ( .A(u2__abc_52138_new_n6415_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11281_));
OAI21X1 OAI21X1_2789 ( .A(u2__abc_52138_new_n11281_), .B(u2__abc_52138_new_n11280_), .C(u2__abc_52138_new_n11282_), .Y(u2__abc_52138_new_n11283_));
OAI21X1 OAI21X1_279 ( .A(u2__abc_52138_new_n3235_), .B(u2__abc_52138_new_n3229_), .C(u2__abc_52138_new_n3232_), .Y(u2__abc_52138_new_n3236_));
OAI21X1 OAI21X1_2790 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_442_), .Y(u2__abc_52138_new_n11285_));
OAI21X1 OAI21X1_2791 ( .A(u2__abc_52138_new_n6414_), .B(u2_remHi_439_), .C(u2__abc_52138_new_n5968_), .Y(u2__abc_52138_new_n11288_));
OAI21X1 OAI21X1_2792 ( .A(u2_o_439_), .B(u2__abc_52138_new_n6415_), .C(u2__abc_52138_new_n11288_), .Y(u2__abc_52138_new_n11289_));
OAI21X1 OAI21X1_2793 ( .A(u2__abc_52138_new_n5975_), .B(u2__abc_52138_new_n5977_), .C(u2__abc_52138_new_n11290_), .Y(u2__abc_52138_new_n11292_));
OAI21X1 OAI21X1_2794 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n11292_), .Y(u2__abc_52138_new_n11293_));
OAI21X1 OAI21X1_2795 ( .A(u2__abc_52138_new_n5974_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11295_));
OAI21X1 OAI21X1_2796 ( .A(u2__abc_52138_new_n11295_), .B(u2__abc_52138_new_n11294_), .C(u2__abc_52138_new_n11296_), .Y(u2__abc_52138_new_n11297_));
OAI21X1 OAI21X1_2797 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_443_), .Y(u2__abc_52138_new_n11299_));
OAI21X1 OAI21X1_2798 ( .A(u2__abc_52138_new_n5977_), .B(u2__abc_52138_new_n11290_), .C(u2__abc_52138_new_n11300_), .Y(u2__abc_52138_new_n11301_));
OAI21X1 OAI21X1_2799 ( .A(u2__abc_52138_new_n5983_), .B(u2__abc_52138_new_n11301_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11302_));
OAI21X1 OAI21X1_28 ( .A(aNan), .B(_abc_65734_new_n911_), .C(_abc_65734_new_n912_), .Y(\o[139] ));
OAI21X1 OAI21X1_280 ( .A(u2__abc_52138_new_n3158_), .B(u2__abc_52138_new_n3217_), .C(u2__abc_52138_new_n3237_), .Y(u2__abc_52138_new_n3238_));
OAI21X1 OAI21X1_2800 ( .A(u2__abc_52138_new_n5981_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11304_));
OAI21X1 OAI21X1_2801 ( .A(u2__abc_52138_new_n11304_), .B(u2__abc_52138_new_n11303_), .C(u2__abc_52138_new_n11305_), .Y(u2__abc_52138_new_n11306_));
OAI21X1 OAI21X1_2802 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_444_), .Y(u2__abc_52138_new_n11308_));
OAI21X1 OAI21X1_2803 ( .A(u2__abc_52138_new_n5980_), .B(u2__abc_52138_new_n11300_), .C(u2__abc_52138_new_n11309_), .Y(u2__abc_52138_new_n11310_));
OAI21X1 OAI21X1_2804 ( .A(u2__abc_52138_new_n5964_), .B(u2__abc_52138_new_n11313_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11316_));
OAI21X1 OAI21X1_2805 ( .A(u2__abc_52138_new_n5960_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11318_));
OAI21X1 OAI21X1_2806 ( .A(u2__abc_52138_new_n11318_), .B(u2__abc_52138_new_n11317_), .C(u2__abc_52138_new_n11319_), .Y(u2__abc_52138_new_n11320_));
OAI21X1 OAI21X1_2807 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_445_), .Y(u2__abc_52138_new_n11322_));
OAI21X1 OAI21X1_2808 ( .A(u2_o_442_), .B(u2__abc_52138_new_n5960_), .C(u2__abc_52138_new_n11314_), .Y(u2__abc_52138_new_n11323_));
OAI21X1 OAI21X1_2809 ( .A(u2__abc_52138_new_n5957_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11326_));
OAI21X1 OAI21X1_281 ( .A(u2__abc_52138_new_n3433_), .B(u2__abc_52138_new_n3436_), .C(u2__abc_52138_new_n3440_), .Y(u2__abc_52138_new_n3441_));
OAI21X1 OAI21X1_2810 ( .A(u2__abc_52138_new_n11326_), .B(u2__abc_52138_new_n11325_), .C(u2__abc_52138_new_n11327_), .Y(u2__abc_52138_new_n11328_));
OAI21X1 OAI21X1_2811 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_446_), .Y(u2__abc_52138_new_n11330_));
OAI21X1 OAI21X1_2812 ( .A(u2__abc_52138_new_n11333_), .B(u2__abc_52138_new_n11315_), .C(u2__abc_52138_new_n11331_), .Y(u2__abc_52138_new_n11334_));
OAI21X1 OAI21X1_2813 ( .A(u2__abc_52138_new_n5948_), .B(u2__abc_52138_new_n11335_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11336_));
OAI21X1 OAI21X1_2814 ( .A(u2__abc_52138_new_n5944_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11338_));
OAI21X1 OAI21X1_2815 ( .A(u2__abc_52138_new_n11338_), .B(u2__abc_52138_new_n11337_), .C(u2__abc_52138_new_n11339_), .Y(u2__abc_52138_new_n11340_));
OAI21X1 OAI21X1_2816 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_447_), .Y(u2__abc_52138_new_n11342_));
OAI21X1 OAI21X1_2817 ( .A(u2__abc_52138_new_n5947_), .B(u2__abc_52138_new_n11334_), .C(u2__abc_52138_new_n11343_), .Y(u2__abc_52138_new_n11344_));
OAI21X1 OAI21X1_2818 ( .A(u2__abc_52138_new_n5953_), .B(u2__abc_52138_new_n11344_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11345_));
OAI21X1 OAI21X1_2819 ( .A(u2__abc_52138_new_n5951_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11347_));
OAI21X1 OAI21X1_282 ( .A(u2__abc_52138_new_n3429_), .B(u2__abc_52138_new_n3446_), .C(u2__abc_52138_new_n3449_), .Y(u2__abc_52138_new_n3450_));
OAI21X1 OAI21X1_2820 ( .A(u2__abc_52138_new_n11347_), .B(u2__abc_52138_new_n11346_), .C(u2__abc_52138_new_n11348_), .Y(u2__abc_52138_new_n11349_));
OAI21X1 OAI21X1_2821 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_448_), .Y(u2__abc_52138_new_n11351_));
OAI21X1 OAI21X1_2822 ( .A(u2__abc_52138_new_n5950_), .B(u2__abc_52138_new_n11343_), .C(u2__abc_52138_new_n6424_), .Y(u2__abc_52138_new_n11354_));
OAI21X1 OAI21X1_2823 ( .A(u2__abc_52138_new_n11353_), .B(u2__abc_52138_new_n11311_), .C(u2__abc_52138_new_n11356_), .Y(u2__abc_52138_new_n11357_));
OAI21X1 OAI21X1_2824 ( .A(u2__abc_52138_new_n6035_), .B(u2__abc_52138_new_n11184_), .C(u2__abc_52138_new_n11358_), .Y(u2__abc_52138_new_n11359_));
OAI21X1 OAI21X1_2825 ( .A(u2__abc_52138_new_n3012_), .B(u2__abc_52138_new_n11361_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11362_));
OAI21X1 OAI21X1_2826 ( .A(u2__abc_52138_new_n3008_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11364_));
OAI21X1 OAI21X1_2827 ( .A(u2__abc_52138_new_n11364_), .B(u2__abc_52138_new_n11363_), .C(u2__abc_52138_new_n11365_), .Y(u2__abc_52138_new_n11366_));
OAI21X1 OAI21X1_2828 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_449_), .Y(u2__abc_52138_new_n11368_));
OAI21X1 OAI21X1_2829 ( .A(u2__abc_52138_new_n3011_), .B(u2__abc_52138_new_n11360_), .C(u2__abc_52138_new_n11369_), .Y(u2__abc_52138_new_n11370_));
OAI21X1 OAI21X1_283 ( .A(u2__abc_52138_new_n3338_), .B(u2__abc_52138_new_n3456_), .C(u2__abc_52138_new_n3343_), .Y(u2__abc_52138_new_n3457_));
OAI21X1 OAI21X1_2830 ( .A(u2__abc_52138_new_n3007_), .B(u2__abc_52138_new_n11370_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n11371_));
OAI21X1 OAI21X1_2831 ( .A(u2__abc_52138_new_n3003_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n11373_));
OAI21X1 OAI21X1_2832 ( .A(u2__abc_52138_new_n11373_), .B(u2__abc_52138_new_n11372_), .C(u2__abc_52138_new_n11374_), .Y(u2__abc_52138_new_n11375_));
OAI21X1 OAI21X1_2833 ( .A(u2__abc_52138_new_n2962_), .B(u2__abc_52138_new_n2963_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11378_));
OAI21X1 OAI21X1_2834 ( .A(u2__abc_52138_new_n11378_), .B(u2__abc_52138_new_n2991_), .C(u2__abc_52138_new_n11377_), .Y(u2__abc_52138_new_n11379_));
OAI21X1 OAI21X1_2835 ( .A(rst), .B(ce), .C(u2_cnt_0_), .Y(u2__abc_52138_new_n11380_));
OAI21X1 OAI21X1_2836 ( .A(u2__abc_52138_new_n2962_), .B(u2__abc_52138_new_n2963_), .C(u2__abc_52138_new_n11388_), .Y(u2__abc_52138_new_n11389_));
OAI21X1 OAI21X1_2837 ( .A(u2_cnt_3_), .B(u2__abc_52138_new_n11391_), .C(u2__abc_52138_new_n11395_), .Y(u2__abc_52138_new_n11396_));
OAI21X1 OAI21X1_2838 ( .A(u2_cnt_4_), .B(u2__abc_52138_new_n11393_), .C(u2__abc_52138_new_n11395_), .Y(u2__abc_52138_new_n11399_));
OAI21X1 OAI21X1_2839 ( .A(u2_cnt_5_), .B(u2__abc_52138_new_n11398_), .C(u2__abc_52138_new_n11395_), .Y(u2__abc_52138_new_n11403_));
OAI21X1 OAI21X1_284 ( .A(u2__abc_52138_new_n3455_), .B(u2__abc_52138_new_n3452_), .C(u2__abc_52138_new_n3458_), .Y(u2__abc_52138_new_n3459_));
OAI21X1 OAI21X1_2840 ( .A(u2__abc_52138_new_n11406_), .B(u2__abc_52138_new_n11401_), .C(u2__abc_52138_new_n2965_), .Y(u2__abc_52138_new_n11407_));
OAI21X1 OAI21X1_2841 ( .A(u2__abc_52138_new_n11407_), .B(u2__abc_52138_new_n11405_), .C(u2__abc_52138_new_n7779_), .Y(u2__0cnt_7_0__6_));
OAI21X1 OAI21X1_2842 ( .A(u2__abc_52138_new_n11394_), .B(u2__abc_52138_new_n11410_), .C(u2__abc_52138_new_n7779_), .Y(u2__0cnt_7_0__7_));
OAI21X1 OAI21X1_2843 ( .A(ld), .B(u2__abc_52138_new_n2963_), .C(u2__abc_52138_new_n2992_), .Y(u2__abc_52138_new_n11412_));
OAI21X1 OAI21X1_2844 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_0_), .Y(u2__abc_52138_new_n11413_));
OAI21X1 OAI21X1_2845 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_1_), .Y(u2__abc_52138_new_n11415_));
OAI21X1 OAI21X1_2846 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_2_), .Y(u2__abc_52138_new_n11417_));
OAI21X1 OAI21X1_2847 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_3_), .Y(u2__abc_52138_new_n11420_));
OAI21X1 OAI21X1_2848 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_4_), .Y(u2__abc_52138_new_n11423_));
OAI21X1 OAI21X1_2849 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_5_), .Y(u2__abc_52138_new_n11426_));
OAI21X1 OAI21X1_285 ( .A(u2__abc_52138_new_n3377_), .B(u2__abc_52138_new_n3460_), .C(u2__abc_52138_new_n3372_), .Y(u2__abc_52138_new_n3461_));
OAI21X1 OAI21X1_2850 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_6_), .Y(u2__abc_52138_new_n11429_));
OAI21X1 OAI21X1_2851 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_7_), .Y(u2__abc_52138_new_n11432_));
OAI21X1 OAI21X1_2852 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_8_), .Y(u2__abc_52138_new_n11435_));
OAI21X1 OAI21X1_2853 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_9_), .Y(u2__abc_52138_new_n11438_));
OAI21X1 OAI21X1_2854 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_10_), .Y(u2__abc_52138_new_n11441_));
OAI21X1 OAI21X1_2855 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_11_), .Y(u2__abc_52138_new_n11444_));
OAI21X1 OAI21X1_2856 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_12_), .Y(u2__abc_52138_new_n11447_));
OAI21X1 OAI21X1_2857 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_13_), .Y(u2__abc_52138_new_n11450_));
OAI21X1 OAI21X1_2858 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_14_), .Y(u2__abc_52138_new_n11453_));
OAI21X1 OAI21X1_2859 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_15_), .Y(u2__abc_52138_new_n11456_));
OAI21X1 OAI21X1_286 ( .A(u2__abc_52138_new_n3361_), .B(u2__abc_52138_new_n3463_), .C(u2__abc_52138_new_n3366_), .Y(u2__abc_52138_new_n3464_));
OAI21X1 OAI21X1_2860 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_16_), .Y(u2__abc_52138_new_n11459_));
OAI21X1 OAI21X1_2861 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_17_), .Y(u2__abc_52138_new_n11462_));
OAI21X1 OAI21X1_2862 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_18_), .Y(u2__abc_52138_new_n11465_));
OAI21X1 OAI21X1_2863 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_19_), .Y(u2__abc_52138_new_n11468_));
OAI21X1 OAI21X1_2864 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_20_), .Y(u2__abc_52138_new_n11471_));
OAI21X1 OAI21X1_2865 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_21_), .Y(u2__abc_52138_new_n11474_));
OAI21X1 OAI21X1_2866 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_22_), .Y(u2__abc_52138_new_n11477_));
OAI21X1 OAI21X1_2867 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_23_), .Y(u2__abc_52138_new_n11480_));
OAI21X1 OAI21X1_2868 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_24_), .Y(u2__abc_52138_new_n11483_));
OAI21X1 OAI21X1_2869 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_25_), .Y(u2__abc_52138_new_n11486_));
OAI21X1 OAI21X1_287 ( .A(u2__abc_52138_new_n3427_), .B(u2__abc_52138_new_n3451_), .C(u2__abc_52138_new_n3467_), .Y(u2__abc_52138_new_n3468_));
OAI21X1 OAI21X1_2870 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_26_), .Y(u2__abc_52138_new_n11489_));
OAI21X1 OAI21X1_2871 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_27_), .Y(u2__abc_52138_new_n11492_));
OAI21X1 OAI21X1_2872 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_28_), .Y(u2__abc_52138_new_n11495_));
OAI21X1 OAI21X1_2873 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_29_), .Y(u2__abc_52138_new_n11498_));
OAI21X1 OAI21X1_2874 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_30_), .Y(u2__abc_52138_new_n11501_));
OAI21X1 OAI21X1_2875 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_31_), .Y(u2__abc_52138_new_n11504_));
OAI21X1 OAI21X1_2876 ( .A(u2__abc_52138_new_n11515_), .B(u2__abc_52138_new_n11513_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11516_));
OAI21X1 OAI21X1_2877 ( .A(u2__abc_52138_new_n11512_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11516_), .Y(u2__0remLo_451_0__33_));
OAI21X1 OAI21X1_2878 ( .A(u2__abc_52138_new_n11527_), .B(u2__abc_52138_new_n11525_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11528_));
OAI21X1 OAI21X1_2879 ( .A(u2__abc_52138_new_n11524_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11528_), .Y(u2__0remLo_451_0__36_));
OAI21X1 OAI21X1_288 ( .A(u2__abc_52138_new_n3472_), .B(u2__abc_52138_new_n3293_), .C(u2__abc_52138_new_n3473_), .Y(u2__abc_52138_new_n3474_));
OAI21X1 OAI21X1_2880 ( .A(u2__abc_52138_new_n11566_), .B(u2__abc_52138_new_n11564_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11567_));
OAI21X1 OAI21X1_2881 ( .A(u2__abc_52138_new_n11563_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11567_), .Y(u2__0remLo_451_0__48_));
OAI21X1 OAI21X1_2882 ( .A(u2__abc_52138_new_n11626_), .B(u2__abc_52138_new_n11624_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11627_));
OAI21X1 OAI21X1_2883 ( .A(u2__abc_52138_new_n11623_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11627_), .Y(u2__0remLo_451_0__67_));
OAI21X1 OAI21X1_2884 ( .A(u2__abc_52138_new_n11656_), .B(u2__abc_52138_new_n11654_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11657_));
OAI21X1 OAI21X1_2885 ( .A(u2__abc_52138_new_n11653_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11657_), .Y(u2__0remLo_451_0__76_));
OAI21X1 OAI21X1_2886 ( .A(u2__abc_52138_new_n11716_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11719_), .Y(u2__0remLo_451_0__96_));
OAI21X1 OAI21X1_2887 ( .A(u2__abc_52138_new_n11724_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11726_), .Y(u2__0remLo_451_0__98_));
OAI21X1 OAI21X1_2888 ( .A(u2__abc_52138_new_n11731_), .B(u2__abc_52138_new_n11729_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11732_));
OAI21X1 OAI21X1_2889 ( .A(u2__abc_52138_new_n11728_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11732_), .Y(u2__0remLo_451_0__99_));
OAI21X1 OAI21X1_289 ( .A(u2__abc_52138_new_n3471_), .B(u2__abc_52138_new_n3297_), .C(u2__abc_52138_new_n3475_), .Y(u2__abc_52138_new_n3476_));
OAI21X1 OAI21X1_2890 ( .A(u2__abc_52138_new_n11785_), .B(u2__abc_52138_new_n11783_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11786_));
OAI21X1 OAI21X1_2891 ( .A(u2__abc_52138_new_n11782_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11786_), .Y(u2__0remLo_451_0__116_));
OAI21X1 OAI21X1_2892 ( .A(u2__abc_52138_new_n11833_), .B(u2__abc_52138_new_n11831_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11834_));
OAI21X1 OAI21X1_2893 ( .A(u2__abc_52138_new_n11830_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11834_), .Y(u2__0remLo_451_0__131_));
OAI21X1 OAI21X1_2894 ( .A(u2__abc_52138_new_n11839_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11841_), .Y(u2__0remLo_451_0__133_));
OAI21X1 OAI21X1_2895 ( .A(u2__abc_52138_new_n11933_), .B(u2__abc_52138_new_n11931_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n11934_));
OAI21X1 OAI21X1_2896 ( .A(u2__abc_52138_new_n11930_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11934_), .Y(u2__0remLo_451_0__163_));
OAI21X1 OAI21X1_2897 ( .A(u2__abc_52138_new_n11966_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n11968_), .Y(u2__0remLo_451_0__174_));
OAI21X1 OAI21X1_2898 ( .A(u2__abc_52138_new_n12033_), .B(u2__abc_52138_new_n12031_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n12034_));
OAI21X1 OAI21X1_2899 ( .A(u2__abc_52138_new_n12030_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n12034_), .Y(u2__0remLo_451_0__195_));
OAI21X1 OAI21X1_29 ( .A(aNan), .B(_abc_65734_new_n914_), .C(_abc_65734_new_n915_), .Y(\o[140] ));
OAI21X1 OAI21X1_290 ( .A(u2__abc_52138_new_n3330_), .B(u2__abc_52138_new_n3478_), .C(u2__abc_52138_new_n3325_), .Y(u2__abc_52138_new_n3479_));
OAI21X1 OAI21X1_2900 ( .A(u2__abc_52138_new_n12063_), .B(u2__abc_52138_new_n12061_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n12064_));
OAI21X1 OAI21X1_2901 ( .A(u2__abc_52138_new_n12060_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n12064_), .Y(u2__0remLo_451_0__204_));
OAI21X1 OAI21X1_2902 ( .A(u2__abc_52138_new_n12069_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n12071_), .Y(u2__0remLo_451_0__206_));
OAI21X1 OAI21X1_2903 ( .A(u2__abc_52138_new_n12136_), .B(u2__abc_52138_new_n12134_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n12137_));
OAI21X1 OAI21X1_2904 ( .A(u2__abc_52138_new_n12133_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n12137_), .Y(u2__0remLo_451_0__227_));
OAI21X1 OAI21X1_2905 ( .A(u2__abc_52138_new_n12142_), .B(u2__abc_52138_new_n12140_), .C(u2__abc_52138_new_n2981_), .Y(u2__abc_52138_new_n12143_));
OAI21X1 OAI21X1_2906 ( .A(u2__abc_52138_new_n12139_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n12143_), .Y(u2__0remLo_451_0__228_));
OAI21X1 OAI21X1_2907 ( .A(u2__abc_52138_new_n12160_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n12162_), .Y(u2__0remLo_451_0__234_));
OAI21X1 OAI21X1_2908 ( .A(u2__abc_52138_new_n12227_), .B(u2__abc_52138_new_n11508_), .C(u2__abc_52138_new_n12229_), .Y(u2__0remLo_451_0__256_));
OAI21X1 OAI21X1_2909 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_258_), .Y(u2__abc_52138_new_n12234_));
OAI21X1 OAI21X1_291 ( .A(u2__abc_52138_new_n3480_), .B(u2__abc_52138_new_n3477_), .C(u2__abc_52138_new_n3483_), .Y(u2__abc_52138_new_n3484_));
OAI21X1 OAI21X1_2910 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_259_), .Y(u2__abc_52138_new_n12237_));
OAI21X1 OAI21X1_2911 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_260_), .Y(u2__abc_52138_new_n12240_));
OAI21X1 OAI21X1_2912 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_261_), .Y(u2__abc_52138_new_n12243_));
OAI21X1 OAI21X1_2913 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_262_), .Y(u2__abc_52138_new_n12246_));
OAI21X1 OAI21X1_2914 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_263_), .Y(u2__abc_52138_new_n12249_));
OAI21X1 OAI21X1_2915 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_264_), .Y(u2__abc_52138_new_n12252_));
OAI21X1 OAI21X1_2916 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_265_), .Y(u2__abc_52138_new_n12255_));
OAI21X1 OAI21X1_2917 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_266_), .Y(u2__abc_52138_new_n12258_));
OAI21X1 OAI21X1_2918 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_267_), .Y(u2__abc_52138_new_n12261_));
OAI21X1 OAI21X1_2919 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_268_), .Y(u2__abc_52138_new_n12264_));
OAI21X1 OAI21X1_292 ( .A(u2__abc_52138_new_n3243_), .B(u2__abc_52138_new_n3249_), .C(u2__abc_52138_new_n3248_), .Y(u2__abc_52138_new_n3491_));
OAI21X1 OAI21X1_2920 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_269_), .Y(u2__abc_52138_new_n12267_));
OAI21X1 OAI21X1_2921 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_270_), .Y(u2__abc_52138_new_n12270_));
OAI21X1 OAI21X1_2922 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_271_), .Y(u2__abc_52138_new_n12273_));
OAI21X1 OAI21X1_2923 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_272_), .Y(u2__abc_52138_new_n12276_));
OAI21X1 OAI21X1_2924 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_273_), .Y(u2__abc_52138_new_n12279_));
OAI21X1 OAI21X1_2925 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_274_), .Y(u2__abc_52138_new_n12282_));
OAI21X1 OAI21X1_2926 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_275_), .Y(u2__abc_52138_new_n12285_));
OAI21X1 OAI21X1_2927 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_276_), .Y(u2__abc_52138_new_n12288_));
OAI21X1 OAI21X1_2928 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_277_), .Y(u2__abc_52138_new_n12291_));
OAI21X1 OAI21X1_2929 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_278_), .Y(u2__abc_52138_new_n12294_));
OAI21X1 OAI21X1_293 ( .A(u2__abc_52138_new_n3490_), .B(u2__abc_52138_new_n3487_), .C(u2__abc_52138_new_n3492_), .Y(u2__abc_52138_new_n3493_));
OAI21X1 OAI21X1_2930 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_279_), .Y(u2__abc_52138_new_n12297_));
OAI21X1 OAI21X1_2931 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_280_), .Y(u2__abc_52138_new_n12300_));
OAI21X1 OAI21X1_2932 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_281_), .Y(u2__abc_52138_new_n12303_));
OAI21X1 OAI21X1_2933 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_282_), .Y(u2__abc_52138_new_n12306_));
OAI21X1 OAI21X1_2934 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_283_), .Y(u2__abc_52138_new_n12309_));
OAI21X1 OAI21X1_2935 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_284_), .Y(u2__abc_52138_new_n12312_));
OAI21X1 OAI21X1_2936 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_285_), .Y(u2__abc_52138_new_n12315_));
OAI21X1 OAI21X1_2937 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_286_), .Y(u2__abc_52138_new_n12318_));
OAI21X1 OAI21X1_2938 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_287_), .Y(u2__abc_52138_new_n12321_));
OAI21X1 OAI21X1_2939 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_288_), .Y(u2__abc_52138_new_n12324_));
OAI21X1 OAI21X1_294 ( .A(u2__abc_52138_new_n3282_), .B(u2__abc_52138_new_n3494_), .C(u2__abc_52138_new_n3277_), .Y(u2__abc_52138_new_n3495_));
OAI21X1 OAI21X1_2940 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_289_), .Y(u2__abc_52138_new_n12327_));
OAI21X1 OAI21X1_2941 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_290_), .Y(u2__abc_52138_new_n12330_));
OAI21X1 OAI21X1_2942 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_291_), .Y(u2__abc_52138_new_n12333_));
OAI21X1 OAI21X1_2943 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_292_), .Y(u2__abc_52138_new_n12336_));
OAI21X1 OAI21X1_2944 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_293_), .Y(u2__abc_52138_new_n12339_));
OAI21X1 OAI21X1_2945 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_294_), .Y(u2__abc_52138_new_n12342_));
OAI21X1 OAI21X1_2946 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_295_), .Y(u2__abc_52138_new_n12345_));
OAI21X1 OAI21X1_2947 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_296_), .Y(u2__abc_52138_new_n12348_));
OAI21X1 OAI21X1_2948 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_297_), .Y(u2__abc_52138_new_n12351_));
OAI21X1 OAI21X1_2949 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_298_), .Y(u2__abc_52138_new_n12354_));
OAI21X1 OAI21X1_295 ( .A(u2__abc_52138_new_n3422_), .B(u2__abc_52138_new_n3485_), .C(u2__abc_52138_new_n3499_), .Y(u2__abc_52138_new_n3500_));
OAI21X1 OAI21X1_2950 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_299_), .Y(u2__abc_52138_new_n12357_));
OAI21X1 OAI21X1_2951 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_300_), .Y(u2__abc_52138_new_n12360_));
OAI21X1 OAI21X1_2952 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_301_), .Y(u2__abc_52138_new_n12363_));
OAI21X1 OAI21X1_2953 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_302_), .Y(u2__abc_52138_new_n12366_));
OAI21X1 OAI21X1_2954 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_303_), .Y(u2__abc_52138_new_n12369_));
OAI21X1 OAI21X1_2955 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_304_), .Y(u2__abc_52138_new_n12372_));
OAI21X1 OAI21X1_2956 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_305_), .Y(u2__abc_52138_new_n12375_));
OAI21X1 OAI21X1_2957 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_306_), .Y(u2__abc_52138_new_n12378_));
OAI21X1 OAI21X1_2958 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_307_), .Y(u2__abc_52138_new_n12381_));
OAI21X1 OAI21X1_2959 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_308_), .Y(u2__abc_52138_new_n12384_));
OAI21X1 OAI21X1_296 ( .A(u2__abc_52138_new_n3421_), .B(u2__abc_52138_new_n3239_), .C(u2__abc_52138_new_n3501_), .Y(u2__abc_52138_new_n3502_));
OAI21X1 OAI21X1_2960 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_309_), .Y(u2__abc_52138_new_n12387_));
OAI21X1 OAI21X1_2961 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_310_), .Y(u2__abc_52138_new_n12390_));
OAI21X1 OAI21X1_2962 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_311_), .Y(u2__abc_52138_new_n12393_));
OAI21X1 OAI21X1_2963 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_312_), .Y(u2__abc_52138_new_n12396_));
OAI21X1 OAI21X1_2964 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_313_), .Y(u2__abc_52138_new_n12399_));
OAI21X1 OAI21X1_2965 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_314_), .Y(u2__abc_52138_new_n12402_));
OAI21X1 OAI21X1_2966 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_315_), .Y(u2__abc_52138_new_n12405_));
OAI21X1 OAI21X1_2967 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_316_), .Y(u2__abc_52138_new_n12408_));
OAI21X1 OAI21X1_2968 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_317_), .Y(u2__abc_52138_new_n12411_));
OAI21X1 OAI21X1_2969 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_318_), .Y(u2__abc_52138_new_n12414_));
OAI21X1 OAI21X1_297 ( .A(u2__abc_52138_new_n3873_), .B(u2__abc_52138_new_n3876_), .C(u2__abc_52138_new_n3879_), .Y(u2__abc_52138_new_n3880_));
OAI21X1 OAI21X1_2970 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_319_), .Y(u2__abc_52138_new_n12417_));
OAI21X1 OAI21X1_2971 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_320_), .Y(u2__abc_52138_new_n12420_));
OAI21X1 OAI21X1_2972 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_321_), .Y(u2__abc_52138_new_n12423_));
OAI21X1 OAI21X1_2973 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_322_), .Y(u2__abc_52138_new_n12426_));
OAI21X1 OAI21X1_2974 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_323_), .Y(u2__abc_52138_new_n12429_));
OAI21X1 OAI21X1_2975 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_324_), .Y(u2__abc_52138_new_n12432_));
OAI21X1 OAI21X1_2976 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_325_), .Y(u2__abc_52138_new_n12435_));
OAI21X1 OAI21X1_2977 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_326_), .Y(u2__abc_52138_new_n12438_));
OAI21X1 OAI21X1_2978 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_327_), .Y(u2__abc_52138_new_n12441_));
OAI21X1 OAI21X1_2979 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_328_), .Y(u2__abc_52138_new_n12444_));
OAI21X1 OAI21X1_298 ( .A(u2__abc_52138_new_n3889_), .B(u2__abc_52138_new_n3890_), .C(u2__abc_52138_new_n3859_), .Y(u2__abc_52138_new_n3891_));
OAI21X1 OAI21X1_2980 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_329_), .Y(u2__abc_52138_new_n12447_));
OAI21X1 OAI21X1_2981 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_330_), .Y(u2__abc_52138_new_n12450_));
OAI21X1 OAI21X1_2982 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_331_), .Y(u2__abc_52138_new_n12453_));
OAI21X1 OAI21X1_2983 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_332_), .Y(u2__abc_52138_new_n12456_));
OAI21X1 OAI21X1_2984 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_333_), .Y(u2__abc_52138_new_n12459_));
OAI21X1 OAI21X1_2985 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_334_), .Y(u2__abc_52138_new_n12462_));
OAI21X1 OAI21X1_2986 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_335_), .Y(u2__abc_52138_new_n12465_));
OAI21X1 OAI21X1_2987 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_336_), .Y(u2__abc_52138_new_n12468_));
OAI21X1 OAI21X1_2988 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_337_), .Y(u2__abc_52138_new_n12471_));
OAI21X1 OAI21X1_2989 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_338_), .Y(u2__abc_52138_new_n12474_));
OAI21X1 OAI21X1_299 ( .A(u2__abc_52138_new_n3860_), .B(u2__abc_52138_new_n3887_), .C(u2__abc_52138_new_n3892_), .Y(u2__abc_52138_new_n3893_));
OAI21X1 OAI21X1_2990 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_339_), .Y(u2__abc_52138_new_n12477_));
OAI21X1 OAI21X1_2991 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_340_), .Y(u2__abc_52138_new_n12480_));
OAI21X1 OAI21X1_2992 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_341_), .Y(u2__abc_52138_new_n12483_));
OAI21X1 OAI21X1_2993 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_342_), .Y(u2__abc_52138_new_n12486_));
OAI21X1 OAI21X1_2994 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_343_), .Y(u2__abc_52138_new_n12489_));
OAI21X1 OAI21X1_2995 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_344_), .Y(u2__abc_52138_new_n12492_));
OAI21X1 OAI21X1_2996 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_345_), .Y(u2__abc_52138_new_n12495_));
OAI21X1 OAI21X1_2997 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_346_), .Y(u2__abc_52138_new_n12498_));
OAI21X1 OAI21X1_2998 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_347_), .Y(u2__abc_52138_new_n12501_));
OAI21X1 OAI21X1_2999 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_348_), .Y(u2__abc_52138_new_n12504_));
OAI21X1 OAI21X1_3 ( .A(aNan), .B(_abc_65734_new_n836_), .C(_abc_65734_new_n837_), .Y(\o[114] ));
OAI21X1 OAI21X1_30 ( .A(aNan), .B(_abc_65734_new_n917_), .C(_abc_65734_new_n918_), .Y(\o[141] ));
OAI21X1 OAI21X1_300 ( .A(u2__abc_52138_new_n3896_), .B(u2__abc_52138_new_n3806_), .C(u2__abc_52138_new_n3899_), .Y(u2__abc_52138_new_n3900_));
OAI21X1 OAI21X1_3000 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_349_), .Y(u2__abc_52138_new_n12507_));
OAI21X1 OAI21X1_3001 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_350_), .Y(u2__abc_52138_new_n12510_));
OAI21X1 OAI21X1_3002 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_351_), .Y(u2__abc_52138_new_n12513_));
OAI21X1 OAI21X1_3003 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_352_), .Y(u2__abc_52138_new_n12516_));
OAI21X1 OAI21X1_3004 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_353_), .Y(u2__abc_52138_new_n12519_));
OAI21X1 OAI21X1_3005 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_354_), .Y(u2__abc_52138_new_n12522_));
OAI21X1 OAI21X1_3006 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_355_), .Y(u2__abc_52138_new_n12525_));
OAI21X1 OAI21X1_3007 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_356_), .Y(u2__abc_52138_new_n12528_));
OAI21X1 OAI21X1_3008 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_357_), .Y(u2__abc_52138_new_n12531_));
OAI21X1 OAI21X1_3009 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_358_), .Y(u2__abc_52138_new_n12534_));
OAI21X1 OAI21X1_301 ( .A(u2__abc_52138_new_n3902_), .B(u2__abc_52138_new_n3818_), .C(u2__abc_52138_new_n3904_), .Y(u2__abc_52138_new_n3905_));
OAI21X1 OAI21X1_3010 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_359_), .Y(u2__abc_52138_new_n12537_));
OAI21X1 OAI21X1_3011 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_360_), .Y(u2__abc_52138_new_n12540_));
OAI21X1 OAI21X1_3012 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_361_), .Y(u2__abc_52138_new_n12543_));
OAI21X1 OAI21X1_3013 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_362_), .Y(u2__abc_52138_new_n12546_));
OAI21X1 OAI21X1_3014 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_363_), .Y(u2__abc_52138_new_n12549_));
OAI21X1 OAI21X1_3015 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_364_), .Y(u2__abc_52138_new_n12552_));
OAI21X1 OAI21X1_3016 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_365_), .Y(u2__abc_52138_new_n12555_));
OAI21X1 OAI21X1_3017 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_366_), .Y(u2__abc_52138_new_n12558_));
OAI21X1 OAI21X1_3018 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_367_), .Y(u2__abc_52138_new_n12561_));
OAI21X1 OAI21X1_3019 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_368_), .Y(u2__abc_52138_new_n12564_));
OAI21X1 OAI21X1_302 ( .A(u2__abc_52138_new_n3831_), .B(u2__abc_52138_new_n3894_), .C(u2__abc_52138_new_n3906_), .Y(u2__abc_52138_new_n3907_));
OAI21X1 OAI21X1_3020 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_369_), .Y(u2__abc_52138_new_n12567_));
OAI21X1 OAI21X1_3021 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_370_), .Y(u2__abc_52138_new_n12570_));
OAI21X1 OAI21X1_3022 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_371_), .Y(u2__abc_52138_new_n12573_));
OAI21X1 OAI21X1_3023 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_372_), .Y(u2__abc_52138_new_n12576_));
OAI21X1 OAI21X1_3024 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_373_), .Y(u2__abc_52138_new_n12579_));
OAI21X1 OAI21X1_3025 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_374_), .Y(u2__abc_52138_new_n12582_));
OAI21X1 OAI21X1_3026 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_375_), .Y(u2__abc_52138_new_n12585_));
OAI21X1 OAI21X1_3027 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_376_), .Y(u2__abc_52138_new_n12588_));
OAI21X1 OAI21X1_3028 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_377_), .Y(u2__abc_52138_new_n12591_));
OAI21X1 OAI21X1_3029 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_378_), .Y(u2__abc_52138_new_n12594_));
OAI21X1 OAI21X1_303 ( .A(u2__abc_52138_new_n3910_), .B(u2__abc_52138_new_n3759_), .C(u2__abc_52138_new_n3913_), .Y(u2__abc_52138_new_n3914_));
OAI21X1 OAI21X1_3030 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_379_), .Y(u2__abc_52138_new_n12597_));
OAI21X1 OAI21X1_3031 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_380_), .Y(u2__abc_52138_new_n12600_));
OAI21X1 OAI21X1_3032 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_381_), .Y(u2__abc_52138_new_n12603_));
OAI21X1 OAI21X1_3033 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_382_), .Y(u2__abc_52138_new_n12606_));
OAI21X1 OAI21X1_3034 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_383_), .Y(u2__abc_52138_new_n12609_));
OAI21X1 OAI21X1_3035 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_384_), .Y(u2__abc_52138_new_n12612_));
OAI21X1 OAI21X1_3036 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_385_), .Y(u2__abc_52138_new_n12615_));
OAI21X1 OAI21X1_3037 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_386_), .Y(u2__abc_52138_new_n12618_));
OAI21X1 OAI21X1_3038 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_387_), .Y(u2__abc_52138_new_n12621_));
OAI21X1 OAI21X1_3039 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_388_), .Y(u2__abc_52138_new_n12624_));
OAI21X1 OAI21X1_304 ( .A(u2__abc_52138_new_n3764_), .B(u2__abc_52138_new_n3918_), .C(u2__abc_52138_new_n3769_), .Y(u2__abc_52138_new_n3919_));
OAI21X1 OAI21X1_3040 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_389_), .Y(u2__abc_52138_new_n12627_));
OAI21X1 OAI21X1_3041 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_390_), .Y(u2__abc_52138_new_n12630_));
OAI21X1 OAI21X1_3042 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_391_), .Y(u2__abc_52138_new_n12633_));
OAI21X1 OAI21X1_3043 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_392_), .Y(u2__abc_52138_new_n12636_));
OAI21X1 OAI21X1_3044 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_393_), .Y(u2__abc_52138_new_n12639_));
OAI21X1 OAI21X1_3045 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_394_), .Y(u2__abc_52138_new_n12642_));
OAI21X1 OAI21X1_3046 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_395_), .Y(u2__abc_52138_new_n12645_));
OAI21X1 OAI21X1_3047 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_396_), .Y(u2__abc_52138_new_n12648_));
OAI21X1 OAI21X1_3048 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_397_), .Y(u2__abc_52138_new_n12651_));
OAI21X1 OAI21X1_3049 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_398_), .Y(u2__abc_52138_new_n12654_));
OAI21X1 OAI21X1_305 ( .A(u2__abc_52138_new_n3917_), .B(u2__abc_52138_new_n3915_), .C(u2__abc_52138_new_n3920_), .Y(u2__abc_52138_new_n3921_));
OAI21X1 OAI21X1_3050 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_399_), .Y(u2__abc_52138_new_n12657_));
OAI21X1 OAI21X1_3051 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_400_), .Y(u2__abc_52138_new_n12660_));
OAI21X1 OAI21X1_3052 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_401_), .Y(u2__abc_52138_new_n12663_));
OAI21X1 OAI21X1_3053 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_402_), .Y(u2__abc_52138_new_n12666_));
OAI21X1 OAI21X1_3054 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_403_), .Y(u2__abc_52138_new_n12669_));
OAI21X1 OAI21X1_3055 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_404_), .Y(u2__abc_52138_new_n12672_));
OAI21X1 OAI21X1_3056 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_405_), .Y(u2__abc_52138_new_n12675_));
OAI21X1 OAI21X1_3057 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_406_), .Y(u2__abc_52138_new_n12678_));
OAI21X1 OAI21X1_3058 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_407_), .Y(u2__abc_52138_new_n12681_));
OAI21X1 OAI21X1_3059 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_408_), .Y(u2__abc_52138_new_n12684_));
OAI21X1 OAI21X1_306 ( .A(u2__abc_52138_new_n3718_), .B(u2_remHi_89_), .C(u2__abc_52138_new_n3924_), .Y(u2__abc_52138_new_n3925_));
OAI21X1 OAI21X1_3060 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_409_), .Y(u2__abc_52138_new_n12687_));
OAI21X1 OAI21X1_3061 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_410_), .Y(u2__abc_52138_new_n12690_));
OAI21X1 OAI21X1_3062 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_411_), .Y(u2__abc_52138_new_n12693_));
OAI21X1 OAI21X1_3063 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_412_), .Y(u2__abc_52138_new_n12696_));
OAI21X1 OAI21X1_3064 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_413_), .Y(u2__abc_52138_new_n12699_));
OAI21X1 OAI21X1_3065 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_414_), .Y(u2__abc_52138_new_n12702_));
OAI21X1 OAI21X1_3066 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_415_), .Y(u2__abc_52138_new_n12705_));
OAI21X1 OAI21X1_3067 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_416_), .Y(u2__abc_52138_new_n12708_));
OAI21X1 OAI21X1_3068 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_417_), .Y(u2__abc_52138_new_n12711_));
OAI21X1 OAI21X1_3069 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_418_), .Y(u2__abc_52138_new_n12714_));
OAI21X1 OAI21X1_307 ( .A(u2__abc_52138_new_n3923_), .B(u2__abc_52138_new_n3723_), .C(u2__abc_52138_new_n3926_), .Y(u2__abc_52138_new_n3927_));
OAI21X1 OAI21X1_3070 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_419_), .Y(u2__abc_52138_new_n12717_));
OAI21X1 OAI21X1_3071 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_420_), .Y(u2__abc_52138_new_n12720_));
OAI21X1 OAI21X1_3072 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_421_), .Y(u2__abc_52138_new_n12723_));
OAI21X1 OAI21X1_3073 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_422_), .Y(u2__abc_52138_new_n12726_));
OAI21X1 OAI21X1_3074 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_423_), .Y(u2__abc_52138_new_n12729_));
OAI21X1 OAI21X1_3075 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_424_), .Y(u2__abc_52138_new_n12732_));
OAI21X1 OAI21X1_3076 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_425_), .Y(u2__abc_52138_new_n12735_));
OAI21X1 OAI21X1_3077 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_426_), .Y(u2__abc_52138_new_n12738_));
OAI21X1 OAI21X1_3078 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_427_), .Y(u2__abc_52138_new_n12741_));
OAI21X1 OAI21X1_3079 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_428_), .Y(u2__abc_52138_new_n12744_));
OAI21X1 OAI21X1_308 ( .A(sqrto_91_), .B(u2__abc_52138_new_n3704_), .C(u2__abc_52138_new_n3709_), .Y(u2__abc_52138_new_n3929_));
OAI21X1 OAI21X1_3080 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_429_), .Y(u2__abc_52138_new_n12747_));
OAI21X1 OAI21X1_3081 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_430_), .Y(u2__abc_52138_new_n12750_));
OAI21X1 OAI21X1_3082 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_431_), .Y(u2__abc_52138_new_n12753_));
OAI21X1 OAI21X1_3083 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_432_), .Y(u2__abc_52138_new_n12756_));
OAI21X1 OAI21X1_3084 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_433_), .Y(u2__abc_52138_new_n12759_));
OAI21X1 OAI21X1_3085 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_434_), .Y(u2__abc_52138_new_n12762_));
OAI21X1 OAI21X1_3086 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_435_), .Y(u2__abc_52138_new_n12765_));
OAI21X1 OAI21X1_3087 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_436_), .Y(u2__abc_52138_new_n12768_));
OAI21X1 OAI21X1_3088 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_437_), .Y(u2__abc_52138_new_n12771_));
OAI21X1 OAI21X1_3089 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_438_), .Y(u2__abc_52138_new_n12774_));
OAI21X1 OAI21X1_309 ( .A(u2__abc_52138_new_n3702_), .B(u2_remHi_91_), .C(u2__abc_52138_new_n3929_), .Y(u2__abc_52138_new_n3930_));
OAI21X1 OAI21X1_3090 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_439_), .Y(u2__abc_52138_new_n12777_));
OAI21X1 OAI21X1_3091 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_440_), .Y(u2__abc_52138_new_n12780_));
OAI21X1 OAI21X1_3092 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_441_), .Y(u2__abc_52138_new_n12783_));
OAI21X1 OAI21X1_3093 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_442_), .Y(u2__abc_52138_new_n12786_));
OAI21X1 OAI21X1_3094 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_443_), .Y(u2__abc_52138_new_n12789_));
OAI21X1 OAI21X1_3095 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_444_), .Y(u2__abc_52138_new_n12792_));
OAI21X1 OAI21X1_3096 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_445_), .Y(u2__abc_52138_new_n12795_));
OAI21X1 OAI21X1_3097 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_446_), .Y(u2__abc_52138_new_n12798_));
OAI21X1 OAI21X1_3098 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_447_), .Y(u2__abc_52138_new_n12801_));
OAI21X1 OAI21X1_3099 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_448_), .Y(u2__abc_52138_new_n12804_));
OAI21X1 OAI21X1_31 ( .A(aNan), .B(_abc_65734_new_n920_), .C(_abc_65734_new_n921_), .Y(\o[142] ));
OAI21X1 OAI21X1_310 ( .A(u2__abc_52138_new_n3694_), .B(u2__abc_52138_new_n3932_), .C(u2__abc_52138_new_n3699_), .Y(u2__abc_52138_new_n3933_));
OAI21X1 OAI21X1_3100 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remLo_449_), .Y(u2__abc_52138_new_n12807_));
OAI21X1 OAI21X1_3101 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remHiShift_0_), .Y(u2__abc_52138_new_n12810_));
OAI21X1 OAI21X1_3102 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_remHiShift_1_), .Y(u2__abc_52138_new_n12813_));
OAI21X1 OAI21X1_3103 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n11412_), .C(u2_root_0_), .Y(u2__abc_52138_new_n12816_));
OAI21X1 OAI21X1_3104 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_0_), .Y(u2__abc_52138_new_n12818_));
OAI21X1 OAI21X1_3105 ( .A(u2__abc_52138_new_n3063_), .B(u2__abc_52138_new_n6463_), .C(u2__abc_52138_new_n3082_), .Y(u2__abc_52138_new_n12825_));
OAI21X1 OAI21X1_3106 ( .A(u2__abc_52138_new_n3087_), .B(u2__abc_52138_new_n6579_), .C(u2__abc_52138_new_n3055_), .Y(u2__abc_52138_new_n12826_));
OAI21X1 OAI21X1_3107 ( .A(u2__abc_52138_new_n6466_), .B(u2__abc_52138_new_n12824_), .C(u2__abc_52138_new_n12827_), .Y(u2__abc_52138_new_n12828_));
OAI21X1 OAI21X1_3108 ( .A(u2__abc_52138_new_n3048_), .B(u2__abc_52138_new_n6600_), .C(u2__abc_52138_new_n3043_), .Y(u2__abc_52138_new_n12829_));
OAI21X1 OAI21X1_3109 ( .A(u2__abc_52138_new_n3035_), .B(u2_remHi_9_), .C(u2__abc_52138_new_n3098_), .Y(u2__abc_52138_new_n12830_));
OAI21X1 OAI21X1_311 ( .A(u2__abc_52138_new_n3737_), .B(u2__abc_52138_new_n3922_), .C(u2__abc_52138_new_n3936_), .Y(u2__abc_52138_new_n3937_));
OAI21X1 OAI21X1_3110 ( .A(u2__abc_52138_new_n3102_), .B(u2__abc_52138_new_n6653_), .C(u2__abc_52138_new_n3018_), .Y(u2__abc_52138_new_n12832_));
OAI21X1 OAI21X1_3111 ( .A(u2__abc_52138_new_n3030_), .B(u2__abc_52138_new_n12833_), .C(u2__abc_52138_new_n3025_), .Y(u2__abc_52138_new_n12834_));
OAI21X1 OAI21X1_3112 ( .A(u2__abc_52138_new_n12819_), .B(u2__abc_52138_new_n12831_), .C(u2__abc_52138_new_n12835_), .Y(u2__abc_52138_new_n12836_));
OAI21X1 OAI21X1_3113 ( .A(u2__abc_52138_new_n3173_), .B(u2__abc_52138_new_n6692_), .C(u2__abc_52138_new_n3178_), .Y(u2__abc_52138_new_n12841_));
OAI21X1 OAI21X1_3114 ( .A(u2__abc_52138_new_n3162_), .B(u2__abc_52138_new_n6713_), .C(u2__abc_52138_new_n3167_), .Y(u2__abc_52138_new_n12842_));
OAI21X1 OAI21X1_3115 ( .A(u2__abc_52138_new_n3192_), .B(u2__abc_52138_new_n12844_), .C(u2__abc_52138_new_n12845_), .Y(u2__abc_52138_new_n12846_));
OAI21X1 OAI21X1_3116 ( .A(u2__abc_52138_new_n12840_), .B(u2__abc_52138_new_n12843_), .C(u2__abc_52138_new_n12847_), .Y(u2__abc_52138_new_n12848_));
OAI21X1 OAI21X1_3117 ( .A(u2__abc_52138_new_n3131_), .B(u2__abc_52138_new_n3127_), .C(u2__abc_52138_new_n3126_), .Y(u2__abc_52138_new_n12849_));
OAI21X1 OAI21X1_3118 ( .A(u2__abc_52138_new_n3154_), .B(u2__abc_52138_new_n3150_), .C(u2__abc_52138_new_n3149_), .Y(u2__abc_52138_new_n12852_));
OAI21X1 OAI21X1_3119 ( .A(u2__abc_52138_new_n3157_), .B(u2__abc_52138_new_n12850_), .C(u2__abc_52138_new_n12853_), .Y(u2__abc_52138_new_n12854_));
OAI21X1 OAI21X1_312 ( .A(u2__abc_52138_new_n3942_), .B(u2__abc_52138_new_n3648_), .C(u2__abc_52138_new_n3943_), .Y(u2__abc_52138_new_n3944_));
OAI21X1 OAI21X1_3120 ( .A(u2__abc_52138_new_n12839_), .B(u2__abc_52138_new_n12837_), .C(u2__abc_52138_new_n12855_), .Y(u2__abc_52138_new_n12856_));
OAI21X1 OAI21X1_3121 ( .A(u2__abc_52138_new_n3392_), .B(u2__abc_52138_new_n12858_), .C(u2__abc_52138_new_n3397_), .Y(u2__abc_52138_new_n12859_));
OAI21X1 OAI21X1_3122 ( .A(sqrto_33_), .B(u2__abc_52138_new_n3385_), .C(u2__abc_52138_new_n3438_), .Y(u2__abc_52138_new_n12860_));
OAI21X1 OAI21X1_3123 ( .A(u2__abc_52138_new_n3383_), .B(u2_remHi_33_), .C(u2__abc_52138_new_n12860_), .Y(u2__abc_52138_new_n12861_));
OAI21X1 OAI21X1_3124 ( .A(u2__abc_52138_new_n3444_), .B(u2__abc_52138_new_n6895_), .C(u2__abc_52138_new_n3415_), .Y(u2__abc_52138_new_n12863_));
OAI21X1 OAI21X1_3125 ( .A(u2__abc_52138_new_n3404_), .B(u2__abc_52138_new_n3410_), .C(u2__abc_52138_new_n3409_), .Y(u2__abc_52138_new_n12864_));
OAI21X1 OAI21X1_3126 ( .A(u2__abc_52138_new_n3418_), .B(u2__abc_52138_new_n12862_), .C(u2__abc_52138_new_n12865_), .Y(u2__abc_52138_new_n12866_));
OAI21X1 OAI21X1_3127 ( .A(u2__abc_52138_new_n3349_), .B(u2__abc_52138_new_n6947_), .C(u2__abc_52138_new_n3354_), .Y(u2__abc_52138_new_n12867_));
OAI21X1 OAI21X1_3128 ( .A(u2__abc_52138_new_n3380_), .B(u2__abc_52138_new_n12868_), .C(u2__abc_52138_new_n12869_), .Y(u2__abc_52138_new_n12870_));
OAI21X1 OAI21X1_3129 ( .A(u2__abc_52138_new_n3306_), .B(u2__abc_52138_new_n3299_), .C(u2__abc_52138_new_n7030_), .Y(u2__abc_52138_new_n12874_));
OAI21X1 OAI21X1_313 ( .A(u2__abc_52138_new_n3941_), .B(u2__abc_52138_new_n3652_), .C(u2__abc_52138_new_n3945_), .Y(u2__abc_52138_new_n3946_));
OAI21X1 OAI21X1_3130 ( .A(u2__abc_52138_new_n7093_), .B(u2__abc_52138_new_n12875_), .C(u2__abc_52138_new_n12877_), .Y(u2__abc_52138_new_n12878_));
OAI21X1 OAI21X1_3131 ( .A(u2__abc_52138_new_n3254_), .B(u2__abc_52138_new_n3260_), .C(u2__abc_52138_new_n3259_), .Y(u2__abc_52138_new_n12879_));
OAI21X1 OAI21X1_3132 ( .A(u2__abc_52138_new_n3266_), .B(u2__abc_52138_new_n3272_), .C(u2__abc_52138_new_n3269_), .Y(u2__abc_52138_new_n12881_));
OAI21X1 OAI21X1_3133 ( .A(u2__abc_52138_new_n3285_), .B(u2__abc_52138_new_n12880_), .C(u2__abc_52138_new_n12882_), .Y(u2__abc_52138_new_n12883_));
OAI21X1 OAI21X1_3134 ( .A(u2__abc_52138_new_n3334_), .B(u2__abc_52138_new_n12871_), .C(u2__abc_52138_new_n12884_), .Y(u2__abc_52138_new_n12885_));
OAI21X1 OAI21X1_3135 ( .A(u2__abc_52138_new_n3835_), .B(u2__abc_52138_new_n3841_), .C(u2__abc_52138_new_n3840_), .Y(u2__abc_52138_new_n12891_));
OAI21X1 OAI21X1_3136 ( .A(u2__abc_52138_new_n3846_), .B(u2__abc_52138_new_n7212_), .C(u2__abc_52138_new_n3851_), .Y(u2__abc_52138_new_n12892_));
OAI21X1 OAI21X1_3137 ( .A(u2__abc_52138_new_n3865_), .B(u2__abc_52138_new_n12896_), .C(u2__abc_52138_new_n3884_), .Y(u2__abc_52138_new_n12897_));
OAI21X1 OAI21X1_3138 ( .A(u2__abc_52138_new_n12890_), .B(u2__abc_52138_new_n12893_), .C(u2__abc_52138_new_n12898_), .Y(u2__abc_52138_new_n12899_));
OAI21X1 OAI21X1_3139 ( .A(sqrto_71_), .B(u2__abc_52138_new_n3791_), .C(u2__abc_52138_new_n3789_), .Y(u2__abc_52138_new_n12900_));
OAI21X1 OAI21X1_314 ( .A(u2__abc_52138_new_n3950_), .B(u2__abc_52138_new_n3947_), .C(u2__abc_52138_new_n3953_), .Y(u2__abc_52138_new_n3954_));
OAI21X1 OAI21X1_3140 ( .A(u2__abc_52138_new_n3793_), .B(u2_remHi_71_), .C(u2__abc_52138_new_n12900_), .Y(u2__abc_52138_new_n12901_));
OAI21X1 OAI21X1_3141 ( .A(u2__abc_52138_new_n3800_), .B(u2__abc_52138_new_n7298_), .C(u2__abc_52138_new_n3805_), .Y(u2__abc_52138_new_n12902_));
OAI21X1 OAI21X1_3142 ( .A(u2__abc_52138_new_n3820_), .B(u2__abc_52138_new_n12904_), .C(u2__abc_52138_new_n7357_), .Y(u2__abc_52138_new_n12905_));
OAI21X1 OAI21X1_3143 ( .A(u2__abc_52138_new_n7355_), .B(u2__abc_52138_new_n12903_), .C(u2__abc_52138_new_n12907_), .Y(u2__abc_52138_new_n12908_));
OAI21X1 OAI21X1_3144 ( .A(u2__abc_52138_new_n3741_), .B(u2__abc_52138_new_n3747_), .C(u2__abc_52138_new_n3746_), .Y(u2__abc_52138_new_n12910_));
OAI21X1 OAI21X1_3145 ( .A(u2__abc_52138_new_n3752_), .B(u2__abc_52138_new_n7402_), .C(u2__abc_52138_new_n3757_), .Y(u2__abc_52138_new_n12911_));
OAI21X1 OAI21X1_3146 ( .A(u2__abc_52138_new_n3772_), .B(u2_remHi_83_), .C(u2__abc_52138_new_n3916_), .Y(u2__abc_52138_new_n12913_));
OAI21X1 OAI21X1_3147 ( .A(u2__abc_52138_new_n7447_), .B(u2__abc_52138_new_n12912_), .C(u2__abc_52138_new_n12914_), .Y(u2__abc_52138_new_n12915_));
OAI21X1 OAI21X1_3148 ( .A(sqrto_87_), .B(u2__abc_52138_new_n3724_), .C(u2__abc_52138_new_n3733_), .Y(u2__abc_52138_new_n12919_));
OAI21X1 OAI21X1_3149 ( .A(u2__abc_52138_new_n3727_), .B(u2_remHi_87_), .C(u2__abc_52138_new_n12919_), .Y(u2__abc_52138_new_n12920_));
OAI21X1 OAI21X1_315 ( .A(sqrto_103_), .B(u2__abc_52138_new_n3610_), .C(u2__abc_52138_new_n3615_), .Y(u2__abc_52138_new_n3956_));
OAI21X1 OAI21X1_3150 ( .A(u2__abc_52138_new_n12921_), .B(u2__abc_52138_new_n12917_), .C(u2__abc_52138_new_n12922_), .Y(u2__abc_52138_new_n12923_));
OAI21X1 OAI21X1_3151 ( .A(u2__abc_52138_new_n12888_), .B(u2__abc_52138_new_n12909_), .C(u2__abc_52138_new_n12924_), .Y(u2__abc_52138_new_n12925_));
OAI21X1 OAI21X1_3152 ( .A(u2__abc_52138_new_n3661_), .B(u2__abc_52138_new_n3657_), .C(u2__abc_52138_new_n3656_), .Y(u2__abc_52138_new_n12928_));
OAI21X1 OAI21X1_3153 ( .A(u2__abc_52138_new_n3684_), .B(u2__abc_52138_new_n3680_), .C(u2__abc_52138_new_n3679_), .Y(u2__abc_52138_new_n12930_));
OAI21X1 OAI21X1_3154 ( .A(u2__abc_52138_new_n7625_), .B(u2__abc_52138_new_n12929_), .C(u2__abc_52138_new_n12932_), .Y(u2__abc_52138_new_n12933_));
OAI21X1 OAI21X1_3155 ( .A(u2__abc_52138_new_n3608_), .B(u2_remHi_103_), .C(u2__abc_52138_new_n3956_), .Y(u2__abc_52138_new_n12935_));
OAI21X1 OAI21X1_3156 ( .A(u2__abc_52138_new_n3622_), .B(u2__abc_52138_new_n3966_), .C(u2__abc_52138_new_n3627_), .Y(u2__abc_52138_new_n12937_));
OAI21X1 OAI21X1_3157 ( .A(u2__abc_52138_new_n7714_), .B(u2__abc_52138_new_n12936_), .C(u2__abc_52138_new_n12938_), .Y(u2__abc_52138_new_n12939_));
OAI21X1 OAI21X1_3158 ( .A(u2__abc_52138_new_n3553_), .B(u2__abc_52138_new_n3559_), .C(u2__abc_52138_new_n3558_), .Y(u2__abc_52138_new_n12943_));
OAI21X1 OAI21X1_3159 ( .A(u2__abc_52138_new_n12942_), .B(u2__abc_52138_new_n12944_), .C(u2__abc_52138_new_n12945_), .Y(u2__abc_52138_new_n12946_));
OAI21X1 OAI21X1_316 ( .A(u2__abc_52138_new_n3600_), .B(u2__abc_52138_new_n3958_), .C(u2__abc_52138_new_n3605_), .Y(u2__abc_52138_new_n3959_));
OAI21X1 OAI21X1_3160 ( .A(u2__abc_52138_new_n3519_), .B(u2__abc_52138_new_n3525_), .C(u2__abc_52138_new_n3524_), .Y(u2__abc_52138_new_n12947_));
OAI21X1 OAI21X1_3161 ( .A(u2__abc_52138_new_n12948_), .B(u2__abc_52138_new_n6488_), .C(u2__abc_52138_new_n3996_), .Y(u2__abc_52138_new_n12949_));
OAI21X1 OAI21X1_3162 ( .A(u2__abc_52138_new_n7893_), .B(u2__abc_52138_new_n12940_), .C(u2__abc_52138_new_n12950_), .Y(u2__abc_52138_new_n12951_));
OAI21X1 OAI21X1_3163 ( .A(u2__abc_52138_new_n7888_), .B(u2__abc_52138_new_n12886_), .C(u2__abc_52138_new_n12952_), .Y(u2__abc_52138_new_n12953_));
OAI21X1 OAI21X1_3164 ( .A(u2__abc_52138_new_n4716_), .B(u2__abc_52138_new_n12955_), .C(u2__abc_52138_new_n4722_), .Y(u2__abc_52138_new_n12956_));
OAI21X1 OAI21X1_3165 ( .A(sqrto_129_), .B(u2__abc_52138_new_n4729_), .C(u2__abc_52138_new_n4771_), .Y(u2__abc_52138_new_n12957_));
OAI21X1 OAI21X1_3166 ( .A(u2__abc_52138_new_n4727_), .B(u2_remHi_129_), .C(u2__abc_52138_new_n12957_), .Y(u2__abc_52138_new_n12958_));
OAI21X1 OAI21X1_3167 ( .A(u2__abc_52138_new_n4750_), .B(u2__abc_52138_new_n12959_), .C(u2__abc_52138_new_n12960_), .Y(u2__abc_52138_new_n12961_));
OAI21X1 OAI21X1_3168 ( .A(u2__abc_52138_new_n4680_), .B(u2__abc_52138_new_n8007_), .C(u2__abc_52138_new_n4685_), .Y(u2__abc_52138_new_n12962_));
OAI21X1 OAI21X1_3169 ( .A(u2__abc_52138_new_n8070_), .B(u2__abc_52138_new_n12963_), .C(u2__abc_52138_new_n12964_), .Y(u2__abc_52138_new_n12965_));
OAI21X1 OAI21X1_317 ( .A(u2__abc_52138_new_n3957_), .B(u2__abc_52138_new_n3607_), .C(u2__abc_52138_new_n3960_), .Y(u2__abc_52138_new_n3961_));
OAI21X1 OAI21X1_3170 ( .A(sqrto_143_), .B(u2__abc_52138_new_n4652_), .C(u2__abc_52138_new_n4661_), .Y(u2__abc_52138_new_n12969_));
OAI21X1 OAI21X1_3171 ( .A(u2__abc_52138_new_n4655_), .B(u2_remHi_143_), .C(u2__abc_52138_new_n12969_), .Y(u2__abc_52138_new_n12970_));
OAI21X1 OAI21X1_3172 ( .A(u2__abc_52138_new_n4647_), .B(u2_remHi_145_), .C(u2__abc_52138_new_n4803_), .Y(u2__abc_52138_new_n12971_));
OAI21X1 OAI21X1_3173 ( .A(u2__abc_52138_new_n12967_), .B(u2__abc_52138_new_n12972_), .C(u2__abc_52138_new_n12974_), .Y(u2__abc_52138_new_n12975_));
OAI21X1 OAI21X1_3174 ( .A(u2__abc_52138_new_n4617_), .B(u2__abc_52138_new_n12976_), .C(u2__abc_52138_new_n12977_), .Y(u2__abc_52138_new_n12978_));
OAI21X1 OAI21X1_3175 ( .A(u2__abc_52138_new_n4665_), .B(u2__abc_52138_new_n12966_), .C(u2__abc_52138_new_n12979_), .Y(u2__abc_52138_new_n12980_));
OAI21X1 OAI21X1_3176 ( .A(u2__abc_52138_new_n12981_), .B(u2__abc_52138_new_n12983_), .C(u2__abc_52138_new_n12984_), .Y(u2__abc_52138_new_n12985_));
OAI21X1 OAI21X1_3177 ( .A(u2__abc_52138_new_n4481_), .B(u2__abc_52138_new_n8425_), .C(u2__abc_52138_new_n4486_), .Y(u2__abc_52138_new_n12987_));
OAI21X1 OAI21X1_3178 ( .A(u2__abc_52138_new_n4500_), .B(u2__abc_52138_new_n12986_), .C(u2__abc_52138_new_n12988_), .Y(u2__abc_52138_new_n12989_));
OAI21X1 OAI21X1_3179 ( .A(u2__abc_52138_new_n4477_), .B(u2__abc_52138_new_n12990_), .C(u2__abc_52138_new_n12991_), .Y(u2__abc_52138_new_n12992_));
OAI21X1 OAI21X1_318 ( .A(sqrto_107_), .B(u2__abc_52138_new_n3632_), .C(u2__abc_52138_new_n3637_), .Y(u2__abc_52138_new_n3963_));
OAI21X1 OAI21X1_3180 ( .A(sqrto_191_), .B(u2__abc_52138_new_n4369_), .C(u2__abc_52138_new_n4367_), .Y(u2__abc_52138_new_n12995_));
OAI21X1 OAI21X1_3181 ( .A(u2__abc_52138_new_n4372_), .B(u2_remHi_191_), .C(u2__abc_52138_new_n12995_), .Y(u2__abc_52138_new_n12996_));
OAI21X1 OAI21X1_3182 ( .A(u2__abc_52138_new_n6467_), .B(u2__abc_52138_new_n12998_), .C(u2__abc_52138_new_n12999_), .Y(u2__abc_52138_new_n13000_));
OAI21X1 OAI21X1_3183 ( .A(u2__abc_52138_new_n4315_), .B(u2__abc_52138_new_n4909_), .C(u2__abc_52138_new_n4320_), .Y(u2__abc_52138_new_n13002_));
OAI21X1 OAI21X1_3184 ( .A(u2__abc_52138_new_n4329_), .B(u2__abc_52138_new_n13001_), .C(u2__abc_52138_new_n13003_), .Y(u2__abc_52138_new_n13004_));
OAI21X1 OAI21X1_3185 ( .A(u2__abc_52138_new_n4255_), .B(u2__abc_52138_new_n4261_), .C(u2__abc_52138_new_n4260_), .Y(u2__abc_52138_new_n13007_));
OAI21X1 OAI21X1_3186 ( .A(sqrto_211_), .B(u2__abc_52138_new_n4275_), .C(u2__abc_52138_new_n4283_), .Y(u2__abc_52138_new_n13010_));
OAI21X1 OAI21X1_3187 ( .A(u2__abc_52138_new_n4277_), .B(u2_remHi_211_), .C(u2__abc_52138_new_n13010_), .Y(u2__abc_52138_new_n13011_));
OAI21X1 OAI21X1_3188 ( .A(u2__abc_52138_new_n13009_), .B(u2__abc_52138_new_n8854_), .C(u2__abc_52138_new_n13013_), .Y(u2__abc_52138_new_n13014_));
OAI21X1 OAI21X1_3189 ( .A(u2__abc_52138_new_n13015_), .B(u2__abc_52138_new_n8939_), .C(u2__abc_52138_new_n4939_), .Y(u2__abc_52138_new_n13016_));
OAI21X1 OAI21X1_319 ( .A(u2__abc_52138_new_n3630_), .B(u2_remHi_107_), .C(u2__abc_52138_new_n3963_), .Y(u2__abc_52138_new_n3964_));
OAI21X1 OAI21X1_3190 ( .A(u2__abc_52138_new_n12994_), .B(u2__abc_52138_new_n13005_), .C(u2__abc_52138_new_n13017_), .Y(u2__abc_52138_new_n13018_));
OAI21X1 OAI21X1_3191 ( .A(u2__abc_52138_new_n4190_), .B(u2__abc_52138_new_n13020_), .C(u2__abc_52138_new_n13021_), .Y(u2__abc_52138_new_n13022_));
OAI21X1 OAI21X1_3192 ( .A(u2__abc_52138_new_n4974_), .B(u2__abc_52138_new_n13024_), .C(u2__abc_52138_new_n4971_), .Y(u2__abc_52138_new_n13025_));
OAI21X1 OAI21X1_3193 ( .A(u2__abc_52138_new_n9269_), .B(u2__abc_52138_new_n13023_), .C(u2__abc_52138_new_n13027_), .Y(u2__abc_52138_new_n13028_));
OAI21X1 OAI21X1_3194 ( .A(u2__abc_52138_new_n9268_), .B(u2__abc_52138_new_n12993_), .C(u2__abc_52138_new_n13029_), .Y(u2__abc_52138_new_n13030_));
OAI21X1 OAI21X1_3195 ( .A(u2__abc_52138_new_n5546_), .B(u2__abc_52138_new_n13032_), .C(u2__abc_52138_new_n13033_), .Y(u2__abc_52138_new_n13034_));
OAI21X1 OAI21X1_3196 ( .A(u2__abc_52138_new_n10646_), .B(u2__abc_52138_new_n13031_), .C(u2__abc_52138_new_n13038_), .Y(u2__abc_52138_new_n13039_));
OAI21X1 OAI21X1_3197 ( .A(u2__abc_52138_new_n3014_), .B(u2__abc_52138_new_n13042_), .C(u2__abc_52138_new_n6450_), .Y(u2__abc_52138_new_n13043_));
OAI21X1 OAI21X1_3198 ( .A(u2__abc_52138_new_n13044_), .B(u2__abc_52138_new_n13045_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13046_));
OAI21X1 OAI21X1_3199 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_1_), .Y(u2__abc_52138_new_n13050_));
OAI21X1 OAI21X1_32 ( .A(aNan), .B(_abc_65734_new_n923_), .C(_abc_65734_new_n924_), .Y(\o[143] ));
OAI21X1 OAI21X1_320 ( .A(u2__abc_52138_new_n3641_), .B(u2__abc_52138_new_n3955_), .C(u2__abc_52138_new_n3969_), .Y(u2__abc_52138_new_n3970_));
OAI21X1 OAI21X1_3200 ( .A(u2__abc_52138_new_n13051_), .B(u2__abc_52138_new_n13052_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13053_));
OAI21X1 OAI21X1_3201 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_2_), .Y(u2__abc_52138_new_n13057_));
OAI21X1 OAI21X1_3202 ( .A(u2__abc_52138_new_n6541_), .B(u2__abc_52138_new_n6539_), .C(u2_root_0_), .Y(u2__abc_52138_new_n13059_));
OAI21X1 OAI21X1_3203 ( .A(u2__abc_52138_new_n13060_), .B(u2__abc_52138_new_n13058_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13061_));
OAI21X1 OAI21X1_3204 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_3_), .Y(u2__abc_52138_new_n13065_));
OAI21X1 OAI21X1_3205 ( .A(u2__abc_52138_new_n13066_), .B(u2__abc_52138_new_n13068_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13069_));
OAI21X1 OAI21X1_3206 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_4_), .Y(u2__abc_52138_new_n13073_));
OAI21X1 OAI21X1_3207 ( .A(u2__abc_52138_new_n13076_), .B(u2__abc_52138_new_n13074_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13077_));
OAI21X1 OAI21X1_3208 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_5_), .Y(u2__abc_52138_new_n13081_));
OAI21X1 OAI21X1_3209 ( .A(u2__abc_52138_new_n13083_), .B(u2__abc_52138_new_n13082_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13084_));
OAI21X1 OAI21X1_321 ( .A(u2__abc_52138_new_n3564_), .B(u2__abc_52138_new_n3975_), .C(u2__abc_52138_new_n3569_), .Y(u2__abc_52138_new_n3976_));
OAI21X1 OAI21X1_3210 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_6_), .Y(u2__abc_52138_new_n13088_));
OAI21X1 OAI21X1_3211 ( .A(u2__abc_52138_new_n13091_), .B(u2__abc_52138_new_n13089_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13092_));
OAI21X1 OAI21X1_3212 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_7_), .Y(u2__abc_52138_new_n13096_));
OAI21X1 OAI21X1_3213 ( .A(u2__abc_52138_new_n13097_), .B(u2__abc_52138_new_n13099_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13100_));
OAI21X1 OAI21X1_3214 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_8_), .Y(u2__abc_52138_new_n13104_));
OAI21X1 OAI21X1_3215 ( .A(u2__abc_52138_new_n13107_), .B(u2__abc_52138_new_n13105_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13108_));
OAI21X1 OAI21X1_3216 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_9_), .Y(u2__abc_52138_new_n13112_));
OAI21X1 OAI21X1_3217 ( .A(u2__abc_52138_new_n13114_), .B(u2__abc_52138_new_n13113_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13115_));
OAI21X1 OAI21X1_3218 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_10_), .Y(u2__abc_52138_new_n13119_));
OAI21X1 OAI21X1_3219 ( .A(u2__abc_52138_new_n13122_), .B(u2__abc_52138_new_n13120_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13123_));
OAI21X1 OAI21X1_322 ( .A(u2__abc_52138_new_n3974_), .B(u2__abc_52138_new_n3971_), .C(u2__abc_52138_new_n3977_), .Y(u2__abc_52138_new_n3978_));
OAI21X1 OAI21X1_3220 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_11_), .Y(u2__abc_52138_new_n13127_));
OAI21X1 OAI21X1_3221 ( .A(u2__abc_52138_new_n13128_), .B(u2__abc_52138_new_n13130_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13131_));
OAI21X1 OAI21X1_3222 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_12_), .Y(u2__abc_52138_new_n13135_));
OAI21X1 OAI21X1_3223 ( .A(u2__abc_52138_new_n13138_), .B(u2__abc_52138_new_n13136_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13139_));
OAI21X1 OAI21X1_3224 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_13_), .Y(u2__abc_52138_new_n13143_));
OAI21X1 OAI21X1_3225 ( .A(u2__abc_52138_new_n13145_), .B(u2__abc_52138_new_n13144_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13146_));
OAI21X1 OAI21X1_3226 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_14_), .Y(u2__abc_52138_new_n13150_));
OAI21X1 OAI21X1_3227 ( .A(u2__abc_52138_new_n13153_), .B(u2__abc_52138_new_n13151_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13154_));
OAI21X1 OAI21X1_3228 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_15_), .Y(u2__abc_52138_new_n13158_));
OAI21X1 OAI21X1_3229 ( .A(u2__abc_52138_new_n13159_), .B(u2__abc_52138_new_n13161_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13162_));
OAI21X1 OAI21X1_323 ( .A(sqrto_117_), .B(u2__abc_52138_new_n3580_), .C(u2__abc_52138_new_n3576_), .Y(u2__abc_52138_new_n3979_));
OAI21X1 OAI21X1_3230 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_16_), .Y(u2__abc_52138_new_n13166_));
OAI21X1 OAI21X1_3231 ( .A(u2__abc_52138_new_n13169_), .B(u2__abc_52138_new_n13167_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13170_));
OAI21X1 OAI21X1_3232 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_17_), .Y(u2__abc_52138_new_n13174_));
OAI21X1 OAI21X1_3233 ( .A(u2__abc_52138_new_n13176_), .B(u2__abc_52138_new_n13175_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13177_));
OAI21X1 OAI21X1_3234 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_18_), .Y(u2__abc_52138_new_n13181_));
OAI21X1 OAI21X1_3235 ( .A(u2__abc_52138_new_n13184_), .B(u2__abc_52138_new_n13182_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13185_));
OAI21X1 OAI21X1_3236 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_19_), .Y(u2__abc_52138_new_n13189_));
OAI21X1 OAI21X1_3237 ( .A(u2__abc_52138_new_n13190_), .B(u2__abc_52138_new_n13192_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13193_));
OAI21X1 OAI21X1_3238 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_20_), .Y(u2__abc_52138_new_n13197_));
OAI21X1 OAI21X1_3239 ( .A(u2__abc_52138_new_n13200_), .B(u2__abc_52138_new_n13198_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13201_));
OAI21X1 OAI21X1_324 ( .A(u2__abc_52138_new_n3578_), .B(u2_remHi_117_), .C(u2__abc_52138_new_n3979_), .Y(u2__abc_52138_new_n3980_));
OAI21X1 OAI21X1_3240 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_21_), .Y(u2__abc_52138_new_n13205_));
OAI21X1 OAI21X1_3241 ( .A(u2__abc_52138_new_n13207_), .B(u2__abc_52138_new_n13206_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13208_));
OAI21X1 OAI21X1_3242 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_22_), .Y(u2__abc_52138_new_n13212_));
OAI21X1 OAI21X1_3243 ( .A(u2__abc_52138_new_n13215_), .B(u2__abc_52138_new_n13213_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13216_));
OAI21X1 OAI21X1_3244 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_23_), .Y(u2__abc_52138_new_n13220_));
OAI21X1 OAI21X1_3245 ( .A(u2__abc_52138_new_n13221_), .B(u2__abc_52138_new_n13223_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13224_));
OAI21X1 OAI21X1_3246 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_24_), .Y(u2__abc_52138_new_n13228_));
OAI21X1 OAI21X1_3247 ( .A(u2__abc_52138_new_n13231_), .B(u2__abc_52138_new_n13229_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13232_));
OAI21X1 OAI21X1_3248 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_25_), .Y(u2__abc_52138_new_n13236_));
OAI21X1 OAI21X1_3249 ( .A(u2__abc_52138_new_n13238_), .B(u2__abc_52138_new_n13237_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13239_));
OAI21X1 OAI21X1_325 ( .A(u2__abc_52138_new_n3591_), .B(u2__abc_52138_new_n3982_), .C(u2__abc_52138_new_n3586_), .Y(u2__abc_52138_new_n3983_));
OAI21X1 OAI21X1_3250 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_26_), .Y(u2__abc_52138_new_n13243_));
OAI21X1 OAI21X1_3251 ( .A(u2__abc_52138_new_n13246_), .B(u2__abc_52138_new_n13244_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13247_));
OAI21X1 OAI21X1_3252 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_27_), .Y(u2__abc_52138_new_n13251_));
OAI21X1 OAI21X1_3253 ( .A(u2__abc_52138_new_n13252_), .B(u2__abc_52138_new_n13254_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13255_));
OAI21X1 OAI21X1_3254 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_28_), .Y(u2__abc_52138_new_n13259_));
OAI21X1 OAI21X1_3255 ( .A(u2__abc_52138_new_n13262_), .B(u2__abc_52138_new_n13260_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13263_));
OAI21X1 OAI21X1_3256 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_29_), .Y(u2__abc_52138_new_n13267_));
OAI21X1 OAI21X1_3257 ( .A(u2__abc_52138_new_n13269_), .B(u2__abc_52138_new_n13268_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13270_));
OAI21X1 OAI21X1_3258 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_30_), .Y(u2__abc_52138_new_n13274_));
OAI21X1 OAI21X1_3259 ( .A(u2__abc_52138_new_n13277_), .B(u2__abc_52138_new_n13275_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13278_));
OAI21X1 OAI21X1_326 ( .A(u2__abc_52138_new_n3984_), .B(u2__abc_52138_new_n3582_), .C(u2__abc_52138_new_n3981_), .Y(u2__abc_52138_new_n3985_));
OAI21X1 OAI21X1_3260 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_31_), .Y(u2__abc_52138_new_n13282_));
OAI21X1 OAI21X1_3261 ( .A(u2__abc_52138_new_n13283_), .B(u2__abc_52138_new_n13285_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13286_));
OAI21X1 OAI21X1_3262 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_32_), .Y(u2__abc_52138_new_n13290_));
OAI21X1 OAI21X1_3263 ( .A(u2__abc_52138_new_n13293_), .B(u2__abc_52138_new_n13291_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13294_));
OAI21X1 OAI21X1_3264 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_33_), .Y(u2__abc_52138_new_n13298_));
OAI21X1 OAI21X1_3265 ( .A(u2__abc_52138_new_n13300_), .B(u2__abc_52138_new_n13299_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13301_));
OAI21X1 OAI21X1_3266 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_34_), .Y(u2__abc_52138_new_n13305_));
OAI21X1 OAI21X1_3267 ( .A(u2__abc_52138_new_n13308_), .B(u2__abc_52138_new_n13306_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13309_));
OAI21X1 OAI21X1_3268 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_35_), .Y(u2__abc_52138_new_n13314_));
OAI21X1 OAI21X1_3269 ( .A(u2__abc_52138_new_n13315_), .B(u2__abc_52138_new_n13317_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13318_));
OAI21X1 OAI21X1_327 ( .A(u2__abc_52138_new_n3506_), .B(u2__abc_52138_new_n3509_), .C(u2__abc_52138_new_n3513_), .Y(u2__abc_52138_new_n3987_));
OAI21X1 OAI21X1_3270 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_36_), .Y(u2__abc_52138_new_n13322_));
OAI21X1 OAI21X1_3271 ( .A(u2__abc_52138_new_n13325_), .B(u2__abc_52138_new_n13323_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13326_));
OAI21X1 OAI21X1_3272 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_37_), .Y(u2__abc_52138_new_n13330_));
OAI21X1 OAI21X1_3273 ( .A(u2__abc_52138_new_n13332_), .B(u2__abc_52138_new_n13331_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13333_));
OAI21X1 OAI21X1_3274 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_38_), .Y(u2__abc_52138_new_n13337_));
OAI21X1 OAI21X1_3275 ( .A(u2__abc_52138_new_n13340_), .B(u2__abc_52138_new_n13338_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13341_));
OAI21X1 OAI21X1_3276 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_39_), .Y(u2__abc_52138_new_n13345_));
OAI21X1 OAI21X1_3277 ( .A(u2__abc_52138_new_n13346_), .B(u2__abc_52138_new_n13348_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13349_));
OAI21X1 OAI21X1_3278 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_40_), .Y(u2__abc_52138_new_n13353_));
OAI21X1 OAI21X1_3279 ( .A(u2__abc_52138_new_n13356_), .B(u2__abc_52138_new_n13354_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13357_));
OAI21X1 OAI21X1_328 ( .A(u2__abc_52138_new_n3530_), .B(u2__abc_52138_new_n3992_), .C(u2__abc_52138_new_n3533_), .Y(u2__abc_52138_new_n3993_));
OAI21X1 OAI21X1_3280 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_41_), .Y(u2__abc_52138_new_n13361_));
OAI21X1 OAI21X1_3281 ( .A(u2__abc_52138_new_n13363_), .B(u2__abc_52138_new_n13362_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13364_));
OAI21X1 OAI21X1_3282 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_42_), .Y(u2__abc_52138_new_n13368_));
OAI21X1 OAI21X1_3283 ( .A(u2__abc_52138_new_n13371_), .B(u2__abc_52138_new_n13369_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13372_));
OAI21X1 OAI21X1_3284 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_43_), .Y(u2__abc_52138_new_n13376_));
OAI21X1 OAI21X1_3285 ( .A(u2__abc_52138_new_n13377_), .B(u2__abc_52138_new_n13379_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13380_));
OAI21X1 OAI21X1_3286 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_44_), .Y(u2__abc_52138_new_n13384_));
OAI21X1 OAI21X1_3287 ( .A(u2__abc_52138_new_n13387_), .B(u2__abc_52138_new_n13385_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13388_));
OAI21X1 OAI21X1_3288 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_45_), .Y(u2__abc_52138_new_n13392_));
OAI21X1 OAI21X1_3289 ( .A(u2__abc_52138_new_n13394_), .B(u2__abc_52138_new_n13393_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13395_));
OAI21X1 OAI21X1_329 ( .A(sqrto_123_), .B(u2__abc_52138_new_n3540_), .C(u2__abc_52138_new_n3545_), .Y(u2__abc_52138_new_n3994_));
OAI21X1 OAI21X1_3290 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_46_), .Y(u2__abc_52138_new_n13399_));
OAI21X1 OAI21X1_3291 ( .A(u2__abc_52138_new_n13402_), .B(u2__abc_52138_new_n13400_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13403_));
OAI21X1 OAI21X1_3292 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_47_), .Y(u2__abc_52138_new_n13407_));
OAI21X1 OAI21X1_3293 ( .A(u2__abc_52138_new_n13408_), .B(u2__abc_52138_new_n13410_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13411_));
OAI21X1 OAI21X1_3294 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_48_), .Y(u2__abc_52138_new_n13415_));
OAI21X1 OAI21X1_3295 ( .A(u2__abc_52138_new_n13418_), .B(u2__abc_52138_new_n13416_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13419_));
OAI21X1 OAI21X1_3296 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_49_), .Y(u2__abc_52138_new_n13423_));
OAI21X1 OAI21X1_3297 ( .A(u2__abc_52138_new_n13425_), .B(u2__abc_52138_new_n13424_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13426_));
OAI21X1 OAI21X1_3298 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_50_), .Y(u2__abc_52138_new_n13430_));
OAI21X1 OAI21X1_3299 ( .A(u2__abc_52138_new_n13433_), .B(u2__abc_52138_new_n13431_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13434_));
OAI21X1 OAI21X1_33 ( .A(aNan), .B(_abc_65734_new_n926_), .C(_abc_65734_new_n927_), .Y(\o[144] ));
OAI21X1 OAI21X1_330 ( .A(u2__abc_52138_new_n3538_), .B(u2_remHi_123_), .C(u2__abc_52138_new_n3994_), .Y(u2__abc_52138_new_n3995_));
OAI21X1 OAI21X1_3300 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_51_), .Y(u2__abc_52138_new_n13438_));
OAI21X1 OAI21X1_3301 ( .A(u2__abc_52138_new_n13439_), .B(u2__abc_52138_new_n13441_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13442_));
OAI21X1 OAI21X1_3302 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_52_), .Y(u2__abc_52138_new_n13446_));
OAI21X1 OAI21X1_3303 ( .A(u2__abc_52138_new_n13449_), .B(u2__abc_52138_new_n13447_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13450_));
OAI21X1 OAI21X1_3304 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_53_), .Y(u2__abc_52138_new_n13454_));
OAI21X1 OAI21X1_3305 ( .A(u2__abc_52138_new_n13456_), .B(u2__abc_52138_new_n13455_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13457_));
OAI21X1 OAI21X1_3306 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_54_), .Y(u2__abc_52138_new_n13461_));
OAI21X1 OAI21X1_3307 ( .A(u2__abc_52138_new_n13464_), .B(u2__abc_52138_new_n13462_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13465_));
OAI21X1 OAI21X1_3308 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_55_), .Y(u2__abc_52138_new_n13469_));
OAI21X1 OAI21X1_3309 ( .A(u2__abc_52138_new_n13470_), .B(u2__abc_52138_new_n13472_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13473_));
OAI21X1 OAI21X1_331 ( .A(u2__abc_52138_new_n3549_), .B(u2__abc_52138_new_n3986_), .C(u2__abc_52138_new_n3998_), .Y(u2__abc_52138_new_n3999_));
OAI21X1 OAI21X1_3310 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_56_), .Y(u2__abc_52138_new_n13477_));
OAI21X1 OAI21X1_3311 ( .A(u2__abc_52138_new_n13480_), .B(u2__abc_52138_new_n13478_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13481_));
OAI21X1 OAI21X1_3312 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_57_), .Y(u2__abc_52138_new_n13485_));
OAI21X1 OAI21X1_3313 ( .A(u2__abc_52138_new_n13487_), .B(u2__abc_52138_new_n13486_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13488_));
OAI21X1 OAI21X1_3314 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_58_), .Y(u2__abc_52138_new_n13492_));
OAI21X1 OAI21X1_3315 ( .A(u2__abc_52138_new_n13495_), .B(u2__abc_52138_new_n13493_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13496_));
OAI21X1 OAI21X1_3316 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_59_), .Y(u2__abc_52138_new_n13500_));
OAI21X1 OAI21X1_3317 ( .A(u2__abc_52138_new_n13501_), .B(u2__abc_52138_new_n13503_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13504_));
OAI21X1 OAI21X1_3318 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_60_), .Y(u2__abc_52138_new_n13508_));
OAI21X1 OAI21X1_3319 ( .A(u2__abc_52138_new_n13511_), .B(u2__abc_52138_new_n13509_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13512_));
OAI21X1 OAI21X1_332 ( .A(u2__abc_52138_new_n3690_), .B(u2__abc_52138_new_n3938_), .C(u2__abc_52138_new_n4000_), .Y(u2__abc_52138_new_n4001_));
OAI21X1 OAI21X1_3320 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_61_), .Y(u2__abc_52138_new_n13516_));
OAI21X1 OAI21X1_3321 ( .A(u2__abc_52138_new_n13518_), .B(u2__abc_52138_new_n13517_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13519_));
OAI21X1 OAI21X1_3322 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_62_), .Y(u2__abc_52138_new_n13523_));
OAI21X1 OAI21X1_3323 ( .A(u2__abc_52138_new_n13526_), .B(u2__abc_52138_new_n13524_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13527_));
OAI21X1 OAI21X1_3324 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_63_), .Y(u2__abc_52138_new_n13531_));
OAI21X1 OAI21X1_3325 ( .A(u2__abc_52138_new_n13532_), .B(u2__abc_52138_new_n13534_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13535_));
OAI21X1 OAI21X1_3326 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_64_), .Y(u2__abc_52138_new_n13539_));
OAI21X1 OAI21X1_3327 ( .A(u2__abc_52138_new_n13542_), .B(u2__abc_52138_new_n13540_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13543_));
OAI21X1 OAI21X1_3328 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_65_), .Y(u2__abc_52138_new_n13547_));
OAI21X1 OAI21X1_3329 ( .A(u2__abc_52138_new_n13549_), .B(u2__abc_52138_new_n13548_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13550_));
OAI21X1 OAI21X1_333 ( .A(u2__abc_52138_new_n4731_), .B(u2__abc_52138_new_n4769_), .C(u2__abc_52138_new_n4773_), .Y(u2__abc_52138_new_n4774_));
OAI21X1 OAI21X1_3330 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_66_), .Y(u2__abc_52138_new_n13554_));
OAI21X1 OAI21X1_3331 ( .A(u2__abc_52138_new_n13557_), .B(u2__abc_52138_new_n13555_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13558_));
OAI21X1 OAI21X1_3332 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_67_), .Y(u2__abc_52138_new_n13562_));
OAI21X1 OAI21X1_3333 ( .A(u2__abc_52138_new_n13563_), .B(u2__abc_52138_new_n13565_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13566_));
OAI21X1 OAI21X1_3334 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_68_), .Y(u2__abc_52138_new_n13570_));
OAI21X1 OAI21X1_3335 ( .A(u2__abc_52138_new_n13573_), .B(u2__abc_52138_new_n13571_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13574_));
OAI21X1 OAI21X1_3336 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_69_), .Y(u2__abc_52138_new_n13578_));
OAI21X1 OAI21X1_3337 ( .A(u2__abc_52138_new_n13580_), .B(u2__abc_52138_new_n13579_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13581_));
OAI21X1 OAI21X1_3338 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_70_), .Y(u2__abc_52138_new_n13585_));
OAI21X1 OAI21X1_3339 ( .A(u2__abc_52138_new_n13588_), .B(u2__abc_52138_new_n13586_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13589_));
OAI21X1 OAI21X1_334 ( .A(u2__abc_52138_new_n4777_), .B(u2__abc_52138_new_n4775_), .C(u2__abc_52138_new_n4747_), .Y(u2__abc_52138_new_n4778_));
OAI21X1 OAI21X1_3340 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_71_), .Y(u2__abc_52138_new_n13593_));
OAI21X1 OAI21X1_3341 ( .A(u2__abc_52138_new_n13594_), .B(u2__abc_52138_new_n13596_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13597_));
OAI21X1 OAI21X1_3342 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_72_), .Y(u2__abc_52138_new_n13601_));
OAI21X1 OAI21X1_3343 ( .A(u2__abc_52138_new_n13604_), .B(u2__abc_52138_new_n13602_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13605_));
OAI21X1 OAI21X1_3344 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_73_), .Y(u2__abc_52138_new_n13609_));
OAI21X1 OAI21X1_3345 ( .A(u2__abc_52138_new_n13611_), .B(u2__abc_52138_new_n13610_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13612_));
OAI21X1 OAI21X1_3346 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_74_), .Y(u2__abc_52138_new_n13616_));
OAI21X1 OAI21X1_3347 ( .A(u2__abc_52138_new_n13619_), .B(u2__abc_52138_new_n13617_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13620_));
OAI21X1 OAI21X1_3348 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_75_), .Y(u2__abc_52138_new_n13624_));
OAI21X1 OAI21X1_3349 ( .A(u2__abc_52138_new_n13625_), .B(u2__abc_52138_new_n13627_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13628_));
OAI21X1 OAI21X1_335 ( .A(u2__abc_52138_new_n4736_), .B(u2__abc_52138_new_n4780_), .C(u2__abc_52138_new_n4741_), .Y(u2__abc_52138_new_n4781_));
OAI21X1 OAI21X1_3350 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_76_), .Y(u2__abc_52138_new_n13632_));
OAI21X1 OAI21X1_3351 ( .A(u2__abc_52138_new_n13635_), .B(u2__abc_52138_new_n13633_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13636_));
OAI21X1 OAI21X1_3352 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_77_), .Y(u2__abc_52138_new_n13640_));
OAI21X1 OAI21X1_3353 ( .A(u2__abc_52138_new_n13642_), .B(u2__abc_52138_new_n13641_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13643_));
OAI21X1 OAI21X1_3354 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_78_), .Y(u2__abc_52138_new_n13647_));
OAI21X1 OAI21X1_3355 ( .A(u2__abc_52138_new_n13650_), .B(u2__abc_52138_new_n13648_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13651_));
OAI21X1 OAI21X1_3356 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_79_), .Y(u2__abc_52138_new_n13655_));
OAI21X1 OAI21X1_3357 ( .A(u2__abc_52138_new_n13656_), .B(u2__abc_52138_new_n13658_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13659_));
OAI21X1 OAI21X1_3358 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_80_), .Y(u2__abc_52138_new_n13663_));
OAI21X1 OAI21X1_3359 ( .A(u2__abc_52138_new_n13665_), .B(u2__abc_52138_new_n13666_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13667_));
OAI21X1 OAI21X1_336 ( .A(u2__abc_52138_new_n4764_), .B(u2__abc_52138_new_n4779_), .C(u2__abc_52138_new_n4782_), .Y(u2__abc_52138_new_n4783_));
OAI21X1 OAI21X1_3360 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_81_), .Y(u2__abc_52138_new_n13671_));
OAI21X1 OAI21X1_3361 ( .A(u2__abc_52138_new_n13673_), .B(u2__abc_52138_new_n13672_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13674_));
OAI21X1 OAI21X1_3362 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_82_), .Y(u2__abc_52138_new_n13678_));
OAI21X1 OAI21X1_3363 ( .A(u2__abc_52138_new_n13681_), .B(u2__abc_52138_new_n13679_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13682_));
OAI21X1 OAI21X1_3364 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_83_), .Y(u2__abc_52138_new_n13686_));
OAI21X1 OAI21X1_3365 ( .A(u2__abc_52138_new_n13687_), .B(u2__abc_52138_new_n13689_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13690_));
OAI21X1 OAI21X1_3366 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_84_), .Y(u2__abc_52138_new_n13694_));
OAI21X1 OAI21X1_3367 ( .A(u2__abc_52138_new_n13697_), .B(u2__abc_52138_new_n13695_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13698_));
OAI21X1 OAI21X1_3368 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_85_), .Y(u2__abc_52138_new_n13702_));
OAI21X1 OAI21X1_3369 ( .A(u2__abc_52138_new_n13704_), .B(u2__abc_52138_new_n13703_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13705_));
OAI21X1 OAI21X1_337 ( .A(u2__abc_52138_new_n4669_), .B(u2__abc_52138_new_n4789_), .C(u2__abc_52138_new_n4674_), .Y(u2__abc_52138_new_n4790_));
OAI21X1 OAI21X1_3370 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_86_), .Y(u2__abc_52138_new_n13709_));
OAI21X1 OAI21X1_3371 ( .A(u2__abc_52138_new_n13712_), .B(u2__abc_52138_new_n13710_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13713_));
OAI21X1 OAI21X1_3372 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_87_), .Y(u2__abc_52138_new_n13717_));
OAI21X1 OAI21X1_3373 ( .A(u2__abc_52138_new_n13718_), .B(u2__abc_52138_new_n13720_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13721_));
OAI21X1 OAI21X1_3374 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_88_), .Y(u2__abc_52138_new_n13725_));
OAI21X1 OAI21X1_3375 ( .A(u2__abc_52138_new_n13727_), .B(u2__abc_52138_new_n13728_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13729_));
OAI21X1 OAI21X1_3376 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_89_), .Y(u2__abc_52138_new_n13733_));
OAI21X1 OAI21X1_3377 ( .A(u2__abc_52138_new_n13735_), .B(u2__abc_52138_new_n13734_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13736_));
OAI21X1 OAI21X1_3378 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_90_), .Y(u2__abc_52138_new_n13740_));
OAI21X1 OAI21X1_3379 ( .A(u2__abc_52138_new_n13743_), .B(u2__abc_52138_new_n13741_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13744_));
OAI21X1 OAI21X1_338 ( .A(u2__abc_52138_new_n4788_), .B(u2__abc_52138_new_n4785_), .C(u2__abc_52138_new_n4791_), .Y(u2__abc_52138_new_n4792_));
OAI21X1 OAI21X1_3380 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_91_), .Y(u2__abc_52138_new_n13748_));
OAI21X1 OAI21X1_3381 ( .A(u2__abc_52138_new_n13749_), .B(u2__abc_52138_new_n13751_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13752_));
OAI21X1 OAI21X1_3382 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_92_), .Y(u2__abc_52138_new_n13756_));
OAI21X1 OAI21X1_3383 ( .A(u2__abc_52138_new_n13758_), .B(u2__abc_52138_new_n13759_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13760_));
OAI21X1 OAI21X1_3384 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_93_), .Y(u2__abc_52138_new_n13764_));
OAI21X1 OAI21X1_3385 ( .A(u2__abc_52138_new_n13766_), .B(u2__abc_52138_new_n13765_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13767_));
OAI21X1 OAI21X1_3386 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_94_), .Y(u2__abc_52138_new_n13771_));
OAI21X1 OAI21X1_3387 ( .A(u2__abc_52138_new_n13773_), .B(u2__abc_52138_new_n13774_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13775_));
OAI21X1 OAI21X1_3388 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_95_), .Y(u2__abc_52138_new_n13779_));
OAI21X1 OAI21X1_3389 ( .A(u2__abc_52138_new_n13780_), .B(u2__abc_52138_new_n13782_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13783_));
OAI21X1 OAI21X1_339 ( .A(u2__abc_52138_new_n4708_), .B(u2__abc_52138_new_n4793_), .C(u2__abc_52138_new_n4703_), .Y(u2__abc_52138_new_n4794_));
OAI21X1 OAI21X1_3390 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_96_), .Y(u2__abc_52138_new_n13787_));
OAI21X1 OAI21X1_3391 ( .A(u2__abc_52138_new_n13790_), .B(u2__abc_52138_new_n13788_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13791_));
OAI21X1 OAI21X1_3392 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_97_), .Y(u2__abc_52138_new_n13795_));
OAI21X1 OAI21X1_3393 ( .A(u2__abc_52138_new_n13797_), .B(u2__abc_52138_new_n13796_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13798_));
OAI21X1 OAI21X1_3394 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_98_), .Y(u2__abc_52138_new_n13802_));
OAI21X1 OAI21X1_3395 ( .A(u2__abc_52138_new_n13805_), .B(u2__abc_52138_new_n13803_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13806_));
OAI21X1 OAI21X1_3396 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_99_), .Y(u2__abc_52138_new_n13810_));
OAI21X1 OAI21X1_3397 ( .A(u2__abc_52138_new_n13811_), .B(u2__abc_52138_new_n13813_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13814_));
OAI21X1 OAI21X1_3398 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_100_), .Y(u2__abc_52138_new_n13818_));
OAI21X1 OAI21X1_3399 ( .A(u2__abc_52138_new_n13821_), .B(u2__abc_52138_new_n13819_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13822_));
OAI21X1 OAI21X1_34 ( .A(aNan), .B(_abc_65734_new_n929_), .C(_abc_65734_new_n930_), .Y(\o[145] ));
OAI21X1 OAI21X1_340 ( .A(u2__abc_52138_new_n4692_), .B(u2__abc_52138_new_n4698_), .C(u2__abc_52138_new_n4697_), .Y(u2__abc_52138_new_n4796_));
OAI21X1 OAI21X1_3400 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_101_), .Y(u2__abc_52138_new_n13826_));
OAI21X1 OAI21X1_3401 ( .A(u2__abc_52138_new_n13828_), .B(u2__abc_52138_new_n13827_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13829_));
OAI21X1 OAI21X1_3402 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_102_), .Y(u2__abc_52138_new_n13833_));
OAI21X1 OAI21X1_3403 ( .A(u2__abc_52138_new_n13836_), .B(u2__abc_52138_new_n13834_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13837_));
OAI21X1 OAI21X1_3404 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_103_), .Y(u2__abc_52138_new_n13841_));
OAI21X1 OAI21X1_3405 ( .A(u2__abc_52138_new_n13842_), .B(u2__abc_52138_new_n13844_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13845_));
OAI21X1 OAI21X1_3406 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_104_), .Y(u2__abc_52138_new_n13849_));
OAI21X1 OAI21X1_3407 ( .A(u2__abc_52138_new_n13851_), .B(u2__abc_52138_new_n13852_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13853_));
OAI21X1 OAI21X1_3408 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_105_), .Y(u2__abc_52138_new_n13857_));
OAI21X1 OAI21X1_3409 ( .A(u2__abc_52138_new_n13859_), .B(u2__abc_52138_new_n13858_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13860_));
OAI21X1 OAI21X1_341 ( .A(u2__abc_52138_new_n4712_), .B(u2__abc_52138_new_n4784_), .C(u2__abc_52138_new_n4799_), .Y(u2__abc_52138_new_n4800_));
OAI21X1 OAI21X1_3410 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_106_), .Y(u2__abc_52138_new_n13864_));
OAI21X1 OAI21X1_3411 ( .A(u2__abc_52138_new_n13867_), .B(u2__abc_52138_new_n13865_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13868_));
OAI21X1 OAI21X1_3412 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_107_), .Y(u2__abc_52138_new_n13872_));
OAI21X1 OAI21X1_3413 ( .A(u2__abc_52138_new_n13873_), .B(u2__abc_52138_new_n13875_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13876_));
OAI21X1 OAI21X1_3414 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_108_), .Y(u2__abc_52138_new_n13880_));
OAI21X1 OAI21X1_3415 ( .A(u2__abc_52138_new_n13882_), .B(u2__abc_52138_new_n13883_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13884_));
OAI21X1 OAI21X1_3416 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_109_), .Y(u2__abc_52138_new_n13888_));
OAI21X1 OAI21X1_3417 ( .A(u2__abc_52138_new_n13890_), .B(u2__abc_52138_new_n13889_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13891_));
OAI21X1 OAI21X1_3418 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_110_), .Y(u2__abc_52138_new_n13895_));
OAI21X1 OAI21X1_3419 ( .A(u2__abc_52138_new_n13897_), .B(u2__abc_52138_new_n13898_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13899_));
OAI21X1 OAI21X1_342 ( .A(sqrto_145_), .B(u2__abc_52138_new_n4649_), .C(u2__abc_52138_new_n4802_), .Y(u2__abc_52138_new_n4803_));
OAI21X1 OAI21X1_3420 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_111_), .Y(u2__abc_52138_new_n13903_));
OAI21X1 OAI21X1_3421 ( .A(u2__abc_52138_new_n13904_), .B(u2__abc_52138_new_n13906_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13907_));
OAI21X1 OAI21X1_3422 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_112_), .Y(u2__abc_52138_new_n13911_));
OAI21X1 OAI21X1_3423 ( .A(u2__abc_52138_new_n13914_), .B(u2__abc_52138_new_n13912_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13915_));
OAI21X1 OAI21X1_3424 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_113_), .Y(u2__abc_52138_new_n13919_));
OAI21X1 OAI21X1_3425 ( .A(u2__abc_52138_new_n13921_), .B(u2__abc_52138_new_n13920_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13922_));
OAI21X1 OAI21X1_3426 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_114_), .Y(u2__abc_52138_new_n13926_));
OAI21X1 OAI21X1_3427 ( .A(u2__abc_52138_new_n13929_), .B(u2__abc_52138_new_n13927_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13930_));
OAI21X1 OAI21X1_3428 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_115_), .Y(u2__abc_52138_new_n13934_));
OAI21X1 OAI21X1_3429 ( .A(u2__abc_52138_new_n13935_), .B(u2__abc_52138_new_n13937_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13938_));
OAI21X1 OAI21X1_343 ( .A(u2__abc_52138_new_n4801_), .B(u2__abc_52138_new_n4651_), .C(u2__abc_52138_new_n4804_), .Y(u2__abc_52138_new_n4805_));
OAI21X1 OAI21X1_3430 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_116_), .Y(u2__abc_52138_new_n13942_));
OAI21X1 OAI21X1_3431 ( .A(u2__abc_52138_new_n13944_), .B(u2__abc_52138_new_n13945_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13946_));
OAI21X1 OAI21X1_3432 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_117_), .Y(u2__abc_52138_new_n13950_));
OAI21X1 OAI21X1_3433 ( .A(u2__abc_52138_new_n13952_), .B(u2__abc_52138_new_n13951_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13953_));
OAI21X1 OAI21X1_3434 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_118_), .Y(u2__abc_52138_new_n13957_));
OAI21X1 OAI21X1_3435 ( .A(u2__abc_52138_new_n13959_), .B(u2__abc_52138_new_n13960_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13961_));
OAI21X1 OAI21X1_3436 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_119_), .Y(u2__abc_52138_new_n13966_));
OAI21X1 OAI21X1_3437 ( .A(u2__abc_52138_new_n13967_), .B(u2__abc_52138_new_n13969_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13970_));
OAI21X1 OAI21X1_3438 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_120_), .Y(u2__abc_52138_new_n13974_));
OAI21X1 OAI21X1_3439 ( .A(u2__abc_52138_new_n13977_), .B(u2__abc_52138_new_n13975_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13978_));
OAI21X1 OAI21X1_344 ( .A(u2__abc_52138_new_n4638_), .B(u2__abc_52138_new_n4807_), .C(u2__abc_52138_new_n4633_), .Y(u2__abc_52138_new_n4808_));
OAI21X1 OAI21X1_3440 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_121_), .Y(u2__abc_52138_new_n13982_));
OAI21X1 OAI21X1_3441 ( .A(u2__abc_52138_new_n13984_), .B(u2__abc_52138_new_n13983_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13985_));
OAI21X1 OAI21X1_3442 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_122_), .Y(u2__abc_52138_new_n13989_));
OAI21X1 OAI21X1_3443 ( .A(u2__abc_52138_new_n13991_), .B(u2__abc_52138_new_n13992_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n13993_));
OAI21X1 OAI21X1_3444 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_123_), .Y(u2__abc_52138_new_n13997_));
OAI21X1 OAI21X1_3445 ( .A(u2__abc_52138_new_n13998_), .B(u2__abc_52138_new_n14000_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14001_));
OAI21X1 OAI21X1_3446 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_124_), .Y(u2__abc_52138_new_n14005_));
OAI21X1 OAI21X1_3447 ( .A(u2__abc_52138_new_n14008_), .B(u2__abc_52138_new_n14006_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14009_));
OAI21X1 OAI21X1_3448 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_125_), .Y(u2__abc_52138_new_n14013_));
OAI21X1 OAI21X1_3449 ( .A(u2__abc_52138_new_n14015_), .B(u2__abc_52138_new_n14014_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14016_));
OAI21X1 OAI21X1_345 ( .A(u2__abc_52138_new_n4809_), .B(u2__abc_52138_new_n4806_), .C(u2__abc_52138_new_n4812_), .Y(u2__abc_52138_new_n4813_));
OAI21X1 OAI21X1_3450 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_126_), .Y(u2__abc_52138_new_n14020_));
OAI21X1 OAI21X1_3451 ( .A(u2__abc_52138_new_n14022_), .B(u2__abc_52138_new_n14023_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14024_));
OAI21X1 OAI21X1_3452 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_127_), .Y(u2__abc_52138_new_n14028_));
OAI21X1 OAI21X1_3453 ( .A(u2__abc_52138_new_n14029_), .B(u2__abc_52138_new_n14031_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14032_));
OAI21X1 OAI21X1_3454 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_128_), .Y(u2__abc_52138_new_n14036_));
OAI21X1 OAI21X1_3455 ( .A(u2__abc_52138_new_n14039_), .B(u2__abc_52138_new_n14037_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14040_));
OAI21X1 OAI21X1_3456 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_129_), .Y(u2__abc_52138_new_n14044_));
OAI21X1 OAI21X1_3457 ( .A(u2__abc_52138_new_n14046_), .B(u2__abc_52138_new_n14045_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14047_));
OAI21X1 OAI21X1_3458 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_130_), .Y(u2__abc_52138_new_n14051_));
OAI21X1 OAI21X1_3459 ( .A(u2__abc_52138_new_n14054_), .B(u2__abc_52138_new_n14052_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14055_));
OAI21X1 OAI21X1_346 ( .A(u2__abc_52138_new_n4592_), .B(u2__abc_52138_new_n4816_), .C(u2__abc_52138_new_n4587_), .Y(u2__abc_52138_new_n4817_));
OAI21X1 OAI21X1_3460 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_131_), .Y(u2__abc_52138_new_n14060_));
OAI21X1 OAI21X1_3461 ( .A(u2__abc_52138_new_n14061_), .B(u2__abc_52138_new_n14063_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14064_));
OAI21X1 OAI21X1_3462 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_132_), .Y(u2__abc_52138_new_n14068_));
OAI21X1 OAI21X1_3463 ( .A(u2__abc_52138_new_n14071_), .B(u2__abc_52138_new_n14069_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14072_));
OAI21X1 OAI21X1_3464 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_133_), .Y(u2__abc_52138_new_n14076_));
OAI21X1 OAI21X1_3465 ( .A(u2__abc_52138_new_n14078_), .B(u2__abc_52138_new_n14077_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14079_));
OAI21X1 OAI21X1_3466 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_134_), .Y(u2__abc_52138_new_n14083_));
OAI21X1 OAI21X1_3467 ( .A(u2__abc_52138_new_n14086_), .B(u2__abc_52138_new_n14084_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14087_));
OAI21X1 OAI21X1_3468 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_135_), .Y(u2__abc_52138_new_n14091_));
OAI21X1 OAI21X1_3469 ( .A(u2__abc_52138_new_n14092_), .B(u2__abc_52138_new_n14094_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14095_));
OAI21X1 OAI21X1_347 ( .A(u2__abc_52138_new_n4576_), .B(u2__abc_52138_new_n4582_), .C(u2__abc_52138_new_n4581_), .Y(u2__abc_52138_new_n4819_));
OAI21X1 OAI21X1_3470 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_136_), .Y(u2__abc_52138_new_n14099_));
OAI21X1 OAI21X1_3471 ( .A(u2__abc_52138_new_n14101_), .B(u2__abc_52138_new_n14102_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14103_));
OAI21X1 OAI21X1_3472 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_137_), .Y(u2__abc_52138_new_n14107_));
OAI21X1 OAI21X1_3473 ( .A(u2__abc_52138_new_n14109_), .B(u2__abc_52138_new_n14108_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14110_));
OAI21X1 OAI21X1_3474 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_138_), .Y(u2__abc_52138_new_n14114_));
OAI21X1 OAI21X1_3475 ( .A(u2__abc_52138_new_n14117_), .B(u2__abc_52138_new_n14115_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14118_));
OAI21X1 OAI21X1_3476 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_139_), .Y(u2__abc_52138_new_n14122_));
OAI21X1 OAI21X1_3477 ( .A(u2__abc_52138_new_n14123_), .B(u2__abc_52138_new_n14125_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14126_));
OAI21X1 OAI21X1_3478 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_140_), .Y(u2__abc_52138_new_n14130_));
OAI21X1 OAI21X1_3479 ( .A(u2__abc_52138_new_n14132_), .B(u2__abc_52138_new_n14133_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14134_));
OAI21X1 OAI21X1_348 ( .A(sqrto_155_), .B(u2__abc_52138_new_n4607_), .C(u2__abc_52138_new_n4615_), .Y(u2__abc_52138_new_n4822_));
OAI21X1 OAI21X1_3480 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_141_), .Y(u2__abc_52138_new_n14138_));
OAI21X1 OAI21X1_3481 ( .A(u2__abc_52138_new_n14140_), .B(u2__abc_52138_new_n14139_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14141_));
OAI21X1 OAI21X1_3482 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_142_), .Y(u2__abc_52138_new_n14145_));
OAI21X1 OAI21X1_3483 ( .A(u2__abc_52138_new_n14147_), .B(u2__abc_52138_new_n14148_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14149_));
OAI21X1 OAI21X1_3484 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_143_), .Y(u2__abc_52138_new_n14153_));
OAI21X1 OAI21X1_3485 ( .A(u2__abc_52138_new_n14154_), .B(u2__abc_52138_new_n14156_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14157_));
OAI21X1 OAI21X1_3486 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_144_), .Y(u2__abc_52138_new_n14161_));
OAI21X1 OAI21X1_3487 ( .A(u2__abc_52138_new_n14164_), .B(u2__abc_52138_new_n14162_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14165_));
OAI21X1 OAI21X1_3488 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_145_), .Y(u2__abc_52138_new_n14169_));
OAI21X1 OAI21X1_3489 ( .A(u2__abc_52138_new_n14171_), .B(u2__abc_52138_new_n14170_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14172_));
OAI21X1 OAI21X1_349 ( .A(u2__abc_52138_new_n4609_), .B(u2_remHi_155_), .C(u2__abc_52138_new_n4822_), .Y(u2__abc_52138_new_n4823_));
OAI21X1 OAI21X1_3490 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_146_), .Y(u2__abc_52138_new_n14176_));
OAI21X1 OAI21X1_3491 ( .A(u2__abc_52138_new_n14179_), .B(u2__abc_52138_new_n14177_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14180_));
OAI21X1 OAI21X1_3492 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_147_), .Y(u2__abc_52138_new_n14184_));
OAI21X1 OAI21X1_3493 ( .A(u2__abc_52138_new_n14185_), .B(u2__abc_52138_new_n14187_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14188_));
OAI21X1 OAI21X1_3494 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_148_), .Y(u2__abc_52138_new_n14192_));
OAI21X1 OAI21X1_3495 ( .A(u2__abc_52138_new_n14194_), .B(u2__abc_52138_new_n14195_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14196_));
OAI21X1 OAI21X1_3496 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_149_), .Y(u2__abc_52138_new_n14200_));
OAI21X1 OAI21X1_3497 ( .A(u2__abc_52138_new_n14202_), .B(u2__abc_52138_new_n14201_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14203_));
OAI21X1 OAI21X1_3498 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_150_), .Y(u2__abc_52138_new_n14207_));
OAI21X1 OAI21X1_3499 ( .A(u2__abc_52138_new_n14209_), .B(u2__abc_52138_new_n14210_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14211_));
OAI21X1 OAI21X1_35 ( .A(aNan), .B(_abc_65734_new_n932_), .C(_abc_65734_new_n933_), .Y(\o[146] ));
OAI21X1 OAI21X1_350 ( .A(u2__abc_52138_new_n4599_), .B(u2__abc_52138_new_n4605_), .C(u2__abc_52138_new_n4604_), .Y(u2__abc_52138_new_n4825_));
OAI21X1 OAI21X1_3500 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_151_), .Y(u2__abc_52138_new_n14215_));
OAI21X1 OAI21X1_3501 ( .A(u2__abc_52138_new_n14216_), .B(u2__abc_52138_new_n14218_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14219_));
OAI21X1 OAI21X1_3502 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_152_), .Y(u2__abc_52138_new_n14223_));
OAI21X1 OAI21X1_3503 ( .A(u2__abc_52138_new_n14226_), .B(u2__abc_52138_new_n14224_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14227_));
OAI21X1 OAI21X1_3504 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_153_), .Y(u2__abc_52138_new_n14231_));
OAI21X1 OAI21X1_3505 ( .A(u2__abc_52138_new_n14233_), .B(u2__abc_52138_new_n14232_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14234_));
OAI21X1 OAI21X1_3506 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_154_), .Y(u2__abc_52138_new_n14238_));
OAI21X1 OAI21X1_3507 ( .A(u2__abc_52138_new_n14240_), .B(u2__abc_52138_new_n14241_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14242_));
OAI21X1 OAI21X1_3508 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_155_), .Y(u2__abc_52138_new_n14246_));
OAI21X1 OAI21X1_3509 ( .A(u2__abc_52138_new_n14247_), .B(u2__abc_52138_new_n14249_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14250_));
OAI21X1 OAI21X1_351 ( .A(u2__abc_52138_new_n4760_), .B(u2__abc_52138_new_n4814_), .C(u2__abc_52138_new_n4828_), .Y(u2__abc_52138_new_n4829_));
OAI21X1 OAI21X1_3510 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_156_), .Y(u2__abc_52138_new_n14254_));
OAI21X1 OAI21X1_3511 ( .A(u2__abc_52138_new_n14257_), .B(u2__abc_52138_new_n14255_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14258_));
OAI21X1 OAI21X1_3512 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_157_), .Y(u2__abc_52138_new_n14262_));
OAI21X1 OAI21X1_3513 ( .A(u2__abc_52138_new_n14264_), .B(u2__abc_52138_new_n14263_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14265_));
OAI21X1 OAI21X1_3514 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_158_), .Y(u2__abc_52138_new_n14269_));
OAI21X1 OAI21X1_3515 ( .A(u2__abc_52138_new_n14271_), .B(u2__abc_52138_new_n14272_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14273_));
OAI21X1 OAI21X1_3516 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_159_), .Y(u2__abc_52138_new_n14277_));
OAI21X1 OAI21X1_3517 ( .A(u2__abc_52138_new_n14278_), .B(u2__abc_52138_new_n14280_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14281_));
OAI21X1 OAI21X1_3518 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_160_), .Y(u2__abc_52138_new_n14285_));
OAI21X1 OAI21X1_3519 ( .A(u2__abc_52138_new_n14288_), .B(u2__abc_52138_new_n14286_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14289_));
OAI21X1 OAI21X1_352 ( .A(u2__abc_52138_new_n4528_), .B(u2__abc_52138_new_n4833_), .C(u2__abc_52138_new_n4533_), .Y(u2__abc_52138_new_n4834_));
OAI21X1 OAI21X1_3520 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_161_), .Y(u2__abc_52138_new_n14293_));
OAI21X1 OAI21X1_3521 ( .A(u2__abc_52138_new_n14295_), .B(u2__abc_52138_new_n14294_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14296_));
OAI21X1 OAI21X1_3522 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_162_), .Y(u2__abc_52138_new_n14300_));
OAI21X1 OAI21X1_3523 ( .A(u2__abc_52138_new_n14303_), .B(u2__abc_52138_new_n14301_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14304_));
OAI21X1 OAI21X1_3524 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_163_), .Y(u2__abc_52138_new_n14308_));
OAI21X1 OAI21X1_3525 ( .A(u2__abc_52138_new_n14309_), .B(u2__abc_52138_new_n14311_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14312_));
OAI21X1 OAI21X1_3526 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_164_), .Y(u2__abc_52138_new_n14316_));
OAI21X1 OAI21X1_3527 ( .A(u2__abc_52138_new_n14318_), .B(u2__abc_52138_new_n14319_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14320_));
OAI21X1 OAI21X1_3528 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_165_), .Y(u2__abc_52138_new_n14324_));
OAI21X1 OAI21X1_3529 ( .A(u2__abc_52138_new_n14326_), .B(u2__abc_52138_new_n14325_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14327_));
OAI21X1 OAI21X1_353 ( .A(u2__abc_52138_new_n4832_), .B(u2__abc_52138_new_n4831_), .C(u2__abc_52138_new_n4835_), .Y(u2__abc_52138_new_n4836_));
OAI21X1 OAI21X1_3530 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_166_), .Y(u2__abc_52138_new_n14331_));
OAI21X1 OAI21X1_3531 ( .A(u2__abc_52138_new_n14333_), .B(u2__abc_52138_new_n14334_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14335_));
OAI21X1 OAI21X1_3532 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_167_), .Y(u2__abc_52138_new_n14339_));
OAI21X1 OAI21X1_3533 ( .A(u2__abc_52138_new_n14340_), .B(u2__abc_52138_new_n14342_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14343_));
OAI21X1 OAI21X1_3534 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_168_), .Y(u2__abc_52138_new_n14347_));
OAI21X1 OAI21X1_3535 ( .A(u2__abc_52138_new_n14350_), .B(u2__abc_52138_new_n14348_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14351_));
OAI21X1 OAI21X1_3536 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_169_), .Y(u2__abc_52138_new_n14355_));
OAI21X1 OAI21X1_3537 ( .A(u2__abc_52138_new_n14357_), .B(u2__abc_52138_new_n14356_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14358_));
OAI21X1 OAI21X1_3538 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_170_), .Y(u2__abc_52138_new_n14362_));
OAI21X1 OAI21X1_3539 ( .A(u2__abc_52138_new_n14364_), .B(u2__abc_52138_new_n14365_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14366_));
OAI21X1 OAI21X1_354 ( .A(u2__abc_52138_new_n4567_), .B(u2__abc_52138_new_n4838_), .C(u2__abc_52138_new_n4562_), .Y(u2__abc_52138_new_n4839_));
OAI21X1 OAI21X1_3540 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_171_), .Y(u2__abc_52138_new_n14370_));
OAI21X1 OAI21X1_3541 ( .A(u2__abc_52138_new_n14371_), .B(u2__abc_52138_new_n14373_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14374_));
OAI21X1 OAI21X1_3542 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_172_), .Y(u2__abc_52138_new_n14378_));
OAI21X1 OAI21X1_3543 ( .A(u2__abc_52138_new_n14381_), .B(u2__abc_52138_new_n14379_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14382_));
OAI21X1 OAI21X1_3544 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_173_), .Y(u2__abc_52138_new_n14386_));
OAI21X1 OAI21X1_3545 ( .A(u2__abc_52138_new_n14388_), .B(u2__abc_52138_new_n14387_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14389_));
OAI21X1 OAI21X1_3546 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_174_), .Y(u2__abc_52138_new_n14393_));
OAI21X1 OAI21X1_3547 ( .A(u2__abc_52138_new_n14395_), .B(u2__abc_52138_new_n14396_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14397_));
OAI21X1 OAI21X1_3548 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_175_), .Y(u2__abc_52138_new_n14401_));
OAI21X1 OAI21X1_3549 ( .A(u2__abc_52138_new_n14402_), .B(u2__abc_52138_new_n14404_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14405_));
OAI21X1 OAI21X1_355 ( .A(u2__abc_52138_new_n4551_), .B(u2__abc_52138_new_n4557_), .C(u2__abc_52138_new_n4556_), .Y(u2__abc_52138_new_n4841_));
OAI21X1 OAI21X1_3550 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_176_), .Y(u2__abc_52138_new_n14409_));
OAI21X1 OAI21X1_3551 ( .A(u2__abc_52138_new_n14412_), .B(u2__abc_52138_new_n14410_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14413_));
OAI21X1 OAI21X1_3552 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_177_), .Y(u2__abc_52138_new_n14417_));
OAI21X1 OAI21X1_3553 ( .A(u2__abc_52138_new_n14419_), .B(u2__abc_52138_new_n14418_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14420_));
OAI21X1 OAI21X1_3554 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_178_), .Y(u2__abc_52138_new_n14424_));
OAI21X1 OAI21X1_3555 ( .A(u2__abc_52138_new_n14426_), .B(u2__abc_52138_new_n14427_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14428_));
OAI21X1 OAI21X1_3556 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_179_), .Y(u2__abc_52138_new_n14432_));
OAI21X1 OAI21X1_3557 ( .A(u2__abc_52138_new_n14433_), .B(u2__abc_52138_new_n14435_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14436_));
OAI21X1 OAI21X1_3558 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_180_), .Y(u2__abc_52138_new_n14440_));
OAI21X1 OAI21X1_3559 ( .A(u2__abc_52138_new_n14443_), .B(u2__abc_52138_new_n14441_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14444_));
OAI21X1 OAI21X1_356 ( .A(u2__abc_52138_new_n4840_), .B(u2__abc_52138_new_n4837_), .C(u2__abc_52138_new_n4842_), .Y(u2__abc_52138_new_n4843_));
OAI21X1 OAI21X1_3560 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_181_), .Y(u2__abc_52138_new_n14448_));
OAI21X1 OAI21X1_3561 ( .A(u2__abc_52138_new_n14450_), .B(u2__abc_52138_new_n14449_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14451_));
OAI21X1 OAI21X1_3562 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_182_), .Y(u2__abc_52138_new_n14455_));
OAI21X1 OAI21X1_3563 ( .A(u2__abc_52138_new_n14457_), .B(u2__abc_52138_new_n14458_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14459_));
OAI21X1 OAI21X1_3564 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_183_), .Y(u2__abc_52138_new_n14463_));
OAI21X1 OAI21X1_3565 ( .A(u2__abc_52138_new_n14464_), .B(u2__abc_52138_new_n14466_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14467_));
OAI21X1 OAI21X1_3566 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_184_), .Y(u2__abc_52138_new_n14471_));
OAI21X1 OAI21X1_3567 ( .A(u2__abc_52138_new_n14474_), .B(u2__abc_52138_new_n14472_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14475_));
OAI21X1 OAI21X1_3568 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_185_), .Y(u2__abc_52138_new_n14479_));
OAI21X1 OAI21X1_3569 ( .A(u2__abc_52138_new_n14481_), .B(u2__abc_52138_new_n14480_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14482_));
OAI21X1 OAI21X1_357 ( .A(sqrto_167_), .B(u2__abc_52138_new_n4514_), .C(u2__abc_52138_new_n4520_), .Y(u2__abc_52138_new_n4845_));
OAI21X1 OAI21X1_3570 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_186_), .Y(u2__abc_52138_new_n14486_));
OAI21X1 OAI21X1_3571 ( .A(u2__abc_52138_new_n14488_), .B(u2__abc_52138_new_n14489_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14490_));
OAI21X1 OAI21X1_3572 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_187_), .Y(u2__abc_52138_new_n14494_));
OAI21X1 OAI21X1_3573 ( .A(u2__abc_52138_new_n14495_), .B(u2__abc_52138_new_n14497_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14498_));
OAI21X1 OAI21X1_3574 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_188_), .Y(u2__abc_52138_new_n14502_));
OAI21X1 OAI21X1_3575 ( .A(u2__abc_52138_new_n14505_), .B(u2__abc_52138_new_n14503_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14506_));
OAI21X1 OAI21X1_3576 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_189_), .Y(u2__abc_52138_new_n14510_));
OAI21X1 OAI21X1_3577 ( .A(u2__abc_52138_new_n14512_), .B(u2__abc_52138_new_n14511_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14513_));
OAI21X1 OAI21X1_3578 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_190_), .Y(u2__abc_52138_new_n14517_));
OAI21X1 OAI21X1_3579 ( .A(u2__abc_52138_new_n14519_), .B(u2__abc_52138_new_n14520_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14521_));
OAI21X1 OAI21X1_358 ( .A(u2__abc_52138_new_n4512_), .B(u2_remHi_167_), .C(u2__abc_52138_new_n4845_), .Y(u2__abc_52138_new_n4846_));
OAI21X1 OAI21X1_3580 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_191_), .Y(u2__abc_52138_new_n14525_));
OAI21X1 OAI21X1_3581 ( .A(u2__abc_52138_new_n14526_), .B(u2__abc_52138_new_n14528_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14529_));
OAI21X1 OAI21X1_3582 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_192_), .Y(u2__abc_52138_new_n14533_));
OAI21X1 OAI21X1_3583 ( .A(u2__abc_52138_new_n14535_), .B(u2__abc_52138_new_n14536_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14537_));
OAI21X1 OAI21X1_3584 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_193_), .Y(u2__abc_52138_new_n14541_));
OAI21X1 OAI21X1_3585 ( .A(u2__abc_52138_new_n14543_), .B(u2__abc_52138_new_n14542_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14544_));
OAI21X1 OAI21X1_3586 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_194_), .Y(u2__abc_52138_new_n14548_));
OAI21X1 OAI21X1_3587 ( .A(u2__abc_52138_new_n14551_), .B(u2__abc_52138_new_n14549_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14552_));
OAI21X1 OAI21X1_3588 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_195_), .Y(u2__abc_52138_new_n14556_));
OAI21X1 OAI21X1_3589 ( .A(u2__abc_52138_new_n14557_), .B(u2__abc_52138_new_n14559_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14560_));
OAI21X1 OAI21X1_359 ( .A(u2__abc_52138_new_n4504_), .B(u2__abc_52138_new_n4510_), .C(u2__abc_52138_new_n4509_), .Y(u2__abc_52138_new_n4848_));
OAI21X1 OAI21X1_3590 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_196_), .Y(u2__abc_52138_new_n14564_));
OAI21X1 OAI21X1_3591 ( .A(u2__abc_52138_new_n14566_), .B(u2__abc_52138_new_n14567_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14568_));
OAI21X1 OAI21X1_3592 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_197_), .Y(u2__abc_52138_new_n14572_));
OAI21X1 OAI21X1_3593 ( .A(u2__abc_52138_new_n14574_), .B(u2__abc_52138_new_n14573_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14575_));
OAI21X1 OAI21X1_3594 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_198_), .Y(u2__abc_52138_new_n14579_));
OAI21X1 OAI21X1_3595 ( .A(u2__abc_52138_new_n14581_), .B(u2__abc_52138_new_n14582_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14583_));
OAI21X1 OAI21X1_3596 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_199_), .Y(u2__abc_52138_new_n14587_));
OAI21X1 OAI21X1_3597 ( .A(u2__abc_52138_new_n14588_), .B(u2__abc_52138_new_n14590_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14591_));
OAI21X1 OAI21X1_3598 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_200_), .Y(u2__abc_52138_new_n14595_));
OAI21X1 OAI21X1_3599 ( .A(u2__abc_52138_new_n14598_), .B(u2__abc_52138_new_n14596_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14599_));
OAI21X1 OAI21X1_36 ( .A(aNan), .B(_abc_65734_new_n935_), .C(_abc_65734_new_n936_), .Y(\o[147] ));
OAI21X1 OAI21X1_360 ( .A(u2__abc_52138_new_n4497_), .B(u2__abc_52138_new_n4493_), .C(u2__abc_52138_new_n4492_), .Y(u2__abc_52138_new_n4851_));
OAI21X1 OAI21X1_3600 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_201_), .Y(u2__abc_52138_new_n14603_));
OAI21X1 OAI21X1_3601 ( .A(u2__abc_52138_new_n14605_), .B(u2__abc_52138_new_n14604_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14606_));
OAI21X1 OAI21X1_3602 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_202_), .Y(u2__abc_52138_new_n14610_));
OAI21X1 OAI21X1_3603 ( .A(u2__abc_52138_new_n14612_), .B(u2__abc_52138_new_n14613_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14614_));
OAI21X1 OAI21X1_3604 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_203_), .Y(u2__abc_52138_new_n14619_));
OAI21X1 OAI21X1_3605 ( .A(u2__abc_52138_new_n14620_), .B(u2__abc_52138_new_n14622_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14623_));
OAI21X1 OAI21X1_3606 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_204_), .Y(u2__abc_52138_new_n14627_));
OAI21X1 OAI21X1_3607 ( .A(u2__abc_52138_new_n14630_), .B(u2__abc_52138_new_n14628_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14631_));
OAI21X1 OAI21X1_3608 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_205_), .Y(u2__abc_52138_new_n14635_));
OAI21X1 OAI21X1_3609 ( .A(u2__abc_52138_new_n14637_), .B(u2__abc_52138_new_n14636_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14638_));
OAI21X1 OAI21X1_361 ( .A(sqrto_173_), .B(u2__abc_52138_new_n4485_), .C(u2__abc_52138_new_n4853_), .Y(u2__abc_52138_new_n4854_));
OAI21X1 OAI21X1_3610 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_206_), .Y(u2__abc_52138_new_n14642_));
OAI21X1 OAI21X1_3611 ( .A(u2__abc_52138_new_n14644_), .B(u2__abc_52138_new_n14645_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14646_));
OAI21X1 OAI21X1_3612 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_207_), .Y(u2__abc_52138_new_n14650_));
OAI21X1 OAI21X1_3613 ( .A(u2__abc_52138_new_n14651_), .B(u2__abc_52138_new_n14653_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14654_));
OAI21X1 OAI21X1_3614 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_208_), .Y(u2__abc_52138_new_n14658_));
OAI21X1 OAI21X1_3615 ( .A(u2__abc_52138_new_n14661_), .B(u2__abc_52138_new_n14659_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14662_));
OAI21X1 OAI21X1_3616 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_209_), .Y(u2__abc_52138_new_n14666_));
OAI21X1 OAI21X1_3617 ( .A(u2__abc_52138_new_n14668_), .B(u2__abc_52138_new_n14667_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14669_));
OAI21X1 OAI21X1_3618 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_210_), .Y(u2__abc_52138_new_n14673_));
OAI21X1 OAI21X1_3619 ( .A(u2__abc_52138_new_n14675_), .B(u2__abc_52138_new_n14676_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14677_));
OAI21X1 OAI21X1_362 ( .A(u2__abc_52138_new_n4756_), .B(u2__abc_52138_new_n4844_), .C(u2__abc_52138_new_n4856_), .Y(u2__abc_52138_new_n4857_));
OAI21X1 OAI21X1_3620 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_211_), .Y(u2__abc_52138_new_n14681_));
OAI21X1 OAI21X1_3621 ( .A(u2__abc_52138_new_n14682_), .B(u2__abc_52138_new_n14684_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14685_));
OAI21X1 OAI21X1_3622 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_212_), .Y(u2__abc_52138_new_n14689_));
OAI21X1 OAI21X1_3623 ( .A(u2__abc_52138_new_n14692_), .B(u2__abc_52138_new_n14690_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14693_));
OAI21X1 OAI21X1_3624 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_213_), .Y(u2__abc_52138_new_n14697_));
OAI21X1 OAI21X1_3625 ( .A(u2__abc_52138_new_n14699_), .B(u2__abc_52138_new_n14698_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14700_));
OAI21X1 OAI21X1_3626 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_214_), .Y(u2__abc_52138_new_n14704_));
OAI21X1 OAI21X1_3627 ( .A(u2__abc_52138_new_n14706_), .B(u2__abc_52138_new_n14707_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14708_));
OAI21X1 OAI21X1_3628 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_215_), .Y(u2__abc_52138_new_n14712_));
OAI21X1 OAI21X1_3629 ( .A(u2__abc_52138_new_n14713_), .B(u2__abc_52138_new_n14715_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14716_));
OAI21X1 OAI21X1_363 ( .A(u2__abc_52138_new_n4466_), .B(u2__abc_52138_new_n4858_), .C(u2__abc_52138_new_n4472_), .Y(u2__abc_52138_new_n4859_));
OAI21X1 OAI21X1_3630 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_216_), .Y(u2__abc_52138_new_n14720_));
OAI21X1 OAI21X1_3631 ( .A(u2__abc_52138_new_n14723_), .B(u2__abc_52138_new_n14721_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14724_));
OAI21X1 OAI21X1_3632 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_217_), .Y(u2__abc_52138_new_n14728_));
OAI21X1 OAI21X1_3633 ( .A(u2__abc_52138_new_n14730_), .B(u2__abc_52138_new_n14729_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14731_));
OAI21X1 OAI21X1_3634 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_218_), .Y(u2__abc_52138_new_n14735_));
OAI21X1 OAI21X1_3635 ( .A(u2__abc_52138_new_n14737_), .B(u2__abc_52138_new_n14738_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14739_));
OAI21X1 OAI21X1_3636 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_219_), .Y(u2__abc_52138_new_n14743_));
OAI21X1 OAI21X1_3637 ( .A(u2__abc_52138_new_n14744_), .B(u2__abc_52138_new_n14746_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14747_));
OAI21X1 OAI21X1_3638 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_220_), .Y(u2__abc_52138_new_n14751_));
OAI21X1 OAI21X1_3639 ( .A(u2__abc_52138_new_n14754_), .B(u2__abc_52138_new_n14752_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14755_));
OAI21X1 OAI21X1_364 ( .A(u2__abc_52138_new_n4455_), .B(u2__abc_52138_new_n4461_), .C(u2__abc_52138_new_n4460_), .Y(u2__abc_52138_new_n4860_));
OAI21X1 OAI21X1_3640 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_221_), .Y(u2__abc_52138_new_n14759_));
OAI21X1 OAI21X1_3641 ( .A(u2__abc_52138_new_n14761_), .B(u2__abc_52138_new_n14760_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14762_));
OAI21X1 OAI21X1_3642 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_222_), .Y(u2__abc_52138_new_n14766_));
OAI21X1 OAI21X1_3643 ( .A(u2__abc_52138_new_n14768_), .B(u2__abc_52138_new_n14769_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14770_));
OAI21X1 OAI21X1_3644 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_223_), .Y(u2__abc_52138_new_n14774_));
OAI21X1 OAI21X1_3645 ( .A(u2__abc_52138_new_n14775_), .B(u2__abc_52138_new_n14777_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14778_));
OAI21X1 OAI21X1_3646 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_224_), .Y(u2__abc_52138_new_n14782_));
OAI21X1 OAI21X1_3647 ( .A(u2__abc_52138_new_n14784_), .B(u2__abc_52138_new_n14785_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14786_));
OAI21X1 OAI21X1_3648 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(sqrto_225_), .Y(u2__abc_52138_new_n14790_));
OAI21X1 OAI21X1_3649 ( .A(u2__abc_52138_new_n14792_), .B(u2__abc_52138_new_n14791_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14793_));
OAI21X1 OAI21X1_365 ( .A(u2__abc_52138_new_n4432_), .B(u2__abc_52138_new_n4862_), .C(u2__abc_52138_new_n4437_), .Y(u2__abc_52138_new_n4863_));
OAI21X1 OAI21X1_3650 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_226_), .Y(u2__abc_52138_new_n14797_));
OAI21X1 OAI21X1_3651 ( .A(u2__abc_52138_new_n14799_), .B(u2__abc_52138_new_n14800_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14801_));
OAI21X1 OAI21X1_3652 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_227_), .Y(u2__abc_52138_new_n14805_));
OAI21X1 OAI21X1_3653 ( .A(u2__abc_52138_new_n14806_), .B(u2__abc_52138_new_n14808_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14809_));
OAI21X1 OAI21X1_3654 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_228_), .Y(u2__abc_52138_new_n14813_));
OAI21X1 OAI21X1_3655 ( .A(u2__abc_52138_new_n14816_), .B(u2__abc_52138_new_n14814_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14817_));
OAI21X1 OAI21X1_3656 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_229_), .Y(u2__abc_52138_new_n14821_));
OAI21X1 OAI21X1_3657 ( .A(u2__abc_52138_new_n14823_), .B(u2__abc_52138_new_n14822_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14824_));
OAI21X1 OAI21X1_3658 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_230_), .Y(u2__abc_52138_new_n14828_));
OAI21X1 OAI21X1_3659 ( .A(u2__abc_52138_new_n14830_), .B(u2__abc_52138_new_n14831_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14832_));
OAI21X1 OAI21X1_366 ( .A(u2__abc_52138_new_n4448_), .B(u2__abc_52138_new_n4444_), .C(u2__abc_52138_new_n4443_), .Y(u2__abc_52138_new_n4864_));
OAI21X1 OAI21X1_3660 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_231_), .Y(u2__abc_52138_new_n14836_));
OAI21X1 OAI21X1_3661 ( .A(u2__abc_52138_new_n14837_), .B(u2__abc_52138_new_n14839_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14840_));
OAI21X1 OAI21X1_3662 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_232_), .Y(u2__abc_52138_new_n14844_));
OAI21X1 OAI21X1_3663 ( .A(u2__abc_52138_new_n14847_), .B(u2__abc_52138_new_n14845_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14848_));
OAI21X1 OAI21X1_3664 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_233_), .Y(u2__abc_52138_new_n14852_));
OAI21X1 OAI21X1_3665 ( .A(u2__abc_52138_new_n14854_), .B(u2__abc_52138_new_n14853_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14855_));
OAI21X1 OAI21X1_3666 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_234_), .Y(u2__abc_52138_new_n14859_));
OAI21X1 OAI21X1_3667 ( .A(u2__abc_52138_new_n14861_), .B(u2__abc_52138_new_n14862_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14863_));
OAI21X1 OAI21X1_3668 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_235_), .Y(u2__abc_52138_new_n14867_));
OAI21X1 OAI21X1_3669 ( .A(u2__abc_52138_new_n14868_), .B(u2__abc_52138_new_n14870_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14871_));
OAI21X1 OAI21X1_367 ( .A(u2__abc_52138_new_n4451_), .B(u2__abc_52138_new_n4861_), .C(u2__abc_52138_new_n4865_), .Y(u2__abc_52138_new_n4866_));
OAI21X1 OAI21X1_3670 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_236_), .Y(u2__abc_52138_new_n14875_));
OAI21X1 OAI21X1_3671 ( .A(u2__abc_52138_new_n14878_), .B(u2__abc_52138_new_n14876_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14879_));
OAI21X1 OAI21X1_3672 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_237_), .Y(u2__abc_52138_new_n14883_));
OAI21X1 OAI21X1_3673 ( .A(u2__abc_52138_new_n14885_), .B(u2__abc_52138_new_n14884_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14886_));
OAI21X1 OAI21X1_3674 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_238_), .Y(u2__abc_52138_new_n14890_));
OAI21X1 OAI21X1_3675 ( .A(u2__abc_52138_new_n14892_), .B(u2__abc_52138_new_n14893_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14894_));
OAI21X1 OAI21X1_3676 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_239_), .Y(u2__abc_52138_new_n14898_));
OAI21X1 OAI21X1_3677 ( .A(u2__abc_52138_new_n14899_), .B(u2__abc_52138_new_n14901_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14902_));
OAI21X1 OAI21X1_3678 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_240_), .Y(u2__abc_52138_new_n14906_));
OAI21X1 OAI21X1_3679 ( .A(u2__abc_52138_new_n14908_), .B(u2__abc_52138_new_n14909_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14910_));
OAI21X1 OAI21X1_368 ( .A(u2__abc_52138_new_n4385_), .B(u2__abc_52138_new_n4391_), .C(u2__abc_52138_new_n4390_), .Y(u2__abc_52138_new_n4868_));
OAI21X1 OAI21X1_3680 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_241_), .Y(u2__abc_52138_new_n14914_));
OAI21X1 OAI21X1_3681 ( .A(u2__abc_52138_new_n14916_), .B(u2__abc_52138_new_n14915_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14917_));
OAI21X1 OAI21X1_3682 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_242_), .Y(u2__abc_52138_new_n14921_));
OAI21X1 OAI21X1_3683 ( .A(u2__abc_52138_new_n14923_), .B(u2__abc_52138_new_n14924_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14925_));
OAI21X1 OAI21X1_3684 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_243_), .Y(u2__abc_52138_new_n14929_));
OAI21X1 OAI21X1_3685 ( .A(u2__abc_52138_new_n14930_), .B(u2__abc_52138_new_n14932_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14933_));
OAI21X1 OAI21X1_3686 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_244_), .Y(u2__abc_52138_new_n14937_));
OAI21X1 OAI21X1_3687 ( .A(u2__abc_52138_new_n14940_), .B(u2__abc_52138_new_n14938_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14941_));
OAI21X1 OAI21X1_3688 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_245_), .Y(u2__abc_52138_new_n14945_));
OAI21X1 OAI21X1_3689 ( .A(u2__abc_52138_new_n14947_), .B(u2__abc_52138_new_n14946_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14948_));
OAI21X1 OAI21X1_369 ( .A(u2__abc_52138_new_n4396_), .B(u2__abc_52138_new_n4402_), .C(u2__abc_52138_new_n4401_), .Y(u2__abc_52138_new_n4869_));
OAI21X1 OAI21X1_3690 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_246_), .Y(u2__abc_52138_new_n14952_));
OAI21X1 OAI21X1_3691 ( .A(u2__abc_52138_new_n14954_), .B(u2__abc_52138_new_n14955_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14956_));
OAI21X1 OAI21X1_3692 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_247_), .Y(u2__abc_52138_new_n14960_));
OAI21X1 OAI21X1_3693 ( .A(u2__abc_52138_new_n14961_), .B(u2__abc_52138_new_n14963_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14964_));
OAI21X1 OAI21X1_3694 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_248_), .Y(u2__abc_52138_new_n14968_));
OAI21X1 OAI21X1_3695 ( .A(u2__abc_52138_new_n14970_), .B(u2__abc_52138_new_n14971_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14972_));
OAI21X1 OAI21X1_3696 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_249_), .Y(u2__abc_52138_new_n14976_));
OAI21X1 OAI21X1_3697 ( .A(u2__abc_52138_new_n14978_), .B(u2__abc_52138_new_n14977_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14979_));
OAI21X1 OAI21X1_3698 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_250_), .Y(u2__abc_52138_new_n14983_));
OAI21X1 OAI21X1_3699 ( .A(u2__abc_52138_new_n14985_), .B(u2__abc_52138_new_n14986_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14987_));
OAI21X1 OAI21X1_37 ( .A(aNan), .B(_abc_65734_new_n938_), .C(_abc_65734_new_n939_), .Y(\o[148] ));
OAI21X1 OAI21X1_370 ( .A(u2__abc_52138_new_n4424_), .B(u2__abc_52138_new_n4420_), .C(u2__abc_52138_new_n4419_), .Y(u2__abc_52138_new_n4871_));
OAI21X1 OAI21X1_3700 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_251_), .Y(u2__abc_52138_new_n14991_));
OAI21X1 OAI21X1_3701 ( .A(u2__abc_52138_new_n14992_), .B(u2__abc_52138_new_n14994_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n14995_));
OAI21X1 OAI21X1_3702 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_252_), .Y(u2__abc_52138_new_n14999_));
OAI21X1 OAI21X1_3703 ( .A(u2__abc_52138_new_n15001_), .B(u2__abc_52138_new_n15002_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15003_));
OAI21X1 OAI21X1_3704 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_253_), .Y(u2__abc_52138_new_n15007_));
OAI21X1 OAI21X1_3705 ( .A(u2__abc_52138_new_n15009_), .B(u2__abc_52138_new_n15008_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15010_));
OAI21X1 OAI21X1_3706 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_254_), .Y(u2__abc_52138_new_n15014_));
OAI21X1 OAI21X1_3707 ( .A(u2__abc_52138_new_n15016_), .B(u2__abc_52138_new_n15017_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15018_));
OAI21X1 OAI21X1_3708 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_255_), .Y(u2__abc_52138_new_n15022_));
OAI21X1 OAI21X1_3709 ( .A(u2__abc_52138_new_n15023_), .B(u2__abc_52138_new_n15025_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15026_));
OAI21X1 OAI21X1_371 ( .A(u2__abc_52138_new_n4408_), .B(u2__abc_52138_new_n4872_), .C(u2__abc_52138_new_n4413_), .Y(u2__abc_52138_new_n4873_));
OAI21X1 OAI21X1_3710 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_256_), .Y(u2__abc_52138_new_n15030_));
OAI21X1 OAI21X1_3711 ( .A(u2__abc_52138_new_n15032_), .B(u2__abc_52138_new_n15033_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15034_));
OAI21X1 OAI21X1_3712 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_257_), .Y(u2__abc_52138_new_n15038_));
OAI21X1 OAI21X1_3713 ( .A(u2__abc_52138_new_n15040_), .B(u2__abc_52138_new_n15039_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15041_));
OAI21X1 OAI21X1_3714 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_258_), .Y(u2__abc_52138_new_n15045_));
OAI21X1 OAI21X1_3715 ( .A(u2__abc_52138_new_n15048_), .B(u2__abc_52138_new_n15046_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15049_));
OAI21X1 OAI21X1_3716 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_259_), .Y(u2__abc_52138_new_n15053_));
OAI21X1 OAI21X1_3717 ( .A(u2__abc_52138_new_n15054_), .B(u2__abc_52138_new_n15056_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15057_));
OAI21X1 OAI21X1_3718 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_260_), .Y(u2__abc_52138_new_n15061_));
OAI21X1 OAI21X1_3719 ( .A(u2__abc_52138_new_n15063_), .B(u2__abc_52138_new_n15064_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15065_));
OAI21X1 OAI21X1_372 ( .A(u2__abc_52138_new_n4427_), .B(u2__abc_52138_new_n4870_), .C(u2__abc_52138_new_n4874_), .Y(u2__abc_52138_new_n4875_));
OAI21X1 OAI21X1_3720 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_261_), .Y(u2__abc_52138_new_n15069_));
OAI21X1 OAI21X1_3721 ( .A(u2__abc_52138_new_n15071_), .B(u2__abc_52138_new_n15070_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15072_));
OAI21X1 OAI21X1_3722 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_262_), .Y(u2__abc_52138_new_n15076_));
OAI21X1 OAI21X1_3723 ( .A(u2__abc_52138_new_n15078_), .B(u2__abc_52138_new_n15079_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15080_));
OAI21X1 OAI21X1_3724 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_263_), .Y(u2__abc_52138_new_n15084_));
OAI21X1 OAI21X1_3725 ( .A(u2__abc_52138_new_n15085_), .B(u2__abc_52138_new_n15087_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15088_));
OAI21X1 OAI21X1_3726 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_264_), .Y(u2__abc_52138_new_n15092_));
OAI21X1 OAI21X1_3727 ( .A(u2__abc_52138_new_n15095_), .B(u2__abc_52138_new_n15093_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15096_));
OAI21X1 OAI21X1_3728 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_265_), .Y(u2__abc_52138_new_n15100_));
OAI21X1 OAI21X1_3729 ( .A(u2__abc_52138_new_n15102_), .B(u2__abc_52138_new_n15101_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15103_));
OAI21X1 OAI21X1_373 ( .A(u2__abc_52138_new_n4759_), .B(u2__abc_52138_new_n4830_), .C(u2__abc_52138_new_n4878_), .Y(u2__abc_52138_new_n4879_));
OAI21X1 OAI21X1_3730 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_266_), .Y(u2__abc_52138_new_n15107_));
OAI21X1 OAI21X1_3731 ( .A(u2__abc_52138_new_n15109_), .B(u2__abc_52138_new_n15110_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15111_));
OAI21X1 OAI21X1_3732 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_267_), .Y(u2__abc_52138_new_n15115_));
OAI21X1 OAI21X1_3733 ( .A(u2__abc_52138_new_n15116_), .B(u2__abc_52138_new_n15118_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15119_));
OAI21X1 OAI21X1_3734 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_268_), .Y(u2__abc_52138_new_n15123_));
OAI21X1 OAI21X1_3735 ( .A(u2__abc_52138_new_n15126_), .B(u2__abc_52138_new_n15124_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15127_));
OAI21X1 OAI21X1_3736 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_269_), .Y(u2__abc_52138_new_n15131_));
OAI21X1 OAI21X1_3737 ( .A(u2__abc_52138_new_n15133_), .B(u2__abc_52138_new_n15132_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15134_));
OAI21X1 OAI21X1_3738 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_270_), .Y(u2__abc_52138_new_n15138_));
OAI21X1 OAI21X1_3739 ( .A(u2__abc_52138_new_n15140_), .B(u2__abc_52138_new_n15141_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15142_));
OAI21X1 OAI21X1_374 ( .A(u2__abc_52138_new_n4885_), .B(u2__abc_52138_new_n4884_), .C(u2__abc_52138_new_n4886_), .Y(u2__abc_52138_new_n4887_));
OAI21X1 OAI21X1_3740 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_271_), .Y(u2__abc_52138_new_n15146_));
OAI21X1 OAI21X1_3741 ( .A(u2__abc_52138_new_n15147_), .B(u2__abc_52138_new_n15149_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15150_));
OAI21X1 OAI21X1_3742 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_272_), .Y(u2__abc_52138_new_n15154_));
OAI21X1 OAI21X1_3743 ( .A(u2__abc_52138_new_n15157_), .B(u2__abc_52138_new_n15155_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15158_));
OAI21X1 OAI21X1_3744 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_273_), .Y(u2__abc_52138_new_n15162_));
OAI21X1 OAI21X1_3745 ( .A(u2__abc_52138_new_n15164_), .B(u2__abc_52138_new_n15163_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15165_));
OAI21X1 OAI21X1_3746 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_274_), .Y(u2__abc_52138_new_n15169_));
OAI21X1 OAI21X1_3747 ( .A(u2__abc_52138_new_n15171_), .B(u2__abc_52138_new_n15172_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15173_));
OAI21X1 OAI21X1_3748 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_275_), .Y(u2__abc_52138_new_n15177_));
OAI21X1 OAI21X1_3749 ( .A(u2__abc_52138_new_n15178_), .B(u2__abc_52138_new_n15180_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15181_));
OAI21X1 OAI21X1_375 ( .A(u2__abc_52138_new_n4350_), .B(u2__abc_52138_new_n4889_), .C(u2__abc_52138_new_n4345_), .Y(u2__abc_52138_new_n4890_));
OAI21X1 OAI21X1_3750 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_276_), .Y(u2__abc_52138_new_n15185_));
OAI21X1 OAI21X1_3751 ( .A(u2__abc_52138_new_n15188_), .B(u2__abc_52138_new_n15186_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15189_));
OAI21X1 OAI21X1_3752 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_277_), .Y(u2__abc_52138_new_n15193_));
OAI21X1 OAI21X1_3753 ( .A(u2__abc_52138_new_n15195_), .B(u2__abc_52138_new_n15194_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15196_));
OAI21X1 OAI21X1_3754 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_278_), .Y(u2__abc_52138_new_n15200_));
OAI21X1 OAI21X1_3755 ( .A(u2__abc_52138_new_n15202_), .B(u2__abc_52138_new_n15203_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15204_));
OAI21X1 OAI21X1_3756 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_279_), .Y(u2__abc_52138_new_n15208_));
OAI21X1 OAI21X1_3757 ( .A(u2__abc_52138_new_n15209_), .B(u2__abc_52138_new_n15211_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15212_));
OAI21X1 OAI21X1_3758 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_280_), .Y(u2__abc_52138_new_n15216_));
OAI21X1 OAI21X1_3759 ( .A(u2__abc_52138_new_n15219_), .B(u2__abc_52138_new_n15217_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15220_));
OAI21X1 OAI21X1_376 ( .A(u2__abc_52138_new_n4334_), .B(u2__abc_52138_new_n4892_), .C(u2__abc_52138_new_n4339_), .Y(u2__abc_52138_new_n4893_));
OAI21X1 OAI21X1_3760 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_281_), .Y(u2__abc_52138_new_n15224_));
OAI21X1 OAI21X1_3761 ( .A(u2__abc_52138_new_n15226_), .B(u2__abc_52138_new_n15225_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15227_));
OAI21X1 OAI21X1_3762 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_282_), .Y(u2__abc_52138_new_n15231_));
OAI21X1 OAI21X1_3763 ( .A(u2__abc_52138_new_n15233_), .B(u2__abc_52138_new_n15234_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15235_));
OAI21X1 OAI21X1_3764 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_283_), .Y(u2__abc_52138_new_n15239_));
OAI21X1 OAI21X1_3765 ( .A(u2__abc_52138_new_n15240_), .B(u2__abc_52138_new_n15242_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15243_));
OAI21X1 OAI21X1_3766 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_284_), .Y(u2__abc_52138_new_n15247_));
OAI21X1 OAI21X1_3767 ( .A(u2__abc_52138_new_n15250_), .B(u2__abc_52138_new_n15248_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15251_));
OAI21X1 OAI21X1_3768 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_285_), .Y(u2__abc_52138_new_n15255_));
OAI21X1 OAI21X1_3769 ( .A(u2__abc_52138_new_n15257_), .B(u2__abc_52138_new_n15256_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15258_));
OAI21X1 OAI21X1_377 ( .A(u2__abc_52138_new_n4891_), .B(u2__abc_52138_new_n4888_), .C(u2__abc_52138_new_n4894_), .Y(u2__abc_52138_new_n4895_));
OAI21X1 OAI21X1_3770 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_286_), .Y(u2__abc_52138_new_n15262_));
OAI21X1 OAI21X1_3771 ( .A(u2__abc_52138_new_n15264_), .B(u2__abc_52138_new_n15265_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15266_));
OAI21X1 OAI21X1_3772 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_287_), .Y(u2__abc_52138_new_n15270_));
OAI21X1 OAI21X1_3773 ( .A(u2__abc_52138_new_n15271_), .B(u2__abc_52138_new_n15273_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15274_));
OAI21X1 OAI21X1_3774 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_288_), .Y(u2__abc_52138_new_n15278_));
OAI21X1 OAI21X1_3775 ( .A(u2__abc_52138_new_n15280_), .B(u2__abc_52138_new_n15281_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15282_));
OAI21X1 OAI21X1_3776 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_289_), .Y(u2__abc_52138_new_n15286_));
OAI21X1 OAI21X1_3777 ( .A(u2__abc_52138_new_n15288_), .B(u2__abc_52138_new_n15287_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15289_));
OAI21X1 OAI21X1_3778 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_290_), .Y(u2__abc_52138_new_n15293_));
OAI21X1 OAI21X1_3779 ( .A(u2__abc_52138_new_n15295_), .B(u2__abc_52138_new_n15296_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15297_));
OAI21X1 OAI21X1_378 ( .A(u2__abc_52138_new_n4308_), .B(u2__abc_52138_new_n4898_), .C(u2__abc_52138_new_n4303_), .Y(u2__abc_52138_new_n4899_));
OAI21X1 OAI21X1_3780 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_291_), .Y(u2__abc_52138_new_n15301_));
OAI21X1 OAI21X1_3781 ( .A(u2__abc_52138_new_n15302_), .B(u2__abc_52138_new_n15304_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15305_));
OAI21X1 OAI21X1_3782 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_292_), .Y(u2__abc_52138_new_n15309_));
OAI21X1 OAI21X1_3783 ( .A(u2__abc_52138_new_n15312_), .B(u2__abc_52138_new_n15310_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15313_));
OAI21X1 OAI21X1_3784 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_293_), .Y(u2__abc_52138_new_n15317_));
OAI21X1 OAI21X1_3785 ( .A(u2__abc_52138_new_n15319_), .B(u2__abc_52138_new_n15318_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15320_));
OAI21X1 OAI21X1_3786 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_294_), .Y(u2__abc_52138_new_n15324_));
OAI21X1 OAI21X1_3787 ( .A(u2__abc_52138_new_n15326_), .B(u2__abc_52138_new_n15327_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15328_));
OAI21X1 OAI21X1_3788 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_295_), .Y(u2__abc_52138_new_n15332_));
OAI21X1 OAI21X1_3789 ( .A(u2__abc_52138_new_n15333_), .B(u2__abc_52138_new_n15335_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15336_));
OAI21X1 OAI21X1_379 ( .A(u2__abc_52138_new_n4292_), .B(u2__abc_52138_new_n4298_), .C(u2__abc_52138_new_n4297_), .Y(u2__abc_52138_new_n4901_));
OAI21X1 OAI21X1_3790 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_296_), .Y(u2__abc_52138_new_n15340_));
OAI21X1 OAI21X1_3791 ( .A(u2__abc_52138_new_n15343_), .B(u2__abc_52138_new_n15341_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15344_));
OAI21X1 OAI21X1_3792 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_297_), .Y(u2__abc_52138_new_n15348_));
OAI21X1 OAI21X1_3793 ( .A(u2__abc_52138_new_n15350_), .B(u2__abc_52138_new_n15349_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15351_));
OAI21X1 OAI21X1_3794 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_298_), .Y(u2__abc_52138_new_n15355_));
OAI21X1 OAI21X1_3795 ( .A(u2__abc_52138_new_n15357_), .B(u2__abc_52138_new_n15358_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15359_));
OAI21X1 OAI21X1_3796 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_299_), .Y(u2__abc_52138_new_n15363_));
OAI21X1 OAI21X1_3797 ( .A(u2__abc_52138_new_n15364_), .B(u2__abc_52138_new_n15366_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15367_));
OAI21X1 OAI21X1_3798 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_300_), .Y(u2__abc_52138_new_n15371_));
OAI21X1 OAI21X1_3799 ( .A(u2__abc_52138_new_n15374_), .B(u2__abc_52138_new_n15372_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15375_));
OAI21X1 OAI21X1_38 ( .A(aNan), .B(_abc_65734_new_n941_), .C(_abc_65734_new_n942_), .Y(\o[149] ));
OAI21X1 OAI21X1_380 ( .A(u2__abc_52138_new_n4906_), .B(u2__abc_52138_new_n4324_), .C(u2__abc_52138_new_n4904_), .Y(u2__abc_52138_new_n4907_));
OAI21X1 OAI21X1_3800 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_301_), .Y(u2__abc_52138_new_n15379_));
OAI21X1 OAI21X1_3801 ( .A(u2__abc_52138_new_n15381_), .B(u2__abc_52138_new_n15380_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15382_));
OAI21X1 OAI21X1_3802 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_302_), .Y(u2__abc_52138_new_n15386_));
OAI21X1 OAI21X1_3803 ( .A(u2__abc_52138_new_n15388_), .B(u2__abc_52138_new_n15389_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15390_));
OAI21X1 OAI21X1_3804 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_303_), .Y(u2__abc_52138_new_n15394_));
OAI21X1 OAI21X1_3805 ( .A(u2__abc_52138_new_n15395_), .B(u2__abc_52138_new_n15397_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15398_));
OAI21X1 OAI21X1_3806 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_304_), .Y(u2__abc_52138_new_n15402_));
OAI21X1 OAI21X1_3807 ( .A(u2__abc_52138_new_n15404_), .B(u2__abc_52138_new_n15405_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15406_));
OAI21X1 OAI21X1_3808 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_305_), .Y(u2__abc_52138_new_n15410_));
OAI21X1 OAI21X1_3809 ( .A(u2__abc_52138_new_n15412_), .B(u2__abc_52138_new_n15411_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15413_));
OAI21X1 OAI21X1_381 ( .A(u2__abc_52138_new_n4330_), .B(u2__abc_52138_new_n4896_), .C(u2__abc_52138_new_n4912_), .Y(u2__abc_52138_new_n4913_));
OAI21X1 OAI21X1_3810 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_306_), .Y(u2__abc_52138_new_n15417_));
OAI21X1 OAI21X1_3811 ( .A(u2__abc_52138_new_n15419_), .B(u2__abc_52138_new_n15420_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15421_));
OAI21X1 OAI21X1_3812 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_307_), .Y(u2__abc_52138_new_n15425_));
OAI21X1 OAI21X1_3813 ( .A(u2__abc_52138_new_n15426_), .B(u2__abc_52138_new_n15428_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15429_));
OAI21X1 OAI21X1_3814 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_308_), .Y(u2__abc_52138_new_n15433_));
OAI21X1 OAI21X1_3815 ( .A(u2__abc_52138_new_n15436_), .B(u2__abc_52138_new_n15434_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15437_));
OAI21X1 OAI21X1_3816 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_309_), .Y(u2__abc_52138_new_n15441_));
OAI21X1 OAI21X1_3817 ( .A(u2__abc_52138_new_n15443_), .B(u2__abc_52138_new_n15442_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15444_));
OAI21X1 OAI21X1_3818 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_310_), .Y(u2__abc_52138_new_n15448_));
OAI21X1 OAI21X1_3819 ( .A(u2__abc_52138_new_n15450_), .B(u2__abc_52138_new_n15451_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15452_));
OAI21X1 OAI21X1_382 ( .A(u2__abc_52138_new_n4916_), .B(u2__abc_52138_new_n4251_), .C(u2__abc_52138_new_n4919_), .Y(u2__abc_52138_new_n4920_));
OAI21X1 OAI21X1_3820 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_311_), .Y(u2__abc_52138_new_n15456_));
OAI21X1 OAI21X1_3821 ( .A(u2__abc_52138_new_n15457_), .B(u2__abc_52138_new_n15459_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15460_));
OAI21X1 OAI21X1_3822 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_312_), .Y(u2__abc_52138_new_n15464_));
OAI21X1 OAI21X1_3823 ( .A(u2__abc_52138_new_n15466_), .B(u2__abc_52138_new_n15467_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15468_));
OAI21X1 OAI21X1_3824 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_313_), .Y(u2__abc_52138_new_n15472_));
OAI21X1 OAI21X1_3825 ( .A(u2__abc_52138_new_n15474_), .B(u2__abc_52138_new_n15473_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15475_));
OAI21X1 OAI21X1_3826 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_314_), .Y(u2__abc_52138_new_n15479_));
OAI21X1 OAI21X1_3827 ( .A(u2__abc_52138_new_n15481_), .B(u2__abc_52138_new_n15482_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15483_));
OAI21X1 OAI21X1_3828 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_315_), .Y(u2__abc_52138_new_n15488_));
OAI21X1 OAI21X1_3829 ( .A(u2__abc_52138_new_n15489_), .B(u2__abc_52138_new_n15491_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15492_));
OAI21X1 OAI21X1_383 ( .A(sqrto_213_), .B(u2__abc_52138_new_n4269_), .C(u2__abc_52138_new_n4267_), .Y(u2__abc_52138_new_n4924_));
OAI21X1 OAI21X1_3830 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_316_), .Y(u2__abc_52138_new_n15496_));
OAI21X1 OAI21X1_3831 ( .A(u2__abc_52138_new_n15498_), .B(u2__abc_52138_new_n15499_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15500_));
OAI21X1 OAI21X1_3832 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_317_), .Y(u2__abc_52138_new_n15504_));
OAI21X1 OAI21X1_3833 ( .A(u2__abc_52138_new_n15506_), .B(u2__abc_52138_new_n15505_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15507_));
OAI21X1 OAI21X1_3834 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_318_), .Y(u2__abc_52138_new_n15511_));
OAI21X1 OAI21X1_3835 ( .A(u2__abc_52138_new_n15513_), .B(u2__abc_52138_new_n15514_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15515_));
OAI21X1 OAI21X1_3836 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_319_), .Y(u2__abc_52138_new_n15519_));
OAI21X1 OAI21X1_3837 ( .A(u2__abc_52138_new_n15520_), .B(u2__abc_52138_new_n15522_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15523_));
OAI21X1 OAI21X1_3838 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_320_), .Y(u2__abc_52138_new_n15527_));
OAI21X1 OAI21X1_3839 ( .A(u2__abc_52138_new_n15529_), .B(u2__abc_52138_new_n15530_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15531_));
OAI21X1 OAI21X1_384 ( .A(u2__abc_52138_new_n4922_), .B(u2__abc_52138_new_n4274_), .C(u2__abc_52138_new_n4925_), .Y(u2__abc_52138_new_n4926_));
OAI21X1 OAI21X1_3840 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_321_), .Y(u2__abc_52138_new_n15535_));
OAI21X1 OAI21X1_3841 ( .A(u2__abc_52138_new_n15537_), .B(u2__abc_52138_new_n15536_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15538_));
OAI21X1 OAI21X1_3842 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_322_), .Y(u2__abc_52138_new_n15542_));
OAI21X1 OAI21X1_3843 ( .A(u2__abc_52138_new_n15544_), .B(u2__abc_52138_new_n15545_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15546_));
OAI21X1 OAI21X1_3844 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_323_), .Y(u2__abc_52138_new_n15550_));
OAI21X1 OAI21X1_3845 ( .A(u2__abc_52138_new_n15551_), .B(u2__abc_52138_new_n15553_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15554_));
OAI21X1 OAI21X1_3846 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_324_), .Y(u2__abc_52138_new_n15558_));
OAI21X1 OAI21X1_3847 ( .A(u2__abc_52138_new_n15561_), .B(u2__abc_52138_new_n15559_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15562_));
OAI21X1 OAI21X1_3848 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_325_), .Y(u2__abc_52138_new_n15566_));
OAI21X1 OAI21X1_3849 ( .A(u2__abc_52138_new_n15568_), .B(u2__abc_52138_new_n15567_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15569_));
OAI21X1 OAI21X1_385 ( .A(u2__abc_52138_new_n4208_), .B(u2__abc_52138_new_n4214_), .C(u2__abc_52138_new_n4213_), .Y(u2__abc_52138_new_n4929_));
OAI21X1 OAI21X1_3850 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_326_), .Y(u2__abc_52138_new_n15573_));
OAI21X1 OAI21X1_3851 ( .A(u2__abc_52138_new_n15575_), .B(u2__abc_52138_new_n15576_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15577_));
OAI21X1 OAI21X1_3852 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_327_), .Y(u2__abc_52138_new_n15581_));
OAI21X1 OAI21X1_3853 ( .A(u2__abc_52138_new_n15582_), .B(u2__abc_52138_new_n15584_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15585_));
OAI21X1 OAI21X1_3854 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_328_), .Y(u2__abc_52138_new_n15589_));
OAI21X1 OAI21X1_3855 ( .A(u2__abc_52138_new_n15592_), .B(u2__abc_52138_new_n15590_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15593_));
OAI21X1 OAI21X1_3856 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_329_), .Y(u2__abc_52138_new_n15597_));
OAI21X1 OAI21X1_3857 ( .A(u2__abc_52138_new_n15599_), .B(u2__abc_52138_new_n15598_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15600_));
OAI21X1 OAI21X1_3858 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_330_), .Y(u2__abc_52138_new_n15604_));
OAI21X1 OAI21X1_3859 ( .A(u2__abc_52138_new_n15606_), .B(u2__abc_52138_new_n15607_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15608_));
OAI21X1 OAI21X1_386 ( .A(u2__abc_52138_new_n4197_), .B(u2__abc_52138_new_n4203_), .C(u2__abc_52138_new_n4202_), .Y(u2__abc_52138_new_n4931_));
OAI21X1 OAI21X1_3860 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_331_), .Y(u2__abc_52138_new_n15612_));
OAI21X1 OAI21X1_3861 ( .A(u2__abc_52138_new_n15613_), .B(u2__abc_52138_new_n15615_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15616_));
OAI21X1 OAI21X1_3862 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_332_), .Y(u2__abc_52138_new_n15620_));
OAI21X1 OAI21X1_3863 ( .A(u2__abc_52138_new_n15623_), .B(u2__abc_52138_new_n15621_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15624_));
OAI21X1 OAI21X1_3864 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_333_), .Y(u2__abc_52138_new_n15628_));
OAI21X1 OAI21X1_3865 ( .A(u2__abc_52138_new_n15630_), .B(u2__abc_52138_new_n15629_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15631_));
OAI21X1 OAI21X1_3866 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_334_), .Y(u2__abc_52138_new_n15635_));
OAI21X1 OAI21X1_3867 ( .A(u2__abc_52138_new_n15637_), .B(u2__abc_52138_new_n15638_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15639_));
OAI21X1 OAI21X1_3868 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_335_), .Y(u2__abc_52138_new_n15644_));
OAI21X1 OAI21X1_3869 ( .A(u2__abc_52138_new_n15645_), .B(u2__abc_52138_new_n15647_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15648_));
OAI21X1 OAI21X1_387 ( .A(u2__abc_52138_new_n4220_), .B(u2__abc_52138_new_n4935_), .C(u2__abc_52138_new_n4225_), .Y(u2__abc_52138_new_n4936_));
OAI21X1 OAI21X1_3870 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_336_), .Y(u2__abc_52138_new_n15652_));
OAI21X1 OAI21X1_3871 ( .A(u2__abc_52138_new_n15654_), .B(u2__abc_52138_new_n15655_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15656_));
OAI21X1 OAI21X1_3872 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_337_), .Y(u2__abc_52138_new_n15660_));
OAI21X1 OAI21X1_3873 ( .A(u2__abc_52138_new_n15662_), .B(u2__abc_52138_new_n15661_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15663_));
OAI21X1 OAI21X1_3874 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_338_), .Y(u2__abc_52138_new_n15667_));
OAI21X1 OAI21X1_3875 ( .A(u2__abc_52138_new_n15669_), .B(u2__abc_52138_new_n15670_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15671_));
OAI21X1 OAI21X1_3876 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_339_), .Y(u2__abc_52138_new_n15676_));
OAI21X1 OAI21X1_3877 ( .A(u2__abc_52138_new_n15677_), .B(u2__abc_52138_new_n15679_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15680_));
OAI21X1 OAI21X1_3878 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_340_), .Y(u2__abc_52138_new_n15684_));
OAI21X1 OAI21X1_3879 ( .A(u2__abc_52138_new_n15687_), .B(u2__abc_52138_new_n15685_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15688_));
OAI21X1 OAI21X1_388 ( .A(u2__abc_52138_new_n4236_), .B(u2__abc_52138_new_n4229_), .C(u2__abc_52138_new_n4937_), .Y(u2__abc_52138_new_n4938_));
OAI21X1 OAI21X1_3880 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_341_), .Y(u2__abc_52138_new_n15692_));
OAI21X1 OAI21X1_3881 ( .A(u2__abc_52138_new_n15694_), .B(u2__abc_52138_new_n15693_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15695_));
OAI21X1 OAI21X1_3882 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_342_), .Y(u2__abc_52138_new_n15699_));
OAI21X1 OAI21X1_3883 ( .A(u2__abc_52138_new_n15701_), .B(u2__abc_52138_new_n15702_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15703_));
OAI21X1 OAI21X1_3884 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_343_), .Y(u2__abc_52138_new_n15707_));
OAI21X1 OAI21X1_3885 ( .A(u2__abc_52138_new_n15708_), .B(u2__abc_52138_new_n15710_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15711_));
OAI21X1 OAI21X1_3886 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_344_), .Y(u2__abc_52138_new_n15715_));
OAI21X1 OAI21X1_3887 ( .A(u2__abc_52138_new_n15717_), .B(u2__abc_52138_new_n15718_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15719_));
OAI21X1 OAI21X1_3888 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_345_), .Y(u2__abc_52138_new_n15723_));
OAI21X1 OAI21X1_3889 ( .A(u2__abc_52138_new_n15725_), .B(u2__abc_52138_new_n15724_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15726_));
OAI21X1 OAI21X1_389 ( .A(u2__abc_52138_new_n4240_), .B(u2__abc_52138_new_n4927_), .C(u2__abc_52138_new_n4941_), .Y(u2__abc_52138_new_n4942_));
OAI21X1 OAI21X1_3890 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_346_), .Y(u2__abc_52138_new_n15730_));
OAI21X1 OAI21X1_3891 ( .A(u2__abc_52138_new_n15732_), .B(u2__abc_52138_new_n15733_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15734_));
OAI21X1 OAI21X1_3892 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_347_), .Y(u2__abc_52138_new_n15738_));
OAI21X1 OAI21X1_3893 ( .A(u2__abc_52138_new_n15739_), .B(u2__abc_52138_new_n15741_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15742_));
OAI21X1 OAI21X1_3894 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_348_), .Y(u2__abc_52138_new_n15746_));
OAI21X1 OAI21X1_3895 ( .A(u2__abc_52138_new_n15748_), .B(u2__abc_52138_new_n15749_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15750_));
OAI21X1 OAI21X1_3896 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_349_), .Y(u2__abc_52138_new_n15754_));
OAI21X1 OAI21X1_3897 ( .A(u2__abc_52138_new_n15756_), .B(u2__abc_52138_new_n15755_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15757_));
OAI21X1 OAI21X1_3898 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_350_), .Y(u2__abc_52138_new_n15761_));
OAI21X1 OAI21X1_3899 ( .A(u2__abc_52138_new_n15763_), .B(u2__abc_52138_new_n15764_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15765_));
OAI21X1 OAI21X1_39 ( .A(aNan), .B(_abc_65734_new_n944_), .C(_abc_65734_new_n945_), .Y(\o[150] ));
OAI21X1 OAI21X1_390 ( .A(u2__abc_52138_new_n4165_), .B(u2__abc_52138_new_n4945_), .C(u2__abc_52138_new_n4160_), .Y(u2__abc_52138_new_n4946_));
OAI21X1 OAI21X1_3900 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_351_), .Y(u2__abc_52138_new_n15769_));
OAI21X1 OAI21X1_3901 ( .A(u2__abc_52138_new_n15770_), .B(u2__abc_52138_new_n15772_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15773_));
OAI21X1 OAI21X1_3902 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_352_), .Y(u2__abc_52138_new_n15777_));
OAI21X1 OAI21X1_3903 ( .A(u2__abc_52138_new_n15779_), .B(u2__abc_52138_new_n15780_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15781_));
OAI21X1 OAI21X1_3904 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_353_), .Y(u2__abc_52138_new_n15785_));
OAI21X1 OAI21X1_3905 ( .A(u2__abc_52138_new_n15787_), .B(u2__abc_52138_new_n15786_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15788_));
OAI21X1 OAI21X1_3906 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_354_), .Y(u2__abc_52138_new_n15792_));
OAI21X1 OAI21X1_3907 ( .A(u2__abc_52138_new_n15794_), .B(u2__abc_52138_new_n15795_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15796_));
OAI21X1 OAI21X1_3908 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_355_), .Y(u2__abc_52138_new_n15800_));
OAI21X1 OAI21X1_3909 ( .A(u2__abc_52138_new_n15801_), .B(u2__abc_52138_new_n15803_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15804_));
OAI21X1 OAI21X1_391 ( .A(u2__abc_52138_new_n4149_), .B(u2__abc_52138_new_n4155_), .C(u2__abc_52138_new_n4154_), .Y(u2__abc_52138_new_n4948_));
OAI21X1 OAI21X1_3910 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_356_), .Y(u2__abc_52138_new_n15808_));
OAI21X1 OAI21X1_3911 ( .A(u2__abc_52138_new_n15811_), .B(u2__abc_52138_new_n15809_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15812_));
OAI21X1 OAI21X1_3912 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_357_), .Y(u2__abc_52138_new_n15816_));
OAI21X1 OAI21X1_3913 ( .A(u2__abc_52138_new_n15818_), .B(u2__abc_52138_new_n15817_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15819_));
OAI21X1 OAI21X1_3914 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_358_), .Y(u2__abc_52138_new_n15823_));
OAI21X1 OAI21X1_3915 ( .A(u2__abc_52138_new_n15825_), .B(u2__abc_52138_new_n15826_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15827_));
OAI21X1 OAI21X1_3916 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_359_), .Y(u2__abc_52138_new_n15831_));
OAI21X1 OAI21X1_3917 ( .A(u2__abc_52138_new_n15832_), .B(u2__abc_52138_new_n15834_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15835_));
OAI21X1 OAI21X1_3918 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_360_), .Y(u2__abc_52138_new_n15839_));
OAI21X1 OAI21X1_3919 ( .A(u2__abc_52138_new_n15841_), .B(u2__abc_52138_new_n15842_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15843_));
OAI21X1 OAI21X1_392 ( .A(u2_o_227_), .B(u2__abc_52138_new_n4180_), .C(u2__abc_52138_new_n4188_), .Y(u2__abc_52138_new_n4951_));
OAI21X1 OAI21X1_3920 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_361_), .Y(u2__abc_52138_new_n15847_));
OAI21X1 OAI21X1_3921 ( .A(u2__abc_52138_new_n15849_), .B(u2__abc_52138_new_n15848_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15850_));
OAI21X1 OAI21X1_3922 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_362_), .Y(u2__abc_52138_new_n15854_));
OAI21X1 OAI21X1_3923 ( .A(u2__abc_52138_new_n15856_), .B(u2__abc_52138_new_n15857_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15858_));
OAI21X1 OAI21X1_3924 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_363_), .Y(u2__abc_52138_new_n15862_));
OAI21X1 OAI21X1_3925 ( .A(u2__abc_52138_new_n15863_), .B(u2__abc_52138_new_n15865_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15866_));
OAI21X1 OAI21X1_3926 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_364_), .Y(u2__abc_52138_new_n15870_));
OAI21X1 OAI21X1_3927 ( .A(u2__abc_52138_new_n15872_), .B(u2__abc_52138_new_n15873_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15874_));
OAI21X1 OAI21X1_3928 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_365_), .Y(u2__abc_52138_new_n15878_));
OAI21X1 OAI21X1_3929 ( .A(u2__abc_52138_new_n15880_), .B(u2__abc_52138_new_n15879_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15881_));
OAI21X1 OAI21X1_393 ( .A(u2__abc_52138_new_n4182_), .B(u2_remHi_227_), .C(u2__abc_52138_new_n4951_), .Y(u2__abc_52138_new_n4952_));
OAI21X1 OAI21X1_3930 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_366_), .Y(u2__abc_52138_new_n15885_));
OAI21X1 OAI21X1_3931 ( .A(u2__abc_52138_new_n15887_), .B(u2__abc_52138_new_n15888_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15889_));
OAI21X1 OAI21X1_3932 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_367_), .Y(u2__abc_52138_new_n15893_));
OAI21X1 OAI21X1_3933 ( .A(u2__abc_52138_new_n15894_), .B(u2__abc_52138_new_n15896_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15897_));
OAI21X1 OAI21X1_3934 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_368_), .Y(u2__abc_52138_new_n15901_));
OAI21X1 OAI21X1_3935 ( .A(u2__abc_52138_new_n15903_), .B(u2__abc_52138_new_n15904_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15905_));
OAI21X1 OAI21X1_3936 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_369_), .Y(u2__abc_52138_new_n15909_));
OAI21X1 OAI21X1_3937 ( .A(u2__abc_52138_new_n15911_), .B(u2__abc_52138_new_n15910_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15912_));
OAI21X1 OAI21X1_3938 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_370_), .Y(u2__abc_52138_new_n15917_));
OAI21X1 OAI21X1_3939 ( .A(u2__abc_52138_new_n15919_), .B(u2__abc_52138_new_n15920_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15921_));
OAI21X1 OAI21X1_394 ( .A(u2__abc_52138_new_n4172_), .B(u2__abc_52138_new_n4954_), .C(u2__abc_52138_new_n4177_), .Y(u2__abc_52138_new_n4955_));
OAI21X1 OAI21X1_3940 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_371_), .Y(u2__abc_52138_new_n15925_));
OAI21X1 OAI21X1_3941 ( .A(u2__abc_52138_new_n15926_), .B(u2__abc_52138_new_n15928_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15929_));
OAI21X1 OAI21X1_3942 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_372_), .Y(u2__abc_52138_new_n15933_));
OAI21X1 OAI21X1_3943 ( .A(u2__abc_52138_new_n15935_), .B(u2__abc_52138_new_n15936_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15937_));
OAI21X1 OAI21X1_3944 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_373_), .Y(u2__abc_52138_new_n15941_));
OAI21X1 OAI21X1_3945 ( .A(u2__abc_52138_new_n15943_), .B(u2__abc_52138_new_n15942_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15944_));
OAI21X1 OAI21X1_3946 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_374_), .Y(u2__abc_52138_new_n15948_));
OAI21X1 OAI21X1_3947 ( .A(u2__abc_52138_new_n15950_), .B(u2__abc_52138_new_n15951_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15952_));
OAI21X1 OAI21X1_3948 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_375_), .Y(u2__abc_52138_new_n15956_));
OAI21X1 OAI21X1_3949 ( .A(u2__abc_52138_new_n15957_), .B(u2__abc_52138_new_n15959_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15960_));
OAI21X1 OAI21X1_395 ( .A(u2_o_231_), .B(u2__abc_52138_new_n4134_), .C(u2__abc_52138_new_n4141_), .Y(u2__abc_52138_new_n4961_));
OAI21X1 OAI21X1_3950 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_376_), .Y(u2__abc_52138_new_n15964_));
OAI21X1 OAI21X1_3951 ( .A(u2__abc_52138_new_n15966_), .B(u2__abc_52138_new_n15967_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15968_));
OAI21X1 OAI21X1_3952 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_377_), .Y(u2__abc_52138_new_n15972_));
OAI21X1 OAI21X1_3953 ( .A(u2__abc_52138_new_n15974_), .B(u2__abc_52138_new_n15973_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15975_));
OAI21X1 OAI21X1_3954 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_378_), .Y(u2__abc_52138_new_n15979_));
OAI21X1 OAI21X1_3955 ( .A(u2__abc_52138_new_n15981_), .B(u2__abc_52138_new_n15982_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15983_));
OAI21X1 OAI21X1_3956 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_379_), .Y(u2__abc_52138_new_n15987_));
OAI21X1 OAI21X1_3957 ( .A(u2__abc_52138_new_n15988_), .B(u2__abc_52138_new_n15990_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15991_));
OAI21X1 OAI21X1_3958 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_380_), .Y(u2__abc_52138_new_n15995_));
OAI21X1 OAI21X1_3959 ( .A(u2__abc_52138_new_n15997_), .B(u2__abc_52138_new_n15998_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n15999_));
OAI21X1 OAI21X1_396 ( .A(u2__abc_52138_new_n4960_), .B(u2_remHi_231_), .C(u2__abc_52138_new_n4961_), .Y(u2__abc_52138_new_n4962_));
OAI21X1 OAI21X1_3960 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_381_), .Y(u2__abc_52138_new_n16003_));
OAI21X1 OAI21X1_3961 ( .A(u2__abc_52138_new_n16005_), .B(u2__abc_52138_new_n16004_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16006_));
OAI21X1 OAI21X1_3962 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_382_), .Y(u2__abc_52138_new_n16010_));
OAI21X1 OAI21X1_3963 ( .A(u2__abc_52138_new_n16012_), .B(u2__abc_52138_new_n16013_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16014_));
OAI21X1 OAI21X1_3964 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_383_), .Y(u2__abc_52138_new_n16018_));
OAI21X1 OAI21X1_3965 ( .A(u2__abc_52138_new_n16019_), .B(u2__abc_52138_new_n16021_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16022_));
OAI21X1 OAI21X1_3966 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_384_), .Y(u2__abc_52138_new_n16026_));
OAI21X1 OAI21X1_3967 ( .A(u2__abc_52138_new_n16028_), .B(u2__abc_52138_new_n16029_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16030_));
OAI21X1 OAI21X1_3968 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_385_), .Y(u2__abc_52138_new_n16034_));
OAI21X1 OAI21X1_3969 ( .A(u2__abc_52138_new_n16036_), .B(u2__abc_52138_new_n16035_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16037_));
OAI21X1 OAI21X1_397 ( .A(u2__abc_52138_new_n4126_), .B(u2__abc_52138_new_n4132_), .C(u2__abc_52138_new_n4131_), .Y(u2__abc_52138_new_n4963_));
OAI21X1 OAI21X1_3970 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_386_), .Y(u2__abc_52138_new_n16041_));
OAI21X1 OAI21X1_3971 ( .A(u2__abc_52138_new_n16043_), .B(u2__abc_52138_new_n16044_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16045_));
OAI21X1 OAI21X1_3972 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_387_), .Y(u2__abc_52138_new_n16049_));
OAI21X1 OAI21X1_3973 ( .A(u2__abc_52138_new_n16050_), .B(u2__abc_52138_new_n16052_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16053_));
OAI21X1 OAI21X1_3974 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_388_), .Y(u2__abc_52138_new_n16057_));
OAI21X1 OAI21X1_3975 ( .A(u2__abc_52138_new_n16060_), .B(u2__abc_52138_new_n16058_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16061_));
OAI21X1 OAI21X1_3976 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_389_), .Y(u2__abc_52138_new_n16065_));
OAI21X1 OAI21X1_3977 ( .A(u2__abc_52138_new_n16067_), .B(u2__abc_52138_new_n16066_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16068_));
OAI21X1 OAI21X1_3978 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_390_), .Y(u2__abc_52138_new_n16072_));
OAI21X1 OAI21X1_3979 ( .A(u2__abc_52138_new_n16074_), .B(u2__abc_52138_new_n16075_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16076_));
OAI21X1 OAI21X1_398 ( .A(u2__abc_52138_new_n4118_), .B(u2__abc_52138_new_n4114_), .C(u2__abc_52138_new_n4113_), .Y(u2__abc_52138_new_n4965_));
OAI21X1 OAI21X1_3980 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_391_), .Y(u2__abc_52138_new_n16081_));
OAI21X1 OAI21X1_3981 ( .A(u2__abc_52138_new_n16082_), .B(u2__abc_52138_new_n16084_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16085_));
OAI21X1 OAI21X1_3982 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_392_), .Y(u2__abc_52138_new_n16090_));
OAI21X1 OAI21X1_3983 ( .A(u2__abc_52138_new_n16093_), .B(u2__abc_52138_new_n16091_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16094_));
OAI21X1 OAI21X1_3984 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_393_), .Y(u2__abc_52138_new_n16098_));
OAI21X1 OAI21X1_3985 ( .A(u2__abc_52138_new_n16100_), .B(u2__abc_52138_new_n16099_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16101_));
OAI21X1 OAI21X1_3986 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_394_), .Y(u2__abc_52138_new_n16105_));
OAI21X1 OAI21X1_3987 ( .A(u2__abc_52138_new_n16107_), .B(u2__abc_52138_new_n16108_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16109_));
OAI21X1 OAI21X1_3988 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_395_), .Y(u2__abc_52138_new_n16114_));
OAI21X1 OAI21X1_3989 ( .A(u2__abc_52138_new_n16115_), .B(u2__abc_52138_new_n16117_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16118_));
OAI21X1 OAI21X1_399 ( .A(u2__abc_52138_new_n4102_), .B(u2__abc_52138_new_n4108_), .C(u2__abc_52138_new_n4107_), .Y(u2__abc_52138_new_n4966_));
OAI21X1 OAI21X1_3990 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_396_), .Y(u2__abc_52138_new_n16122_));
OAI21X1 OAI21X1_3991 ( .A(u2__abc_52138_new_n16125_), .B(u2__abc_52138_new_n16123_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16126_));
OAI21X1 OAI21X1_3992 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_397_), .Y(u2__abc_52138_new_n16130_));
OAI21X1 OAI21X1_3993 ( .A(u2__abc_52138_new_n16132_), .B(u2__abc_52138_new_n16131_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16133_));
OAI21X1 OAI21X1_3994 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_398_), .Y(u2__abc_52138_new_n16137_));
OAI21X1 OAI21X1_3995 ( .A(u2__abc_52138_new_n16139_), .B(u2__abc_52138_new_n16140_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16141_));
OAI21X1 OAI21X1_3996 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_399_), .Y(u2__abc_52138_new_n16145_));
OAI21X1 OAI21X1_3997 ( .A(u2__abc_52138_new_n16146_), .B(u2__abc_52138_new_n16148_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16149_));
OAI21X1 OAI21X1_3998 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_400_), .Y(u2__abc_52138_new_n16153_));
OAI21X1 OAI21X1_3999 ( .A(u2__abc_52138_new_n16155_), .B(u2__abc_52138_new_n16156_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16157_));
OAI21X1 OAI21X1_4 ( .A(aNan), .B(_abc_65734_new_n839_), .C(_abc_65734_new_n840_), .Y(\o[115] ));
OAI21X1 OAI21X1_40 ( .A(aNan), .B(_abc_65734_new_n947_), .C(_abc_65734_new_n948_), .Y(\o[151] ));
OAI21X1 OAI21X1_400 ( .A(u2__abc_52138_new_n4121_), .B(u2__abc_52138_new_n4964_), .C(u2__abc_52138_new_n4967_), .Y(u2__abc_52138_new_n4968_));
OAI21X1 OAI21X1_4000 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_401_), .Y(u2__abc_52138_new_n16161_));
OAI21X1 OAI21X1_4001 ( .A(u2__abc_52138_new_n16163_), .B(u2__abc_52138_new_n16162_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16164_));
OAI21X1 OAI21X1_4002 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_402_), .Y(u2__abc_52138_new_n16168_));
OAI21X1 OAI21X1_4003 ( .A(u2__abc_52138_new_n16170_), .B(u2__abc_52138_new_n16171_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16172_));
OAI21X1 OAI21X1_4004 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_403_), .Y(u2__abc_52138_new_n16176_));
OAI21X1 OAI21X1_4005 ( .A(u2__abc_52138_new_n16177_), .B(u2__abc_52138_new_n16179_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16180_));
OAI21X1 OAI21X1_4006 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_404_), .Y(u2__abc_52138_new_n16184_));
OAI21X1 OAI21X1_4007 ( .A(u2__abc_52138_new_n16187_), .B(u2__abc_52138_new_n16185_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16188_));
OAI21X1 OAI21X1_4008 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_405_), .Y(u2__abc_52138_new_n16192_));
OAI21X1 OAI21X1_4009 ( .A(u2__abc_52138_new_n16194_), .B(u2__abc_52138_new_n16193_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16195_));
OAI21X1 OAI21X1_401 ( .A(u2__abc_52138_new_n4145_), .B(u2__abc_52138_new_n4958_), .C(u2__abc_52138_new_n4969_), .Y(u2__abc_52138_new_n4970_));
OAI21X1 OAI21X1_4010 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_406_), .Y(u2__abc_52138_new_n16199_));
OAI21X1 OAI21X1_4011 ( .A(u2__abc_52138_new_n16201_), .B(u2__abc_52138_new_n16202_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16203_));
OAI21X1 OAI21X1_4012 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_407_), .Y(u2__abc_52138_new_n16207_));
OAI21X1 OAI21X1_4013 ( .A(u2__abc_52138_new_n16208_), .B(u2__abc_52138_new_n16210_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16211_));
OAI21X1 OAI21X1_4014 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_408_), .Y(u2__abc_52138_new_n16215_));
OAI21X1 OAI21X1_4015 ( .A(u2__abc_52138_new_n16217_), .B(u2__abc_52138_new_n16218_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16219_));
OAI21X1 OAI21X1_4016 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_409_), .Y(u2__abc_52138_new_n16223_));
OAI21X1 OAI21X1_4017 ( .A(u2__abc_52138_new_n16225_), .B(u2__abc_52138_new_n16224_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16226_));
OAI21X1 OAI21X1_4018 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_410_), .Y(u2__abc_52138_new_n16230_));
OAI21X1 OAI21X1_4019 ( .A(u2__abc_52138_new_n16232_), .B(u2__abc_52138_new_n16233_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16234_));
OAI21X1 OAI21X1_402 ( .A(u2__abc_52138_new_n4006_), .B(u2__abc_52138_new_n4012_), .C(u2__abc_52138_new_n4011_), .Y(u2__abc_52138_new_n4972_));
OAI21X1 OAI21X1_4020 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_411_), .Y(u2__abc_52138_new_n16238_));
OAI21X1 OAI21X1_4021 ( .A(u2__abc_52138_new_n16239_), .B(u2__abc_52138_new_n16241_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16242_));
OAI21X1 OAI21X1_4022 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_412_), .Y(u2__abc_52138_new_n16246_));
OAI21X1 OAI21X1_4023 ( .A(u2__abc_52138_new_n16248_), .B(u2__abc_52138_new_n16249_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16250_));
OAI21X1 OAI21X1_4024 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_413_), .Y(u2__abc_52138_new_n16254_));
OAI21X1 OAI21X1_4025 ( .A(u2__abc_52138_new_n16256_), .B(u2__abc_52138_new_n16255_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16257_));
OAI21X1 OAI21X1_4026 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_414_), .Y(u2__abc_52138_new_n16261_));
OAI21X1 OAI21X1_4027 ( .A(u2__abc_52138_new_n16263_), .B(u2__abc_52138_new_n16264_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16265_));
OAI21X1 OAI21X1_4028 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_415_), .Y(u2__abc_52138_new_n16269_));
OAI21X1 OAI21X1_4029 ( .A(u2__abc_52138_new_n16270_), .B(u2__abc_52138_new_n16272_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16273_));
OAI21X1 OAI21X1_403 ( .A(u2__abc_52138_new_n4017_), .B(u2__abc_52138_new_n4023_), .C(u2__abc_52138_new_n4022_), .Y(u2__abc_52138_new_n4974_));
OAI21X1 OAI21X1_4030 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_416_), .Y(u2__abc_52138_new_n16277_));
OAI21X1 OAI21X1_4031 ( .A(u2__abc_52138_new_n16279_), .B(u2__abc_52138_new_n16280_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16281_));
OAI21X1 OAI21X1_4032 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_417_), .Y(u2__abc_52138_new_n16285_));
OAI21X1 OAI21X1_4033 ( .A(u2__abc_52138_new_n16287_), .B(u2__abc_52138_new_n16286_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16288_));
OAI21X1 OAI21X1_4034 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_418_), .Y(u2__abc_52138_new_n16292_));
OAI21X1 OAI21X1_4035 ( .A(u2__abc_52138_new_n16294_), .B(u2__abc_52138_new_n16295_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16296_));
OAI21X1 OAI21X1_4036 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_419_), .Y(u2__abc_52138_new_n16300_));
OAI21X1 OAI21X1_4037 ( .A(u2__abc_52138_new_n16301_), .B(u2__abc_52138_new_n16303_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16304_));
OAI21X1 OAI21X1_4038 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_420_), .Y(u2__abc_52138_new_n16308_));
OAI21X1 OAI21X1_4039 ( .A(u2__abc_52138_new_n16311_), .B(u2__abc_52138_new_n16309_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16312_));
OAI21X1 OAI21X1_404 ( .A(u2__abc_52138_new_n4029_), .B(u2__abc_52138_new_n4035_), .C(u2__abc_52138_new_n4032_), .Y(u2__abc_52138_new_n4977_));
OAI21X1 OAI21X1_4040 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_421_), .Y(u2__abc_52138_new_n16316_));
OAI21X1 OAI21X1_4041 ( .A(u2__abc_52138_new_n16318_), .B(u2__abc_52138_new_n16317_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16319_));
OAI21X1 OAI21X1_4042 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_422_), .Y(u2__abc_52138_new_n16323_));
OAI21X1 OAI21X1_4043 ( .A(u2__abc_52138_new_n16325_), .B(u2__abc_52138_new_n16326_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16327_));
OAI21X1 OAI21X1_4044 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_423_), .Y(u2__abc_52138_new_n16331_));
OAI21X1 OAI21X1_4045 ( .A(u2__abc_52138_new_n16332_), .B(u2__abc_52138_new_n16334_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16335_));
OAI21X1 OAI21X1_4046 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_424_), .Y(u2__abc_52138_new_n16339_));
OAI21X1 OAI21X1_4047 ( .A(u2__abc_52138_new_n16341_), .B(u2__abc_52138_new_n16342_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16343_));
OAI21X1 OAI21X1_4048 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_425_), .Y(u2__abc_52138_new_n16347_));
OAI21X1 OAI21X1_4049 ( .A(u2__abc_52138_new_n16349_), .B(u2__abc_52138_new_n16348_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16350_));
OAI21X1 OAI21X1_405 ( .A(u2__abc_52138_new_n4045_), .B(u2__abc_52138_new_n4041_), .C(u2__abc_52138_new_n4040_), .Y(u2__abc_52138_new_n4978_));
OAI21X1 OAI21X1_4050 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_426_), .Y(u2__abc_52138_new_n16354_));
OAI21X1 OAI21X1_4051 ( .A(u2__abc_52138_new_n16356_), .B(u2__abc_52138_new_n16357_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16358_));
OAI21X1 OAI21X1_4052 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_427_), .Y(u2__abc_52138_new_n16362_));
OAI21X1 OAI21X1_4053 ( .A(u2__abc_52138_new_n16363_), .B(u2__abc_52138_new_n16365_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16366_));
OAI21X1 OAI21X1_4054 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_428_), .Y(u2__abc_52138_new_n16370_));
OAI21X1 OAI21X1_4055 ( .A(u2__abc_52138_new_n16372_), .B(u2__abc_52138_new_n16373_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16374_));
OAI21X1 OAI21X1_4056 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_429_), .Y(u2__abc_52138_new_n16378_));
OAI21X1 OAI21X1_4057 ( .A(u2__abc_52138_new_n16380_), .B(u2__abc_52138_new_n16379_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16381_));
OAI21X1 OAI21X1_4058 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_430_), .Y(u2__abc_52138_new_n16385_));
OAI21X1 OAI21X1_4059 ( .A(u2__abc_52138_new_n16387_), .B(u2__abc_52138_new_n16388_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16389_));
OAI21X1 OAI21X1_406 ( .A(u2__abc_52138_new_n4053_), .B(u2__abc_52138_new_n4059_), .C(u2__abc_52138_new_n4058_), .Y(u2__abc_52138_new_n4984_));
OAI21X1 OAI21X1_4060 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_431_), .Y(u2__abc_52138_new_n16393_));
OAI21X1 OAI21X1_4061 ( .A(u2__abc_52138_new_n16394_), .B(u2__abc_52138_new_n16396_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16397_));
OAI21X1 OAI21X1_4062 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_432_), .Y(u2__abc_52138_new_n16401_));
OAI21X1 OAI21X1_4063 ( .A(u2__abc_52138_new_n16403_), .B(u2__abc_52138_new_n16404_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16405_));
OAI21X1 OAI21X1_4064 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_433_), .Y(u2__abc_52138_new_n16409_));
OAI21X1 OAI21X1_4065 ( .A(u2__abc_52138_new_n16411_), .B(u2__abc_52138_new_n16410_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16412_));
OAI21X1 OAI21X1_4066 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_434_), .Y(u2__abc_52138_new_n16416_));
OAI21X1 OAI21X1_4067 ( .A(u2__abc_52138_new_n16418_), .B(u2__abc_52138_new_n16419_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16420_));
OAI21X1 OAI21X1_4068 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_435_), .Y(u2__abc_52138_new_n16424_));
OAI21X1 OAI21X1_4069 ( .A(u2__abc_52138_new_n16425_), .B(u2__abc_52138_new_n16427_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16428_));
OAI21X1 OAI21X1_407 ( .A(u2__abc_52138_new_n4064_), .B(u2__abc_52138_new_n4070_), .C(u2__abc_52138_new_n4069_), .Y(u2__abc_52138_new_n4985_));
OAI21X1 OAI21X1_4070 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_436_), .Y(u2__abc_52138_new_n16432_));
OAI21X1 OAI21X1_4071 ( .A(u2__abc_52138_new_n16434_), .B(u2__abc_52138_new_n16435_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16436_));
OAI21X1 OAI21X1_4072 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_437_), .Y(u2__abc_52138_new_n16440_));
OAI21X1 OAI21X1_4073 ( .A(u2__abc_52138_new_n16442_), .B(u2__abc_52138_new_n16441_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16443_));
OAI21X1 OAI21X1_4074 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_438_), .Y(u2__abc_52138_new_n16447_));
OAI21X1 OAI21X1_4075 ( .A(u2__abc_52138_new_n16449_), .B(u2__abc_52138_new_n16450_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16451_));
OAI21X1 OAI21X1_4076 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_439_), .Y(u2__abc_52138_new_n16455_));
OAI21X1 OAI21X1_4077 ( .A(u2__abc_52138_new_n16456_), .B(u2__abc_52138_new_n16458_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16459_));
OAI21X1 OAI21X1_4078 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_440_), .Y(u2__abc_52138_new_n16463_));
OAI21X1 OAI21X1_4079 ( .A(u2__abc_52138_new_n16465_), .B(u2__abc_52138_new_n16466_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16467_));
OAI21X1 OAI21X1_408 ( .A(u2__abc_52138_new_n4077_), .B(u2__abc_52138_new_n4987_), .C(u2__abc_52138_new_n4082_), .Y(u2__abc_52138_new_n4988_));
OAI21X1 OAI21X1_4080 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_441_), .Y(u2__abc_52138_new_n16471_));
OAI21X1 OAI21X1_4081 ( .A(u2__abc_52138_new_n16473_), .B(u2__abc_52138_new_n16472_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16474_));
OAI21X1 OAI21X1_4082 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_442_), .Y(u2__abc_52138_new_n16478_));
OAI21X1 OAI21X1_4083 ( .A(u2__abc_52138_new_n16480_), .B(u2__abc_52138_new_n16481_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16482_));
OAI21X1 OAI21X1_4084 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_443_), .Y(u2__abc_52138_new_n16486_));
OAI21X1 OAI21X1_4085 ( .A(u2__abc_52138_new_n16487_), .B(u2__abc_52138_new_n16489_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16490_));
OAI21X1 OAI21X1_4086 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_444_), .Y(u2__abc_52138_new_n16494_));
OAI21X1 OAI21X1_4087 ( .A(u2__abc_52138_new_n16496_), .B(u2__abc_52138_new_n16497_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16498_));
OAI21X1 OAI21X1_4088 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_445_), .Y(u2__abc_52138_new_n16502_));
OAI21X1 OAI21X1_4089 ( .A(u2__abc_52138_new_n16504_), .B(u2__abc_52138_new_n16503_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16505_));
OAI21X1 OAI21X1_409 ( .A(u2__abc_52138_new_n4093_), .B(u2__abc_52138_new_n4086_), .C(u2__abc_52138_new_n4989_), .Y(u2__abc_52138_new_n4990_));
OAI21X1 OAI21X1_4090 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_446_), .Y(u2__abc_52138_new_n16509_));
OAI21X1 OAI21X1_4091 ( .A(u2__abc_52138_new_n16511_), .B(u2__abc_52138_new_n16512_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16513_));
OAI21X1 OAI21X1_4092 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_447_), .Y(u2__abc_52138_new_n16517_));
OAI21X1 OAI21X1_4093 ( .A(u2__abc_52138_new_n16518_), .B(u2__abc_52138_new_n16520_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16521_));
OAI21X1 OAI21X1_4094 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_448_), .Y(u2__abc_52138_new_n16525_));
OAI21X1 OAI21X1_4095 ( .A(u2__abc_52138_new_n16528_), .B(u2__abc_52138_new_n16526_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n16529_));
OAI21X1 OAI21X1_4096 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_o_449_), .Y(u2__abc_52138_new_n16533_));
OAI21X1 OAI21X1_4097 ( .A(u2__abc_52138_new_n16535_), .B(u2__abc_52138_new_n16534_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n16536_));
OAI21X1 OAI21X1_41 ( .A(aNan), .B(_abc_65734_new_n950_), .C(_abc_65734_new_n951_), .Y(\o[152] ));
OAI21X1 OAI21X1_410 ( .A(u2__abc_52138_new_n4986_), .B(u2__abc_52138_new_n4983_), .C(u2__abc_52138_new_n4991_), .Y(u2__abc_52138_new_n4992_));
OAI21X1 OAI21X1_411 ( .A(u2__abc_52138_new_n4193_), .B(u2__abc_52138_new_n4943_), .C(u2__abc_52138_new_n4995_), .Y(u2__abc_52138_new_n4996_));
OAI21X1 OAI21X1_412 ( .A(u2__abc_52138_new_n4753_), .B(u2__abc_52138_new_n4002_), .C(u2__abc_52138_new_n4997_), .Y(u2__abc_52138_new_n4998_));
OAI21X1 OAI21X1_413 ( .A(u2_remHi_254_), .B(u2__abc_52138_new_n5687_), .C(u2__abc_52138_new_n5689_), .Y(u2__abc_52138_new_n5690_));
OAI21X1 OAI21X1_414 ( .A(u2__abc_52138_new_n5691_), .B(u2_o_254_), .C(u2__abc_52138_new_n5693_), .Y(u2__abc_52138_new_n5694_));
OAI21X1 OAI21X1_415 ( .A(u2__abc_52138_new_n5688_), .B(u2_o_255_), .C(u2__abc_52138_new_n5690_), .Y(u2__abc_52138_new_n5737_));
OAI21X1 OAI21X1_416 ( .A(u2__abc_52138_new_n5737_), .B(u2__abc_52138_new_n5707_), .C(u2__abc_52138_new_n5739_), .Y(u2__abc_52138_new_n5740_));
OAI21X1 OAI21X1_417 ( .A(u2__abc_52138_new_n5723_), .B(u2__abc_52138_new_n5728_), .C(u2__abc_52138_new_n5741_), .Y(u2__abc_52138_new_n5742_));
OAI21X1 OAI21X1_418 ( .A(u2__abc_52138_new_n5742_), .B(u2__abc_52138_new_n5719_), .C(u2__abc_52138_new_n5743_), .Y(u2__abc_52138_new_n5744_));
OAI21X1 OAI21X1_419 ( .A(u2__abc_52138_new_n5673_), .B(u2__abc_52138_new_n5747_), .C(u2__abc_52138_new_n5748_), .Y(u2__abc_52138_new_n5749_));
OAI21X1 OAI21X1_42 ( .A(aNan), .B(_abc_65734_new_n953_), .C(_abc_65734_new_n954_), .Y(\o[153] ));
OAI21X1 OAI21X1_420 ( .A(u2__abc_52138_new_n5754_), .B(u2__abc_52138_new_n5746_), .C(u2__abc_52138_new_n5638_), .Y(u2__abc_52138_new_n5755_));
OAI21X1 OAI21X1_421 ( .A(u2__abc_52138_new_n5609_), .B(u2__abc_52138_new_n5614_), .C(u2__abc_52138_new_n5756_), .Y(u2__abc_52138_new_n5757_));
OAI21X1 OAI21X1_422 ( .A(u2__abc_52138_new_n5757_), .B(u2__abc_52138_new_n5605_), .C(u2__abc_52138_new_n5758_), .Y(u2__abc_52138_new_n5759_));
OAI21X1 OAI21X1_423 ( .A(u2_remHi_274_), .B(u2__abc_52138_new_n5761_), .C(u2__abc_52138_new_n5762_), .Y(u2__abc_52138_new_n5763_));
OAI21X1 OAI21X1_424 ( .A(u2__abc_52138_new_n5630_), .B(u2_o_275_), .C(u2__abc_52138_new_n5763_), .Y(u2__abc_52138_new_n5764_));
OAI21X1 OAI21X1_425 ( .A(u2__abc_52138_new_n5764_), .B(u2__abc_52138_new_n5628_), .C(u2__abc_52138_new_n5760_), .Y(u2__abc_52138_new_n5765_));
OAI21X1 OAI21X1_426 ( .A(u2__abc_52138_new_n5562_), .B(u2__abc_52138_new_n5567_), .C(u2__abc_52138_new_n5768_), .Y(u2__abc_52138_new_n5769_));
OAI21X1 OAI21X1_427 ( .A(u2__abc_52138_new_n5769_), .B(u2__abc_52138_new_n5558_), .C(u2__abc_52138_new_n5771_), .Y(u2__abc_52138_new_n5772_));
OAI21X1 OAI21X1_428 ( .A(u2__abc_52138_new_n5590_), .B(u2__abc_52138_new_n5775_), .C(u2__abc_52138_new_n5774_), .Y(u2__abc_52138_new_n5776_));
OAI21X1 OAI21X1_429 ( .A(u2__abc_52138_new_n5574_), .B(u2__abc_52138_new_n5579_), .C(u2__abc_52138_new_n5777_), .Y(u2__abc_52138_new_n5778_));
OAI21X1 OAI21X1_43 ( .A(aNan), .B(_abc_65734_new_n956_), .C(_abc_65734_new_n957_), .Y(\o[154] ));
OAI21X1 OAI21X1_430 ( .A(u2__abc_52138_new_n5505_), .B(u2__abc_52138_new_n5510_), .C(u2__abc_52138_new_n5782_), .Y(u2__abc_52138_new_n5783_));
OAI21X1 OAI21X1_431 ( .A(u2__abc_52138_new_n5516_), .B(u2__abc_52138_new_n5521_), .C(u2__abc_52138_new_n5784_), .Y(u2__abc_52138_new_n5785_));
OAI21X1 OAI21X1_432 ( .A(u2__abc_52138_new_n5785_), .B(u2__abc_52138_new_n5512_), .C(u2__abc_52138_new_n5783_), .Y(u2__abc_52138_new_n5786_));
OAI21X1 OAI21X1_433 ( .A(u2_remHi_290_), .B(u2__abc_52138_new_n5787_), .C(u2__abc_52138_new_n5788_), .Y(u2__abc_52138_new_n5789_));
OAI21X1 OAI21X1_434 ( .A(u2__abc_52138_new_n5537_), .B(u2_o_291_), .C(u2__abc_52138_new_n5789_), .Y(u2__abc_52138_new_n5790_));
OAI21X1 OAI21X1_435 ( .A(u2__abc_52138_new_n5535_), .B(u2__abc_52138_new_n5790_), .C(u2__abc_52138_new_n5791_), .Y(u2__abc_52138_new_n5792_));
OAI21X1 OAI21X1_436 ( .A(u2_remHi_294_), .B(u2__abc_52138_new_n5455_), .C(u2__abc_52138_new_n5461_), .Y(u2__abc_52138_new_n5795_));
OAI21X1 OAI21X1_437 ( .A(u2__abc_52138_new_n5460_), .B(u2_o_295_), .C(u2__abc_52138_new_n5795_), .Y(u2__abc_52138_new_n5796_));
OAI21X1 OAI21X1_438 ( .A(u2__abc_52138_new_n5796_), .B(u2__abc_52138_new_n5476_), .C(u2__abc_52138_new_n5798_), .Y(u2__abc_52138_new_n5799_));
OAI21X1 OAI21X1_439 ( .A(u2_remHi_299_), .B(u2__abc_52138_new_n5496_), .C(u2__abc_52138_new_n5802_), .Y(u2__abc_52138_new_n5803_));
OAI21X1 OAI21X1_44 ( .A(aNan), .B(_abc_65734_new_n959_), .C(_abc_65734_new_n960_), .Y(\o[155] ));
OAI21X1 OAI21X1_440 ( .A(u2__abc_52138_new_n5806_), .B(u2__abc_52138_new_n5794_), .C(u2__abc_52138_new_n5454_), .Y(u2__abc_52138_new_n5807_));
OAI21X1 OAI21X1_441 ( .A(u2_remHi_310_), .B(u2__abc_52138_new_n5811_), .C(u2__abc_52138_new_n5812_), .Y(u2__abc_52138_new_n5813_));
OAI21X1 OAI21X1_442 ( .A(u2__abc_52138_new_n5374_), .B(u2__abc_52138_new_n5815_), .C(u2__abc_52138_new_n5810_), .Y(u2__abc_52138_new_n5816_));
OAI21X1 OAI21X1_443 ( .A(u2__abc_52138_new_n5399_), .B(u2_o_315_), .C(u2__abc_52138_new_n5821_), .Y(u2__abc_52138_new_n5822_));
OAI21X1 OAI21X1_444 ( .A(u2__abc_52138_new_n5428_), .B(u2__abc_52138_new_n5824_), .C(u2__abc_52138_new_n5826_), .Y(u2__abc_52138_new_n5827_));
OAI21X1 OAI21X1_445 ( .A(u2__abc_52138_new_n5440_), .B(u2__abc_52138_new_n5828_), .C(u2__abc_52138_new_n5829_), .Y(u2__abc_52138_new_n5830_));
OAI21X1 OAI21X1_446 ( .A(u2_remHi_318_), .B(u2__abc_52138_new_n5341_), .C(u2__abc_52138_new_n5347_), .Y(u2__abc_52138_new_n5836_));
OAI21X1 OAI21X1_447 ( .A(u2__abc_52138_new_n5346_), .B(u2_o_319_), .C(u2__abc_52138_new_n5836_), .Y(u2__abc_52138_new_n5837_));
OAI21X1 OAI21X1_448 ( .A(u2__abc_52138_new_n5837_), .B(u2__abc_52138_new_n5362_), .C(u2__abc_52138_new_n5839_), .Y(u2__abc_52138_new_n5840_));
OAI21X1 OAI21X1_449 ( .A(u2_remHi_322_), .B(u2__abc_52138_new_n5844_), .C(u2__abc_52138_new_n5336_), .Y(u2__abc_52138_new_n5845_));
OAI21X1 OAI21X1_45 ( .A(aNan), .B(_abc_65734_new_n962_), .C(_abc_65734_new_n963_), .Y(\o[156] ));
OAI21X1 OAI21X1_450 ( .A(u2_remHi_326_), .B(u2__abc_52138_new_n5274_), .C(u2__abc_52138_new_n5280_), .Y(u2__abc_52138_new_n5848_));
OAI21X1 OAI21X1_451 ( .A(u2__abc_52138_new_n5279_), .B(u2_o_327_), .C(u2__abc_52138_new_n5848_), .Y(u2__abc_52138_new_n5849_));
OAI21X1 OAI21X1_452 ( .A(u2__abc_52138_new_n5849_), .B(u2__abc_52138_new_n5295_), .C(u2__abc_52138_new_n5851_), .Y(u2__abc_52138_new_n5852_));
OAI21X1 OAI21X1_453 ( .A(u2__abc_52138_new_n5316_), .B(u2__abc_52138_new_n5855_), .C(u2__abc_52138_new_n5854_), .Y(u2__abc_52138_new_n5856_));
OAI21X1 OAI21X1_454 ( .A(u2_remHi_343_), .B(u2__abc_52138_new_n5202_), .C(u2__abc_52138_new_n5860_), .Y(u2__abc_52138_new_n5861_));
OAI21X1 OAI21X1_455 ( .A(u2__abc_52138_new_n5186_), .B(u2__abc_52138_new_n5189_), .C(u2__abc_52138_new_n5862_), .Y(u2__abc_52138_new_n5863_));
OAI21X1 OAI21X1_456 ( .A(u2__abc_52138_new_n5209_), .B(u2__abc_52138_new_n5211_), .C(u2__abc_52138_new_n5868_), .Y(u2__abc_52138_new_n5869_));
OAI21X1 OAI21X1_457 ( .A(u2__abc_52138_new_n5227_), .B(u2__abc_52138_new_n5864_), .C(u2__abc_52138_new_n5870_), .Y(u2__abc_52138_new_n5871_));
OAI21X1 OAI21X1_458 ( .A(u2__abc_52138_new_n5875_), .B(u2__abc_52138_new_n5246_), .C(u2__abc_52138_new_n5245_), .Y(u2__abc_52138_new_n5876_));
OAI21X1 OAI21X1_459 ( .A(u2__abc_52138_new_n5252_), .B(u2__abc_52138_new_n5255_), .C(u2__abc_52138_new_n5878_), .Y(u2__abc_52138_new_n5879_));
OAI21X1 OAI21X1_46 ( .A(aNan), .B(_abc_65734_new_n965_), .C(_abc_65734_new_n966_), .Y(\o[157] ));
OAI21X1 OAI21X1_460 ( .A(u2__abc_52138_new_n5264_), .B(u2__abc_52138_new_n5267_), .C(u2__abc_52138_new_n5880_), .Y(u2__abc_52138_new_n5881_));
OAI21X1 OAI21X1_461 ( .A(u2__abc_52138_new_n5271_), .B(u2__abc_52138_new_n5877_), .C(u2__abc_52138_new_n5882_), .Y(u2__abc_52138_new_n5883_));
OAI21X1 OAI21X1_462 ( .A(u2__abc_52138_new_n5273_), .B(u2__abc_52138_new_n5859_), .C(u2__abc_52138_new_n5884_), .Y(u2__abc_52138_new_n5885_));
OAI21X1 OAI21X1_463 ( .A(u2_remHi_368_), .B(u2__abc_52138_new_n5047_), .C(u2__abc_52138_new_n5887_), .Y(u2__abc_52138_new_n5888_));
OAI21X1 OAI21X1_464 ( .A(u2__abc_52138_new_n5886_), .B(u2_o_369_), .C(u2__abc_52138_new_n5888_), .Y(u2__abc_52138_new_n5889_));
OAI21X1 OAI21X1_465 ( .A(u2_remHi_366_), .B(u2__abc_52138_new_n5890_), .C(u2__abc_52138_new_n5060_), .Y(u2__abc_52138_new_n5891_));
OAI21X1 OAI21X1_466 ( .A(u2__abc_52138_new_n5059_), .B(u2_o_367_), .C(u2__abc_52138_new_n5891_), .Y(u2__abc_52138_new_n5892_));
OAI21X1 OAI21X1_467 ( .A(u2__abc_52138_new_n5892_), .B(u2__abc_52138_new_n5051_), .C(u2__abc_52138_new_n5889_), .Y(u2__abc_52138_new_n5893_));
OAI21X1 OAI21X1_468 ( .A(u2__abc_52138_new_n5085_), .B(u2__abc_52138_new_n5080_), .C(u2__abc_52138_new_n5079_), .Y(u2__abc_52138_new_n5896_));
OAI21X1 OAI21X1_469 ( .A(u2__abc_52138_new_n5070_), .B(u2_o_373_), .C(u2__abc_52138_new_n5068_), .Y(u2__abc_52138_new_n5898_));
OAI21X1 OAI21X1_47 ( .A(aNan), .B(_abc_65734_new_n968_), .C(_abc_65734_new_n969_), .Y(\o[158] ));
OAI21X1 OAI21X1_470 ( .A(u2__abc_52138_new_n5105_), .B(u2__abc_52138_new_n5903_), .C(u2__abc_52138_new_n5108_), .Y(u2__abc_52138_new_n5904_));
OAI21X1 OAI21X1_471 ( .A(u2_remHi_358_), .B(u2__abc_52138_new_n5091_), .C(u2__abc_52138_new_n5097_), .Y(u2__abc_52138_new_n5905_));
OAI21X1 OAI21X1_472 ( .A(u2__abc_52138_new_n5096_), .B(u2_o_359_), .C(u2__abc_52138_new_n5905_), .Y(u2__abc_52138_new_n5906_));
OAI21X1 OAI21X1_473 ( .A(u2__abc_52138_new_n5906_), .B(u2__abc_52138_new_n5112_), .C(u2__abc_52138_new_n5904_), .Y(u2__abc_52138_new_n5907_));
OAI21X1 OAI21X1_474 ( .A(u2_remHi_362_), .B(u2__abc_52138_new_n5911_), .C(u2__abc_52138_new_n5912_), .Y(u2__abc_52138_new_n5913_));
OAI21X1 OAI21X1_475 ( .A(u2__abc_52138_new_n5137_), .B(u2__abc_52138_new_n5142_), .C(u2__abc_52138_new_n5918_), .Y(u2__abc_52138_new_n5919_));
OAI21X1 OAI21X1_476 ( .A(u2__abc_52138_new_n5148_), .B(u2__abc_52138_new_n5153_), .C(u2__abc_52138_new_n5920_), .Y(u2__abc_52138_new_n5921_));
OAI21X1 OAI21X1_477 ( .A(u2__abc_52138_new_n5921_), .B(u2__abc_52138_new_n5144_), .C(u2__abc_52138_new_n5919_), .Y(u2__abc_52138_new_n5922_));
OAI21X1 OAI21X1_478 ( .A(u2__abc_52138_new_n5167_), .B(u2__abc_52138_new_n5924_), .C(u2__abc_52138_new_n5923_), .Y(u2__abc_52138_new_n5925_));
OAI21X1 OAI21X1_479 ( .A(u2__abc_52138_new_n5927_), .B(u2__abc_52138_new_n5917_), .C(u2__abc_52138_new_n5090_), .Y(u2__abc_52138_new_n5928_));
OAI21X1 OAI21X1_48 ( .A(aNan), .B(_abc_65734_new_n971_), .C(_abc_65734_new_n972_), .Y(\o[159] ));
OAI21X1 OAI21X1_480 ( .A(u2__abc_52138_new_n5033_), .B(u2__abc_52138_new_n5039_), .C(u2__abc_52138_new_n5037_), .Y(u2__abc_52138_new_n5929_));
OAI21X1 OAI21X1_481 ( .A(u2_remHi_374_), .B(u2__abc_52138_new_n5018_), .C(u2__abc_52138_new_n5024_), .Y(u2__abc_52138_new_n5930_));
OAI21X1 OAI21X1_482 ( .A(u2__abc_52138_new_n5023_), .B(u2_o_375_), .C(u2__abc_52138_new_n5930_), .Y(u2__abc_52138_new_n5931_));
OAI21X1 OAI21X1_483 ( .A(u2__abc_52138_new_n5931_), .B(u2__abc_52138_new_n5042_), .C(u2__abc_52138_new_n5929_), .Y(u2__abc_52138_new_n5932_));
OAI21X1 OAI21X1_484 ( .A(u2_remHi_378_), .B(u2__abc_52138_new_n5933_), .C(u2__abc_52138_new_n5934_), .Y(u2__abc_52138_new_n5935_));
OAI21X1 OAI21X1_485 ( .A(u2__abc_52138_new_n5011_), .B(u2_o_379_), .C(u2__abc_52138_new_n5935_), .Y(u2__abc_52138_new_n5936_));
OAI21X1 OAI21X1_486 ( .A(u2__abc_52138_new_n5009_), .B(u2__abc_52138_new_n5936_), .C(u2__abc_52138_new_n5937_), .Y(u2__abc_52138_new_n5938_));
OAI21X1 OAI21X1_487 ( .A(u2__abc_52138_new_n5367_), .B(u2__abc_52138_new_n5835_), .C(u2__abc_52138_new_n5941_), .Y(u2__abc_52138_new_n5942_));
OAI21X1 OAI21X1_488 ( .A(u2__abc_52138_new_n6335_), .B(u2__abc_52138_new_n6170_), .C(u2__abc_52138_new_n6337_), .Y(u2__abc_52138_new_n6338_));
OAI21X1 OAI21X1_489 ( .A(u2__abc_52138_new_n6340_), .B(u2__abc_52138_new_n6146_), .C(u2__abc_52138_new_n6341_), .Y(u2__abc_52138_new_n6342_));
OAI21X1 OAI21X1_49 ( .A(aNan), .B(_abc_65734_new_n974_), .C(_abc_65734_new_n975_), .Y(\o[160] ));
OAI21X1 OAI21X1_490 ( .A(u2__abc_52138_new_n6323_), .B(u2__abc_52138_new_n6318_), .C(u2__abc_52138_new_n6346_), .Y(u2__abc_52138_new_n6347_));
OAI21X1 OAI21X1_491 ( .A(u2__abc_52138_new_n6352_), .B(u2_o_393_), .C(u2__abc_52138_new_n6283_), .Y(u2__abc_52138_new_n6353_));
OAI21X1 OAI21X1_492 ( .A(u2__abc_52138_new_n6351_), .B(u2__abc_52138_new_n6291_), .C(u2__abc_52138_new_n6353_), .Y(u2__abc_52138_new_n6354_));
OAI21X1 OAI21X1_493 ( .A(u2__abc_52138_new_n6286_), .B(u2__abc_52138_new_n6354_), .C(u2__abc_52138_new_n6326_), .Y(u2__abc_52138_new_n6355_));
OAI21X1 OAI21X1_494 ( .A(u2__abc_52138_new_n6344_), .B(u2__abc_52138_new_n6356_), .C(u2__abc_52138_new_n6279_), .Y(u2__abc_52138_new_n6357_));
OAI21X1 OAI21X1_495 ( .A(u2__abc_52138_new_n6359_), .B(u2__abc_52138_new_n6195_), .C(u2__abc_52138_new_n6361_), .Y(u2__abc_52138_new_n6362_));
OAI21X1 OAI21X1_496 ( .A(u2__abc_52138_new_n6222_), .B(u2__abc_52138_new_n6366_), .C(u2__abc_52138_new_n6365_), .Y(u2__abc_52138_new_n6367_));
OAI21X1 OAI21X1_497 ( .A(u2__abc_52138_new_n6374_), .B(u2__abc_52138_new_n6253_), .C(u2__abc_52138_new_n6376_), .Y(u2__abc_52138_new_n6377_));
OAI21X1 OAI21X1_498 ( .A(u2__abc_52138_new_n6379_), .B(u2__abc_52138_new_n6265_), .C(u2__abc_52138_new_n6381_), .Y(u2__abc_52138_new_n6382_));
OAI21X1 OAI21X1_499 ( .A(u2__abc_52138_new_n6123_), .B(u2__abc_52138_new_n6389_), .C(u2__abc_52138_new_n6388_), .Y(u2__abc_52138_new_n6390_));
OAI21X1 OAI21X1_5 ( .A(aNan), .B(_abc_65734_new_n842_), .C(_abc_65734_new_n843_), .Y(\o[116] ));
OAI21X1 OAI21X1_50 ( .A(aNan), .B(_abc_65734_new_n977_), .C(_abc_65734_new_n978_), .Y(\o[161] ));
OAI21X1 OAI21X1_500 ( .A(u2__abc_52138_new_n6111_), .B(u2__abc_52138_new_n6117_), .C(u2__abc_52138_new_n6114_), .Y(u2__abc_52138_new_n6391_));
OAI21X1 OAI21X1_501 ( .A(u2__abc_52138_new_n6099_), .B(u2__abc_52138_new_n6394_), .C(u2__abc_52138_new_n6393_), .Y(u2__abc_52138_new_n6395_));
OAI21X1 OAI21X1_502 ( .A(u2__abc_52138_new_n6087_), .B(u2__abc_52138_new_n6093_), .C(u2__abc_52138_new_n6092_), .Y(u2__abc_52138_new_n6396_));
OAI21X1 OAI21X1_503 ( .A(u2__abc_52138_new_n6392_), .B(u2__abc_52138_new_n6387_), .C(u2__abc_52138_new_n6397_), .Y(u2__abc_52138_new_n6398_));
OAI21X1 OAI21X1_504 ( .A(u2__abc_52138_new_n6039_), .B(u2__abc_52138_new_n6045_), .C(u2__abc_52138_new_n6042_), .Y(u2__abc_52138_new_n6404_));
OAI21X1 OAI21X1_505 ( .A(u2__abc_52138_new_n6404_), .B(u2__abc_52138_new_n6403_), .C(u2__abc_52138_new_n6081_), .Y(u2__abc_52138_new_n6405_));
OAI21X1 OAI21X1_506 ( .A(u2__abc_52138_new_n6073_), .B(u2__abc_52138_new_n6407_), .C(u2__abc_52138_new_n6406_), .Y(u2__abc_52138_new_n6408_));
OAI21X1 OAI21X1_507 ( .A(u2__abc_52138_new_n6061_), .B(u2__abc_52138_new_n6067_), .C(u2__abc_52138_new_n6066_), .Y(u2__abc_52138_new_n6409_));
OAI21X1 OAI21X1_508 ( .A(u2__abc_52138_new_n6411_), .B(u2__abc_52138_new_n6399_), .C(u2__abc_52138_new_n6034_), .Y(u2__abc_52138_new_n6412_));
OAI21X1 OAI21X1_509 ( .A(u2_o_439_), .B(u2__abc_52138_new_n6415_), .C(u2__abc_52138_new_n5970_), .Y(u2__abc_52138_new_n6416_));
OAI21X1 OAI21X1_51 ( .A(aNan), .B(_abc_65734_new_n980_), .C(_abc_65734_new_n981_), .Y(\o[162] ));
OAI21X1 OAI21X1_510 ( .A(u2__abc_52138_new_n6414_), .B(u2_remHi_439_), .C(u2__abc_52138_new_n6416_), .Y(u2__abc_52138_new_n6417_));
OAI21X1 OAI21X1_511 ( .A(u2__abc_52138_new_n5981_), .B(u2_o_441_), .C(u2__abc_52138_new_n5977_), .Y(u2__abc_52138_new_n6419_));
OAI21X1 OAI21X1_512 ( .A(u2_remHi_441_), .B(u2__abc_52138_new_n5979_), .C(u2__abc_52138_new_n6419_), .Y(u2__abc_52138_new_n6420_));
OAI21X1 OAI21X1_513 ( .A(u2__abc_52138_new_n6420_), .B(u2__abc_52138_new_n6418_), .C(u2__abc_52138_new_n5966_), .Y(u2__abc_52138_new_n6421_));
OAI21X1 OAI21X1_514 ( .A(u2__abc_52138_new_n6428_), .B(u2__abc_52138_new_n6031_), .C(u2__abc_52138_new_n6429_), .Y(u2__abc_52138_new_n6430_));
OAI21X1 OAI21X1_515 ( .A(u2__abc_52138_new_n6432_), .B(u2__abc_52138_new_n5997_), .C(u2__abc_52138_new_n6434_), .Y(u2__abc_52138_new_n6435_));
OAI21X1 OAI21X1_516 ( .A(u2__abc_52138_new_n6332_), .B(u2__abc_52138_new_n5943_), .C(u2__abc_52138_new_n6440_), .Y(u2__abc_52138_new_n6441_));
OAI21X1 OAI21X1_517 ( .A(u2__abc_52138_new_n3003_), .B(u2_o_447_), .C(u2__abc_52138_new_n3002_), .Y(u2__abc_52138_new_n6444_));
OAI21X1 OAI21X1_518 ( .A(u2_o_449_), .B(u2__abc_52138_new_n6447_), .C(u2__abc_52138_new_n2998_), .Y(u2__abc_52138_new_n6448_));
OAI21X1 OAI21X1_519 ( .A(u2__abc_52138_new_n6446_), .B(u2_remHi_449_), .C(u2__abc_52138_new_n6448_), .Y(u2__abc_52138_new_n6449_));
OAI21X1 OAI21X1_52 ( .A(aNan), .B(_abc_65734_new_n983_), .C(_abc_65734_new_n984_), .Y(\o[163] ));
OAI21X1 OAI21X1_520 ( .A(u2_remHiShift_0_), .B(u2__abc_52138_new_n6498_), .C(u2__abc_52138_new_n2990_), .Y(u2__abc_52138_new_n6501_));
OAI21X1 OAI21X1_521 ( .A(u2__abc_52138_new_n6501_), .B(u2__abc_52138_new_n6500_), .C(u2__abc_52138_new_n6506_), .Y(u2__abc_52138_new_n6507_));
OAI21X1 OAI21X1_522 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_1_), .Y(u2__abc_52138_new_n6509_));
OAI21X1 OAI21X1_523 ( .A(u2__abc_52138_new_n6454_), .B(u2__abc_52138_new_n3071_), .C(u2__abc_52138_new_n2996_), .Y(u2__abc_52138_new_n6511_));
OAI21X1 OAI21X1_524 ( .A(u2__abc_52138_new_n6498_), .B(u2__abc_52138_new_n6512_), .C(u2__abc_52138_new_n6513_), .Y(u2__abc_52138_new_n6514_));
OAI21X1 OAI21X1_525 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6514_), .C(u2__abc_52138_new_n6516_), .Y(u2__abc_52138_new_n6517_));
OAI21X1 OAI21X1_526 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_2_), .Y(u2__abc_52138_new_n6519_));
OAI21X1 OAI21X1_527 ( .A(u2__abc_52138_new_n2996_), .B(u2__abc_52138_new_n6454_), .C(u2__abc_52138_new_n3070_), .Y(u2__abc_52138_new_n6520_));
OAI21X1 OAI21X1_528 ( .A(u2__abc_52138_new_n6502_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6523_), .Y(u2__abc_52138_new_n6524_));
OAI21X1 OAI21X1_529 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6524_), .C(u2__abc_52138_new_n6525_), .Y(u2__abc_52138_new_n6526_));
OAI21X1 OAI21X1_53 ( .A(aNan), .B(_abc_65734_new_n986_), .C(_abc_65734_new_n987_), .Y(\o[164] ));
OAI21X1 OAI21X1_530 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_3_), .Y(u2__abc_52138_new_n6528_));
OAI21X1 OAI21X1_531 ( .A(u2__abc_52138_new_n6502_), .B(sqrto_0_), .C(u2__abc_52138_new_n6521_), .Y(u2__abc_52138_new_n6529_));
OAI21X1 OAI21X1_532 ( .A(u2__abc_52138_new_n6515_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6532_), .Y(u2__abc_52138_new_n6533_));
OAI21X1 OAI21X1_533 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6533_), .C(u2__abc_52138_new_n6534_), .Y(u2__abc_52138_new_n6535_));
OAI21X1 OAI21X1_534 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_4_), .Y(u2__abc_52138_new_n6537_));
OAI21X1 OAI21X1_535 ( .A(sqrto_1_), .B(u2__abc_52138_new_n6515_), .C(u2__abc_52138_new_n6531_), .Y(u2__abc_52138_new_n6542_));
OAI21X1 OAI21X1_536 ( .A(u2__abc_52138_new_n6541_), .B(u2__abc_52138_new_n6539_), .C(u2__abc_52138_new_n6543_), .Y(u2__abc_52138_new_n6544_));
OAI21X1 OAI21X1_537 ( .A(u2__abc_52138_new_n3062_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6544_), .Y(u2__abc_52138_new_n6545_));
OAI21X1 OAI21X1_538 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6545_), .C(u2__abc_52138_new_n6546_), .Y(u2__abc_52138_new_n6547_));
OAI21X1 OAI21X1_539 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_5_), .Y(u2__abc_52138_new_n6549_));
OAI21X1 OAI21X1_54 ( .A(aNan), .B(_abc_65734_new_n989_), .C(_abc_65734_new_n990_), .Y(\o[165] ));
OAI21X1 OAI21X1_540 ( .A(u2__abc_52138_new_n3084_), .B(u2__abc_52138_new_n6550_), .C(u2__abc_52138_new_n3061_), .Y(u2__abc_52138_new_n6551_));
OAI21X1 OAI21X1_541 ( .A(u2__abc_52138_new_n6541_), .B(u2__abc_52138_new_n6539_), .C(u2__abc_52138_new_n6552_), .Y(u2__abc_52138_new_n6553_));
OAI21X1 OAI21X1_542 ( .A(u2__abc_52138_new_n3081_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6553_), .Y(u2__abc_52138_new_n6554_));
OAI21X1 OAI21X1_543 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6554_), .C(u2__abc_52138_new_n6555_), .Y(u2__abc_52138_new_n6556_));
OAI21X1 OAI21X1_544 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_6_), .Y(u2__abc_52138_new_n6558_));
OAI21X1 OAI21X1_545 ( .A(sqrto_2_), .B(u2__abc_52138_new_n3062_), .C(u2__abc_52138_new_n3080_), .Y(u2__abc_52138_new_n6559_));
OAI21X1 OAI21X1_546 ( .A(u2__abc_52138_new_n6541_), .B(u2__abc_52138_new_n6539_), .C(u2__abc_52138_new_n6561_), .Y(u2__abc_52138_new_n6562_));
OAI21X1 OAI21X1_547 ( .A(u2__abc_52138_new_n3086_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6562_), .Y(u2__abc_52138_new_n6563_));
OAI21X1 OAI21X1_548 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6563_), .C(u2__abc_52138_new_n6564_), .Y(u2__abc_52138_new_n6565_));
OAI21X1 OAI21X1_549 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_7_), .Y(u2__abc_52138_new_n6567_));
OAI21X1 OAI21X1_55 ( .A(aNan), .B(_abc_65734_new_n992_), .C(_abc_65734_new_n993_), .Y(\o[166] ));
OAI21X1 OAI21X1_550 ( .A(u2__abc_52138_new_n3088_), .B(u2__abc_52138_new_n6560_), .C(u2__abc_52138_new_n6459_), .Y(u2__abc_52138_new_n6568_));
OAI21X1 OAI21X1_551 ( .A(u2__abc_52138_new_n6541_), .B(u2__abc_52138_new_n6539_), .C(u2__abc_52138_new_n6569_), .Y(u2__abc_52138_new_n6570_));
OAI21X1 OAI21X1_552 ( .A(u2__abc_52138_new_n3054_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6570_), .Y(u2__abc_52138_new_n6571_));
OAI21X1 OAI21X1_553 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6571_), .C(u2__abc_52138_new_n6572_), .Y(u2__abc_52138_new_n6573_));
OAI21X1 OAI21X1_554 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_8_), .Y(u2__abc_52138_new_n6575_));
OAI21X1 OAI21X1_555 ( .A(u2__abc_52138_new_n3079_), .B(u2_remHi_3_), .C(u2__abc_52138_new_n6559_), .Y(u2__abc_52138_new_n6577_));
OAI21X1 OAI21X1_556 ( .A(u2__abc_52138_new_n3058_), .B(u2__abc_52138_new_n6577_), .C(u2__abc_52138_new_n6580_), .Y(u2__abc_52138_new_n6581_));
OAI21X1 OAI21X1_557 ( .A(u2__abc_52138_new_n6541_), .B(u2__abc_52138_new_n6539_), .C(u2__abc_52138_new_n6583_), .Y(u2__abc_52138_new_n6584_));
OAI21X1 OAI21X1_558 ( .A(u2__abc_52138_new_n3047_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6584_), .Y(u2__abc_52138_new_n6585_));
OAI21X1 OAI21X1_559 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6585_), .C(u2__abc_52138_new_n6587_), .Y(u2__abc_52138_new_n6588_));
OAI21X1 OAI21X1_56 ( .A(aNan), .B(_abc_65734_new_n995_), .C(_abc_65734_new_n996_), .Y(\o[167] ));
OAI21X1 OAI21X1_560 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_9_), .Y(u2__abc_52138_new_n6590_));
OAI21X1 OAI21X1_561 ( .A(u2__abc_52138_new_n3094_), .B(u2__abc_52138_new_n6582_), .C(u2__abc_52138_new_n3046_), .Y(u2__abc_52138_new_n6591_));
OAI21X1 OAI21X1_562 ( .A(u2__abc_52138_new_n3042_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6594_));
OAI21X1 OAI21X1_563 ( .A(u2__abc_52138_new_n6593_), .B(u2__abc_52138_new_n6594_), .C(u2__abc_52138_new_n6595_), .Y(u2__abc_52138_new_n6596_));
OAI21X1 OAI21X1_564 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_10_), .Y(u2__abc_52138_new_n6598_));
OAI21X1 OAI21X1_565 ( .A(u2__abc_52138_new_n6600_), .B(u2__abc_52138_new_n6601_), .C(u2__abc_52138_new_n3043_), .Y(u2__abc_52138_new_n6602_));
OAI21X1 OAI21X1_566 ( .A(u2__abc_52138_new_n3050_), .B(u2__abc_52138_new_n6582_), .C(u2__abc_52138_new_n6602_), .Y(u2__abc_52138_new_n6603_));
OAI21X1 OAI21X1_567 ( .A(u2__abc_52138_new_n6586_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6608_), .Y(u2__abc_52138_new_n6609_));
OAI21X1 OAI21X1_568 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6609_), .C(u2__abc_52138_new_n6610_), .Y(u2__abc_52138_new_n6611_));
OAI21X1 OAI21X1_569 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_11_), .Y(u2__abc_52138_new_n6613_));
OAI21X1 OAI21X1_57 ( .A(aNan), .B(_abc_65734_new_n998_), .C(_abc_65734_new_n999_), .Y(\o[168] ));
OAI21X1 OAI21X1_570 ( .A(u2__abc_52138_new_n3097_), .B(u2__abc_52138_new_n6604_), .C(u2__abc_52138_new_n6615_), .Y(u2__abc_52138_new_n6616_));
OAI21X1 OAI21X1_571 ( .A(u2__abc_52138_new_n6541_), .B(u2__abc_52138_new_n6539_), .C(u2__abc_52138_new_n6617_), .Y(u2__abc_52138_new_n6618_));
OAI21X1 OAI21X1_572 ( .A(u2__abc_52138_new_n3037_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6618_), .Y(u2__abc_52138_new_n6619_));
OAI21X1 OAI21X1_573 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6619_), .C(u2__abc_52138_new_n6620_), .Y(u2__abc_52138_new_n6621_));
OAI21X1 OAI21X1_574 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_12_), .Y(u2__abc_52138_new_n6623_));
OAI21X1 OAI21X1_575 ( .A(sqrto_9_), .B(u2__abc_52138_new_n3037_), .C(u2__abc_52138_new_n6615_), .Y(u2__abc_52138_new_n6624_));
OAI21X1 OAI21X1_576 ( .A(u2__abc_52138_new_n3035_), .B(u2_remHi_9_), .C(u2__abc_52138_new_n6624_), .Y(u2__abc_52138_new_n6625_));
OAI21X1 OAI21X1_577 ( .A(u2__abc_52138_new_n3039_), .B(u2__abc_52138_new_n6604_), .C(u2__abc_52138_new_n6625_), .Y(u2__abc_52138_new_n6626_));
OAI21X1 OAI21X1_578 ( .A(u2__abc_52138_new_n3029_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6629_), .Y(u2__abc_52138_new_n6630_));
OAI21X1 OAI21X1_579 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6630_), .C(u2__abc_52138_new_n6631_), .Y(u2__abc_52138_new_n6632_));
OAI21X1 OAI21X1_58 ( .A(aNan), .B(_abc_65734_new_n1001_), .C(_abc_65734_new_n1002_), .Y(\o[169] ));
OAI21X1 OAI21X1_580 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_13_), .Y(u2__abc_52138_new_n6634_));
OAI21X1 OAI21X1_581 ( .A(sqrto_10_), .B(u2__abc_52138_new_n3029_), .C(u2__abc_52138_new_n6628_), .Y(u2__abc_52138_new_n6635_));
OAI21X1 OAI21X1_582 ( .A(u2__abc_52138_new_n3024_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6638_));
OAI21X1 OAI21X1_583 ( .A(u2__abc_52138_new_n6637_), .B(u2__abc_52138_new_n6638_), .C(u2__abc_52138_new_n6639_), .Y(u2__abc_52138_new_n6640_));
OAI21X1 OAI21X1_584 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_14_), .Y(u2__abc_52138_new_n6642_));
OAI21X1 OAI21X1_585 ( .A(sqrto_10_), .B(u2__abc_52138_new_n3029_), .C(u2__abc_52138_new_n3023_), .Y(u2__abc_52138_new_n6644_));
OAI21X1 OAI21X1_586 ( .A(u2__abc_52138_new_n6644_), .B(u2__abc_52138_new_n6643_), .C(u2__abc_52138_new_n3025_), .Y(u2__abc_52138_new_n6645_));
OAI21X1 OAI21X1_587 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6646_), .Y(u2__abc_52138_new_n6647_));
OAI21X1 OAI21X1_588 ( .A(u2__abc_52138_new_n3101_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6647_), .Y(u2__abc_52138_new_n6648_));
OAI21X1 OAI21X1_589 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6648_), .C(u2__abc_52138_new_n6649_), .Y(u2__abc_52138_new_n6650_));
OAI21X1 OAI21X1_59 ( .A(aNan), .B(_abc_65734_new_n1004_), .C(_abc_65734_new_n1005_), .Y(\o[170] ));
OAI21X1 OAI21X1_590 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_15_), .Y(u2__abc_52138_new_n6652_));
OAI21X1 OAI21X1_591 ( .A(u2__abc_52138_new_n3103_), .B(u2__abc_52138_new_n6645_), .C(u2__abc_52138_new_n6655_), .Y(u2__abc_52138_new_n6656_));
OAI21X1 OAI21X1_592 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6657_), .Y(u2__abc_52138_new_n6658_));
OAI21X1 OAI21X1_593 ( .A(u2__abc_52138_new_n3017_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6658_), .Y(u2__abc_52138_new_n6659_));
OAI21X1 OAI21X1_594 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6659_), .C(u2__abc_52138_new_n6660_), .Y(u2__abc_52138_new_n6661_));
OAI21X1 OAI21X1_595 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_16_), .Y(u2__abc_52138_new_n6663_));
OAI21X1 OAI21X1_596 ( .A(u2__abc_52138_new_n3039_), .B(u2__abc_52138_new_n6602_), .C(u2__abc_52138_new_n6625_), .Y(u2__abc_52138_new_n6665_));
OAI21X1 OAI21X1_597 ( .A(u2__abc_52138_new_n3028_), .B(u2__abc_52138_new_n3106_), .C(u2__abc_52138_new_n3023_), .Y(u2__abc_52138_new_n6669_));
OAI21X1 OAI21X1_598 ( .A(u2__abc_52138_new_n6655_), .B(u2__abc_52138_new_n3104_), .C(u2__abc_52138_new_n3020_), .Y(u2__abc_52138_new_n6670_));
OAI21X1 OAI21X1_599 ( .A(u2__abc_52138_new_n3052_), .B(u2__abc_52138_new_n6582_), .C(u2__abc_52138_new_n6672_), .Y(u2__abc_52138_new_n6673_));
OAI21X1 OAI21X1_6 ( .A(aNan), .B(_abc_65734_new_n845_), .C(_abc_65734_new_n846_), .Y(\o[117] ));
OAI21X1 OAI21X1_60 ( .A(aNan), .B(_abc_65734_new_n1007_), .C(_abc_65734_new_n1008_), .Y(\o[171] ));
OAI21X1 OAI21X1_600 ( .A(u2__abc_52138_new_n6664_), .B(u2__abc_52138_new_n3199_), .C(u2__abc_52138_new_n6674_), .Y(u2__abc_52138_new_n6675_));
OAI21X1 OAI21X1_601 ( .A(u2__abc_52138_new_n3172_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6677_), .Y(u2__abc_52138_new_n6678_));
OAI21X1 OAI21X1_602 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6678_), .C(u2__abc_52138_new_n6679_), .Y(u2__abc_52138_new_n6680_));
OAI21X1 OAI21X1_603 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_17_), .Y(u2__abc_52138_new_n6682_));
OAI21X1 OAI21X1_604 ( .A(u2__abc_52138_new_n3199_), .B(u2__abc_52138_new_n6674_), .C(u2__abc_52138_new_n3171_), .Y(u2__abc_52138_new_n6683_));
OAI21X1 OAI21X1_605 ( .A(u2__abc_52138_new_n3177_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6686_));
OAI21X1 OAI21X1_606 ( .A(u2__abc_52138_new_n6685_), .B(u2__abc_52138_new_n6686_), .C(u2__abc_52138_new_n6687_), .Y(u2__abc_52138_new_n6688_));
OAI21X1 OAI21X1_607 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_18_), .Y(u2__abc_52138_new_n6690_));
OAI21X1 OAI21X1_608 ( .A(u2__abc_52138_new_n6691_), .B(u2__abc_52138_new_n3202_), .C(u2__abc_52138_new_n6693_), .Y(u2__abc_52138_new_n6694_));
OAI21X1 OAI21X1_609 ( .A(u2__abc_52138_new_n3161_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6696_), .Y(u2__abc_52138_new_n6697_));
OAI21X1 OAI21X1_61 ( .A(aNan), .B(_abc_65734_new_n1010_), .C(_abc_65734_new_n1011_), .Y(\o[172] ));
OAI21X1 OAI21X1_610 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6697_), .C(u2__abc_52138_new_n6698_), .Y(u2__abc_52138_new_n6699_));
OAI21X1 OAI21X1_611 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_19_), .Y(u2__abc_52138_new_n6701_));
OAI21X1 OAI21X1_612 ( .A(u2__abc_52138_new_n3202_), .B(u2__abc_52138_new_n6693_), .C(u2__abc_52138_new_n3160_), .Y(u2__abc_52138_new_n6702_));
OAI21X1 OAI21X1_613 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6703_), .Y(u2__abc_52138_new_n6704_));
OAI21X1 OAI21X1_614 ( .A(u2__abc_52138_new_n3166_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6704_), .Y(u2__abc_52138_new_n6705_));
OAI21X1 OAI21X1_615 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6705_), .C(u2__abc_52138_new_n6707_), .Y(u2__abc_52138_new_n6708_));
OAI21X1 OAI21X1_616 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_20_), .Y(u2__abc_52138_new_n6710_));
OAI21X1 OAI21X1_617 ( .A(u2__abc_52138_new_n6664_), .B(u2__abc_52138_new_n6692_), .C(u2__abc_52138_new_n3178_), .Y(u2__abc_52138_new_n6712_));
OAI21X1 OAI21X1_618 ( .A(u2__abc_52138_new_n3198_), .B(u2__abc_52138_new_n6712_), .C(u2__abc_52138_new_n6714_), .Y(u2__abc_52138_new_n6715_));
OAI21X1 OAI21X1_619 ( .A(u2__abc_52138_new_n3191_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6719_), .Y(u2__abc_52138_new_n6720_));
OAI21X1 OAI21X1_62 ( .A(aNan), .B(_abc_65734_new_n1013_), .C(_abc_65734_new_n1014_), .Y(\o[173] ));
OAI21X1 OAI21X1_620 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6720_), .C(u2__abc_52138_new_n6721_), .Y(u2__abc_52138_new_n6722_));
OAI21X1 OAI21X1_621 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_21_), .Y(u2__abc_52138_new_n6724_));
OAI21X1 OAI21X1_622 ( .A(u2__abc_52138_new_n3209_), .B(u2__abc_52138_new_n6716_), .C(u2__abc_52138_new_n3190_), .Y(u2__abc_52138_new_n6725_));
OAI21X1 OAI21X1_623 ( .A(u2__abc_52138_new_n6541_), .B(u2__abc_52138_new_n6539_), .C(u2__abc_52138_new_n6726_), .Y(u2__abc_52138_new_n6727_));
OAI21X1 OAI21X1_624 ( .A(u2__abc_52138_new_n6706_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6727_), .Y(u2__abc_52138_new_n6728_));
OAI21X1 OAI21X1_625 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6728_), .C(u2__abc_52138_new_n6729_), .Y(u2__abc_52138_new_n6730_));
OAI21X1 OAI21X1_626 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_22_), .Y(u2__abc_52138_new_n6732_));
OAI21X1 OAI21X1_627 ( .A(u2__abc_52138_new_n3190_), .B(u2__abc_52138_new_n3208_), .C(u2__abc_52138_new_n3207_), .Y(u2__abc_52138_new_n6737_));
OAI21X1 OAI21X1_628 ( .A(u2__abc_52138_new_n6737_), .B(u2__abc_52138_new_n6736_), .C(u2__abc_52138_new_n3182_), .Y(u2__abc_52138_new_n6740_));
OAI21X1 OAI21X1_629 ( .A(u2__abc_52138_new_n3211_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6741_), .Y(u2__abc_52138_new_n6742_));
OAI21X1 OAI21X1_63 ( .A(aNan), .B(_abc_65734_new_n1016_), .C(_abc_65734_new_n1017_), .Y(\o[174] ));
OAI21X1 OAI21X1_630 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6742_), .C(u2__abc_52138_new_n6743_), .Y(u2__abc_52138_new_n6744_));
OAI21X1 OAI21X1_631 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_23_), .Y(u2__abc_52138_new_n6746_));
OAI21X1 OAI21X1_632 ( .A(sqrto_20_), .B(u2__abc_52138_new_n3211_), .C(u2__abc_52138_new_n6740_), .Y(u2__abc_52138_new_n6748_));
OAI21X1 OAI21X1_633 ( .A(u2__abc_52138_new_n3185_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6751_));
OAI21X1 OAI21X1_634 ( .A(u2__abc_52138_new_n6750_), .B(u2__abc_52138_new_n6751_), .C(u2__abc_52138_new_n6752_), .Y(u2__abc_52138_new_n6753_));
OAI21X1 OAI21X1_635 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_24_), .Y(u2__abc_52138_new_n6755_));
OAI21X1 OAI21X1_636 ( .A(u2__abc_52138_new_n6762_), .B(u2__abc_52138_new_n6756_), .C(u2__abc_52138_new_n6765_), .Y(u2__abc_52138_new_n6766_));
OAI21X1 OAI21X1_637 ( .A(u2__abc_52138_new_n3130_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6767_), .Y(u2__abc_52138_new_n6768_));
OAI21X1 OAI21X1_638 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6768_), .C(u2__abc_52138_new_n6769_), .Y(u2__abc_52138_new_n6770_));
OAI21X1 OAI21X1_639 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_25_), .Y(u2__abc_52138_new_n6772_));
OAI21X1 OAI21X1_64 ( .A(aNan), .B(_abc_65734_new_n1019_), .C(_abc_65734_new_n1020_), .Y(\o[175] ));
OAI21X1 OAI21X1_640 ( .A(sqrto_22_), .B(u2__abc_52138_new_n3130_), .C(u2__abc_52138_new_n6766_), .Y(u2__abc_52138_new_n6773_));
OAI21X1 OAI21X1_641 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6774_), .Y(u2__abc_52138_new_n6775_));
OAI21X1 OAI21X1_642 ( .A(u2__abc_52138_new_n3125_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6775_), .Y(u2__abc_52138_new_n6776_));
OAI21X1 OAI21X1_643 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6776_), .C(u2__abc_52138_new_n6777_), .Y(u2__abc_52138_new_n6778_));
OAI21X1 OAI21X1_644 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_26_), .Y(u2__abc_52138_new_n6780_));
OAI21X1 OAI21X1_645 ( .A(sqrto_22_), .B(u2__abc_52138_new_n3130_), .C(u2__abc_52138_new_n3124_), .Y(u2__abc_52138_new_n6781_));
OAI21X1 OAI21X1_646 ( .A(u2__abc_52138_new_n3123_), .B(u2_remHi_23_), .C(u2__abc_52138_new_n6781_), .Y(u2__abc_52138_new_n6782_));
OAI21X1 OAI21X1_647 ( .A(u2__abc_52138_new_n6762_), .B(u2__abc_52138_new_n6756_), .C(u2__abc_52138_new_n3133_), .Y(u2__abc_52138_new_n6783_));
OAI21X1 OAI21X1_648 ( .A(u2__abc_52138_new_n3114_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6787_), .Y(u2__abc_52138_new_n6788_));
OAI21X1 OAI21X1_649 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6788_), .C(u2__abc_52138_new_n6789_), .Y(u2__abc_52138_new_n6790_));
OAI21X1 OAI21X1_65 ( .A(aNan), .B(_abc_65734_new_n1022_), .C(_abc_65734_new_n1023_), .Y(\o[176] ));
OAI21X1 OAI21X1_650 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_27_), .Y(u2__abc_52138_new_n6792_));
OAI21X1 OAI21X1_651 ( .A(sqrto_24_), .B(u2__abc_52138_new_n3114_), .C(u2__abc_52138_new_n6786_), .Y(u2__abc_52138_new_n6793_));
OAI21X1 OAI21X1_652 ( .A(u2__abc_52138_new_n3119_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6796_));
OAI21X1 OAI21X1_653 ( .A(u2__abc_52138_new_n6796_), .B(u2__abc_52138_new_n6795_), .C(u2__abc_52138_new_n6797_), .Y(u2__abc_52138_new_n6798_));
OAI21X1 OAI21X1_654 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_28_), .Y(u2__abc_52138_new_n6800_));
OAI21X1 OAI21X1_655 ( .A(u2__abc_52138_new_n3113_), .B(u2__abc_52138_new_n3121_), .C(u2__abc_52138_new_n3118_), .Y(u2__abc_52138_new_n6801_));
OAI21X1 OAI21X1_656 ( .A(u2__abc_52138_new_n6782_), .B(u2__abc_52138_new_n3221_), .C(u2__abc_52138_new_n6802_), .Y(u2__abc_52138_new_n6803_));
OAI21X1 OAI21X1_657 ( .A(u2__abc_52138_new_n3134_), .B(u2__abc_52138_new_n6763_), .C(u2__abc_52138_new_n6804_), .Y(u2__abc_52138_new_n6805_));
OAI21X1 OAI21X1_658 ( .A(u2__abc_52138_new_n3153_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6810_), .Y(u2__abc_52138_new_n6811_));
OAI21X1 OAI21X1_659 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6811_), .C(u2__abc_52138_new_n6812_), .Y(u2__abc_52138_new_n6813_));
OAI21X1 OAI21X1_66 ( .A(aNan), .B(_abc_65734_new_n1025_), .C(_abc_65734_new_n1026_), .Y(\o[177] ));
OAI21X1 OAI21X1_660 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_29_), .Y(u2__abc_52138_new_n6815_));
OAI21X1 OAI21X1_661 ( .A(u2__abc_52138_new_n3234_), .B(u2__abc_52138_new_n6806_), .C(u2__abc_52138_new_n3152_), .Y(u2__abc_52138_new_n6816_));
OAI21X1 OAI21X1_662 ( .A(u2__abc_52138_new_n3148_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6819_));
OAI21X1 OAI21X1_663 ( .A(u2__abc_52138_new_n6819_), .B(u2__abc_52138_new_n6818_), .C(u2__abc_52138_new_n6820_), .Y(u2__abc_52138_new_n6821_));
OAI21X1 OAI21X1_664 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_30_), .Y(u2__abc_52138_new_n6823_));
OAI21X1 OAI21X1_665 ( .A(sqrto_26_), .B(u2__abc_52138_new_n3153_), .C(u2__abc_52138_new_n3147_), .Y(u2__abc_52138_new_n6824_));
OAI21X1 OAI21X1_666 ( .A(u2__abc_52138_new_n6824_), .B(u2__abc_52138_new_n6808_), .C(u2__abc_52138_new_n3149_), .Y(u2__abc_52138_new_n6825_));
OAI21X1 OAI21X1_667 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6826_), .Y(u2__abc_52138_new_n6827_));
OAI21X1 OAI21X1_668 ( .A(u2__abc_52138_new_n3137_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6827_), .Y(u2__abc_52138_new_n6828_));
OAI21X1 OAI21X1_669 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6828_), .C(u2__abc_52138_new_n6829_), .Y(u2__abc_52138_new_n6830_));
OAI21X1 OAI21X1_67 ( .A(aNan), .B(_abc_65734_new_n1028_), .C(_abc_65734_new_n1029_), .Y(\o[178] ));
OAI21X1 OAI21X1_670 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_31_), .Y(u2__abc_52138_new_n6832_));
OAI21X1 OAI21X1_671 ( .A(u2__abc_52138_new_n3230_), .B(u2__abc_52138_new_n6825_), .C(u2__abc_52138_new_n3136_), .Y(u2__abc_52138_new_n6833_));
OAI21X1 OAI21X1_672 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6834_), .Y(u2__abc_52138_new_n6835_));
OAI21X1 OAI21X1_673 ( .A(u2__abc_52138_new_n3140_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6835_), .Y(u2__abc_52138_new_n6836_));
OAI21X1 OAI21X1_674 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6836_), .C(u2__abc_52138_new_n6837_), .Y(u2__abc_52138_new_n6838_));
OAI21X1 OAI21X1_675 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_32_), .Y(u2__abc_52138_new_n6840_));
OAI21X1 OAI21X1_676 ( .A(u2__abc_52138_new_n3136_), .B(u2__abc_52138_new_n3231_), .C(u2__abc_52138_new_n3143_), .Y(u2__abc_52138_new_n6842_));
OAI21X1 OAI21X1_677 ( .A(u2__abc_52138_new_n3157_), .B(u2__abc_52138_new_n6806_), .C(u2__abc_52138_new_n6843_), .Y(u2__abc_52138_new_n6844_));
OAI21X1 OAI21X1_678 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6845_), .Y(u2__abc_52138_new_n6846_));
OAI21X1 OAI21X1_679 ( .A(u2__abc_52138_new_n3391_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6846_), .Y(u2__abc_52138_new_n6847_));
OAI21X1 OAI21X1_68 ( .A(aNan), .B(_abc_65734_new_n1031_), .C(_abc_65734_new_n1032_), .Y(\o[179] ));
OAI21X1 OAI21X1_680 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6847_), .C(u2__abc_52138_new_n6849_), .Y(u2__abc_52138_new_n6850_));
OAI21X1 OAI21X1_681 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_33_), .Y(u2__abc_52138_new_n6852_));
OAI21X1 OAI21X1_682 ( .A(u2__abc_52138_new_n3434_), .B(u2__abc_52138_new_n6853_), .C(u2__abc_52138_new_n3390_), .Y(u2__abc_52138_new_n6854_));
OAI21X1 OAI21X1_683 ( .A(u2__abc_52138_new_n3396_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6857_));
OAI21X1 OAI21X1_684 ( .A(u2__abc_52138_new_n6857_), .B(u2__abc_52138_new_n6856_), .C(u2__abc_52138_new_n6858_), .Y(u2__abc_52138_new_n6859_));
OAI21X1 OAI21X1_685 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_34_), .Y(u2__abc_52138_new_n6861_));
OAI21X1 OAI21X1_686 ( .A(u2__abc_52138_new_n3435_), .B(u2__abc_52138_new_n6862_), .C(u2__abc_52138_new_n3395_), .Y(u2__abc_52138_new_n6863_));
OAI21X1 OAI21X1_687 ( .A(u2__abc_52138_new_n6848_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6866_), .Y(u2__abc_52138_new_n6867_));
OAI21X1 OAI21X1_688 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6867_), .C(u2__abc_52138_new_n6868_), .Y(u2__abc_52138_new_n6869_));
OAI21X1 OAI21X1_689 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_35_), .Y(u2__abc_52138_new_n6871_));
OAI21X1 OAI21X1_69 ( .A(aNan), .B(_abc_65734_new_n1034_), .C(_abc_65734_new_n1035_), .Y(\o[180] ));
OAI21X1 OAI21X1_690 ( .A(sqrto_32_), .B(u2__abc_52138_new_n6848_), .C(u2__abc_52138_new_n6865_), .Y(u2__abc_52138_new_n6872_));
OAI21X1 OAI21X1_691 ( .A(u2__abc_52138_new_n6873_), .B(u2__abc_52138_new_n6874_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6875_));
OAI21X1 OAI21X1_692 ( .A(u2__abc_52138_new_n3385_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6875_), .Y(u2__abc_52138_new_n6876_));
OAI21X1 OAI21X1_693 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6876_), .C(u2__abc_52138_new_n6877_), .Y(u2__abc_52138_new_n6878_));
OAI21X1 OAI21X1_694 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_36_), .Y(u2__abc_52138_new_n6880_));
OAI21X1 OAI21X1_695 ( .A(u2__abc_52138_new_n3390_), .B(u2__abc_52138_new_n3398_), .C(u2__abc_52138_new_n3395_), .Y(u2__abc_52138_new_n6881_));
OAI21X1 OAI21X1_696 ( .A(u2__abc_52138_new_n6882_), .B(u2__abc_52138_new_n3439_), .C(u2__abc_52138_new_n3384_), .Y(u2__abc_52138_new_n6883_));
OAI21X1 OAI21X1_697 ( .A(u2__abc_52138_new_n3400_), .B(u2__abc_52138_new_n6853_), .C(u2__abc_52138_new_n6884_), .Y(u2__abc_52138_new_n6885_));
OAI21X1 OAI21X1_698 ( .A(u2__abc_52138_new_n6886_), .B(u2__abc_52138_new_n6888_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6889_));
OAI21X1 OAI21X1_699 ( .A(u2_remHi_34_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6889_), .Y(u2__abc_52138_new_n6890_));
OAI21X1 OAI21X1_7 ( .A(aNan), .B(_abc_65734_new_n848_), .C(_abc_65734_new_n849_), .Y(\o[118] ));
OAI21X1 OAI21X1_70 ( .A(aNan), .B(_abc_65734_new_n1037_), .C(_abc_65734_new_n1038_), .Y(\o[181] ));
OAI21X1 OAI21X1_700 ( .A(u2_remHi_36_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6891_), .Y(u2__abc_52138_new_n6892_));
OAI21X1 OAI21X1_701 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_37_), .Y(u2__abc_52138_new_n6894_));
OAI21X1 OAI21X1_702 ( .A(sqrto_34_), .B(u2__abc_52138_new_n3443_), .C(u2__abc_52138_new_n6887_), .Y(u2__abc_52138_new_n6896_));
OAI21X1 OAI21X1_703 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6897_), .Y(u2__abc_52138_new_n6898_));
OAI21X1 OAI21X1_704 ( .A(u2__abc_52138_new_n3414_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6898_), .Y(u2__abc_52138_new_n6899_));
OAI21X1 OAI21X1_705 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6899_), .C(u2__abc_52138_new_n6900_), .Y(u2__abc_52138_new_n6901_));
OAI21X1 OAI21X1_706 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_38_), .Y(u2__abc_52138_new_n6903_));
OAI21X1 OAI21X1_707 ( .A(sqrto_34_), .B(u2__abc_52138_new_n3443_), .C(u2__abc_52138_new_n3413_), .Y(u2__abc_52138_new_n6905_));
OAI21X1 OAI21X1_708 ( .A(u2__abc_52138_new_n6905_), .B(u2__abc_52138_new_n6888_), .C(u2__abc_52138_new_n3415_), .Y(u2__abc_52138_new_n6906_));
OAI21X1 OAI21X1_709 ( .A(u2__abc_52138_new_n6904_), .B(u2__abc_52138_new_n3447_), .C(u2__abc_52138_new_n6906_), .Y(u2__abc_52138_new_n6907_));
OAI21X1 OAI21X1_71 ( .A(aNan), .B(_abc_65734_new_n1040_), .C(_abc_65734_new_n1041_), .Y(\o[182] ));
OAI21X1 OAI21X1_710 ( .A(u2__abc_52138_new_n3403_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6909_), .Y(u2__abc_52138_new_n6910_));
OAI21X1 OAI21X1_711 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6910_), .C(u2__abc_52138_new_n6911_), .Y(u2__abc_52138_new_n6912_));
OAI21X1 OAI21X1_712 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_39_), .Y(u2__abc_52138_new_n6914_));
OAI21X1 OAI21X1_713 ( .A(u2__abc_52138_new_n3447_), .B(u2__abc_52138_new_n6906_), .C(u2__abc_52138_new_n3402_), .Y(u2__abc_52138_new_n6915_));
OAI21X1 OAI21X1_714 ( .A(u2__abc_52138_new_n3408_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6918_));
OAI21X1 OAI21X1_715 ( .A(u2__abc_52138_new_n6918_), .B(u2__abc_52138_new_n6917_), .C(u2__abc_52138_new_n6919_), .Y(u2__abc_52138_new_n6920_));
OAI21X1 OAI21X1_716 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_40_), .Y(u2__abc_52138_new_n6922_));
OAI21X1 OAI21X1_717 ( .A(u2__abc_52138_new_n3412_), .B(u2_remHi_35_), .C(u2__abc_52138_new_n6905_), .Y(u2__abc_52138_new_n6925_));
OAI21X1 OAI21X1_718 ( .A(u2__abc_52138_new_n3429_), .B(u2__abc_52138_new_n6925_), .C(u2__abc_52138_new_n3407_), .Y(u2__abc_52138_new_n6926_));
OAI21X1 OAI21X1_719 ( .A(u2__abc_52138_new_n6930_), .B(u2__abc_52138_new_n6932_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6933_));
OAI21X1 OAI21X1_72 ( .A(aNan), .B(_abc_65734_new_n1043_), .C(_abc_65734_new_n1044_), .Y(\o[183] ));
OAI21X1 OAI21X1_720 ( .A(u2_remHi_38_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6933_), .Y(u2__abc_52138_new_n6934_));
OAI21X1 OAI21X1_721 ( .A(u2_remHi_40_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n6935_), .Y(u2__abc_52138_new_n6936_));
OAI21X1 OAI21X1_722 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_41_), .Y(u2__abc_52138_new_n6938_));
OAI21X1 OAI21X1_723 ( .A(sqrto_38_), .B(u2__abc_52138_new_n3348_), .C(u2__abc_52138_new_n6931_), .Y(u2__abc_52138_new_n6939_));
OAI21X1 OAI21X1_724 ( .A(u2__abc_52138_new_n3353_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6942_));
OAI21X1 OAI21X1_725 ( .A(u2__abc_52138_new_n6942_), .B(u2__abc_52138_new_n6941_), .C(u2__abc_52138_new_n6943_), .Y(u2__abc_52138_new_n6944_));
OAI21X1 OAI21X1_726 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_42_), .Y(u2__abc_52138_new_n6946_));
OAI21X1 OAI21X1_727 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n6949_), .Y(u2__abc_52138_new_n6950_));
OAI21X1 OAI21X1_728 ( .A(u2__abc_52138_new_n3337_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6950_), .Y(u2__abc_52138_new_n6951_));
OAI21X1 OAI21X1_729 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6951_), .C(u2__abc_52138_new_n6952_), .Y(u2__abc_52138_new_n6953_));
OAI21X1 OAI21X1_73 ( .A(aNan), .B(_abc_65734_new_n1046_), .C(_abc_65734_new_n1047_), .Y(\o[184] ));
OAI21X1 OAI21X1_730 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_43_), .Y(u2__abc_52138_new_n6955_));
OAI21X1 OAI21X1_731 ( .A(u2__abc_52138_new_n3339_), .B(u2__abc_52138_new_n6948_), .C(u2__abc_52138_new_n3336_), .Y(u2__abc_52138_new_n6958_));
OAI21X1 OAI21X1_732 ( .A(u2__abc_52138_new_n6957_), .B(u2__abc_52138_new_n6958_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n6959_));
OAI21X1 OAI21X1_733 ( .A(u2__abc_52138_new_n3342_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6961_));
OAI21X1 OAI21X1_734 ( .A(u2__abc_52138_new_n6961_), .B(u2__abc_52138_new_n6960_), .C(u2__abc_52138_new_n6962_), .Y(u2__abc_52138_new_n6963_));
OAI21X1 OAI21X1_735 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_44_), .Y(u2__abc_52138_new_n6965_));
OAI21X1 OAI21X1_736 ( .A(u2__abc_52138_new_n6966_), .B(u2__abc_52138_new_n6947_), .C(u2__abc_52138_new_n3354_), .Y(u2__abc_52138_new_n6967_));
OAI21X1 OAI21X1_737 ( .A(u2__abc_52138_new_n6967_), .B(u2__abc_52138_new_n3452_), .C(u2__abc_52138_new_n6969_), .Y(u2__abc_52138_new_n6970_));
OAI21X1 OAI21X1_738 ( .A(u2__abc_52138_new_n3376_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n6974_), .Y(u2__abc_52138_new_n6975_));
OAI21X1 OAI21X1_739 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n6975_), .C(u2__abc_52138_new_n6976_), .Y(u2__abc_52138_new_n6977_));
OAI21X1 OAI21X1_74 ( .A(aNan), .B(_abc_65734_new_n1049_), .C(_abc_65734_new_n1050_), .Y(\o[185] ));
OAI21X1 OAI21X1_740 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_45_), .Y(u2__abc_52138_new_n6979_));
OAI21X1 OAI21X1_741 ( .A(u2__abc_52138_new_n3378_), .B(u2__abc_52138_new_n6971_), .C(u2__abc_52138_new_n3375_), .Y(u2__abc_52138_new_n6980_));
OAI21X1 OAI21X1_742 ( .A(u2__abc_52138_new_n3371_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6983_));
OAI21X1 OAI21X1_743 ( .A(u2__abc_52138_new_n6983_), .B(u2__abc_52138_new_n6982_), .C(u2__abc_52138_new_n6984_), .Y(u2__abc_52138_new_n6985_));
OAI21X1 OAI21X1_744 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_46_), .Y(u2__abc_52138_new_n6987_));
OAI21X1 OAI21X1_745 ( .A(u2__abc_52138_new_n3360_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n6993_));
OAI21X1 OAI21X1_746 ( .A(u2__abc_52138_new_n6993_), .B(u2__abc_52138_new_n6992_), .C(u2__abc_52138_new_n6994_), .Y(u2__abc_52138_new_n6995_));
OAI21X1 OAI21X1_747 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_47_), .Y(u2__abc_52138_new_n6997_));
OAI21X1 OAI21X1_748 ( .A(u2__abc_52138_new_n3365_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7002_));
OAI21X1 OAI21X1_749 ( .A(u2__abc_52138_new_n7002_), .B(u2__abc_52138_new_n7001_), .C(u2__abc_52138_new_n7003_), .Y(u2__abc_52138_new_n7004_));
OAI21X1 OAI21X1_75 ( .A(aNan), .B(_abc_65734_new_n1052_), .C(_abc_65734_new_n1053_), .Y(\o[186] ));
OAI21X1 OAI21X1_750 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_48_), .Y(u2__abc_52138_new_n7006_));
OAI21X1 OAI21X1_751 ( .A(u2__abc_52138_new_n3375_), .B(u2__abc_52138_new_n6988_), .C(u2__abc_52138_new_n3370_), .Y(u2__abc_52138_new_n7007_));
OAI21X1 OAI21X1_752 ( .A(u2__abc_52138_new_n3359_), .B(u2__abc_52138_new_n3367_), .C(u2__abc_52138_new_n3364_), .Y(u2__abc_52138_new_n7008_));
OAI21X1 OAI21X1_753 ( .A(u2__abc_52138_new_n3427_), .B(u2__abc_52138_new_n6927_), .C(u2__abc_52138_new_n7009_), .Y(u2__abc_52138_new_n7010_));
OAI21X1 OAI21X1_754 ( .A(u2__abc_52138_new_n3420_), .B(u2__abc_52138_new_n6853_), .C(u2__abc_52138_new_n7011_), .Y(u2__abc_52138_new_n7012_));
OAI21X1 OAI21X1_755 ( .A(u2__abc_52138_new_n7013_), .B(u2__abc_52138_new_n7015_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7016_));
OAI21X1 OAI21X1_756 ( .A(u2_remHi_46_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7016_), .Y(u2__abc_52138_new_n7017_));
OAI21X1 OAI21X1_757 ( .A(u2_remHi_48_), .B(u2__abc_52138_new_n2978_), .C(u2__abc_52138_new_n7018_), .Y(u2__abc_52138_new_n7019_));
OAI21X1 OAI21X1_758 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_49_), .Y(u2__abc_52138_new_n7021_));
OAI21X1 OAI21X1_759 ( .A(u2__abc_52138_new_n3470_), .B(u2__abc_52138_new_n7014_), .C(u2__abc_52138_new_n3304_), .Y(u2__abc_52138_new_n7022_));
OAI21X1 OAI21X1_76 ( .A(aNan), .B(_abc_65734_new_n1055_), .C(_abc_65734_new_n1056_), .Y(\o[187] ));
OAI21X1 OAI21X1_760 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7023_), .Y(u2__abc_52138_new_n7024_));
OAI21X1 OAI21X1_761 ( .A(u2__abc_52138_new_n3298_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7024_), .Y(u2__abc_52138_new_n7025_));
OAI21X1 OAI21X1_762 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7025_), .C(u2__abc_52138_new_n7026_), .Y(u2__abc_52138_new_n7027_));
OAI21X1 OAI21X1_763 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_50_), .Y(u2__abc_52138_new_n7029_));
OAI21X1 OAI21X1_764 ( .A(sqrto_47_), .B(u2__abc_52138_new_n3298_), .C(u2__abc_52138_new_n3304_), .Y(u2__abc_52138_new_n7031_));
OAI21X1 OAI21X1_765 ( .A(u2__abc_52138_new_n7031_), .B(u2__abc_52138_new_n7015_), .C(u2__abc_52138_new_n7030_), .Y(u2__abc_52138_new_n7032_));
OAI21X1 OAI21X1_766 ( .A(u2__abc_52138_new_n3288_), .B(u2__abc_52138_new_n3290_), .C(u2__abc_52138_new_n7032_), .Y(u2__abc_52138_new_n7033_));
OAI21X1 OAI21X1_767 ( .A(u2__abc_52138_new_n3287_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7037_), .Y(u2__abc_52138_new_n7038_));
OAI21X1 OAI21X1_768 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7038_), .C(u2__abc_52138_new_n7039_), .Y(u2__abc_52138_new_n7040_));
OAI21X1 OAI21X1_769 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_51_), .Y(u2__abc_52138_new_n7042_));
OAI21X1 OAI21X1_77 ( .A(aNan), .B(_abc_65734_new_n1058_), .C(_abc_65734_new_n1059_), .Y(\o[188] ));
OAI21X1 OAI21X1_770 ( .A(u2__abc_52138_new_n3290_), .B(u2__abc_52138_new_n7032_), .C(u2__abc_52138_new_n7034_), .Y(u2__abc_52138_new_n7043_));
OAI21X1 OAI21X1_771 ( .A(u2__abc_52138_new_n3296_), .B(u2__abc_52138_new_n7043_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7044_));
OAI21X1 OAI21X1_772 ( .A(u2__abc_52138_new_n3292_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7046_));
OAI21X1 OAI21X1_773 ( .A(u2__abc_52138_new_n7046_), .B(u2__abc_52138_new_n7045_), .C(u2__abc_52138_new_n7047_), .Y(u2__abc_52138_new_n7048_));
OAI21X1 OAI21X1_774 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_52_), .Y(u2__abc_52138_new_n7050_));
OAI21X1 OAI21X1_775 ( .A(u2__abc_52138_new_n3300_), .B(u2_remHi_47_), .C(u2__abc_52138_new_n7031_), .Y(u2__abc_52138_new_n7051_));
OAI21X1 OAI21X1_776 ( .A(u2__abc_52138_new_n7034_), .B(u2__abc_52138_new_n3295_), .C(u2__abc_52138_new_n7052_), .Y(u2__abc_52138_new_n7053_));
OAI21X1 OAI21X1_777 ( .A(u2__abc_52138_new_n7051_), .B(u2__abc_52138_new_n3297_), .C(u2__abc_52138_new_n7054_), .Y(u2__abc_52138_new_n7055_));
OAI21X1 OAI21X1_778 ( .A(u2__abc_52138_new_n3329_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7059_), .Y(u2__abc_52138_new_n7060_));
OAI21X1 OAI21X1_779 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7060_), .C(u2__abc_52138_new_n7061_), .Y(u2__abc_52138_new_n7062_));
OAI21X1 OAI21X1_78 ( .A(aNan), .B(_abc_65734_new_n1061_), .C(_abc_65734_new_n1062_), .Y(\o[189] ));
OAI21X1 OAI21X1_780 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_53_), .Y(u2__abc_52138_new_n7064_));
OAI21X1 OAI21X1_781 ( .A(u2__abc_52138_new_n3331_), .B(u2__abc_52138_new_n7056_), .C(u2__abc_52138_new_n3328_), .Y(u2__abc_52138_new_n7065_));
OAI21X1 OAI21X1_782 ( .A(u2__abc_52138_new_n3324_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7068_));
OAI21X1 OAI21X1_783 ( .A(u2__abc_52138_new_n7068_), .B(u2__abc_52138_new_n7067_), .C(u2__abc_52138_new_n7069_), .Y(u2__abc_52138_new_n7070_));
OAI21X1 OAI21X1_784 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_54_), .Y(u2__abc_52138_new_n7072_));
OAI21X1 OAI21X1_785 ( .A(sqrto_51_), .B(u2__abc_52138_new_n3324_), .C(u2__abc_52138_new_n3328_), .Y(u2__abc_52138_new_n7074_));
OAI21X1 OAI21X1_786 ( .A(u2__abc_52138_new_n3313_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7079_));
OAI21X1 OAI21X1_787 ( .A(u2__abc_52138_new_n7079_), .B(u2__abc_52138_new_n7078_), .C(u2__abc_52138_new_n7080_), .Y(u2__abc_52138_new_n7081_));
OAI21X1 OAI21X1_788 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_55_), .Y(u2__abc_52138_new_n7083_));
OAI21X1 OAI21X1_789 ( .A(sqrto_52_), .B(u2__abc_52138_new_n3313_), .C(u2__abc_52138_new_n7084_), .Y(u2__abc_52138_new_n7085_));
OAI21X1 OAI21X1_79 ( .A(aNan), .B(_abc_65734_new_n1064_), .C(_abc_65734_new_n1065_), .Y(\o[190] ));
OAI21X1 OAI21X1_790 ( .A(u2__abc_52138_new_n3318_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7088_));
OAI21X1 OAI21X1_791 ( .A(u2__abc_52138_new_n7088_), .B(u2__abc_52138_new_n7087_), .C(u2__abc_52138_new_n7089_), .Y(u2__abc_52138_new_n7090_));
OAI21X1 OAI21X1_792 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_56_), .Y(u2__abc_52138_new_n7092_));
OAI21X1 OAI21X1_793 ( .A(u2__abc_52138_new_n3328_), .B(u2__abc_52138_new_n7073_), .C(u2__abc_52138_new_n3323_), .Y(u2__abc_52138_new_n7095_));
OAI21X1 OAI21X1_794 ( .A(u2__abc_52138_new_n3312_), .B(u2__abc_52138_new_n3482_), .C(u2__abc_52138_new_n3317_), .Y(u2__abc_52138_new_n7096_));
OAI21X1 OAI21X1_795 ( .A(u2__abc_52138_new_n7093_), .B(u2__abc_52138_new_n7094_), .C(u2__abc_52138_new_n7097_), .Y(u2__abc_52138_new_n7098_));
OAI21X1 OAI21X1_796 ( .A(u2__abc_52138_new_n3253_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7103_), .Y(u2__abc_52138_new_n7104_));
OAI21X1 OAI21X1_797 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7104_), .C(u2__abc_52138_new_n7105_), .Y(u2__abc_52138_new_n7106_));
OAI21X1 OAI21X1_798 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_57_), .Y(u2__abc_52138_new_n7108_));
OAI21X1 OAI21X1_799 ( .A(u2__abc_52138_new_n3258_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7109_));
OAI21X1 OAI21X1_8 ( .A(aNan), .B(_abc_65734_new_n851_), .C(_abc_65734_new_n852_), .Y(\o[119] ));
OAI21X1 OAI21X1_80 ( .A(aNan), .B(_abc_65734_new_n1067_), .C(_abc_65734_new_n1068_), .Y(\o[191] ));
OAI21X1 OAI21X1_800 ( .A(u2__abc_52138_new_n3488_), .B(u2__abc_52138_new_n7100_), .C(u2__abc_52138_new_n3252_), .Y(u2__abc_52138_new_n7110_));
OAI21X1 OAI21X1_801 ( .A(u2__abc_52138_new_n7109_), .B(u2__abc_52138_new_n7112_), .C(u2__abc_52138_new_n7113_), .Y(u2__abc_52138_new_n7114_));
OAI21X1 OAI21X1_802 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_58_), .Y(u2__abc_52138_new_n7116_));
OAI21X1 OAI21X1_803 ( .A(u2__abc_52138_new_n3489_), .B(u2__abc_52138_new_n7117_), .C(u2__abc_52138_new_n3257_), .Y(u2__abc_52138_new_n7118_));
OAI21X1 OAI21X1_804 ( .A(u2__abc_52138_new_n3242_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7121_));
OAI21X1 OAI21X1_805 ( .A(u2__abc_52138_new_n7121_), .B(u2__abc_52138_new_n7120_), .C(u2__abc_52138_new_n7122_), .Y(u2__abc_52138_new_n7123_));
OAI21X1 OAI21X1_806 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_59_), .Y(u2__abc_52138_new_n7125_));
OAI21X1 OAI21X1_807 ( .A(sqrto_56_), .B(u2__abc_52138_new_n3242_), .C(u2__abc_52138_new_n7126_), .Y(u2__abc_52138_new_n7127_));
OAI21X1 OAI21X1_808 ( .A(u2__abc_52138_new_n3247_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7130_));
OAI21X1 OAI21X1_809 ( .A(u2__abc_52138_new_n7130_), .B(u2__abc_52138_new_n7129_), .C(u2__abc_52138_new_n7131_), .Y(u2__abc_52138_new_n7132_));
OAI21X1 OAI21X1_81 ( .A(aNan), .B(_abc_65734_new_n1070_), .C(_abc_65734_new_n1071_), .Y(\o[192] ));
OAI21X1 OAI21X1_810 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_60_), .Y(u2__abc_52138_new_n7134_));
OAI21X1 OAI21X1_811 ( .A(u2__abc_52138_new_n3252_), .B(u2__abc_52138_new_n3260_), .C(u2__abc_52138_new_n3257_), .Y(u2__abc_52138_new_n7136_));
OAI21X1 OAI21X1_812 ( .A(u2__abc_52138_new_n3241_), .B(u2__abc_52138_new_n3249_), .C(u2__abc_52138_new_n3246_), .Y(u2__abc_52138_new_n7137_));
OAI21X1 OAI21X1_813 ( .A(u2__abc_52138_new_n3262_), .B(u2__abc_52138_new_n7100_), .C(u2__abc_52138_new_n7138_), .Y(u2__abc_52138_new_n7139_));
OAI21X1 OAI21X1_814 ( .A(u2__abc_52138_new_n7142_), .B(u2__abc_52138_new_n7141_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7143_));
OAI21X1 OAI21X1_815 ( .A(u2_remHi_58_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7143_), .Y(u2__abc_52138_new_n7144_));
OAI21X1 OAI21X1_816 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_61_), .Y(u2__abc_52138_new_n7149_));
OAI21X1 OAI21X1_817 ( .A(sqrto_58_), .B(u2__abc_52138_new_n3281_), .C(u2__abc_52138_new_n7140_), .Y(u2__abc_52138_new_n7150_));
OAI21X1 OAI21X1_818 ( .A(u2__abc_52138_new_n7152_), .B(u2__abc_52138_new_n7151_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7153_));
OAI21X1 OAI21X1_819 ( .A(u2_remHi_59_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7153_), .Y(u2__abc_52138_new_n7154_));
OAI21X1 OAI21X1_82 ( .A(aNan), .B(_abc_65734_new_n1073_), .C(_abc_65734_new_n1074_), .Y(\o[193] ));
OAI21X1 OAI21X1_820 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_62_), .Y(u2__abc_52138_new_n7159_));
OAI21X1 OAI21X1_821 ( .A(u2__abc_52138_new_n3265_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7164_));
OAI21X1 OAI21X1_822 ( .A(u2__abc_52138_new_n7164_), .B(u2__abc_52138_new_n7163_), .C(u2__abc_52138_new_n7165_), .Y(u2__abc_52138_new_n7166_));
OAI21X1 OAI21X1_823 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_63_), .Y(u2__abc_52138_new_n7168_));
OAI21X1 OAI21X1_824 ( .A(u2__abc_52138_new_n3267_), .B(u2__abc_52138_new_n7160_), .C(u2__abc_52138_new_n3264_), .Y(u2__abc_52138_new_n7169_));
OAI21X1 OAI21X1_825 ( .A(u2__abc_52138_new_n3268_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7172_));
OAI21X1 OAI21X1_826 ( .A(u2__abc_52138_new_n7172_), .B(u2__abc_52138_new_n7171_), .C(u2__abc_52138_new_n7173_), .Y(u2__abc_52138_new_n7174_));
OAI21X1 OAI21X1_827 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_64_), .Y(u2__abc_52138_new_n7176_));
OAI21X1 OAI21X1_828 ( .A(u2__abc_52138_new_n3280_), .B(u2__abc_52138_new_n3278_), .C(u2__abc_52138_new_n3275_), .Y(u2__abc_52138_new_n7178_));
OAI21X1 OAI21X1_829 ( .A(u2__abc_52138_new_n3264_), .B(u2__abc_52138_new_n3272_), .C(u2__abc_52138_new_n3271_), .Y(u2__abc_52138_new_n7179_));
OAI21X1 OAI21X1_83 ( .A(aNan), .B(_abc_65734_new_n1076_), .C(_abc_65734_new_n1077_), .Y(\o[194] ));
OAI21X1 OAI21X1_830 ( .A(u2__abc_52138_new_n3285_), .B(u2__abc_52138_new_n7138_), .C(u2__abc_52138_new_n7180_), .Y(u2__abc_52138_new_n7181_));
OAI21X1 OAI21X1_831 ( .A(u2__abc_52138_new_n3421_), .B(u2__abc_52138_new_n6853_), .C(u2__abc_52138_new_n7184_), .Y(u2__abc_52138_new_n7185_));
OAI21X1 OAI21X1_832 ( .A(u2__abc_52138_new_n3834_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7189_), .Y(u2__abc_52138_new_n7190_));
OAI21X1 OAI21X1_833 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7190_), .C(u2__abc_52138_new_n7191_), .Y(u2__abc_52138_new_n7192_));
OAI21X1 OAI21X1_834 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_65_), .Y(u2__abc_52138_new_n7194_));
OAI21X1 OAI21X1_835 ( .A(u2__abc_52138_new_n3841_), .B(u2__abc_52138_new_n7195_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7196_));
OAI21X1 OAI21X1_836 ( .A(u2__abc_52138_new_n3839_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7198_));
OAI21X1 OAI21X1_837 ( .A(u2__abc_52138_new_n7198_), .B(u2__abc_52138_new_n7197_), .C(u2__abc_52138_new_n7199_), .Y(u2__abc_52138_new_n7200_));
OAI21X1 OAI21X1_838 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_66_), .Y(u2__abc_52138_new_n7202_));
OAI21X1 OAI21X1_839 ( .A(u2__abc_52138_new_n3833_), .B(u2__abc_52138_new_n3875_), .C(u2__abc_52138_new_n3838_), .Y(u2__abc_52138_new_n7203_));
OAI21X1 OAI21X1_84 ( .A(aNan), .B(_abc_65734_new_n1079_), .C(_abc_65734_new_n1080_), .Y(\o[195] ));
OAI21X1 OAI21X1_840 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7205_), .Y(u2__abc_52138_new_n7206_));
OAI21X1 OAI21X1_841 ( .A(u2__abc_52138_new_n3845_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7206_), .Y(u2__abc_52138_new_n7207_));
OAI21X1 OAI21X1_842 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7207_), .C(u2__abc_52138_new_n7208_), .Y(u2__abc_52138_new_n7209_));
OAI21X1 OAI21X1_843 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_67_), .Y(u2__abc_52138_new_n7211_));
OAI21X1 OAI21X1_844 ( .A(u2__abc_52138_new_n3877_), .B(u2__abc_52138_new_n7204_), .C(u2__abc_52138_new_n3844_), .Y(u2__abc_52138_new_n7214_));
OAI21X1 OAI21X1_845 ( .A(u2__abc_52138_new_n7213_), .B(u2__abc_52138_new_n7214_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7215_));
OAI21X1 OAI21X1_846 ( .A(u2__abc_52138_new_n3850_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7217_));
OAI21X1 OAI21X1_847 ( .A(u2__abc_52138_new_n7217_), .B(u2__abc_52138_new_n7216_), .C(u2__abc_52138_new_n7218_), .Y(u2__abc_52138_new_n7219_));
OAI21X1 OAI21X1_848 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_68_), .Y(u2__abc_52138_new_n7221_));
OAI21X1 OAI21X1_849 ( .A(u2__abc_52138_new_n3873_), .B(u2__abc_52138_new_n7223_), .C(u2__abc_52138_new_n7225_), .Y(u2__abc_52138_new_n7226_));
OAI21X1 OAI21X1_85 ( .A(aNan), .B(_abc_65734_new_n1082_), .C(_abc_65734_new_n1083_), .Y(\o[196] ));
OAI21X1 OAI21X1_850 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7228_), .Y(u2__abc_52138_new_n7229_));
OAI21X1 OAI21X1_851 ( .A(u2__abc_52138_new_n3864_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7229_), .Y(u2__abc_52138_new_n7230_));
OAI21X1 OAI21X1_852 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7230_), .C(u2__abc_52138_new_n7231_), .Y(u2__abc_52138_new_n7232_));
OAI21X1 OAI21X1_853 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_69_), .Y(u2__abc_52138_new_n7234_));
OAI21X1 OAI21X1_854 ( .A(u2__abc_52138_new_n3886_), .B(u2__abc_52138_new_n7227_), .C(u2__abc_52138_new_n3863_), .Y(u2__abc_52138_new_n7235_));
OAI21X1 OAI21X1_855 ( .A(u2__abc_52138_new_n3883_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7238_));
OAI21X1 OAI21X1_856 ( .A(u2__abc_52138_new_n7238_), .B(u2__abc_52138_new_n7237_), .C(u2__abc_52138_new_n7239_), .Y(u2__abc_52138_new_n7240_));
OAI21X1 OAI21X1_857 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_70_), .Y(u2__abc_52138_new_n7242_));
OAI21X1 OAI21X1_858 ( .A(sqrto_67_), .B(u2__abc_52138_new_n3883_), .C(u2__abc_52138_new_n7243_), .Y(u2__abc_52138_new_n7244_));
OAI21X1 OAI21X1_859 ( .A(u2__abc_52138_new_n3855_), .B(u2__abc_52138_new_n7244_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7245_));
OAI21X1 OAI21X1_86 ( .A(aNan), .B(_abc_65734_new_n1085_), .C(_abc_65734_new_n1086_), .Y(\o[197] ));
OAI21X1 OAI21X1_860 ( .A(u2__abc_52138_new_n3888_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7247_));
OAI21X1 OAI21X1_861 ( .A(u2__abc_52138_new_n7247_), .B(u2__abc_52138_new_n7246_), .C(u2__abc_52138_new_n7248_), .Y(u2__abc_52138_new_n7249_));
OAI21X1 OAI21X1_862 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_71_), .Y(u2__abc_52138_new_n7251_));
OAI21X1 OAI21X1_863 ( .A(sqrto_68_), .B(u2__abc_52138_new_n3888_), .C(u2__abc_52138_new_n7253_), .Y(u2__abc_52138_new_n7254_));
OAI21X1 OAI21X1_864 ( .A(u2__abc_52138_new_n3858_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7257_));
OAI21X1 OAI21X1_865 ( .A(u2__abc_52138_new_n7257_), .B(u2__abc_52138_new_n7256_), .C(u2__abc_52138_new_n7258_), .Y(u2__abc_52138_new_n7259_));
OAI21X1 OAI21X1_866 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_72_), .Y(u2__abc_52138_new_n7261_));
OAI21X1 OAI21X1_867 ( .A(sqrto_66_), .B(u2__abc_52138_new_n3864_), .C(u2__abc_52138_new_n3882_), .Y(u2__abc_52138_new_n7262_));
OAI21X1 OAI21X1_868 ( .A(u2__abc_52138_new_n3881_), .B(u2_remHi_67_), .C(u2__abc_52138_new_n7262_), .Y(u2__abc_52138_new_n7263_));
OAI21X1 OAI21X1_869 ( .A(u2__abc_52138_new_n7265_), .B(u2__abc_52138_new_n7252_), .C(u2__abc_52138_new_n3857_), .Y(u2__abc_52138_new_n7266_));
OAI21X1 OAI21X1_87 ( .A(aNan), .B(_abc_65734_new_n1088_), .C(_abc_65734_new_n1089_), .Y(\o[198] ));
OAI21X1 OAI21X1_870 ( .A(u2__abc_52138_new_n3860_), .B(u2__abc_52138_new_n7263_), .C(u2__abc_52138_new_n7267_), .Y(u2__abc_52138_new_n7268_));
OAI21X1 OAI21X1_871 ( .A(u2__abc_52138_new_n3868_), .B(u2__abc_52138_new_n7186_), .C(u2__abc_52138_new_n7269_), .Y(u2__abc_52138_new_n7270_));
OAI21X1 OAI21X1_872 ( .A(u2__abc_52138_new_n3787_), .B(u2__abc_52138_new_n3789_), .C(u2__abc_52138_new_n7271_), .Y(u2__abc_52138_new_n7272_));
OAI21X1 OAI21X1_873 ( .A(u2__abc_52138_new_n3786_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7274_), .Y(u2__abc_52138_new_n7275_));
OAI21X1 OAI21X1_874 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7275_), .C(u2__abc_52138_new_n7276_), .Y(u2__abc_52138_new_n7277_));
OAI21X1 OAI21X1_875 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_73_), .Y(u2__abc_52138_new_n7279_));
OAI21X1 OAI21X1_876 ( .A(sqrto_70_), .B(u2__abc_52138_new_n3786_), .C(u2__abc_52138_new_n7273_), .Y(u2__abc_52138_new_n7280_));
OAI21X1 OAI21X1_877 ( .A(u2__abc_52138_new_n3795_), .B(u2__abc_52138_new_n7280_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7281_));
OAI21X1 OAI21X1_878 ( .A(u2__abc_52138_new_n3791_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7283_));
OAI21X1 OAI21X1_879 ( .A(u2__abc_52138_new_n7283_), .B(u2__abc_52138_new_n7282_), .C(u2__abc_52138_new_n7284_), .Y(u2__abc_52138_new_n7285_));
OAI21X1 OAI21X1_88 ( .A(aNan), .B(_abc_65734_new_n1091_), .C(_abc_65734_new_n1092_), .Y(\o[199] ));
OAI21X1 OAI21X1_880 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_74_), .Y(u2__abc_52138_new_n7287_));
OAI21X1 OAI21X1_881 ( .A(u2__abc_52138_new_n3793_), .B(u2_remHi_71_), .C(u2__abc_52138_new_n3787_), .Y(u2__abc_52138_new_n7288_));
OAI21X1 OAI21X1_882 ( .A(u2__abc_52138_new_n3796_), .B(u2__abc_52138_new_n7271_), .C(u2__abc_52138_new_n7289_), .Y(u2__abc_52138_new_n7290_));
OAI21X1 OAI21X1_883 ( .A(u2__abc_52138_new_n3799_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7293_));
OAI21X1 OAI21X1_884 ( .A(u2__abc_52138_new_n7293_), .B(u2__abc_52138_new_n7292_), .C(u2__abc_52138_new_n7294_), .Y(u2__abc_52138_new_n7295_));
OAI21X1 OAI21X1_885 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_75_), .Y(u2__abc_52138_new_n7297_));
OAI21X1 OAI21X1_886 ( .A(sqrto_72_), .B(u2__abc_52138_new_n3799_), .C(u2__abc_52138_new_n7299_), .Y(u2__abc_52138_new_n7300_));
OAI21X1 OAI21X1_887 ( .A(u2__abc_52138_new_n3804_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7303_));
OAI21X1 OAI21X1_888 ( .A(u2__abc_52138_new_n7303_), .B(u2__abc_52138_new_n7302_), .C(u2__abc_52138_new_n7304_), .Y(u2__abc_52138_new_n7305_));
OAI21X1 OAI21X1_889 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_76_), .Y(u2__abc_52138_new_n7307_));
OAI21X1 OAI21X1_89 ( .A(aNan), .B(_abc_65734_new_n1094_), .C(_abc_65734_new_n1095_), .Y(\o[200] ));
OAI21X1 OAI21X1_890 ( .A(u2__abc_52138_new_n3798_), .B(u2__abc_52138_new_n3898_), .C(u2__abc_52138_new_n3803_), .Y(u2__abc_52138_new_n7312_));
OAI21X1 OAI21X1_891 ( .A(u2__abc_52138_new_n7310_), .B(u2__abc_52138_new_n7271_), .C(u2__abc_52138_new_n7313_), .Y(u2__abc_52138_new_n7314_));
OAI21X1 OAI21X1_892 ( .A(u2__abc_52138_new_n7317_), .B(u2__abc_52138_new_n7316_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7318_));
OAI21X1 OAI21X1_893 ( .A(u2_remHi_74_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7318_), .Y(u2__abc_52138_new_n7319_));
OAI21X1 OAI21X1_894 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_77_), .Y(u2__abc_52138_new_n7324_));
OAI21X1 OAI21X1_895 ( .A(u2__abc_52138_new_n3825_), .B(u2__abc_52138_new_n7316_), .C(u2__abc_52138_new_n3823_), .Y(u2__abc_52138_new_n7325_));
OAI21X1 OAI21X1_896 ( .A(sqrto_74_), .B(u2__abc_52138_new_n3824_), .C(u2__abc_52138_new_n7315_), .Y(u2__abc_52138_new_n7327_));
OAI21X1 OAI21X1_897 ( .A(u2__abc_52138_new_n3823_), .B(u2__abc_52138_new_n7327_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7328_));
OAI21X1 OAI21X1_898 ( .A(u2__abc_52138_new_n3819_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7330_));
OAI21X1 OAI21X1_899 ( .A(u2__abc_52138_new_n7330_), .B(u2__abc_52138_new_n7329_), .C(u2__abc_52138_new_n7331_), .Y(u2__abc_52138_new_n7332_));
OAI21X1 OAI21X1_9 ( .A(aNan), .B(_abc_65734_new_n854_), .C(_abc_65734_new_n855_), .Y(\o[120] ));
OAI21X1 OAI21X1_90 ( .A(aNan), .B(_abc_65734_new_n1097_), .C(_abc_65734_new_n1098_), .Y(\o[201] ));
OAI21X1 OAI21X1_900 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_78_), .Y(u2__abc_52138_new_n7334_));
OAI21X1 OAI21X1_901 ( .A(u2__abc_52138_new_n3820_), .B(u2__abc_52138_new_n7326_), .C(u2__abc_52138_new_n3812_), .Y(u2__abc_52138_new_n7335_));
OAI21X1 OAI21X1_902 ( .A(u2__abc_52138_new_n3809_), .B(u2__abc_52138_new_n3811_), .C(u2__abc_52138_new_n7336_), .Y(u2__abc_52138_new_n7337_));
OAI21X1 OAI21X1_903 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7339_), .C(u2__abc_52138_new_n7340_), .Y(u2__abc_52138_new_n7341_));
OAI21X1 OAI21X1_904 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_79_), .Y(u2__abc_52138_new_n7343_));
OAI21X1 OAI21X1_905 ( .A(sqrto_76_), .B(u2__abc_52138_new_n3808_), .C(u2__abc_52138_new_n7335_), .Y(u2__abc_52138_new_n7344_));
OAI21X1 OAI21X1_906 ( .A(u2__abc_52138_new_n3817_), .B(u2__abc_52138_new_n7344_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7345_));
OAI21X1 OAI21X1_907 ( .A(u2__abc_52138_new_n3813_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7347_));
OAI21X1 OAI21X1_908 ( .A(u2__abc_52138_new_n7347_), .B(u2__abc_52138_new_n7346_), .C(u2__abc_52138_new_n7348_), .Y(u2__abc_52138_new_n7349_));
OAI21X1 OAI21X1_909 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_80_), .Y(u2__abc_52138_new_n7351_));
OAI21X1 OAI21X1_91 ( .A(aNan), .B(_abc_65734_new_n1100_), .C(_abc_65734_new_n1101_), .Y(\o[202] ));
OAI21X1 OAI21X1_910 ( .A(u2__abc_52138_new_n7358_), .B(u2__abc_52138_new_n3818_), .C(u2__abc_52138_new_n7359_), .Y(u2__abc_52138_new_n7360_));
OAI21X1 OAI21X1_911 ( .A(u2__abc_52138_new_n3831_), .B(u2__abc_52138_new_n7269_), .C(u2__abc_52138_new_n7361_), .Y(u2__abc_52138_new_n7362_));
OAI21X1 OAI21X1_912 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7364_), .Y(u2__abc_52138_new_n7365_));
OAI21X1 OAI21X1_913 ( .A(u2__abc_52138_new_n3740_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7365_), .Y(u2__abc_52138_new_n7366_));
OAI21X1 OAI21X1_914 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7366_), .C(u2__abc_52138_new_n7367_), .Y(u2__abc_52138_new_n7368_));
OAI21X1 OAI21X1_915 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_81_), .Y(u2__abc_52138_new_n7370_));
OAI21X1 OAI21X1_916 ( .A(u2__abc_52138_new_n3908_), .B(u2__abc_52138_new_n7363_), .C(u2__abc_52138_new_n3739_), .Y(u2__abc_52138_new_n7372_));
OAI21X1 OAI21X1_917 ( .A(u2__abc_52138_new_n7371_), .B(u2__abc_52138_new_n7372_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7373_));
OAI21X1 OAI21X1_918 ( .A(u2__abc_52138_new_n3745_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7375_));
OAI21X1 OAI21X1_919 ( .A(u2__abc_52138_new_n7375_), .B(u2__abc_52138_new_n7374_), .C(u2__abc_52138_new_n7376_), .Y(u2__abc_52138_new_n7377_));
OAI21X1 OAI21X1_92 ( .A(aNan), .B(_abc_65734_new_n1103_), .C(_abc_65734_new_n1104_), .Y(\o[203] ));
OAI21X1 OAI21X1_920 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_82_), .Y(u2__abc_52138_new_n7379_));
OAI21X1 OAI21X1_921 ( .A(u2__abc_52138_new_n3739_), .B(u2__abc_52138_new_n3909_), .C(u2__abc_52138_new_n3744_), .Y(u2__abc_52138_new_n7380_));
OAI21X1 OAI21X1_922 ( .A(u2__abc_52138_new_n3748_), .B(u2__abc_52138_new_n7363_), .C(u2__abc_52138_new_n7381_), .Y(u2__abc_52138_new_n7382_));
OAI21X1 OAI21X1_923 ( .A(u2__abc_52138_new_n3751_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7385_));
OAI21X1 OAI21X1_924 ( .A(u2__abc_52138_new_n7385_), .B(u2__abc_52138_new_n7384_), .C(u2__abc_52138_new_n7386_), .Y(u2__abc_52138_new_n7387_));
OAI21X1 OAI21X1_925 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_83_), .Y(u2__abc_52138_new_n7389_));
OAI21X1 OAI21X1_926 ( .A(sqrto_80_), .B(u2__abc_52138_new_n3751_), .C(u2__abc_52138_new_n7390_), .Y(u2__abc_52138_new_n7391_));
OAI21X1 OAI21X1_927 ( .A(u2__abc_52138_new_n3758_), .B(u2__abc_52138_new_n7391_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7392_));
OAI21X1 OAI21X1_928 ( .A(u2__abc_52138_new_n3756_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7394_));
OAI21X1 OAI21X1_929 ( .A(u2__abc_52138_new_n7394_), .B(u2__abc_52138_new_n7393_), .C(u2__abc_52138_new_n7395_), .Y(u2__abc_52138_new_n7396_));
OAI21X1 OAI21X1_93 ( .A(aNan), .B(_abc_65734_new_n1106_), .C(_abc_65734_new_n1107_), .Y(\o[204] ));
OAI21X1 OAI21X1_930 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_84_), .Y(u2__abc_52138_new_n7398_));
OAI21X1 OAI21X1_931 ( .A(u2__abc_52138_new_n3750_), .B(u2__abc_52138_new_n3912_), .C(u2__abc_52138_new_n3755_), .Y(u2__abc_52138_new_n7404_));
OAI21X1 OAI21X1_932 ( .A(u2__abc_52138_new_n7400_), .B(u2__abc_52138_new_n7363_), .C(u2__abc_52138_new_n7405_), .Y(u2__abc_52138_new_n7406_));
OAI21X1 OAI21X1_933 ( .A(u2__abc_52138_new_n7409_), .B(u2__abc_52138_new_n7408_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7410_));
OAI21X1 OAI21X1_934 ( .A(u2_remHi_82_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7410_), .Y(u2__abc_52138_new_n7411_));
OAI21X1 OAI21X1_935 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_85_), .Y(u2__abc_52138_new_n7416_));
OAI21X1 OAI21X1_936 ( .A(sqrto_82_), .B(u2__abc_52138_new_n3779_), .C(u2__abc_52138_new_n7407_), .Y(u2__abc_52138_new_n7417_));
OAI21X1 OAI21X1_937 ( .A(u2__abc_52138_new_n3774_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7420_));
OAI21X1 OAI21X1_938 ( .A(u2__abc_52138_new_n7420_), .B(u2__abc_52138_new_n7419_), .C(u2__abc_52138_new_n7421_), .Y(u2__abc_52138_new_n7422_));
OAI21X1 OAI21X1_939 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_86_), .Y(u2__abc_52138_new_n7424_));
OAI21X1 OAI21X1_94 ( .A(aNan), .B(_abc_65734_new_n1109_), .C(_abc_65734_new_n1110_), .Y(\o[205] ));
OAI21X1 OAI21X1_940 ( .A(sqrto_82_), .B(u2__abc_52138_new_n3779_), .C(u2__abc_52138_new_n3773_), .Y(u2__abc_52138_new_n7425_));
OAI21X1 OAI21X1_941 ( .A(u2__abc_52138_new_n7425_), .B(u2__abc_52138_new_n7408_), .C(u2__abc_52138_new_n3775_), .Y(u2__abc_52138_new_n7426_));
OAI21X1 OAI21X1_942 ( .A(u2__abc_52138_new_n6539_), .B(u2__abc_52138_new_n6541_), .C(u2__abc_52138_new_n7428_), .Y(u2__abc_52138_new_n7429_));
OAI21X1 OAI21X1_943 ( .A(u2__abc_52138_new_n3763_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7431_));
OAI21X1 OAI21X1_944 ( .A(u2__abc_52138_new_n7431_), .B(u2__abc_52138_new_n7430_), .C(u2__abc_52138_new_n7432_), .Y(u2__abc_52138_new_n7433_));
OAI21X1 OAI21X1_945 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_87_), .Y(u2__abc_52138_new_n7435_));
OAI21X1 OAI21X1_946 ( .A(u2__abc_52138_new_n3765_), .B(u2__abc_52138_new_n7426_), .C(u2__abc_52138_new_n3762_), .Y(u2__abc_52138_new_n7438_));
OAI21X1 OAI21X1_947 ( .A(u2__abc_52138_new_n7437_), .B(u2__abc_52138_new_n7438_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7439_));
OAI21X1 OAI21X1_948 ( .A(u2__abc_52138_new_n3768_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7441_));
OAI21X1 OAI21X1_949 ( .A(u2__abc_52138_new_n7441_), .B(u2__abc_52138_new_n7440_), .C(u2__abc_52138_new_n7442_), .Y(u2__abc_52138_new_n7443_));
OAI21X1 OAI21X1_95 ( .A(aNan), .B(_abc_65734_new_n1112_), .C(_abc_65734_new_n1113_), .Y(\o[206] ));
OAI21X1 OAI21X1_950 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_88_), .Y(u2__abc_52138_new_n7445_));
OAI21X1 OAI21X1_951 ( .A(u2__abc_52138_new_n3762_), .B(u2__abc_52138_new_n3770_), .C(u2__abc_52138_new_n3767_), .Y(u2__abc_52138_new_n7446_));
OAI21X1 OAI21X1_952 ( .A(u2__abc_52138_new_n3772_), .B(u2_remHi_83_), .C(u2__abc_52138_new_n7425_), .Y(u2__abc_52138_new_n7448_));
OAI21X1 OAI21X1_953 ( .A(u2__abc_52138_new_n3784_), .B(u2__abc_52138_new_n7363_), .C(u2__abc_52138_new_n7450_), .Y(u2__abc_52138_new_n7451_));
OAI21X1 OAI21X1_954 ( .A(u2__abc_52138_new_n7454_), .B(u2__abc_52138_new_n7453_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7455_));
OAI21X1 OAI21X1_955 ( .A(u2_remHi_86_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7455_), .Y(u2__abc_52138_new_n7456_));
OAI21X1 OAI21X1_956 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_89_), .Y(u2__abc_52138_new_n7461_));
OAI21X1 OAI21X1_957 ( .A(sqrto_86_), .B(u2__abc_52138_new_n3730_), .C(u2__abc_52138_new_n7452_), .Y(u2__abc_52138_new_n7463_));
OAI21X1 OAI21X1_958 ( .A(u2__abc_52138_new_n7462_), .B(u2__abc_52138_new_n7464_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7465_));
OAI21X1 OAI21X1_959 ( .A(u2__abc_52138_new_n3724_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7467_));
OAI21X1 OAI21X1_96 ( .A(aNan), .B(_abc_65734_new_n1115_), .C(_abc_65734_new_n1116_), .Y(\o[207] ));
OAI21X1 OAI21X1_960 ( .A(u2__abc_52138_new_n7467_), .B(u2__abc_52138_new_n7466_), .C(u2__abc_52138_new_n7468_), .Y(u2__abc_52138_new_n7469_));
OAI21X1 OAI21X1_961 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_90_), .Y(u2__abc_52138_new_n7471_));
OAI21X1 OAI21X1_962 ( .A(u2__abc_52138_new_n3728_), .B(u2__abc_52138_new_n7464_), .C(u2__abc_52138_new_n3726_), .Y(u2__abc_52138_new_n7473_));
OAI21X1 OAI21X1_963 ( .A(u2__abc_52138_new_n7472_), .B(u2__abc_52138_new_n7473_), .C(u2__abc_52138_new_n6499_), .Y(u2__abc_52138_new_n7476_));
OAI21X1 OAI21X1_964 ( .A(u2__abc_52138_new_n3715_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7478_));
OAI21X1 OAI21X1_965 ( .A(u2__abc_52138_new_n7478_), .B(u2__abc_52138_new_n7477_), .C(u2__abc_52138_new_n7479_), .Y(u2__abc_52138_new_n7480_));
OAI21X1 OAI21X1_966 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_91_), .Y(u2__abc_52138_new_n7482_));
OAI21X1 OAI21X1_967 ( .A(sqrto_88_), .B(u2__abc_52138_new_n3715_), .C(u2__abc_52138_new_n7474_), .Y(u2__abc_52138_new_n7483_));
OAI21X1 OAI21X1_968 ( .A(u2__abc_52138_new_n3720_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7486_));
OAI21X1 OAI21X1_969 ( .A(u2__abc_52138_new_n7486_), .B(u2__abc_52138_new_n7485_), .C(u2__abc_52138_new_n7487_), .Y(u2__abc_52138_new_n7488_));
OAI21X1 OAI21X1_97 ( .A(aNan), .B(_abc_65734_new_n1118_), .C(_abc_65734_new_n1119_), .Y(\o[208] ));
OAI21X1 OAI21X1_970 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_92_), .Y(u2__abc_52138_new_n7490_));
OAI21X1 OAI21X1_971 ( .A(sqrto_89_), .B(u2__abc_52138_new_n3720_), .C(u2__abc_52138_new_n3714_), .Y(u2__abc_52138_new_n7492_));
OAI21X1 OAI21X1_972 ( .A(u2__abc_52138_new_n7492_), .B(u2__abc_52138_new_n7475_), .C(u2__abc_52138_new_n3721_), .Y(u2__abc_52138_new_n7493_));
OAI21X1 OAI21X1_973 ( .A(u2__abc_52138_new_n3707_), .B(u2__abc_52138_new_n3709_), .C(u2__abc_52138_new_n7493_), .Y(u2__abc_52138_new_n7496_));
OAI21X1 OAI21X1_974 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7498_), .C(u2__abc_52138_new_n7499_), .Y(u2__abc_52138_new_n7500_));
OAI21X1 OAI21X1_975 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_93_), .Y(u2__abc_52138_new_n7502_));
OAI21X1 OAI21X1_976 ( .A(sqrto_90_), .B(u2__abc_52138_new_n3706_), .C(u2__abc_52138_new_n7495_), .Y(u2__abc_52138_new_n7504_));
OAI21X1 OAI21X1_977 ( .A(u2__abc_52138_new_n3704_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7507_));
OAI21X1 OAI21X1_978 ( .A(u2__abc_52138_new_n7507_), .B(u2__abc_52138_new_n7506_), .C(u2__abc_52138_new_n7508_), .Y(u2__abc_52138_new_n7509_));
OAI21X1 OAI21X1_979 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_94_), .Y(u2__abc_52138_new_n7511_));
OAI21X1 OAI21X1_98 ( .A(aNan), .B(_abc_65734_new_n1121_), .C(_abc_65734_new_n1122_), .Y(\o[209] ));
OAI21X1 OAI21X1_980 ( .A(sqrto_90_), .B(u2__abc_52138_new_n3706_), .C(u2__abc_52138_new_n3703_), .Y(u2__abc_52138_new_n7512_));
OAI21X1 OAI21X1_981 ( .A(u2__abc_52138_new_n3702_), .B(u2_remHi_91_), .C(u2__abc_52138_new_n7512_), .Y(u2__abc_52138_new_n7513_));
OAI21X1 OAI21X1_982 ( .A(u2__abc_52138_new_n3711_), .B(u2__abc_52138_new_n7493_), .C(u2__abc_52138_new_n7513_), .Y(u2__abc_52138_new_n7514_));
OAI21X1 OAI21X1_983 ( .A(u2__abc_52138_new_n3693_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7517_));
OAI21X1 OAI21X1_984 ( .A(u2__abc_52138_new_n7517_), .B(u2__abc_52138_new_n7516_), .C(u2__abc_52138_new_n7518_), .Y(u2__abc_52138_new_n7519_));
OAI21X1 OAI21X1_985 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_95_), .Y(u2__abc_52138_new_n7521_));
OAI21X1 OAI21X1_986 ( .A(u2__abc_52138_new_n3698_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n2978_), .Y(u2__abc_52138_new_n7526_));
OAI21X1 OAI21X1_987 ( .A(u2__abc_52138_new_n7526_), .B(u2__abc_52138_new_n7525_), .C(u2__abc_52138_new_n7527_), .Y(u2__abc_52138_new_n7528_));
OAI21X1 OAI21X1_988 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_96_), .Y(u2__abc_52138_new_n7530_));
OAI21X1 OAI21X1_989 ( .A(u2__abc_52138_new_n7446_), .B(u2__abc_52138_new_n7449_), .C(u2__abc_52138_new_n6484_), .Y(u2__abc_52138_new_n7532_));
OAI21X1 OAI21X1_99 ( .A(aNan), .B(_abc_65734_new_n1124_), .C(_abc_65734_new_n1125_), .Y(\o[210] ));
OAI21X1 OAI21X1_990 ( .A(u2__abc_52138_new_n3725_), .B(u2__abc_52138_new_n3731_), .C(u2__abc_52138_new_n3729_), .Y(u2__abc_52138_new_n7533_));
OAI21X1 OAI21X1_991 ( .A(u2__abc_52138_new_n3718_), .B(u2_remHi_89_), .C(u2__abc_52138_new_n7492_), .Y(u2__abc_52138_new_n7534_));
OAI21X1 OAI21X1_992 ( .A(u2__abc_52138_new_n7533_), .B(u2__abc_52138_new_n3723_), .C(u2__abc_52138_new_n7534_), .Y(u2__abc_52138_new_n7535_));
OAI21X1 OAI21X1_993 ( .A(u2__abc_52138_new_n7522_), .B(u2__abc_52138_new_n3932_), .C(u2__abc_52138_new_n3699_), .Y(u2__abc_52138_new_n7536_));
OAI21X1 OAI21X1_994 ( .A(u2__abc_52138_new_n7513_), .B(u2__abc_52138_new_n3701_), .C(u2__abc_52138_new_n7536_), .Y(u2__abc_52138_new_n7537_));
OAI21X1 OAI21X1_995 ( .A(u2__abc_52138_new_n7539_), .B(u2__abc_52138_new_n7540_), .C(u2__abc_52138_new_n7543_), .Y(u2__abc_52138_new_n7544_));
OAI21X1 OAI21X1_996 ( .A(u2__abc_52138_new_n3660_), .B(u2__abc_52138_new_n6499_), .C(u2__abc_52138_new_n7545_), .Y(u2__abc_52138_new_n7546_));
OAI21X1 OAI21X1_997 ( .A(u2__abc_52138_new_n6510_), .B(u2__abc_52138_new_n7546_), .C(u2__abc_52138_new_n7547_), .Y(u2__abc_52138_new_n7548_));
OAI21X1 OAI21X1_998 ( .A(u2__abc_52138_new_n2994_), .B(u2__abc_52138_new_n2983_), .C(u2_remHi_97_), .Y(u2__abc_52138_new_n7550_));
OAI21X1 OAI21X1_999 ( .A(sqrto_94_), .B(u2__abc_52138_new_n3660_), .C(u2__abc_52138_new_n7544_), .Y(u2__abc_52138_new_n7551_));
OAI22X1 OAI22X1_1 ( .A(u2__abc_52138_new_n3402_), .B(u2__abc_52138_new_n3448_), .C(u2__abc_52138_new_n3418_), .D(u2__abc_52138_new_n6884_), .Y(u2__abc_52138_new_n6924_));
OAI22X1 OAI22X1_10 ( .A(u2_remHi_351_), .B(u2__abc_52138_new_n5152_), .C(u2__abc_52138_new_n10331_), .D(u2__abc_52138_new_n10315_), .Y(u2__abc_52138_new_n10332_));
OAI22X1 OAI22X1_100 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11828_), .C(u2__abc_52138_new_n11827_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__130_));
OAI22X1 OAI22X1_101 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11837_), .C(u2__abc_52138_new_n11836_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__132_));
OAI22X1 OAI22X1_102 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11844_), .C(u2__abc_52138_new_n11843_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__134_));
OAI22X1 OAI22X1_103 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11847_), .C(u2__abc_52138_new_n11846_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__135_));
OAI22X1 OAI22X1_104 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11850_), .C(u2__abc_52138_new_n11849_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__136_));
OAI22X1 OAI22X1_105 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11853_), .C(u2__abc_52138_new_n11852_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__137_));
OAI22X1 OAI22X1_106 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11856_), .C(u2__abc_52138_new_n11855_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__138_));
OAI22X1 OAI22X1_107 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11859_), .C(u2__abc_52138_new_n11858_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__139_));
OAI22X1 OAI22X1_108 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11862_), .C(u2__abc_52138_new_n11861_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__140_));
OAI22X1 OAI22X1_109 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11865_), .C(u2__abc_52138_new_n11864_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__141_));
OAI22X1 OAI22X1_11 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11510_), .C(u2__abc_52138_new_n11507_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__32_));
OAI22X1 OAI22X1_110 ( .A(rst), .B(u2__abc_52138_new_n11868_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11867_), .Y(u2__0remLo_451_0__142_));
OAI22X1 OAI22X1_111 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11871_), .C(u2__abc_52138_new_n11870_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__143_));
OAI22X1 OAI22X1_112 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11874_), .C(u2__abc_52138_new_n11873_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__144_));
OAI22X1 OAI22X1_113 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11877_), .C(u2__abc_52138_new_n11876_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__145_));
OAI22X1 OAI22X1_114 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11880_), .C(u2__abc_52138_new_n11879_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__146_));
OAI22X1 OAI22X1_115 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11883_), .C(u2__abc_52138_new_n11882_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__147_));
OAI22X1 OAI22X1_116 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11886_), .C(u2__abc_52138_new_n11885_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__148_));
OAI22X1 OAI22X1_117 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11889_), .C(u2__abc_52138_new_n11888_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__149_));
OAI22X1 OAI22X1_118 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11892_), .C(u2__abc_52138_new_n11891_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__150_));
OAI22X1 OAI22X1_119 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11895_), .C(u2__abc_52138_new_n11894_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__151_));
OAI22X1 OAI22X1_12 ( .A(rst), .B(u2__abc_52138_new_n11519_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11518_), .Y(u2__0remLo_451_0__34_));
OAI22X1 OAI22X1_120 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11898_), .C(u2__abc_52138_new_n11897_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__152_));
OAI22X1 OAI22X1_121 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11901_), .C(u2__abc_52138_new_n11900_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__153_));
OAI22X1 OAI22X1_122 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11904_), .C(u2__abc_52138_new_n11903_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__154_));
OAI22X1 OAI22X1_123 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11907_), .C(u2__abc_52138_new_n11906_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__155_));
OAI22X1 OAI22X1_124 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11910_), .C(u2__abc_52138_new_n11909_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__156_));
OAI22X1 OAI22X1_125 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11913_), .C(u2__abc_52138_new_n11912_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__157_));
OAI22X1 OAI22X1_126 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11916_), .C(u2__abc_52138_new_n11915_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__158_));
OAI22X1 OAI22X1_127 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11919_), .C(u2__abc_52138_new_n11918_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__159_));
OAI22X1 OAI22X1_128 ( .A(rst), .B(u2__abc_52138_new_n11922_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11921_), .Y(u2__0remLo_451_0__160_));
OAI22X1 OAI22X1_129 ( .A(rst), .B(u2__abc_52138_new_n11925_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11924_), .Y(u2__0remLo_451_0__161_));
OAI22X1 OAI22X1_13 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11522_), .C(u2__abc_52138_new_n11521_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__35_));
OAI22X1 OAI22X1_130 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11928_), .C(u2__abc_52138_new_n11927_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__162_));
OAI22X1 OAI22X1_131 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11937_), .C(u2__abc_52138_new_n11936_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__164_));
OAI22X1 OAI22X1_132 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11940_), .C(u2__abc_52138_new_n11939_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__165_));
OAI22X1 OAI22X1_133 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11943_), .C(u2__abc_52138_new_n11942_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__166_));
OAI22X1 OAI22X1_134 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11946_), .C(u2__abc_52138_new_n11945_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__167_));
OAI22X1 OAI22X1_135 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11949_), .C(u2__abc_52138_new_n11948_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__168_));
OAI22X1 OAI22X1_136 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11952_), .C(u2__abc_52138_new_n11951_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__169_));
OAI22X1 OAI22X1_137 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11955_), .C(u2__abc_52138_new_n11954_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__170_));
OAI22X1 OAI22X1_138 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11958_), .C(u2__abc_52138_new_n11957_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__171_));
OAI22X1 OAI22X1_139 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11961_), .C(u2__abc_52138_new_n11960_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__172_));
OAI22X1 OAI22X1_14 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11531_), .C(u2__abc_52138_new_n11530_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__37_));
OAI22X1 OAI22X1_140 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11964_), .C(u2__abc_52138_new_n11963_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__173_));
OAI22X1 OAI22X1_141 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11971_), .C(u2__abc_52138_new_n11970_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__175_));
OAI22X1 OAI22X1_142 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11974_), .C(u2__abc_52138_new_n11973_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__176_));
OAI22X1 OAI22X1_143 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11977_), .C(u2__abc_52138_new_n11976_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__177_));
OAI22X1 OAI22X1_144 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11980_), .C(u2__abc_52138_new_n11979_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__178_));
OAI22X1 OAI22X1_145 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11983_), .C(u2__abc_52138_new_n11982_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__179_));
OAI22X1 OAI22X1_146 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11986_), .C(u2__abc_52138_new_n11985_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__180_));
OAI22X1 OAI22X1_147 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11989_), .C(u2__abc_52138_new_n11988_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__181_));
OAI22X1 OAI22X1_148 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11992_), .C(u2__abc_52138_new_n11991_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__182_));
OAI22X1 OAI22X1_149 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11995_), .C(u2__abc_52138_new_n11994_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__183_));
OAI22X1 OAI22X1_15 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11534_), .C(u2__abc_52138_new_n11533_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__38_));
OAI22X1 OAI22X1_150 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11998_), .C(u2__abc_52138_new_n11997_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__184_));
OAI22X1 OAI22X1_151 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12001_), .C(u2__abc_52138_new_n12000_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__185_));
OAI22X1 OAI22X1_152 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12004_), .C(u2__abc_52138_new_n12003_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__186_));
OAI22X1 OAI22X1_153 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12007_), .C(u2__abc_52138_new_n12006_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__187_));
OAI22X1 OAI22X1_154 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12010_), .C(u2__abc_52138_new_n12009_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__188_));
OAI22X1 OAI22X1_155 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12013_), .C(u2__abc_52138_new_n12012_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__189_));
OAI22X1 OAI22X1_156 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12016_), .C(u2__abc_52138_new_n12015_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__190_));
OAI22X1 OAI22X1_157 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12019_), .C(u2__abc_52138_new_n12018_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__191_));
OAI22X1 OAI22X1_158 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12022_), .C(u2__abc_52138_new_n12021_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__192_));
OAI22X1 OAI22X1_159 ( .A(rst), .B(u2__abc_52138_new_n12025_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n12024_), .Y(u2__0remLo_451_0__193_));
OAI22X1 OAI22X1_16 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11537_), .C(u2__abc_52138_new_n11536_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__39_));
OAI22X1 OAI22X1_160 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12028_), .C(u2__abc_52138_new_n12027_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__194_));
OAI22X1 OAI22X1_161 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12037_), .C(u2__abc_52138_new_n12036_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__196_));
OAI22X1 OAI22X1_162 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12040_), .C(u2__abc_52138_new_n12039_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__197_));
OAI22X1 OAI22X1_163 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12043_), .C(u2__abc_52138_new_n12042_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__198_));
OAI22X1 OAI22X1_164 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12046_), .C(u2__abc_52138_new_n12045_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__199_));
OAI22X1 OAI22X1_165 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12049_), .C(u2__abc_52138_new_n12048_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__200_));
OAI22X1 OAI22X1_166 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12052_), .C(u2__abc_52138_new_n12051_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__201_));
OAI22X1 OAI22X1_167 ( .A(rst), .B(u2__abc_52138_new_n12055_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n12054_), .Y(u2__0remLo_451_0__202_));
OAI22X1 OAI22X1_168 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12058_), .C(u2__abc_52138_new_n12057_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__203_));
OAI22X1 OAI22X1_169 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12067_), .C(u2__abc_52138_new_n12066_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__205_));
OAI22X1 OAI22X1_17 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11540_), .C(u2__abc_52138_new_n11539_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__40_));
OAI22X1 OAI22X1_170 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12074_), .C(u2__abc_52138_new_n12073_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__207_));
OAI22X1 OAI22X1_171 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12077_), .C(u2__abc_52138_new_n12076_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__208_));
OAI22X1 OAI22X1_172 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12080_), .C(u2__abc_52138_new_n12079_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__209_));
OAI22X1 OAI22X1_173 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12083_), .C(u2__abc_52138_new_n12082_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__210_));
OAI22X1 OAI22X1_174 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12086_), .C(u2__abc_52138_new_n12085_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__211_));
OAI22X1 OAI22X1_175 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12089_), .C(u2__abc_52138_new_n12088_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__212_));
OAI22X1 OAI22X1_176 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12092_), .C(u2__abc_52138_new_n12091_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__213_));
OAI22X1 OAI22X1_177 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12095_), .C(u2__abc_52138_new_n12094_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__214_));
OAI22X1 OAI22X1_178 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12098_), .C(u2__abc_52138_new_n12097_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__215_));
OAI22X1 OAI22X1_179 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12101_), .C(u2__abc_52138_new_n12100_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__216_));
OAI22X1 OAI22X1_18 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11543_), .C(u2__abc_52138_new_n11542_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__41_));
OAI22X1 OAI22X1_180 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12104_), .C(u2__abc_52138_new_n12103_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__217_));
OAI22X1 OAI22X1_181 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12107_), .C(u2__abc_52138_new_n12106_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__218_));
OAI22X1 OAI22X1_182 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12110_), .C(u2__abc_52138_new_n12109_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__219_));
OAI22X1 OAI22X1_183 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12113_), .C(u2__abc_52138_new_n12112_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__220_));
OAI22X1 OAI22X1_184 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12116_), .C(u2__abc_52138_new_n12115_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__221_));
OAI22X1 OAI22X1_185 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12119_), .C(u2__abc_52138_new_n12118_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__222_));
OAI22X1 OAI22X1_186 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12122_), .C(u2__abc_52138_new_n12121_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__223_));
OAI22X1 OAI22X1_187 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12125_), .C(u2__abc_52138_new_n12124_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__224_));
OAI22X1 OAI22X1_188 ( .A(rst), .B(u2__abc_52138_new_n12128_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n12127_), .Y(u2__0remLo_451_0__225_));
OAI22X1 OAI22X1_189 ( .A(rst), .B(u2__abc_52138_new_n12131_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n12130_), .Y(u2__0remLo_451_0__226_));
OAI22X1 OAI22X1_19 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11546_), .C(u2__abc_52138_new_n11545_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__42_));
OAI22X1 OAI22X1_190 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12146_), .C(u2__abc_52138_new_n12145_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__229_));
OAI22X1 OAI22X1_191 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12149_), .C(u2__abc_52138_new_n12148_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__230_));
OAI22X1 OAI22X1_192 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12152_), .C(u2__abc_52138_new_n12151_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__231_));
OAI22X1 OAI22X1_193 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12155_), .C(u2__abc_52138_new_n12154_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__232_));
OAI22X1 OAI22X1_194 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12158_), .C(u2__abc_52138_new_n12157_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__233_));
OAI22X1 OAI22X1_195 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12165_), .C(u2__abc_52138_new_n12164_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__235_));
OAI22X1 OAI22X1_196 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12168_), .C(u2__abc_52138_new_n12167_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__236_));
OAI22X1 OAI22X1_197 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12171_), .C(u2__abc_52138_new_n12170_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__237_));
OAI22X1 OAI22X1_198 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12174_), .C(u2__abc_52138_new_n12173_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__238_));
OAI22X1 OAI22X1_199 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12177_), .C(u2__abc_52138_new_n12176_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__239_));
OAI22X1 OAI22X1_2 ( .A(u2__abc_52138_new_n3915_), .B(u2__abc_52138_new_n7448_), .C(u2__abc_52138_new_n7447_), .D(u2__abc_52138_new_n7405_), .Y(u2__abc_52138_new_n7449_));
OAI22X1 OAI22X1_20 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11549_), .C(u2__abc_52138_new_n11548_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__43_));
OAI22X1 OAI22X1_200 ( .A(rst), .B(u2__abc_52138_new_n12180_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n12179_), .Y(u2__0remLo_451_0__240_));
OAI22X1 OAI22X1_201 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12183_), .C(u2__abc_52138_new_n12182_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__241_));
OAI22X1 OAI22X1_202 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12186_), .C(u2__abc_52138_new_n12185_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__242_));
OAI22X1 OAI22X1_203 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12189_), .C(u2__abc_52138_new_n12188_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__243_));
OAI22X1 OAI22X1_204 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12192_), .C(u2__abc_52138_new_n12191_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__244_));
OAI22X1 OAI22X1_205 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12195_), .C(u2__abc_52138_new_n12194_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__245_));
OAI22X1 OAI22X1_206 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12198_), .C(u2__abc_52138_new_n12197_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__246_));
OAI22X1 OAI22X1_207 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12201_), .C(u2__abc_52138_new_n12200_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__247_));
OAI22X1 OAI22X1_208 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12204_), .C(u2__abc_52138_new_n12203_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__248_));
OAI22X1 OAI22X1_209 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12207_), .C(u2__abc_52138_new_n12206_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__249_));
OAI22X1 OAI22X1_21 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11552_), .C(u2__abc_52138_new_n11551_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__44_));
OAI22X1 OAI22X1_210 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12210_), .C(u2__abc_52138_new_n12209_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__250_));
OAI22X1 OAI22X1_211 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12213_), .C(u2__abc_52138_new_n12212_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__251_));
OAI22X1 OAI22X1_212 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12216_), .C(u2__abc_52138_new_n12215_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__252_));
OAI22X1 OAI22X1_213 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12219_), .C(u2__abc_52138_new_n12218_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__253_));
OAI22X1 OAI22X1_214 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12222_), .C(u2__abc_52138_new_n12221_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__254_));
OAI22X1 OAI22X1_215 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n12225_), .C(u2__abc_52138_new_n12224_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__255_));
OAI22X1 OAI22X1_216 ( .A(rst), .B(u2__abc_52138_new_n12232_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n12231_), .Y(u2__0remLo_451_0__257_));
OAI22X1 OAI22X1_22 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11555_), .C(u2__abc_52138_new_n11554_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__45_));
OAI22X1 OAI22X1_23 ( .A(rst), .B(u2__abc_52138_new_n11558_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11557_), .Y(u2__0remLo_451_0__46_));
OAI22X1 OAI22X1_24 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11561_), .C(u2__abc_52138_new_n11560_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__47_));
OAI22X1 OAI22X1_25 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11570_), .C(u2__abc_52138_new_n11569_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__49_));
OAI22X1 OAI22X1_26 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11573_), .C(u2__abc_52138_new_n11572_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__50_));
OAI22X1 OAI22X1_27 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11576_), .C(u2__abc_52138_new_n11575_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__51_));
OAI22X1 OAI22X1_28 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11579_), .C(u2__abc_52138_new_n11578_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__52_));
OAI22X1 OAI22X1_29 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11582_), .C(u2__abc_52138_new_n11581_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__53_));
OAI22X1 OAI22X1_3 ( .A(u2__abc_52138_new_n3537_), .B(u2__abc_52138_new_n7894_), .C(u2__abc_52138_new_n7850_), .D(u2__abc_52138_new_n6488_), .Y(u2__abc_52138_new_n7895_));
OAI22X1 OAI22X1_30 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11585_), .C(u2__abc_52138_new_n11584_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__54_));
OAI22X1 OAI22X1_31 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11588_), .C(u2__abc_52138_new_n11587_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__55_));
OAI22X1 OAI22X1_32 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11591_), .C(u2__abc_52138_new_n11590_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__56_));
OAI22X1 OAI22X1_33 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11594_), .C(u2__abc_52138_new_n11593_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__57_));
OAI22X1 OAI22X1_34 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11597_), .C(u2__abc_52138_new_n11596_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__58_));
OAI22X1 OAI22X1_35 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11600_), .C(u2__abc_52138_new_n11599_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__59_));
OAI22X1 OAI22X1_36 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11603_), .C(u2__abc_52138_new_n11602_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__60_));
OAI22X1 OAI22X1_37 ( .A(rst), .B(u2__abc_52138_new_n11606_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11605_), .Y(u2__0remLo_451_0__61_));
OAI22X1 OAI22X1_38 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11609_), .C(u2__abc_52138_new_n11608_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__62_));
OAI22X1 OAI22X1_39 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11612_), .C(u2__abc_52138_new_n11611_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__63_));
OAI22X1 OAI22X1_4 ( .A(u2__abc_52138_new_n4227_), .B(u2__abc_52138_new_n8917_), .C(u2__abc_52138_new_n8897_), .D(u2__abc_52138_new_n8939_), .Y(u2__abc_52138_new_n8940_));
OAI22X1 OAI22X1_40 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11615_), .C(u2__abc_52138_new_n11614_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__64_));
OAI22X1 OAI22X1_41 ( .A(rst), .B(u2__abc_52138_new_n11618_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11617_), .Y(u2__0remLo_451_0__65_));
OAI22X1 OAI22X1_42 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11621_), .C(u2__abc_52138_new_n11620_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__66_));
OAI22X1 OAI22X1_43 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11630_), .C(u2__abc_52138_new_n11629_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__68_));
OAI22X1 OAI22X1_44 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11633_), .C(u2__abc_52138_new_n11632_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__69_));
OAI22X1 OAI22X1_45 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11636_), .C(u2__abc_52138_new_n11635_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__70_));
OAI22X1 OAI22X1_46 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11639_), .C(u2__abc_52138_new_n11638_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__71_));
OAI22X1 OAI22X1_47 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11642_), .C(u2__abc_52138_new_n11641_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__72_));
OAI22X1 OAI22X1_48 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11645_), .C(u2__abc_52138_new_n11644_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__73_));
OAI22X1 OAI22X1_49 ( .A(rst), .B(u2__abc_52138_new_n11648_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11647_), .Y(u2__0remLo_451_0__74_));
OAI22X1 OAI22X1_5 ( .A(u2__abc_52138_new_n5671_), .B(u2__abc_52138_new_n9400_), .C(u2__abc_52138_new_n5673_), .D(u2__abc_52138_new_n9382_), .Y(u2__abc_52138_new_n9439_));
OAI22X1 OAI22X1_50 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11651_), .C(u2__abc_52138_new_n11650_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__75_));
OAI22X1 OAI22X1_51 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11660_), .C(u2__abc_52138_new_n11659_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__77_));
OAI22X1 OAI22X1_52 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11663_), .C(u2__abc_52138_new_n11662_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__78_));
OAI22X1 OAI22X1_53 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11666_), .C(u2__abc_52138_new_n11665_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__79_));
OAI22X1 OAI22X1_54 ( .A(rst), .B(u2__abc_52138_new_n11669_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11668_), .Y(u2__0remLo_451_0__80_));
OAI22X1 OAI22X1_55 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11672_), .C(u2__abc_52138_new_n11671_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__81_));
OAI22X1 OAI22X1_56 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11675_), .C(u2__abc_52138_new_n11674_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__82_));
OAI22X1 OAI22X1_57 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11678_), .C(u2__abc_52138_new_n11677_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__83_));
OAI22X1 OAI22X1_58 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11681_), .C(u2__abc_52138_new_n11680_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__84_));
OAI22X1 OAI22X1_59 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11684_), .C(u2__abc_52138_new_n11683_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__85_));
OAI22X1 OAI22X1_6 ( .A(u2_remHi_271_), .B(u2__abc_52138_new_n5613_), .C(u2__abc_52138_new_n9465_), .D(u2__abc_52138_new_n9447_), .Y(u2__abc_52138_new_n9466_));
OAI22X1 OAI22X1_60 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11687_), .C(u2__abc_52138_new_n11686_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__86_));
OAI22X1 OAI22X1_61 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11690_), .C(u2__abc_52138_new_n11689_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__87_));
OAI22X1 OAI22X1_62 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11693_), .C(u2__abc_52138_new_n11692_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__88_));
OAI22X1 OAI22X1_63 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11696_), .C(u2__abc_52138_new_n11695_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__89_));
OAI22X1 OAI22X1_64 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11699_), .C(u2__abc_52138_new_n11698_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__90_));
OAI22X1 OAI22X1_65 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11702_), .C(u2__abc_52138_new_n11701_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__91_));
OAI22X1 OAI22X1_66 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11705_), .C(u2__abc_52138_new_n11704_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__92_));
OAI22X1 OAI22X1_67 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11708_), .C(u2__abc_52138_new_n11707_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__93_));
OAI22X1 OAI22X1_68 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11711_), .C(u2__abc_52138_new_n11710_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__94_));
OAI22X1 OAI22X1_69 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11714_), .C(u2__abc_52138_new_n11713_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__95_));
OAI22X1 OAI22X1_7 ( .A(u2_remHi_279_), .B(u2__abc_52138_new_n5566_), .C(u2__abc_52138_new_n9550_), .D(u2__abc_52138_new_n9534_), .Y(u2__abc_52138_new_n9551_));
OAI22X1 OAI22X1_70 ( .A(rst), .B(u2__abc_52138_new_n11722_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11721_), .Y(u2__0remLo_451_0__97_));
OAI22X1 OAI22X1_71 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11735_), .C(u2__abc_52138_new_n11734_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__100_));
OAI22X1 OAI22X1_72 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11738_), .C(u2__abc_52138_new_n11737_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__101_));
OAI22X1 OAI22X1_73 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11741_), .C(u2__abc_52138_new_n11740_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__102_));
OAI22X1 OAI22X1_74 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11744_), .C(u2__abc_52138_new_n11743_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__103_));
OAI22X1 OAI22X1_75 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11747_), .C(u2__abc_52138_new_n11746_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__104_));
OAI22X1 OAI22X1_76 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11750_), .C(u2__abc_52138_new_n11749_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__105_));
OAI22X1 OAI22X1_77 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11753_), .C(u2__abc_52138_new_n11752_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__106_));
OAI22X1 OAI22X1_78 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11756_), .C(u2__abc_52138_new_n11755_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__107_));
OAI22X1 OAI22X1_79 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11759_), .C(u2__abc_52138_new_n11758_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__108_));
OAI22X1 OAI22X1_8 ( .A(u2_remHi_287_), .B(u2__abc_52138_new_n5520_), .C(u2__abc_52138_new_n9640_), .D(u2__abc_52138_new_n9622_), .Y(u2__abc_52138_new_n9641_));
OAI22X1 OAI22X1_80 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11762_), .C(u2__abc_52138_new_n11761_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__109_));
OAI22X1 OAI22X1_81 ( .A(rst), .B(u2__abc_52138_new_n11765_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11764_), .Y(u2__0remLo_451_0__110_));
OAI22X1 OAI22X1_82 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11768_), .C(u2__abc_52138_new_n11767_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__111_));
OAI22X1 OAI22X1_83 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11771_), .C(u2__abc_52138_new_n11770_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__112_));
OAI22X1 OAI22X1_84 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11774_), .C(u2__abc_52138_new_n11773_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__113_));
OAI22X1 OAI22X1_85 ( .A(rst), .B(u2__abc_52138_new_n11777_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11776_), .Y(u2__0remLo_451_0__114_));
OAI22X1 OAI22X1_86 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11780_), .C(u2__abc_52138_new_n11779_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__115_));
OAI22X1 OAI22X1_87 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11789_), .C(u2__abc_52138_new_n11788_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__117_));
OAI22X1 OAI22X1_88 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11792_), .C(u2__abc_52138_new_n11791_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__118_));
OAI22X1 OAI22X1_89 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11795_), .C(u2__abc_52138_new_n11794_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__119_));
OAI22X1 OAI22X1_9 ( .A(u2__abc_52138_new_n5207_), .B(u2__abc_52138_new_n5213_), .C(u2__abc_52138_new_n5215_), .D(u2__abc_52138_new_n10306_), .Y(u2__abc_52138_new_n10307_));
OAI22X1 OAI22X1_90 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11798_), .C(u2__abc_52138_new_n11797_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__120_));
OAI22X1 OAI22X1_91 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11801_), .C(u2__abc_52138_new_n11800_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__121_));
OAI22X1 OAI22X1_92 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11804_), .C(u2__abc_52138_new_n11803_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__122_));
OAI22X1 OAI22X1_93 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11807_), .C(u2__abc_52138_new_n11806_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__123_));
OAI22X1 OAI22X1_94 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11810_), .C(u2__abc_52138_new_n11809_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__124_));
OAI22X1 OAI22X1_95 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11813_), .C(u2__abc_52138_new_n11812_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__125_));
OAI22X1 OAI22X1_96 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11816_), .C(u2__abc_52138_new_n11815_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__126_));
OAI22X1 OAI22X1_97 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11819_), .C(u2__abc_52138_new_n11818_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__127_));
OAI22X1 OAI22X1_98 ( .A(u2__abc_52138_new_n2986_), .B(u2__abc_52138_new_n11822_), .C(u2__abc_52138_new_n11821_), .D(u2__abc_52138_new_n11508_), .Y(u2__0remLo_451_0__128_));
OAI22X1 OAI22X1_99 ( .A(rst), .B(u2__abc_52138_new_n11825_), .C(u2__abc_52138_new_n2986_), .D(u2__abc_52138_new_n11824_), .Y(u2__0remLo_451_0__129_));
OR2X2 OR2X2_1 ( .A(aNan), .B(sqrto_188_), .Y(\o[224] ));
OR2X2 OR2X2_10 ( .A(u2__abc_52138_new_n3531_), .B(u2__abc_52138_new_n3536_), .Y(u2__abc_52138_new_n3537_));
OR2X2 OR2X2_100 ( .A(u2__abc_52138_new_n3187_), .B(u2__abc_52138_new_n3193_), .Y(u2__abc_52138_new_n12840_));
OR2X2 OR2X2_101 ( .A(u2__abc_52138_new_n3860_), .B(u2__abc_52138_new_n3866_), .Y(u2__abc_52138_new_n12890_));
OR2X2 OR2X2_102 ( .A(u2__abc_52138_new_n4240_), .B(u2__abc_52138_new_n4287_), .Y(u2__abc_52138_new_n12994_));
OR2X2 OR2X2_11 ( .A(u2__abc_52138_new_n3587_), .B(u2__abc_52138_new_n3592_), .Y(u2__abc_52138_new_n3593_));
OR2X2 OR2X2_12 ( .A(u2__abc_52138_new_n3601_), .B(u2__abc_52138_new_n3606_), .Y(u2__abc_52138_new_n3607_));
OR2X2 OR2X2_13 ( .A(u2__abc_52138_new_n3623_), .B(u2__abc_52138_new_n3628_), .Y(u2__abc_52138_new_n3629_));
OR2X2 OR2X2_14 ( .A(u2__abc_52138_new_n3657_), .B(u2__abc_52138_new_n3662_), .Y(u2__abc_52138_new_n3663_));
OR2X2 OR2X2_15 ( .A(u2__abc_52138_new_n3695_), .B(u2__abc_52138_new_n3700_), .Y(u2__abc_52138_new_n3701_));
OR2X2 OR2X2_16 ( .A(u2__abc_52138_new_n3717_), .B(u2__abc_52138_new_n3722_), .Y(u2__abc_52138_new_n3723_));
OR2X2 OR2X2_17 ( .A(u2__abc_52138_new_n3742_), .B(u2__abc_52138_new_n3747_), .Y(u2__abc_52138_new_n3748_));
OR2X2 OR2X2_18 ( .A(u2__abc_52138_new_n3765_), .B(u2__abc_52138_new_n3770_), .Y(u2__abc_52138_new_n3915_));
OR2X2 OR2X2_19 ( .A(u2__abc_52138_new_n3669_), .B(u2__abc_52138_new_n3674_), .Y(u2__abc_52138_new_n3947_));
OR2X2 OR2X2_2 ( .A(u2__abc_52138_new_n3134_), .B(u2__abc_52138_new_n3157_), .Y(u2__abc_52138_new_n3158_));
OR2X2 OR2X2_20 ( .A(u2__abc_52138_new_n3966_), .B(u2__abc_52138_new_n3622_), .Y(u2__abc_52138_new_n3967_));
OR2X2 OR2X2_21 ( .A(u2__abc_52138_new_n3565_), .B(u2__abc_52138_new_n3570_), .Y(u2__abc_52138_new_n3971_));
OR2X2 OR2X2_22 ( .A(u2__abc_52138_new_n3525_), .B(u2__abc_52138_new_n3519_), .Y(u2__abc_52138_new_n3989_));
OR2X2 OR2X2_23 ( .A(u2__abc_52138_new_n4025_), .B(u2__abc_52138_new_n4048_), .Y(u2__abc_52138_new_n4049_));
OR2X2 OR2X2_24 ( .A(u2__abc_52138_new_n4054_), .B(u2__abc_52138_new_n4059_), .Y(u2__abc_52138_new_n4060_));
OR2X2 OR2X2_25 ( .A(u2__abc_52138_new_n4127_), .B(u2__abc_52138_new_n4132_), .Y(u2__abc_52138_new_n4133_));
OR2X2 OR2X2_26 ( .A(u2__abc_52138_new_n4190_), .B(u2__abc_52138_new_n4168_), .Y(u2__abc_52138_new_n4191_));
OR2X2 OR2X2_27 ( .A(u2__abc_52138_new_n4198_), .B(u2__abc_52138_new_n4203_), .Y(u2__abc_52138_new_n4204_));
OR2X2 OR2X2_28 ( .A(u2__abc_52138_new_n4209_), .B(u2__abc_52138_new_n4214_), .Y(u2__abc_52138_new_n4215_));
OR2X2 OR2X2_29 ( .A(u2__abc_52138_new_n4221_), .B(u2__abc_52138_new_n4226_), .Y(u2__abc_52138_new_n4227_));
OR2X2 OR2X2_3 ( .A(u2__abc_52138_new_n3139_), .B(u2__abc_52138_new_n3144_), .Y(u2__abc_52138_new_n3229_));
OR2X2 OR2X2_30 ( .A(u2__abc_52138_new_n4245_), .B(u2__abc_52138_new_n4250_), .Y(u2__abc_52138_new_n4251_));
OR2X2 OR2X2_31 ( .A(u2__abc_52138_new_n4256_), .B(u2__abc_52138_new_n4261_), .Y(u2__abc_52138_new_n4262_));
OR2X2 OR2X2_32 ( .A(u2__abc_52138_new_n4329_), .B(u2__abc_52138_new_n4311_), .Y(u2__abc_52138_new_n4330_));
OR2X2 OR2X2_33 ( .A(u2__abc_52138_new_n4365_), .B(u2__abc_52138_new_n4367_), .Y(u2__abc_52138_new_n4368_));
OR2X2 OR2X2_34 ( .A(u2__abc_52138_new_n4518_), .B(u2__abc_52138_new_n4520_), .Y(u2__abc_52138_new_n4521_));
OR2X2 OR2X2_35 ( .A(u2__abc_52138_new_n4542_), .B(u2__abc_52138_new_n4544_), .Y(u2__abc_52138_new_n4545_));
OR2X2 OR2X2_36 ( .A(u2__abc_52138_new_n4725_), .B(u2__abc_52138_new_n4731_), .Y(u2__abc_52138_new_n4732_));
OR2X2 OR2X2_37 ( .A(u2__abc_52138_new_n4732_), .B(u2__abc_52138_new_n4750_), .Y(u2__abc_52138_new_n4751_));
OR2X2 OR2X2_38 ( .A(u2__abc_52138_new_n4617_), .B(u2__abc_52138_new_n4595_), .Y(u2__abc_52138_new_n4760_));
OR2X2 OR2X2_39 ( .A(u2__abc_52138_new_n4670_), .B(u2__abc_52138_new_n4675_), .Y(u2__abc_52138_new_n4785_));
OR2X2 OR2X2_4 ( .A(u2__abc_52138_new_n3334_), .B(u2__abc_52138_new_n3420_), .Y(u2__abc_52138_new_n3421_));
OR2X2 OR2X2_40 ( .A(u2__abc_52138_new_n4623_), .B(u2__abc_52138_new_n4628_), .Y(u2__abc_52138_new_n4806_));
OR2X2 OR2X2_41 ( .A(u2__abc_52138_new_n4529_), .B(u2__abc_52138_new_n4534_), .Y(u2__abc_52138_new_n4831_));
OR2X2 OR2X2_42 ( .A(u2__abc_52138_new_n4552_), .B(u2__abc_52138_new_n4557_), .Y(u2__abc_52138_new_n4837_));
OR2X2 OR2X2_43 ( .A(u2__abc_52138_new_n4335_), .B(u2__abc_52138_new_n4340_), .Y(u2__abc_52138_new_n4888_));
OR2X2 OR2X2_44 ( .A(u2__abc_52138_new_n4909_), .B(u2__abc_52138_new_n4315_), .Y(u2__abc_52138_new_n4910_));
OR2X2 OR2X2_45 ( .A(u2__abc_52138_new_n5031_), .B(u2__abc_52138_new_n5033_), .Y(u2__abc_52138_new_n5034_));
OR2X2 OR2X2_46 ( .A(u2__abc_52138_new_n5041_), .B(u2__abc_52138_new_n5034_), .Y(u2__abc_52138_new_n5042_));
OR2X2 OR2X2_47 ( .A(u2__abc_52138_new_n5101_), .B(u2__abc_52138_new_n5112_), .Y(u2__abc_52138_new_n5113_));
OR2X2 OR2X2_48 ( .A(u2__abc_52138_new_n5124_), .B(u2__abc_52138_new_n5131_), .Y(u2__abc_52138_new_n5132_));
OR2X2 OR2X2_49 ( .A(u2__abc_52138_new_n5113_), .B(u2__abc_52138_new_n5132_), .Y(u2__abc_52138_new_n5133_));
OR2X2 OR2X2_5 ( .A(u2__abc_52138_new_n3285_), .B(u2__abc_52138_new_n3262_), .Y(u2__abc_52138_new_n3422_));
OR2X2 OR2X2_50 ( .A(u2__abc_52138_new_n5215_), .B(u2__abc_52138_new_n5226_), .Y(u2__abc_52138_new_n5227_));
OR2X2 OR2X2_51 ( .A(u2__abc_52138_new_n5362_), .B(u2__abc_52138_new_n5351_), .Y(u2__abc_52138_new_n5363_));
OR2X2 OR2X2_52 ( .A(u2__abc_52138_new_n5732_), .B(u2__abc_52138_new_n5686_), .Y(u2__abc_52138_new_n5733_));
OR2X2 OR2X2_53 ( .A(u2__abc_52138_new_n5752_), .B(u2__abc_52138_new_n5650_), .Y(u2__abc_52138_new_n5753_));
OR2X2 OR2X2_54 ( .A(u2__abc_52138_new_n5232_), .B(u2__abc_52138_new_n5237_), .Y(u2__abc_52138_new_n5873_));
OR2X2 OR2X2_55 ( .A(u2__abc_52138_new_n5900_), .B(u2__abc_52138_new_n5044_), .Y(u2__abc_52138_new_n5901_));
OR2X2 OR2X2_56 ( .A(u2__abc_52138_new_n6422_), .B(u2__abc_52138_new_n5954_), .Y(u2__abc_52138_new_n6423_));
OR2X2 OR2X2_57 ( .A(u2__abc_52138_new_n6476_), .B(u2__abc_52138_new_n6475_), .Y(u2__abc_52138_new_n6477_));
OR2X2 OR2X2_58 ( .A(u2__abc_52138_new_n3547_), .B(u2__abc_52138_new_n3537_), .Y(u2__abc_52138_new_n6488_));
OR2X2 OR2X2_59 ( .A(u2__abc_52138_new_n6520_), .B(u2__abc_52138_new_n3066_), .Y(u2__abc_52138_new_n6522_));
OR2X2 OR2X2_6 ( .A(u2__abc_52138_new_n3339_), .B(u2__abc_52138_new_n3344_), .Y(u2__abc_52138_new_n3452_));
OR2X2 OR2X2_60 ( .A(u2__abc_52138_new_n6529_), .B(u2__abc_52138_new_n3067_), .Y(u2__abc_52138_new_n6530_));
OR2X2 OR2X2_61 ( .A(u2__abc_52138_new_n6626_), .B(u2__abc_52138_new_n3031_), .Y(u2__abc_52138_new_n6627_));
OR2X2 OR2X2_62 ( .A(u2__abc_52138_new_n6674_), .B(u2__abc_52138_new_n3174_), .Y(u2__abc_52138_new_n6676_));
OR2X2 OR2X2_63 ( .A(u2__abc_52138_new_n6693_), .B(u2__abc_52138_new_n3163_), .Y(u2__abc_52138_new_n6695_));
OR2X2 OR2X2_64 ( .A(u2__abc_52138_new_n6716_), .B(u2__abc_52138_new_n6711_), .Y(u2__abc_52138_new_n6718_));
OR2X2 OR2X2_65 ( .A(u2__abc_52138_new_n6784_), .B(u2__abc_52138_new_n3219_), .Y(u2__abc_52138_new_n6785_));
OR2X2 OR2X2_66 ( .A(u2__abc_52138_new_n6863_), .B(u2__abc_52138_new_n3432_), .Y(u2__abc_52138_new_n6864_));
OR2X2 OR2X2_67 ( .A(u2__abc_52138_new_n6906_), .B(u2__abc_52138_new_n3405_), .Y(u2__abc_52138_new_n6908_));
OR2X2 OR2X2_68 ( .A(u2__abc_52138_new_n6971_), .B(u2__abc_52138_new_n3378_), .Y(u2__abc_52138_new_n6973_));
OR2X2 OR2X2_69 ( .A(u2__abc_52138_new_n7032_), .B(u2__abc_52138_new_n7035_), .Y(u2__abc_52138_new_n7036_));
OR2X2 OR2X2_7 ( .A(u2__abc_52138_new_n3315_), .B(u2__abc_52138_new_n3320_), .Y(u2__abc_52138_new_n3477_));
OR2X2 OR2X2_70 ( .A(u2__abc_52138_new_n7056_), .B(u2__abc_52138_new_n3331_), .Y(u2__abc_52138_new_n7058_));
OR2X2 OR2X2_71 ( .A(u2__abc_52138_new_n7100_), .B(u2__abc_52138_new_n3255_), .Y(u2__abc_52138_new_n7102_));
OR2X2 OR2X2_72 ( .A(u2__abc_52138_new_n7160_), .B(u2__abc_52138_new_n3267_), .Y(u2__abc_52138_new_n7161_));
OR2X2 OR2X2_73 ( .A(u2__abc_52138_new_n7177_), .B(u2__abc_52138_new_n7181_), .Y(u2__abc_52138_new_n7182_));
OR2X2 OR2X2_74 ( .A(u2__abc_52138_new_n7186_), .B(u2__abc_52138_new_n3836_), .Y(u2__abc_52138_new_n7188_));
OR2X2 OR2X2_75 ( .A(u2__abc_52138_new_n3748_), .B(u2__abc_52138_new_n3759_), .Y(u2__abc_52138_new_n7400_));
OR2X2 OR2X2_76 ( .A(u2__abc_52138_new_n3707_), .B(u2__abc_52138_new_n3709_), .Y(u2__abc_52138_new_n7491_));
OR2X2 OR2X2_77 ( .A(u2__abc_52138_new_n3574_), .B(u2__abc_52138_new_n3576_), .Y(u2__abc_52138_new_n7802_));
OR2X2 OR2X2_78 ( .A(u2__abc_52138_new_n7810_), .B(u2__abc_52138_new_n3507_), .Y(u2__abc_52138_new_n7811_));
OR2X2 OR2X2_79 ( .A(u2__abc_52138_new_n3690_), .B(u2__abc_52138_new_n3870_), .Y(u2__abc_52138_new_n7888_));
OR2X2 OR2X2_8 ( .A(u2__abc_52138_new_n3244_), .B(u2__abc_52138_new_n3249_), .Y(u2__abc_52138_new_n3487_));
OR2X2 OR2X2_80 ( .A(u2__abc_52138_new_n4608_), .B(u2__abc_52138_new_n4613_), .Y(u2__abc_52138_new_n8230_));
OR2X2 OR2X2_81 ( .A(u2__abc_52138_new_n8248_), .B(u2__abc_52138_new_n8252_), .Y(u2__abc_52138_new_n8253_));
OR2X2 OR2X2_82 ( .A(u2__abc_52138_new_n4467_), .B(u2__abc_52138_new_n4473_), .Y(u2__abc_52138_new_n8449_));
OR2X2 OR2X2_83 ( .A(u2__abc_52138_new_n4404_), .B(u2__abc_52138_new_n4427_), .Y(u2__abc_52138_new_n8591_));
OR2X2 OR2X2_84 ( .A(u2__abc_52138_new_n8593_), .B(u2__abc_52138_new_n8598_), .Y(u2__abc_52138_new_n8599_));
OR2X2 OR2X2_85 ( .A(u2__abc_52138_new_n4274_), .B(u2__abc_52138_new_n4285_), .Y(u2__abc_52138_new_n8854_));
OR2X2 OR2X2_86 ( .A(u2__abc_52138_new_n4204_), .B(u2__abc_52138_new_n4215_), .Y(u2__abc_52138_new_n8895_));
OR2X2 OR2X2_87 ( .A(u2__abc_52138_new_n4227_), .B(u2__abc_52138_new_n4238_), .Y(u2__abc_52138_new_n8939_));
OR2X2 OR2X2_88 ( .A(u2__abc_52138_new_n4181_), .B(u2__abc_52138_new_n4186_), .Y(u2__abc_52138_new_n9002_));
OR2X2 OR2X2_89 ( .A(u2__abc_52138_new_n9188_), .B(u2__abc_52138_new_n4007_), .Y(u2__abc_52138_new_n9189_));
OR2X2 OR2X2_9 ( .A(u2__abc_52138_new_n3272_), .B(u2__abc_52138_new_n3266_), .Y(u2__abc_52138_new_n3497_));
OR2X2 OR2X2_90 ( .A(u2__abc_52138_new_n4097_), .B(u2__abc_52138_new_n4049_), .Y(u2__abc_52138_new_n9269_));
OR2X2 OR2X2_91 ( .A(u2__abc_52138_new_n9228_), .B(u2__abc_52138_new_n4048_), .Y(u2__abc_52138_new_n9270_));
OR2X2 OR2X2_92 ( .A(u2__abc_52138_new_n9615_), .B(u2__abc_52138_new_n5577_), .Y(u2__abc_52138_new_n9616_));
OR2X2 OR2X2_93 ( .A(u2__abc_52138_new_n9618_), .B(u2__abc_52138_new_n9613_), .Y(u2__abc_52138_new_n9619_));
OR2X2 OR2X2_94 ( .A(u2__abc_52138_new_n5512_), .B(u2__abc_52138_new_n5523_), .Y(u2__abc_52138_new_n9660_));
OR2X2 OR2X2_95 ( .A(u2__abc_52138_new_n5217_), .B(u2__abc_52138_new_n5222_), .Y(u2__abc_52138_new_n10286_));
OR2X2 OR2X2_96 ( .A(u2__abc_52138_new_n10307_), .B(u2__abc_52138_new_n5211_), .Y(u2__abc_52138_new_n10308_));
OR2X2 OR2X2_97 ( .A(u2__abc_52138_new_n10588_), .B(u2__abc_52138_new_n5034_), .Y(u2__abc_52138_new_n10589_));
OR2X2 OR2X2_98 ( .A(u2__abc_52138_new_n11004_), .B(u2__abc_52138_new_n6214_), .Y(u2__abc_52138_new_n11005_));
OR2X2 OR2X2_99 ( .A(u2__abc_52138_new_n6022_), .B(u2__abc_52138_new_n6029_), .Y(u2__abc_52138_new_n11224_));
XNOR2X1 XNOR2X1_1 ( .A(_abc_65734_new_n1492_), .B(\a[119] ), .Y(_abc_65734_new_n1506_));
XNOR2X1 XNOR2X1_10 ( .A(sqrto_4_), .B(u2_remHi_4_), .Y(u2__abc_52138_new_n3053_));
XNOR2X1 XNOR2X1_100 ( .A(u2__abc_52138_new_n10190_), .B(u2__abc_52138_new_n5270_), .Y(u2__abc_52138_new_n10191_));
XNOR2X1 XNOR2X1_101 ( .A(u2__abc_52138_new_n10234_), .B(u2__abc_52138_new_n5204_), .Y(u2__abc_52138_new_n10235_));
XNOR2X1 XNOR2X1_102 ( .A(u2__abc_52138_new_n10277_), .B(u2__abc_52138_new_n5225_), .Y(u2__abc_52138_new_n10278_));
XNOR2X1 XNOR2X1_103 ( .A(u2__abc_52138_new_n10323_), .B(u2__abc_52138_new_n5154_), .Y(u2__abc_52138_new_n10324_));
XNOR2X1 XNOR2X1_104 ( .A(u2__abc_52138_new_n10366_), .B(u2__abc_52138_new_n5177_), .Y(u2__abc_52138_new_n10367_));
XNOR2X1 XNOR2X1_105 ( .A(u2__abc_52138_new_n10453_), .B(u2__abc_52138_new_n5130_), .Y(u2__abc_52138_new_n10454_));
XNOR2X1 XNOR2X1_106 ( .A(u2__abc_52138_new_n10497_), .B(u2__abc_52138_new_n5062_), .Y(u2__abc_52138_new_n10498_));
XNOR2X1 XNOR2X1_107 ( .A(u2__abc_52138_new_n10618_), .B(u2__abc_52138_new_n5015_), .Y(u2__abc_52138_new_n10619_));
XNOR2X1 XNOR2X1_108 ( .A(u2__abc_52138_new_n10714_), .B(u2__abc_52138_new_n6151_), .Y(u2__abc_52138_new_n10715_));
XNOR2X1 XNOR2X1_109 ( .A(u2__abc_52138_new_n10803_), .B(u2__abc_52138_new_n6319_), .Y(u2__abc_52138_new_n10804_));
XNOR2X1 XNOR2X1_11 ( .A(sqrto_3_), .B(u2_remHi_3_), .Y(u2__abc_52138_new_n3059_));
XNOR2X1 XNOR2X1_110 ( .A(u2__abc_52138_new_n10887_), .B(u2__abc_52138_new_n6270_), .Y(u2__abc_52138_new_n10888_));
XNOR2X1 XNOR2X1_111 ( .A(u2__abc_52138_new_n10931_), .B(u2__abc_52138_new_n6200_), .Y(u2__abc_52138_new_n10932_));
XNOR2X1 XNOR2X1_112 ( .A(u2__abc_52138_new_n10975_), .B(u2__abc_52138_new_n6223_), .Y(u2__abc_52138_new_n10976_));
XNOR2X1 XNOR2X1_113 ( .A(u2__abc_52138_new_n11021_), .B(u2__abc_52138_new_n6124_), .Y(u2__abc_52138_new_n11022_));
XNOR2X1 XNOR2X1_114 ( .A(u2__abc_52138_new_n11066_), .B(u2__abc_52138_new_n6100_), .Y(u2__abc_52138_new_n11067_));
XNOR2X1 XNOR2X1_115 ( .A(u2__abc_52138_new_n11109_), .B(u2__abc_52138_new_n6056_), .Y(u2__abc_52138_new_n11110_));
XNOR2X1 XNOR2X1_116 ( .A(u2__abc_52138_new_n11150_), .B(u2__abc_52138_new_n6074_), .Y(u2__abc_52138_new_n11151_));
XNOR2X1 XNOR2X1_117 ( .A(u2__abc_52138_new_n11323_), .B(u2__abc_52138_new_n5959_), .Y(u2__abc_52138_new_n11324_));
XNOR2X1 XNOR2X1_118 ( .A(u2__abc_52138_new_n11409_), .B(u2_cnt_7_), .Y(u2__abc_52138_new_n11410_));
XNOR2X1 XNOR2X1_12 ( .A(u2_remHi_0_), .B(sqrto_0_), .Y(u2__abc_52138_new_n3066_));
XNOR2X1 XNOR2X1_13 ( .A(sqrto_1_), .B(u2_remHi_1_), .Y(u2__abc_52138_new_n3067_));
XNOR2X1 XNOR2X1_14 ( .A(sqrto_20_), .B(u2_remHi_20_), .Y(u2__abc_52138_new_n3182_));
XNOR2X1 XNOR2X1_15 ( .A(sqrto_19_), .B(u2_remHi_19_), .Y(u2__abc_52138_new_n3188_));
XNOR2X1 XNOR2X1_16 ( .A(sqrto_16_), .B(u2_remHi_16_), .Y(u2__abc_52138_new_n3197_));
XNOR2X1 XNOR2X1_17 ( .A(sqrto_34_), .B(u2_remHi_34_), .Y(u2__abc_52138_new_n3417_));
XNOR2X1 XNOR2X1_18 ( .A(sqrto_36_), .B(u2_remHi_36_), .Y(u2__abc_52138_new_n3428_));
XNOR2X1 XNOR2X1_19 ( .A(sqrto_32_), .B(u2_remHi_32_), .Y(u2__abc_52138_new_n3432_));
XNOR2X1 XNOR2X1_2 ( .A(_abc_65734_new_n1544_), .B(_abc_65734_new_n1550_), .Y(_abc_65734_new_n1551_));
XNOR2X1 XNOR2X1_20 ( .A(sqrto_68_), .B(u2_remHi_68_), .Y(u2__abc_52138_new_n3855_));
XNOR2X1 XNOR2X1_21 ( .A(sqrto_67_), .B(u2_remHi_67_), .Y(u2__abc_52138_new_n3861_));
XNOR2X1 XNOR2X1_22 ( .A(sqrto_64_), .B(u2_remHi_64_), .Y(u2__abc_52138_new_n3872_));
XNOR2X1 XNOR2X1_23 ( .A(sqrto_202_), .B(u2_remHi_202_), .Y(u2__abc_52138_new_n4328_));
XNOR2X1 XNOR2X1_24 ( .A(sqrto_128_), .B(u2_remHi_128_), .Y(u2__abc_52138_new_n4726_));
XNOR2X1 XNOR2X1_25 ( .A(sqrto_130_), .B(u2_remHi_130_), .Y(u2__abc_52138_new_n4749_));
XNOR2X1 XNOR2X1_26 ( .A(sqrto_132_), .B(u2_remHi_132_), .Y(u2__abc_52138_new_n4763_));
XNOR2X1 XNOR2X1_27 ( .A(u2_remHi_378_), .B(u2_o_378_), .Y(u2__abc_52138_new_n5010_));
XNOR2X1 XNOR2X1_28 ( .A(u2_remHi_369_), .B(u2_o_369_), .Y(u2__abc_52138_new_n5050_));
XNOR2X1 XNOR2X1_29 ( .A(u2_remHi_362_), .B(u2_o_362_), .Y(u2__abc_52138_new_n5125_));
XNOR2X1 XNOR2X1_3 ( .A(_abc_65734_new_n1549_), .B(_abc_65734_new_n1555_), .Y(_abc_65734_new_n1556_));
XNOR2X1 XNOR2X1_30 ( .A(u2_remHi_334_), .B(u2_o_334_), .Y(u2__abc_52138_new_n5241_));
XNOR2X1 XNOR2X1_31 ( .A(u2_remHi_322_), .B(u2_o_322_), .Y(u2__abc_52138_new_n5332_));
XNOR2X1 XNOR2X1_32 ( .A(u2_remHi_310_), .B(u2_o_310_), .Y(u2__abc_52138_new_n5379_));
XNOR2X1 XNOR2X1_33 ( .A(u2_remHi_314_), .B(u2_o_314_), .Y(u2__abc_52138_new_n5398_));
XNOR2X1 XNOR2X1_34 ( .A(u2_remHi_290_), .B(u2_o_290_), .Y(u2__abc_52138_new_n5536_));
XNOR2X1 XNOR2X1_35 ( .A(u2_remHi_274_), .B(u2_o_274_), .Y(u2__abc_52138_new_n5629_));
XNOR2X1 XNOR2X1_36 ( .A(u2_o_439_), .B(u2_remHi_439_), .Y(u2__abc_52138_new_n5972_));
XNOR2X1 XNOR2X1_37 ( .A(u2__abc_52138_new_n6542_), .B(u2__abc_52138_new_n6464_), .Y(u2__abc_52138_new_n6543_));
XNOR2X1 XNOR2X1_38 ( .A(u2__abc_52138_new_n6551_), .B(u2__abc_52138_new_n6463_), .Y(u2__abc_52138_new_n6552_));
XNOR2X1 XNOR2X1_39 ( .A(u2__abc_52138_new_n6560_), .B(u2__abc_52138_new_n3053_), .Y(u2__abc_52138_new_n6561_));
XNOR2X1 XNOR2X1_4 ( .A(_abc_65734_new_n1549_), .B(\a[124] ), .Y(_abc_65734_new_n1559_));
XNOR2X1 XNOR2X1_40 ( .A(u2__abc_52138_new_n6568_), .B(u2__abc_52138_new_n6461_), .Y(u2__abc_52138_new_n6569_));
XNOR2X1 XNOR2X1_41 ( .A(u2__abc_52138_new_n6582_), .B(u2__abc_52138_new_n3049_), .Y(u2__abc_52138_new_n6583_));
XNOR2X1 XNOR2X1_42 ( .A(u2__abc_52138_new_n6591_), .B(u2__abc_52138_new_n3044_), .Y(u2__abc_52138_new_n6592_));
XNOR2X1 XNOR2X1_43 ( .A(u2__abc_52138_new_n6616_), .B(u2__abc_52138_new_n6614_), .Y(u2__abc_52138_new_n6617_));
XNOR2X1 XNOR2X1_44 ( .A(u2__abc_52138_new_n6635_), .B(u2__abc_52138_new_n3026_), .Y(u2__abc_52138_new_n6636_));
XNOR2X1 XNOR2X1_45 ( .A(u2__abc_52138_new_n6645_), .B(u2__abc_52138_new_n3016_), .Y(u2__abc_52138_new_n6646_));
XNOR2X1 XNOR2X1_46 ( .A(u2__abc_52138_new_n6656_), .B(u2__abc_52138_new_n6653_), .Y(u2__abc_52138_new_n6657_));
XNOR2X1 XNOR2X1_47 ( .A(u2__abc_52138_new_n6702_), .B(u2__abc_52138_new_n3168_), .Y(u2__abc_52138_new_n6703_));
XNOR2X1 XNOR2X1_48 ( .A(u2__abc_52138_new_n6773_), .B(u2__abc_52138_new_n3127_), .Y(u2__abc_52138_new_n6774_));
XNOR2X1 XNOR2X1_49 ( .A(u2__abc_52138_new_n6793_), .B(u2__abc_52138_new_n3220_), .Y(u2__abc_52138_new_n6794_));
XNOR2X1 XNOR2X1_5 ( .A(_abc_65734_new_n1557_), .B(_abc_65734_new_n1567_), .Y(_abc_65734_new_n1568_));
XNOR2X1 XNOR2X1_50 ( .A(u2__abc_52138_new_n6833_), .B(u2__abc_52138_new_n3144_), .Y(u2__abc_52138_new_n6834_));
XNOR2X1 XNOR2X1_51 ( .A(u2__abc_52138_new_n6844_), .B(u2__abc_52138_new_n3393_), .Y(u2__abc_52138_new_n6845_));
XNOR2X1 XNOR2X1_52 ( .A(u2__abc_52138_new_n6896_), .B(u2__abc_52138_new_n6895_), .Y(u2__abc_52138_new_n6897_));
XNOR2X1 XNOR2X1_53 ( .A(u2__abc_52138_new_n6999_), .B(u2__abc_52138_new_n3367_), .Y(u2__abc_52138_new_n7000_));
XNOR2X1 XNOR2X1_54 ( .A(u2__abc_52138_new_n7204_), .B(u2__abc_52138_new_n3872_), .Y(u2__abc_52138_new_n7205_));
XNOR2X1 XNOR2X1_55 ( .A(u2__abc_52138_new_n7235_), .B(u2__abc_52138_new_n3861_), .Y(u2__abc_52138_new_n7236_));
XNOR2X1 XNOR2X1_56 ( .A(u2__abc_52138_new_n7290_), .B(u2__abc_52138_new_n3801_), .Y(u2__abc_52138_new_n7291_));
XNOR2X1 XNOR2X1_57 ( .A(u2__abc_52138_new_n7382_), .B(u2__abc_52138_new_n3753_), .Y(u2__abc_52138_new_n7383_));
XNOR2X1 XNOR2X1_58 ( .A(u2__abc_52138_new_n7523_), .B(u2__abc_52138_new_n3700_), .Y(u2__abc_52138_new_n7524_));
XNOR2X1 XNOR2X1_59 ( .A(u2__abc_52138_new_n7561_), .B(u2__abc_52138_new_n3646_), .Y(u2__abc_52138_new_n7562_));
XNOR2X1 XNOR2X1_6 ( .A(_abc_65734_new_n1566_), .B(\a[126] ), .Y(_abc_65734_new_n1572_));
XNOR2X1 XNOR2X1_60 ( .A(u2__abc_52138_new_n7571_), .B(u2__abc_52138_new_n7570_), .Y(u2__abc_52138_new_n7572_));
XNOR2X1 XNOR2X1_61 ( .A(u2__abc_52138_new_n7685_), .B(u2__abc_52138_new_n7684_), .Y(u2__abc_52138_new_n7686_));
XNOR2X1 XNOR2X1_62 ( .A(u2__abc_52138_new_n7872_), .B(u2__abc_52138_new_n3531_), .Y(u2__abc_52138_new_n7873_));
XNOR2X1 XNOR2X1_63 ( .A(u2__abc_52138_new_n7920_), .B(u2__abc_52138_new_n4726_), .Y(u2__abc_52138_new_n7921_));
XNOR2X1 XNOR2X1_64 ( .A(u2__abc_52138_new_n7954_), .B(u2__abc_52138_new_n4748_), .Y(u2__abc_52138_new_n7955_));
XNOR2X1 XNOR2X1_65 ( .A(u2__abc_52138_new_n8053_), .B(u2__abc_52138_new_n4693_), .Y(u2__abc_52138_new_n8054_));
XNOR2X1 XNOR2X1_66 ( .A(u2__abc_52138_new_n8093_), .B(u2__abc_52138_new_n8092_), .Y(u2__abc_52138_new_n8094_));
XNOR2X1 XNOR2X1_67 ( .A(u2__abc_52138_new_n8191_), .B(u2__abc_52138_new_n4577_), .Y(u2__abc_52138_new_n8192_));
XNOR2X1 XNOR2X1_68 ( .A(u2__abc_52138_new_n8221_), .B(u2__abc_52138_new_n4611_), .Y(u2__abc_52138_new_n8222_));
XNOR2X1 XNOR2X1_69 ( .A(u2__abc_52138_new_n8231_), .B(u2__abc_52138_new_n4600_), .Y(u2__abc_52138_new_n8232_));
XNOR2X1 XNOR2X1_7 ( .A(u2_o_449_), .B(u2_remHi_449_), .Y(u2__abc_52138_new_n3000_));
XNOR2X1 XNOR2X1_70 ( .A(u2__abc_52138_new_n8332_), .B(u2__abc_52138_new_n4557_), .Y(u2__abc_52138_new_n8333_));
XNOR2X1 XNOR2X1_71 ( .A(u2__abc_52138_new_n8402_), .B(u2__abc_52138_new_n4482_), .Y(u2__abc_52138_new_n8403_));
XNOR2X1 XNOR2X1_72 ( .A(u2__abc_52138_new_n8493_), .B(u2__abc_52138_new_n4433_), .Y(u2__abc_52138_new_n8494_));
XNOR2X1 XNOR2X1_73 ( .A(u2__abc_52138_new_n8515_), .B(u2__abc_52138_new_n4386_), .Y(u2__abc_52138_new_n8516_));
XNOR2X1 XNOR2X1_74 ( .A(u2__abc_52138_new_n8574_), .B(u2__abc_52138_new_n4409_), .Y(u2__abc_52138_new_n8575_));
XNOR2X1 XNOR2X1_75 ( .A(u2__abc_52138_new_n8711_), .B(u2__abc_52138_new_n4293_), .Y(u2__abc_52138_new_n8712_));
XNOR2X1 XNOR2X1_76 ( .A(u2__abc_52138_new_n8741_), .B(u2__abc_52138_new_n4327_), .Y(u2__abc_52138_new_n8742_));
XNOR2X1 XNOR2X1_77 ( .A(u2__abc_52138_new_n8751_), .B(u2__abc_52138_new_n4316_), .Y(u2__abc_52138_new_n8752_));
XNOR2X1 XNOR2X1_78 ( .A(u2__abc_52138_new_n8858_), .B(u2__abc_52138_new_n4209_), .Y(u2__abc_52138_new_n8859_));
XNOR2X1 XNOR2X1_79 ( .A(u2__abc_52138_new_n8908_), .B(u2__abc_52138_new_n4232_), .Y(u2__abc_52138_new_n8909_));
XNOR2X1 XNOR2X1_8 ( .A(sqrto_12_), .B(u2_remHi_12_), .Y(u2__abc_52138_new_n3016_));
XNOR2X1 XNOR2X1_80 ( .A(u2__abc_52138_new_n8927_), .B(u2__abc_52138_new_n4226_), .Y(u2__abc_52138_new_n8928_));
XNOR2X1 XNOR2X1_81 ( .A(u2__abc_52138_new_n8964_), .B(u2__abc_52138_new_n4150_), .Y(u2__abc_52138_new_n8965_));
XNOR2X1 XNOR2X1_82 ( .A(u2__abc_52138_new_n8993_), .B(u2__abc_52138_new_n4184_), .Y(u2__abc_52138_new_n8994_));
XNOR2X1 XNOR2X1_83 ( .A(u2__abc_52138_new_n9003_), .B(u2__abc_52138_new_n4173_), .Y(u2__abc_52138_new_n9004_));
XNOR2X1 XNOR2X1_84 ( .A(u2__abc_52138_new_n9081_), .B(u2__abc_52138_new_n4103_), .Y(u2__abc_52138_new_n9082_));
XNOR2X1 XNOR2X1_85 ( .A(u2__abc_52138_new_n9147_), .B(u2__abc_52138_new_n9143_), .Y(u2__abc_52138_new_n9148_));
XNOR2X1 XNOR2X1_86 ( .A(u2__abc_52138_new_n9174_), .B(u2__abc_52138_new_n4083_), .Y(u2__abc_52138_new_n9175_));
XNOR2X1 XNOR2X1_87 ( .A(u2__abc_52138_new_n9331_), .B(u2__abc_52138_new_n5729_), .Y(u2__abc_52138_new_n9332_));
XNOR2X1 XNOR2X1_88 ( .A(u2__abc_52138_new_n9457_), .B(u2__abc_52138_new_n5615_), .Y(u2__abc_52138_new_n9458_));
XNOR2X1 XNOR2X1_89 ( .A(u2__abc_52138_new_n9500_), .B(u2__abc_52138_new_n5634_), .Y(u2__abc_52138_new_n9501_));
XNOR2X1 XNOR2X1_9 ( .A(sqrto_8_), .B(u2_remHi_8_), .Y(u2__abc_52138_new_n3034_));
XNOR2X1 XNOR2X1_90 ( .A(u2__abc_52138_new_n9542_), .B(u2__abc_52138_new_n5568_), .Y(u2__abc_52138_new_n9543_));
XNOR2X1 XNOR2X1_91 ( .A(u2__abc_52138_new_n9585_), .B(u2__abc_52138_new_n5591_), .Y(u2__abc_52138_new_n9586_));
XNOR2X1 XNOR2X1_92 ( .A(u2__abc_52138_new_n9632_), .B(u2__abc_52138_new_n5522_), .Y(u2__abc_52138_new_n9633_));
XNOR2X1 XNOR2X1_93 ( .A(u2__abc_52138_new_n9676_), .B(u2__abc_52138_new_n5541_), .Y(u2__abc_52138_new_n9677_));
XNOR2X1 XNOR2X1_94 ( .A(u2__abc_52138_new_n9758_), .B(u2__abc_52138_new_n5498_), .Y(u2__abc_52138_new_n9759_));
XNOR2X1 XNOR2X1_95 ( .A(u2__abc_52138_new_n9886_), .B(u2__abc_52138_new_n5384_), .Y(u2__abc_52138_new_n9887_));
XNOR2X1 XNOR2X1_96 ( .A(u2__abc_52138_new_n9929_), .B(u2__abc_52138_new_n5403_), .Y(u2__abc_52138_new_n9930_));
XNOR2X1 XNOR2X1_97 ( .A(u2__abc_52138_new_n10019_), .B(u2__abc_52138_new_n5337_), .Y(u2__abc_52138_new_n10020_));
XNOR2X1 XNOR2X1_98 ( .A(u2__abc_52138_new_n10103_), .B(u2__abc_52138_new_n5317_), .Y(u2__abc_52138_new_n10104_));
XNOR2X1 XNOR2X1_99 ( .A(u2__abc_52138_new_n10147_), .B(u2__abc_52138_new_n5247_), .Y(u2__abc_52138_new_n10148_));
XOR2X1 XOR2X1_1 ( .A(_abc_65734_new_n1566_), .B(\a[126] ), .Y(_abc_65734_new_n1575_));
XOR2X1 XOR2X1_10 ( .A(u2__abc_52138_new_n6915_), .B(u2__abc_52138_new_n3410_), .Y(u2__abc_52138_new_n6916_));
XOR2X1 XOR2X1_11 ( .A(u2__abc_52138_new_n6939_), .B(u2__abc_52138_new_n3355_), .Y(u2__abc_52138_new_n6940_));
XOR2X1 XOR2X1_12 ( .A(u2__abc_52138_new_n6948_), .B(u2__abc_52138_new_n3339_), .Y(u2__abc_52138_new_n6949_));
XOR2X1 XOR2X1_13 ( .A(u2__abc_52138_new_n6980_), .B(u2__abc_52138_new_n3373_), .Y(u2__abc_52138_new_n6981_));
XOR2X1 XOR2X1_14 ( .A(u2__abc_52138_new_n6990_), .B(u2__abc_52138_new_n3362_), .Y(u2__abc_52138_new_n6991_));
XOR2X1 XOR2X1_15 ( .A(u2__abc_52138_new_n7022_), .B(u2__abc_52138_new_n3302_), .Y(u2__abc_52138_new_n7023_));
XOR2X1 XOR2X1_16 ( .A(u2__abc_52138_new_n7065_), .B(u2__abc_52138_new_n3326_), .Y(u2__abc_52138_new_n7066_));
XOR2X1 XOR2X1_17 ( .A(u2__abc_52138_new_n7076_), .B(u2__abc_52138_new_n3315_), .Y(u2__abc_52138_new_n7077_));
XOR2X1 XOR2X1_18 ( .A(u2__abc_52138_new_n7085_), .B(u2__abc_52138_new_n3320_), .Y(u2__abc_52138_new_n7086_));
XOR2X1 XOR2X1_19 ( .A(u2__abc_52138_new_n7110_), .B(u2__abc_52138_new_n3260_), .Y(u2__abc_52138_new_n7111_));
XOR2X1 XOR2X1_2 ( .A(sqrto_32_), .B(u2_remHi_32_), .Y(u2__abc_52138_new_n3382_));
XOR2X1 XOR2X1_20 ( .A(u2__abc_52138_new_n7118_), .B(u2__abc_52138_new_n3244_), .Y(u2__abc_52138_new_n7119_));
XOR2X1 XOR2X1_21 ( .A(u2__abc_52138_new_n7127_), .B(u2__abc_52138_new_n3249_), .Y(u2__abc_52138_new_n7128_));
XOR2X1 XOR2X1_22 ( .A(u2__abc_52138_new_n7169_), .B(u2__abc_52138_new_n3272_), .Y(u2__abc_52138_new_n7170_));
XOR2X1 XOR2X1_23 ( .A(u2__abc_52138_new_n7227_), .B(u2__abc_52138_new_n7222_), .Y(u2__abc_52138_new_n7228_));
XOR2X1 XOR2X1_24 ( .A(u2__abc_52138_new_n7254_), .B(u2__abc_52138_new_n7252_), .Y(u2__abc_52138_new_n7255_));
XOR2X1 XOR2X1_25 ( .A(u2__abc_52138_new_n7300_), .B(u2__abc_52138_new_n7298_), .Y(u2__abc_52138_new_n7301_));
XOR2X1 XOR2X1_26 ( .A(u2__abc_52138_new_n7363_), .B(u2__abc_52138_new_n3742_), .Y(u2__abc_52138_new_n7364_));
XOR2X1 XOR2X1_27 ( .A(u2__abc_52138_new_n7417_), .B(u2__abc_52138_new_n3776_), .Y(u2__abc_52138_new_n7418_));
XOR2X1 XOR2X1_28 ( .A(u2__abc_52138_new_n7483_), .B(u2__abc_52138_new_n3722_), .Y(u2__abc_52138_new_n7484_));
XOR2X1 XOR2X1_29 ( .A(u2__abc_52138_new_n7504_), .B(u2__abc_52138_new_n7503_), .Y(u2__abc_52138_new_n7505_));
XOR2X1 XOR2X1_3 ( .A(sqrto_8_), .B(u2_remHi_8_), .Y(u2__abc_52138_new_n6599_));
XOR2X1 XOR2X1_30 ( .A(u2__abc_52138_new_n7514_), .B(u2__abc_52138_new_n3695_), .Y(u2__abc_52138_new_n7515_));
XOR2X1 XOR2X1_31 ( .A(u2__abc_52138_new_n7551_), .B(u2__abc_52138_new_n3657_), .Y(u2__abc_52138_new_n7552_));
XOR2X1 XOR2X1_32 ( .A(u2__abc_52138_new_n7597_), .B(u2__abc_52138_new_n3680_), .Y(u2__abc_52138_new_n7598_));
XOR2X1 XOR2X1_33 ( .A(u2__abc_52138_new_n7643_), .B(u2__abc_52138_new_n7642_), .Y(u2__abc_52138_new_n7644_));
XOR2X1 XOR2X1_34 ( .A(u2__abc_52138_new_n7662_), .B(u2__abc_52138_new_n3606_), .Y(u2__abc_52138_new_n7663_));
XOR2X1 XOR2X1_35 ( .A(u2__abc_52138_new_n7695_), .B(u2__abc_52138_new_n3623_), .Y(u2__abc_52138_new_n7696_));
XOR2X1 XOR2X1_36 ( .A(u2__abc_52138_new_n7721_), .B(u2__abc_52138_new_n3554_), .Y(u2__abc_52138_new_n7722_));
XOR2X1 XOR2X1_37 ( .A(u2__abc_52138_new_n7730_), .B(u2__abc_52138_new_n3559_), .Y(u2__abc_52138_new_n7731_));
XOR2X1 XOR2X1_38 ( .A(u2__abc_52138_new_n7749_), .B(u2__abc_52138_new_n3570_), .Y(u2__abc_52138_new_n7750_));
XOR2X1 XOR2X1_39 ( .A(u2__abc_52138_new_n7793_), .B(u2__abc_52138_new_n7792_), .Y(u2__abc_52138_new_n7794_));
XOR2X1 XOR2X1_4 ( .A(u2__abc_52138_new_n6683_), .B(u2__abc_52138_new_n3179_), .Y(u2__abc_52138_new_n6684_));
XOR2X1 XOR2X1_40 ( .A(u2__abc_52138_new_n7841_), .B(u2__abc_52138_new_n3525_), .Y(u2__abc_52138_new_n7842_));
XOR2X1 XOR2X1_41 ( .A(u2__abc_52138_new_n7863_), .B(u2__abc_52138_new_n7862_), .Y(u2__abc_52138_new_n7864_));
XOR2X1 XOR2X1_42 ( .A(u2__abc_52138_new_n7880_), .B(u2__abc_52138_new_n3536_), .Y(u2__abc_52138_new_n7881_));
XOR2X1 XOR2X1_43 ( .A(u2__abc_52138_new_n7930_), .B(u2__abc_52138_new_n7928_), .Y(u2__abc_52138_new_n7931_));
XOR2X1 XOR2X1_44 ( .A(sqrto_128_), .B(u2_remHi_128_), .Y(u2__abc_52138_new_n7938_));
XOR2X1 XOR2X1_45 ( .A(u2__abc_52138_new_n7973_), .B(u2__abc_52138_new_n4742_), .Y(u2__abc_52138_new_n7974_));
XOR2X1 XOR2X1_46 ( .A(u2__abc_52138_new_n7999_), .B(u2__abc_52138_new_n4686_), .Y(u2__abc_52138_new_n8000_));
XOR2X1 XOR2X1_47 ( .A(u2__abc_52138_new_n8044_), .B(u2__abc_52138_new_n4704_), .Y(u2__abc_52138_new_n8045_));
XOR2X1 XOR2X1_48 ( .A(u2__abc_52138_new_n8061_), .B(u2__abc_52138_new_n4698_), .Y(u2__abc_52138_new_n8062_));
XOR2X1 XOR2X1_49 ( .A(u2__abc_52138_new_n8113_), .B(u2__abc_52138_new_n8112_), .Y(u2__abc_52138_new_n8114_));
XOR2X1 XOR2X1_5 ( .A(u2__abc_52138_new_n6725_), .B(u2__abc_52138_new_n3188_), .Y(u2__abc_52138_new_n6726_));
XOR2X1 XOR2X1_50 ( .A(u2__abc_52138_new_n8154_), .B(u2__abc_52138_new_n4628_), .Y(u2__abc_52138_new_n8155_));
XOR2X1 XOR2X1_51 ( .A(u2__abc_52138_new_n8181_), .B(u2__abc_52138_new_n4588_), .Y(u2__abc_52138_new_n8182_));
XOR2X1 XOR2X1_52 ( .A(u2__abc_52138_new_n8199_), .B(u2__abc_52138_new_n4582_), .Y(u2__abc_52138_new_n8200_));
XOR2X1 XOR2X1_53 ( .A(u2__abc_52138_new_n8239_), .B(u2__abc_52138_new_n4605_), .Y(u2__abc_52138_new_n8240_));
XOR2X1 XOR2X1_54 ( .A(u2__abc_52138_new_n8268_), .B(u2__abc_52138_new_n4540_), .Y(u2__abc_52138_new_n8269_));
XOR2X1 XOR2X1_55 ( .A(u2__abc_52138_new_n8323_), .B(u2__abc_52138_new_n4552_), .Y(u2__abc_52138_new_n8324_));
XOR2X1 XOR2X1_56 ( .A(u2__abc_52138_new_n8355_), .B(u2__abc_52138_new_n4516_), .Y(u2__abc_52138_new_n8356_));
XOR2X1 XOR2X1_57 ( .A(u2__abc_52138_new_n8374_), .B(u2__abc_52138_new_n4510_), .Y(u2__abc_52138_new_n8375_));
XOR2X1 XOR2X1_58 ( .A(u2__abc_52138_new_n8393_), .B(u2__abc_52138_new_n4493_), .Y(u2__abc_52138_new_n8394_));
XOR2X1 XOR2X1_59 ( .A(u2__abc_52138_new_n8410_), .B(u2__abc_52138_new_n4487_), .Y(u2__abc_52138_new_n8411_));
XOR2X1 XOR2X1_6 ( .A(u2__abc_52138_new_n6748_), .B(u2__abc_52138_new_n6747_), .Y(u2__abc_52138_new_n6749_));
XOR2X1 XOR2X1_60 ( .A(u2__abc_52138_new_n8463_), .B(u2__abc_52138_new_n4461_), .Y(u2__abc_52138_new_n8464_));
XOR2X1 XOR2X1_61 ( .A(u2__abc_52138_new_n8484_), .B(u2__abc_52138_new_n4444_), .Y(u2__abc_52138_new_n8485_));
XOR2X1 XOR2X1_62 ( .A(u2__abc_52138_new_n8501_), .B(u2__abc_52138_new_n4438_), .Y(u2__abc_52138_new_n8502_));
XOR2X1 XOR2X1_63 ( .A(u2__abc_52138_new_n8524_), .B(u2__abc_52138_new_n4391_), .Y(u2__abc_52138_new_n8525_));
XOR2X1 XOR2X1_64 ( .A(u2__abc_52138_new_n8535_), .B(u2__abc_52138_new_n4397_), .Y(u2__abc_52138_new_n8536_));
XOR2X1 XOR2X1_65 ( .A(u2__abc_52138_new_n8544_), .B(u2__abc_52138_new_n4402_), .Y(u2__abc_52138_new_n8545_));
XOR2X1 XOR2X1_66 ( .A(u2__abc_52138_new_n8565_), .B(u2__abc_52138_new_n4420_), .Y(u2__abc_52138_new_n8566_));
XOR2X1 XOR2X1_67 ( .A(u2__abc_52138_new_n8582_), .B(u2__abc_52138_new_n4414_), .Y(u2__abc_52138_new_n8583_));
XOR2X1 XOR2X1_68 ( .A(u2__abc_52138_new_n8615_), .B(u2__abc_52138_new_n4375_), .Y(u2__abc_52138_new_n8616_));
XOR2X1 XOR2X1_69 ( .A(u2__abc_52138_new_n8677_), .B(u2__abc_52138_new_n4340_), .Y(u2__abc_52138_new_n8678_));
XOR2X1 XOR2X1_7 ( .A(u2__abc_52138_new_n6816_), .B(u2__abc_52138_new_n3150_), .Y(u2__abc_52138_new_n6817_));
XOR2X1 XOR2X1_70 ( .A(u2__abc_52138_new_n8701_), .B(u2__abc_52138_new_n4304_), .Y(u2__abc_52138_new_n8702_));
XOR2X1 XOR2X1_71 ( .A(u2__abc_52138_new_n8719_), .B(u2__abc_52138_new_n4298_), .Y(u2__abc_52138_new_n8720_));
XOR2X1 XOR2X1_72 ( .A(u2__abc_52138_new_n8759_), .B(u2__abc_52138_new_n4321_), .Y(u2__abc_52138_new_n8760_));
XOR2X1 XOR2X1_73 ( .A(u2__abc_52138_new_n8785_), .B(u2__abc_52138_new_n4261_), .Y(u2__abc_52138_new_n8786_));
XOR2X1 XOR2X1_74 ( .A(u2__abc_52138_new_n8794_), .B(u2__abc_52138_new_n4245_), .Y(u2__abc_52138_new_n8795_));
XOR2X1 XOR2X1_75 ( .A(u2__abc_52138_new_n8803_), .B(u2__abc_52138_new_n4250_), .Y(u2__abc_52138_new_n8804_));
XOR2X1 XOR2X1_76 ( .A(u2__abc_52138_new_n8843_), .B(u2__abc_52138_new_n4273_), .Y(u2__abc_52138_new_n8844_));
XOR2X1 XOR2X1_77 ( .A(u2__abc_52138_new_n8867_), .B(u2__abc_52138_new_n4214_), .Y(u2__abc_52138_new_n8868_));
XOR2X1 XOR2X1_78 ( .A(u2__abc_52138_new_n8877_), .B(u2__abc_52138_new_n4198_), .Y(u2__abc_52138_new_n8878_));
XOR2X1 XOR2X1_79 ( .A(u2__abc_52138_new_n8886_), .B(u2__abc_52138_new_n4203_), .Y(u2__abc_52138_new_n8887_));
XOR2X1 XOR2X1_8 ( .A(u2__abc_52138_new_n6825_), .B(u2__abc_52138_new_n3139_), .Y(u2__abc_52138_new_n6826_));
XOR2X1 XOR2X1_80 ( .A(u2__abc_52138_new_n8918_), .B(u2__abc_52138_new_n4221_), .Y(u2__abc_52138_new_n8919_));
XOR2X1 XOR2X1_81 ( .A(u2__abc_52138_new_n8955_), .B(u2__abc_52138_new_n4161_), .Y(u2__abc_52138_new_n8956_));
XOR2X1 XOR2X1_82 ( .A(u2__abc_52138_new_n8972_), .B(u2__abc_52138_new_n4155_), .Y(u2__abc_52138_new_n8973_));
XOR2X1 XOR2X1_83 ( .A(u2__abc_52138_new_n9011_), .B(u2__abc_52138_new_n4178_), .Y(u2__abc_52138_new_n9012_));
XOR2X1 XOR2X1_84 ( .A(u2__abc_52138_new_n9035_), .B(u2__abc_52138_new_n9034_), .Y(u2__abc_52138_new_n9036_));
XOR2X1 XOR2X1_85 ( .A(u2__abc_52138_new_n9053_), .B(u2__abc_52138_new_n4132_), .Y(u2__abc_52138_new_n9054_));
XOR2X1 XOR2X1_86 ( .A(u2__abc_52138_new_n9072_), .B(u2__abc_52138_new_n4114_), .Y(u2__abc_52138_new_n9073_));
XOR2X1 XOR2X1_87 ( .A(u2__abc_52138_new_n9089_), .B(u2__abc_52138_new_n4108_), .Y(u2__abc_52138_new_n9090_));
XOR2X1 XOR2X1_88 ( .A(u2__abc_52138_new_n9107_), .B(u2__abc_52138_new_n4054_), .Y(u2__abc_52138_new_n9108_));
XOR2X1 XOR2X1_89 ( .A(u2__abc_52138_new_n9116_), .B(u2__abc_52138_new_n4059_), .Y(u2__abc_52138_new_n9117_));
XOR2X1 XOR2X1_9 ( .A(u2__abc_52138_new_n6854_), .B(u2__abc_52138_new_n3398_), .Y(u2__abc_52138_new_n6855_));
XOR2X1 XOR2X1_90 ( .A(u2__abc_52138_new_n9126_), .B(u2__abc_52138_new_n4065_), .Y(u2__abc_52138_new_n9127_));
XOR2X1 XOR2X1_91 ( .A(u2__abc_52138_new_n9135_), .B(u2__abc_52138_new_n4070_), .Y(u2__abc_52138_new_n9136_));
XOR2X1 XOR2X1_92 ( .A(u2__abc_52138_new_n9197_), .B(u2__abc_52138_new_n4012_), .Y(u2__abc_52138_new_n9198_));
XOR2X1 XOR2X1_93 ( .A(u2__abc_52138_new_n9218_), .B(u2__abc_52138_new_n4023_), .Y(u2__abc_52138_new_n9219_));
XOR2X1 XOR2X1_94 ( .A(u2__abc_52138_new_n9239_), .B(u2__abc_52138_new_n4041_), .Y(u2__abc_52138_new_n9240_));
XOR2X1 XOR2X1_95 ( .A(u2__abc_52138_new_n9248_), .B(u2__abc_52138_new_n4030_), .Y(u2__abc_52138_new_n9249_));
XOR2X1 XOR2X1_96 ( .A(u2__abc_52138_new_n9256_), .B(u2__abc_52138_new_n4035_), .Y(u2__abc_52138_new_n9257_));
XOR2X1 XOR2X1_97 ( .A(u2__abc_52138_new_n9410_), .B(u2__abc_52138_new_n5660_), .Y(u2__abc_52138_new_n9411_));

assign \o[0]  = 1'h0;
assign \o[1]  = 1'h0;
assign \o[2]  = 1'h0;
assign \o[3]  = 1'h0;
assign \o[4]  = 1'h0;
assign \o[5]  = 1'h0;
assign \o[6]  = 1'h0;
assign \o[7]  = 1'h0;
assign \o[8]  = 1'h0;
assign \o[9]  = 1'h0;
assign \o[10]  = 1'h0;
assign \o[11]  = 1'h0;
assign \o[12]  = 1'h0;
assign \o[13]  = 1'h0;
assign \o[14]  = 1'h0;
assign \o[15]  = 1'h0;
assign \o[16]  = 1'h0;
assign \o[17]  = 1'h0;
assign \o[18]  = 1'h0;
assign \o[19]  = 1'h0;
assign \o[20]  = 1'h0;
assign \o[21]  = 1'h0;
assign \o[22]  = 1'h0;
assign \o[23]  = 1'h0;
assign \o[24]  = 1'h0;
assign \o[25]  = 1'h0;
assign \o[26]  = 1'h0;
assign \o[27]  = 1'h0;
assign \o[28]  = 1'h0;
assign \o[29]  = 1'h0;
assign \o[30]  = 1'h0;
assign \o[31]  = 1'h0;
assign \o[32]  = 1'h0;
assign \o[33]  = 1'h0;
assign \o[34]  = 1'h0;
assign \o[35]  = 1'h0;

endmodule