module cpu8080(\data[0] , \data[1] , \data[2] , \data[3] , \data[4] , \data[5] , \data[6] , \data[7] , intr, waitr, reset, clock, \addr[0] , \addr[1] , \addr[2] , \addr[3] , \addr[4] , \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , \addr[10] , \addr[11] , \addr[12] , \addr[13] , \addr[14] , \addr[15] , readmem, writemem, readio, writeio, inta);

wire _0addr_15_0__0_; 
wire _0addr_15_0__10_; 
wire _0addr_15_0__11_; 
wire _0addr_15_0__12_; 
wire _0addr_15_0__13_; 
wire _0addr_15_0__14_; 
wire _0addr_15_0__15_; 
wire _0addr_15_0__1_; 
wire _0addr_15_0__2_; 
wire _0addr_15_0__3_; 
wire _0addr_15_0__4_; 
wire _0addr_15_0__5_; 
wire _0addr_15_0__6_; 
wire _0addr_15_0__7_; 
wire _0addr_15_0__8_; 
wire _0addr_15_0__9_; 
wire _0alucin_0_0_; 
wire _0aluopra_7_0__0_; 
wire _0aluopra_7_0__1_; 
wire _0aluopra_7_0__2_; 
wire _0aluopra_7_0__3_; 
wire _0aluopra_7_0__4_; 
wire _0aluopra_7_0__5_; 
wire _0aluopra_7_0__6_; 
wire _0aluopra_7_0__7_; 
wire _0aluoprb_7_0__0_; 
wire _0aluoprb_7_0__1_; 
wire _0aluoprb_7_0__2_; 
wire _0aluoprb_7_0__3_; 
wire _0aluoprb_7_0__4_; 
wire _0aluoprb_7_0__5_; 
wire _0aluoprb_7_0__6_; 
wire _0aluoprb_7_0__7_; 
wire _0alusel_2_0__0_; 
wire _0alusel_2_0__1_; 
wire _0alusel_2_0__2_; 
wire _0auxcar_0_0_; 
wire _0carry_0_0_; 
wire _0datao_7_0__0_; 
wire _0datao_7_0__1_; 
wire _0datao_7_0__2_; 
wire _0datao_7_0__3_; 
wire _0datao_7_0__4_; 
wire _0datao_7_0__5_; 
wire _0datao_7_0__6_; 
wire _0datao_7_0__7_; 
wire _0ei_0_0_; 
wire _0eienb_0_0_; 
wire _0inta_0_0_; 
wire _0intcyc_0_0_; 
wire _0opcode_7_0__0_; 
wire _0opcode_7_0__1_; 
wire _0opcode_7_0__2_; 
wire _0opcode_7_0__3_; 
wire _0opcode_7_0__4_; 
wire _0opcode_7_0__5_; 
wire _0opcode_7_0__6_; 
wire _0opcode_7_0__7_; 
wire _0parity_0_0_; 
wire _0pc_15_0__0_; 
wire _0pc_15_0__10_; 
wire _0pc_15_0__11_; 
wire _0pc_15_0__12_; 
wire _0pc_15_0__13_; 
wire _0pc_15_0__14_; 
wire _0pc_15_0__15_; 
wire _0pc_15_0__1_; 
wire _0pc_15_0__2_; 
wire _0pc_15_0__3_; 
wire _0pc_15_0__4_; 
wire _0pc_15_0__5_; 
wire _0pc_15_0__6_; 
wire _0pc_15_0__7_; 
wire _0pc_15_0__8_; 
wire _0pc_15_0__9_; 
wire _0popdes_1_0__0_; 
wire _0popdes_1_0__1_; 
wire _0raddrhold_15_0__0_; 
wire _0raddrhold_15_0__10_; 
wire _0raddrhold_15_0__11_; 
wire _0raddrhold_15_0__12_; 
wire _0raddrhold_15_0__13_; 
wire _0raddrhold_15_0__14_; 
wire _0raddrhold_15_0__15_; 
wire _0raddrhold_15_0__1_; 
wire _0raddrhold_15_0__2_; 
wire _0raddrhold_15_0__3_; 
wire _0raddrhold_15_0__4_; 
wire _0raddrhold_15_0__5_; 
wire _0raddrhold_15_0__6_; 
wire _0raddrhold_15_0__7_; 
wire _0raddrhold_15_0__8_; 
wire _0raddrhold_15_0__9_; 
wire _0rdatahold2_7_0__0_; 
wire _0rdatahold2_7_0__1_; 
wire _0rdatahold2_7_0__2_; 
wire _0rdatahold2_7_0__3_; 
wire _0rdatahold2_7_0__4_; 
wire _0rdatahold2_7_0__5_; 
wire _0rdatahold2_7_0__6_; 
wire _0rdatahold2_7_0__7_; 
wire _0rdatahold_7_0__0_; 
wire _0rdatahold_7_0__1_; 
wire _0rdatahold_7_0__2_; 
wire _0rdatahold_7_0__3_; 
wire _0rdatahold_7_0__4_; 
wire _0rdatahold_7_0__5_; 
wire _0rdatahold_7_0__6_; 
wire _0rdatahold_7_0__7_; 
wire _0readio_0_0_; 
wire _0readmem_0_0_; 
wire _0regd_2_0__0_; 
wire _0regd_2_0__1_; 
wire _0regd_2_0__2_; 
wire _0sign_0_0_; 
wire _0sp_15_0__0_; 
wire _0sp_15_0__10_; 
wire _0sp_15_0__11_; 
wire _0sp_15_0__12_; 
wire _0sp_15_0__13_; 
wire _0sp_15_0__14_; 
wire _0sp_15_0__15_; 
wire _0sp_15_0__1_; 
wire _0sp_15_0__2_; 
wire _0sp_15_0__3_; 
wire _0sp_15_0__4_; 
wire _0sp_15_0__5_; 
wire _0sp_15_0__6_; 
wire _0sp_15_0__7_; 
wire _0sp_15_0__8_; 
wire _0sp_15_0__9_; 
wire _0statesel_5_0__0_; 
wire _0statesel_5_0__1_; 
wire _0statesel_5_0__2_; 
wire _0statesel_5_0__3_; 
wire _0statesel_5_0__4_; 
wire _0statesel_5_0__5_; 
wire _0waddrhold_15_0__0_; 
wire _0waddrhold_15_0__10_; 
wire _0waddrhold_15_0__11_; 
wire _0waddrhold_15_0__12_; 
wire _0waddrhold_15_0__13_; 
wire _0waddrhold_15_0__14_; 
wire _0waddrhold_15_0__15_; 
wire _0waddrhold_15_0__1_; 
wire _0waddrhold_15_0__2_; 
wire _0waddrhold_15_0__3_; 
wire _0waddrhold_15_0__4_; 
wire _0waddrhold_15_0__5_; 
wire _0waddrhold_15_0__6_; 
wire _0waddrhold_15_0__7_; 
wire _0waddrhold_15_0__8_; 
wire _0waddrhold_15_0__9_; 
wire _0wdatahold2_7_0__0_; 
wire _0wdatahold2_7_0__1_; 
wire _0wdatahold2_7_0__2_; 
wire _0wdatahold2_7_0__3_; 
wire _0wdatahold2_7_0__4_; 
wire _0wdatahold2_7_0__5_; 
wire _0wdatahold2_7_0__6_; 
wire _0wdatahold2_7_0__7_; 
wire _0wdatahold_7_0__0_; 
wire _0wdatahold_7_0__1_; 
wire _0wdatahold_7_0__2_; 
wire _0wdatahold_7_0__3_; 
wire _0wdatahold_7_0__4_; 
wire _0wdatahold_7_0__5_; 
wire _0wdatahold_7_0__6_; 
wire _0wdatahold_7_0__7_; 
wire _0writeio_0_0_; 
wire _0writemem_0_0_; 
wire _0zero_0_0_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_0_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_1_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_2_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_3_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_4_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_5_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_0_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_1_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_2_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_3_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_4_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_5_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_6_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_7_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_0_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_1_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_2_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_3_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_4_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_5_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_6_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_7_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_0_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_1_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_2_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_3_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_4_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_5_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_6_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_7_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_0_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_1_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_2_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_3_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_4_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_5_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_6_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_7_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_0_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_1_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_2_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_3_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_4_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_5_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_6_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_7_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_0_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_1_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_2_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_3_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_4_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_5_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_6_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_7_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_0_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_1_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_2_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_3_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_4_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_5_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_6_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_7_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_0_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_1_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_2_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_3_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_4_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_5_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_6_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_7_; 
wire _abc_41234_new_n1000_; 
wire _abc_41234_new_n1001_; 
wire _abc_41234_new_n1002_; 
wire _abc_41234_new_n1003_; 
wire _abc_41234_new_n1004_; 
wire _abc_41234_new_n1005_; 
wire _abc_41234_new_n1006_; 
wire _abc_41234_new_n1007_; 
wire _abc_41234_new_n1008_; 
wire _abc_41234_new_n1009_; 
wire _abc_41234_new_n1010_; 
wire _abc_41234_new_n1011_; 
wire _abc_41234_new_n1012_; 
wire _abc_41234_new_n1013_; 
wire _abc_41234_new_n1014_; 
wire _abc_41234_new_n1015_; 
wire _abc_41234_new_n1016_; 
wire _abc_41234_new_n1017_; 
wire _abc_41234_new_n1018_; 
wire _abc_41234_new_n1019_; 
wire _abc_41234_new_n1020_; 
wire _abc_41234_new_n1021_; 
wire _abc_41234_new_n1022_; 
wire _abc_41234_new_n1023_; 
wire _abc_41234_new_n1024_; 
wire _abc_41234_new_n1025_; 
wire _abc_41234_new_n1026_; 
wire _abc_41234_new_n1027_; 
wire _abc_41234_new_n1028_; 
wire _abc_41234_new_n1029_; 
wire _abc_41234_new_n1031_; 
wire _abc_41234_new_n1032_; 
wire _abc_41234_new_n1033_; 
wire _abc_41234_new_n1034_; 
wire _abc_41234_new_n1035_; 
wire _abc_41234_new_n1036_; 
wire _abc_41234_new_n1037_; 
wire _abc_41234_new_n1038_; 
wire _abc_41234_new_n1039_; 
wire _abc_41234_new_n1040_; 
wire _abc_41234_new_n1040__bF_buf0; 
wire _abc_41234_new_n1040__bF_buf1; 
wire _abc_41234_new_n1040__bF_buf2; 
wire _abc_41234_new_n1040__bF_buf3; 
wire _abc_41234_new_n1040__bF_buf4; 
wire _abc_41234_new_n1041_; 
wire _abc_41234_new_n1042_; 
wire _abc_41234_new_n1043_; 
wire _abc_41234_new_n1044_; 
wire _abc_41234_new_n1045_; 
wire _abc_41234_new_n1046_; 
wire _abc_41234_new_n1046__bF_buf0; 
wire _abc_41234_new_n1046__bF_buf1; 
wire _abc_41234_new_n1046__bF_buf2; 
wire _abc_41234_new_n1046__bF_buf3; 
wire _abc_41234_new_n1046__bF_buf4; 
wire _abc_41234_new_n1046__bF_buf5; 
wire _abc_41234_new_n1046__bF_buf6; 
wire _abc_41234_new_n1046__bF_buf7; 
wire _abc_41234_new_n1047_; 
wire _abc_41234_new_n1047__bF_buf0; 
wire _abc_41234_new_n1047__bF_buf1; 
wire _abc_41234_new_n1047__bF_buf2; 
wire _abc_41234_new_n1047__bF_buf3; 
wire _abc_41234_new_n1047__bF_buf4; 
wire _abc_41234_new_n1048_; 
wire _abc_41234_new_n1049_; 
wire _abc_41234_new_n1049__bF_buf0; 
wire _abc_41234_new_n1049__bF_buf1; 
wire _abc_41234_new_n1049__bF_buf2; 
wire _abc_41234_new_n1049__bF_buf3; 
wire _abc_41234_new_n1049__bF_buf4; 
wire _abc_41234_new_n1050_; 
wire _abc_41234_new_n1051_; 
wire _abc_41234_new_n1052_; 
wire _abc_41234_new_n1053_; 
wire _abc_41234_new_n1054_; 
wire _abc_41234_new_n1055_; 
wire _abc_41234_new_n1056_; 
wire _abc_41234_new_n1057_; 
wire _abc_41234_new_n1058_; 
wire _abc_41234_new_n1059_; 
wire _abc_41234_new_n1060_; 
wire _abc_41234_new_n1061_; 
wire _abc_41234_new_n1062_; 
wire _abc_41234_new_n1063_; 
wire _abc_41234_new_n1064_; 
wire _abc_41234_new_n1065_; 
wire _abc_41234_new_n1066_; 
wire _abc_41234_new_n1066__bF_buf0; 
wire _abc_41234_new_n1066__bF_buf1; 
wire _abc_41234_new_n1066__bF_buf2; 
wire _abc_41234_new_n1066__bF_buf3; 
wire _abc_41234_new_n1067_; 
wire _abc_41234_new_n1068_; 
wire _abc_41234_new_n1069_; 
wire _abc_41234_new_n1070_; 
wire _abc_41234_new_n1071_; 
wire _abc_41234_new_n1072_; 
wire _abc_41234_new_n1073_; 
wire _abc_41234_new_n1074_; 
wire _abc_41234_new_n1075_; 
wire _abc_41234_new_n1076_; 
wire _abc_41234_new_n1077_; 
wire _abc_41234_new_n1078_; 
wire _abc_41234_new_n1079_; 
wire _abc_41234_new_n1080_; 
wire _abc_41234_new_n1081_; 
wire _abc_41234_new_n1082_; 
wire _abc_41234_new_n1083_; 
wire _abc_41234_new_n1084_; 
wire _abc_41234_new_n1085_; 
wire _abc_41234_new_n1086_; 
wire _abc_41234_new_n1087_; 
wire _abc_41234_new_n1088_; 
wire _abc_41234_new_n1089_; 
wire _abc_41234_new_n1090_; 
wire _abc_41234_new_n1091_; 
wire _abc_41234_new_n1092_; 
wire _abc_41234_new_n1093_; 
wire _abc_41234_new_n1094_; 
wire _abc_41234_new_n1095_; 
wire _abc_41234_new_n1096_; 
wire _abc_41234_new_n1097_; 
wire _abc_41234_new_n1098_; 
wire _abc_41234_new_n1099_; 
wire _abc_41234_new_n1100_; 
wire _abc_41234_new_n1101_; 
wire _abc_41234_new_n1102_; 
wire _abc_41234_new_n1103_; 
wire _abc_41234_new_n1104_; 
wire _abc_41234_new_n1105_; 
wire _abc_41234_new_n1105__bF_buf0; 
wire _abc_41234_new_n1105__bF_buf1; 
wire _abc_41234_new_n1105__bF_buf2; 
wire _abc_41234_new_n1105__bF_buf3; 
wire _abc_41234_new_n1106_; 
wire _abc_41234_new_n1107_; 
wire _abc_41234_new_n1108_; 
wire _abc_41234_new_n1109_; 
wire _abc_41234_new_n1110_; 
wire _abc_41234_new_n1111_; 
wire _abc_41234_new_n1112_; 
wire _abc_41234_new_n1113_; 
wire _abc_41234_new_n1114_; 
wire _abc_41234_new_n1115_; 
wire _abc_41234_new_n1116_; 
wire _abc_41234_new_n1117_; 
wire _abc_41234_new_n1118_; 
wire _abc_41234_new_n1119_; 
wire _abc_41234_new_n1120_; 
wire _abc_41234_new_n1121_; 
wire _abc_41234_new_n1122_; 
wire _abc_41234_new_n1123_; 
wire _abc_41234_new_n1124_; 
wire _abc_41234_new_n1125_; 
wire _abc_41234_new_n1126_; 
wire _abc_41234_new_n1127_; 
wire _abc_41234_new_n1128_; 
wire _abc_41234_new_n1129_; 
wire _abc_41234_new_n1130_; 
wire _abc_41234_new_n1131_; 
wire _abc_41234_new_n1132_; 
wire _abc_41234_new_n1133_; 
wire _abc_41234_new_n1134_; 
wire _abc_41234_new_n1135_; 
wire _abc_41234_new_n1136_; 
wire _abc_41234_new_n1137_; 
wire _abc_41234_new_n1138_; 
wire _abc_41234_new_n1139_; 
wire _abc_41234_new_n1140_; 
wire _abc_41234_new_n1141_; 
wire _abc_41234_new_n1142_; 
wire _abc_41234_new_n1143_; 
wire _abc_41234_new_n1144_; 
wire _abc_41234_new_n1145_; 
wire _abc_41234_new_n1146_; 
wire _abc_41234_new_n1147_; 
wire _abc_41234_new_n1148_; 
wire _abc_41234_new_n1149_; 
wire _abc_41234_new_n1150_; 
wire _abc_41234_new_n1151_; 
wire _abc_41234_new_n1152_; 
wire _abc_41234_new_n1153_; 
wire _abc_41234_new_n1154_; 
wire _abc_41234_new_n1155_; 
wire _abc_41234_new_n1156_; 
wire _abc_41234_new_n1157_; 
wire _abc_41234_new_n1158_; 
wire _abc_41234_new_n1159_; 
wire _abc_41234_new_n1160_; 
wire _abc_41234_new_n1161_; 
wire _abc_41234_new_n1162_; 
wire _abc_41234_new_n1163_; 
wire _abc_41234_new_n1164_; 
wire _abc_41234_new_n1165_; 
wire _abc_41234_new_n1166_; 
wire _abc_41234_new_n1167_; 
wire _abc_41234_new_n1168_; 
wire _abc_41234_new_n1169_; 
wire _abc_41234_new_n1170_; 
wire _abc_41234_new_n1171_; 
wire _abc_41234_new_n1172_; 
wire _abc_41234_new_n1173_; 
wire _abc_41234_new_n1174_; 
wire _abc_41234_new_n1175_; 
wire _abc_41234_new_n1176_; 
wire _abc_41234_new_n1177_; 
wire _abc_41234_new_n1178_; 
wire _abc_41234_new_n1179_; 
wire _abc_41234_new_n1180_; 
wire _abc_41234_new_n1181_; 
wire _abc_41234_new_n1182_; 
wire _abc_41234_new_n1183_; 
wire _abc_41234_new_n1184_; 
wire _abc_41234_new_n1185_; 
wire _abc_41234_new_n1186_; 
wire _abc_41234_new_n1187_; 
wire _abc_41234_new_n1188_; 
wire _abc_41234_new_n1189_; 
wire _abc_41234_new_n1190_; 
wire _abc_41234_new_n1191_; 
wire _abc_41234_new_n1192_; 
wire _abc_41234_new_n1193_; 
wire _abc_41234_new_n1194_; 
wire _abc_41234_new_n1195_; 
wire _abc_41234_new_n1196_; 
wire _abc_41234_new_n1197_; 
wire _abc_41234_new_n1198_; 
wire _abc_41234_new_n1199_; 
wire _abc_41234_new_n1200_; 
wire _abc_41234_new_n1201_; 
wire _abc_41234_new_n1202_; 
wire _abc_41234_new_n1203_; 
wire _abc_41234_new_n1204_; 
wire _abc_41234_new_n1205_; 
wire _abc_41234_new_n1206_; 
wire _abc_41234_new_n1207_; 
wire _abc_41234_new_n1208_; 
wire _abc_41234_new_n1209_; 
wire _abc_41234_new_n1210_; 
wire _abc_41234_new_n1211_; 
wire _abc_41234_new_n1212_; 
wire _abc_41234_new_n1213_; 
wire _abc_41234_new_n1214_; 
wire _abc_41234_new_n1215_; 
wire _abc_41234_new_n1216_; 
wire _abc_41234_new_n1217_; 
wire _abc_41234_new_n1218_; 
wire _abc_41234_new_n1219_; 
wire _abc_41234_new_n1220_; 
wire _abc_41234_new_n1221_; 
wire _abc_41234_new_n1222_; 
wire _abc_41234_new_n1223_; 
wire _abc_41234_new_n1224_; 
wire _abc_41234_new_n1225_; 
wire _abc_41234_new_n1226_; 
wire _abc_41234_new_n1227_; 
wire _abc_41234_new_n1228_; 
wire _abc_41234_new_n1229_; 
wire _abc_41234_new_n1230_; 
wire _abc_41234_new_n1231_; 
wire _abc_41234_new_n1232_; 
wire _abc_41234_new_n1233_; 
wire _abc_41234_new_n1234_; 
wire _abc_41234_new_n1236_; 
wire _abc_41234_new_n1237_; 
wire _abc_41234_new_n1238_; 
wire _abc_41234_new_n1239_; 
wire _abc_41234_new_n1240_; 
wire _abc_41234_new_n1241_; 
wire _abc_41234_new_n1242_; 
wire _abc_41234_new_n1243_; 
wire _abc_41234_new_n1244_; 
wire _abc_41234_new_n1245_; 
wire _abc_41234_new_n1246_; 
wire _abc_41234_new_n1247_; 
wire _abc_41234_new_n1248_; 
wire _abc_41234_new_n1249_; 
wire _abc_41234_new_n1250_; 
wire _abc_41234_new_n1251_; 
wire _abc_41234_new_n1252_; 
wire _abc_41234_new_n1253_; 
wire _abc_41234_new_n1254_; 
wire _abc_41234_new_n1255_; 
wire _abc_41234_new_n1256_; 
wire _abc_41234_new_n1257_; 
wire _abc_41234_new_n1258_; 
wire _abc_41234_new_n1259_; 
wire _abc_41234_new_n1260_; 
wire _abc_41234_new_n1261_; 
wire _abc_41234_new_n1262_; 
wire _abc_41234_new_n1263_; 
wire _abc_41234_new_n1264_; 
wire _abc_41234_new_n1265_; 
wire _abc_41234_new_n1266_; 
wire _abc_41234_new_n1267_; 
wire _abc_41234_new_n1268_; 
wire _abc_41234_new_n1269_; 
wire _abc_41234_new_n1270_; 
wire _abc_41234_new_n1271_; 
wire _abc_41234_new_n1272_; 
wire _abc_41234_new_n1273_; 
wire _abc_41234_new_n1274_; 
wire _abc_41234_new_n1275_; 
wire _abc_41234_new_n1276_; 
wire _abc_41234_new_n1277_; 
wire _abc_41234_new_n1278_; 
wire _abc_41234_new_n1279_; 
wire _abc_41234_new_n1280_; 
wire _abc_41234_new_n1281_; 
wire _abc_41234_new_n1282_; 
wire _abc_41234_new_n1283_; 
wire _abc_41234_new_n1284_; 
wire _abc_41234_new_n1285_; 
wire _abc_41234_new_n1287_; 
wire _abc_41234_new_n1288_; 
wire _abc_41234_new_n1289_; 
wire _abc_41234_new_n1290_; 
wire _abc_41234_new_n1291_; 
wire _abc_41234_new_n1292_; 
wire _abc_41234_new_n1293_; 
wire _abc_41234_new_n1294_; 
wire _abc_41234_new_n1295_; 
wire _abc_41234_new_n1296_; 
wire _abc_41234_new_n1297_; 
wire _abc_41234_new_n1298_; 
wire _abc_41234_new_n1299_; 
wire _abc_41234_new_n1300_; 
wire _abc_41234_new_n1301_; 
wire _abc_41234_new_n1302_; 
wire _abc_41234_new_n1303_; 
wire _abc_41234_new_n1304_; 
wire _abc_41234_new_n1305_; 
wire _abc_41234_new_n1306_; 
wire _abc_41234_new_n1307_; 
wire _abc_41234_new_n1308_; 
wire _abc_41234_new_n1309_; 
wire _abc_41234_new_n1310_; 
wire _abc_41234_new_n1311_; 
wire _abc_41234_new_n1312_; 
wire _abc_41234_new_n1313_; 
wire _abc_41234_new_n1314_; 
wire _abc_41234_new_n1315_; 
wire _abc_41234_new_n1316_; 
wire _abc_41234_new_n1317_; 
wire _abc_41234_new_n1318_; 
wire _abc_41234_new_n1319_; 
wire _abc_41234_new_n1320_; 
wire _abc_41234_new_n1321_; 
wire _abc_41234_new_n1322_; 
wire _abc_41234_new_n1323_; 
wire _abc_41234_new_n1324_; 
wire _abc_41234_new_n1325_; 
wire _abc_41234_new_n1326_; 
wire _abc_41234_new_n1327_; 
wire _abc_41234_new_n1328_; 
wire _abc_41234_new_n1329_; 
wire _abc_41234_new_n1330_; 
wire _abc_41234_new_n1331_; 
wire _abc_41234_new_n1332_; 
wire _abc_41234_new_n1333_; 
wire _abc_41234_new_n1334_; 
wire _abc_41234_new_n1335_; 
wire _abc_41234_new_n1336_; 
wire _abc_41234_new_n1337_; 
wire _abc_41234_new_n1338_; 
wire _abc_41234_new_n1339_; 
wire _abc_41234_new_n1340_; 
wire _abc_41234_new_n1341_; 
wire _abc_41234_new_n1343_; 
wire _abc_41234_new_n1344_; 
wire _abc_41234_new_n1345_; 
wire _abc_41234_new_n1346_; 
wire _abc_41234_new_n1347_; 
wire _abc_41234_new_n1348_; 
wire _abc_41234_new_n1349_; 
wire _abc_41234_new_n1350_; 
wire _abc_41234_new_n1351_; 
wire _abc_41234_new_n1352_; 
wire _abc_41234_new_n1353_; 
wire _abc_41234_new_n1354_; 
wire _abc_41234_new_n1355_; 
wire _abc_41234_new_n1356_; 
wire _abc_41234_new_n1357_; 
wire _abc_41234_new_n1358_; 
wire _abc_41234_new_n1359_; 
wire _abc_41234_new_n1360_; 
wire _abc_41234_new_n1361_; 
wire _abc_41234_new_n1362_; 
wire _abc_41234_new_n1363_; 
wire _abc_41234_new_n1364_; 
wire _abc_41234_new_n1365_; 
wire _abc_41234_new_n1366_; 
wire _abc_41234_new_n1367_; 
wire _abc_41234_new_n1368_; 
wire _abc_41234_new_n1369_; 
wire _abc_41234_new_n1370_; 
wire _abc_41234_new_n1371_; 
wire _abc_41234_new_n1372_; 
wire _abc_41234_new_n1373_; 
wire _abc_41234_new_n1374_; 
wire _abc_41234_new_n1375_; 
wire _abc_41234_new_n1376_; 
wire _abc_41234_new_n1377_; 
wire _abc_41234_new_n1378_; 
wire _abc_41234_new_n1379_; 
wire _abc_41234_new_n1380_; 
wire _abc_41234_new_n1381_; 
wire _abc_41234_new_n1382_; 
wire _abc_41234_new_n1383_; 
wire _abc_41234_new_n1384_; 
wire _abc_41234_new_n1386_; 
wire _abc_41234_new_n1387_; 
wire _abc_41234_new_n1388_; 
wire _abc_41234_new_n1389_; 
wire _abc_41234_new_n1390_; 
wire _abc_41234_new_n1391_; 
wire _abc_41234_new_n1392_; 
wire _abc_41234_new_n1393_; 
wire _abc_41234_new_n1394_; 
wire _abc_41234_new_n1395_; 
wire _abc_41234_new_n1396_; 
wire _abc_41234_new_n1397_; 
wire _abc_41234_new_n1398_; 
wire _abc_41234_new_n1399_; 
wire _abc_41234_new_n1400_; 
wire _abc_41234_new_n1401_; 
wire _abc_41234_new_n1402_; 
wire _abc_41234_new_n1403_; 
wire _abc_41234_new_n1404_; 
wire _abc_41234_new_n1405_; 
wire _abc_41234_new_n1406_; 
wire _abc_41234_new_n1407_; 
wire _abc_41234_new_n1408_; 
wire _abc_41234_new_n1409_; 
wire _abc_41234_new_n1410_; 
wire _abc_41234_new_n1411_; 
wire _abc_41234_new_n1412_; 
wire _abc_41234_new_n1413_; 
wire _abc_41234_new_n1414_; 
wire _abc_41234_new_n1415_; 
wire _abc_41234_new_n1416_; 
wire _abc_41234_new_n1417_; 
wire _abc_41234_new_n1418_; 
wire _abc_41234_new_n1419_; 
wire _abc_41234_new_n1420_; 
wire _abc_41234_new_n1421_; 
wire _abc_41234_new_n1422_; 
wire _abc_41234_new_n1423_; 
wire _abc_41234_new_n1424_; 
wire _abc_41234_new_n1425_; 
wire _abc_41234_new_n1426_; 
wire _abc_41234_new_n1427_; 
wire _abc_41234_new_n1428_; 
wire _abc_41234_new_n1429_; 
wire _abc_41234_new_n1430_; 
wire _abc_41234_new_n1431_; 
wire _abc_41234_new_n1432_; 
wire _abc_41234_new_n1433_; 
wire _abc_41234_new_n1434_; 
wire _abc_41234_new_n1435_; 
wire _abc_41234_new_n1436_; 
wire _abc_41234_new_n1437_; 
wire _abc_41234_new_n1438_; 
wire _abc_41234_new_n1439_; 
wire _abc_41234_new_n1440_; 
wire _abc_41234_new_n1441_; 
wire _abc_41234_new_n1443_; 
wire _abc_41234_new_n1444_; 
wire _abc_41234_new_n1445_; 
wire _abc_41234_new_n1446_; 
wire _abc_41234_new_n1447_; 
wire _abc_41234_new_n1448_; 
wire _abc_41234_new_n1449_; 
wire _abc_41234_new_n1450_; 
wire _abc_41234_new_n1451_; 
wire _abc_41234_new_n1452_; 
wire _abc_41234_new_n1453_; 
wire _abc_41234_new_n1454_; 
wire _abc_41234_new_n1455_; 
wire _abc_41234_new_n1456_; 
wire _abc_41234_new_n1457_; 
wire _abc_41234_new_n1458_; 
wire _abc_41234_new_n1459_; 
wire _abc_41234_new_n1460_; 
wire _abc_41234_new_n1461_; 
wire _abc_41234_new_n1462_; 
wire _abc_41234_new_n1463_; 
wire _abc_41234_new_n1464_; 
wire _abc_41234_new_n1465_; 
wire _abc_41234_new_n1466_; 
wire _abc_41234_new_n1467_; 
wire _abc_41234_new_n1468_; 
wire _abc_41234_new_n1469_; 
wire _abc_41234_new_n1470_; 
wire _abc_41234_new_n1471_; 
wire _abc_41234_new_n1472_; 
wire _abc_41234_new_n1473_; 
wire _abc_41234_new_n1474_; 
wire _abc_41234_new_n1475_; 
wire _abc_41234_new_n1476_; 
wire _abc_41234_new_n1477_; 
wire _abc_41234_new_n1478_; 
wire _abc_41234_new_n1479_; 
wire _abc_41234_new_n1480_; 
wire _abc_41234_new_n1481_; 
wire _abc_41234_new_n1482_; 
wire _abc_41234_new_n1483_; 
wire _abc_41234_new_n1484_; 
wire _abc_41234_new_n1485_; 
wire _abc_41234_new_n1486_; 
wire _abc_41234_new_n1487_; 
wire _abc_41234_new_n1488_; 
wire _abc_41234_new_n1489_; 
wire _abc_41234_new_n1490_; 
wire _abc_41234_new_n1491_; 
wire _abc_41234_new_n1492_; 
wire _abc_41234_new_n1493_; 
wire _abc_41234_new_n1494_; 
wire _abc_41234_new_n1495_; 
wire _abc_41234_new_n1496_; 
wire _abc_41234_new_n1497_; 
wire _abc_41234_new_n1498_; 
wire _abc_41234_new_n1499_; 
wire _abc_41234_new_n1500_; 
wire _abc_41234_new_n1501_; 
wire _abc_41234_new_n1502_; 
wire _abc_41234_new_n1503_; 
wire _abc_41234_new_n1504_; 
wire _abc_41234_new_n1505_; 
wire _abc_41234_new_n1507_; 
wire _abc_41234_new_n1508_; 
wire _abc_41234_new_n1509_; 
wire _abc_41234_new_n1510_; 
wire _abc_41234_new_n1511_; 
wire _abc_41234_new_n1512_; 
wire _abc_41234_new_n1513_; 
wire _abc_41234_new_n1514_; 
wire _abc_41234_new_n1515_; 
wire _abc_41234_new_n1516_; 
wire _abc_41234_new_n1517_; 
wire _abc_41234_new_n1518_; 
wire _abc_41234_new_n1519_; 
wire _abc_41234_new_n1520_; 
wire _abc_41234_new_n1521_; 
wire _abc_41234_new_n1522_; 
wire _abc_41234_new_n1523_; 
wire _abc_41234_new_n1524_; 
wire _abc_41234_new_n1525_; 
wire _abc_41234_new_n1526_; 
wire _abc_41234_new_n1527_; 
wire _abc_41234_new_n1528_; 
wire _abc_41234_new_n1529_; 
wire _abc_41234_new_n1530_; 
wire _abc_41234_new_n1531_; 
wire _abc_41234_new_n1532_; 
wire _abc_41234_new_n1533_; 
wire _abc_41234_new_n1534_; 
wire _abc_41234_new_n1535_; 
wire _abc_41234_new_n1536_; 
wire _abc_41234_new_n1537_; 
wire _abc_41234_new_n1538_; 
wire _abc_41234_new_n1539_; 
wire _abc_41234_new_n1540_; 
wire _abc_41234_new_n1541_; 
wire _abc_41234_new_n1542_; 
wire _abc_41234_new_n1543_; 
wire _abc_41234_new_n1544_; 
wire _abc_41234_new_n1545_; 
wire _abc_41234_new_n1546_; 
wire _abc_41234_new_n1547_; 
wire _abc_41234_new_n1548_; 
wire _abc_41234_new_n1549_; 
wire _abc_41234_new_n1550_; 
wire _abc_41234_new_n1551_; 
wire _abc_41234_new_n1552_; 
wire _abc_41234_new_n1553_; 
wire _abc_41234_new_n1554_; 
wire _abc_41234_new_n1555_; 
wire _abc_41234_new_n1556_; 
wire _abc_41234_new_n1558_; 
wire _abc_41234_new_n1559_; 
wire _abc_41234_new_n1560_; 
wire _abc_41234_new_n1561_; 
wire _abc_41234_new_n1562_; 
wire _abc_41234_new_n1563_; 
wire _abc_41234_new_n1564_; 
wire _abc_41234_new_n1565_; 
wire _abc_41234_new_n1566_; 
wire _abc_41234_new_n1567_; 
wire _abc_41234_new_n1568_; 
wire _abc_41234_new_n1569_; 
wire _abc_41234_new_n1570_; 
wire _abc_41234_new_n1571_; 
wire _abc_41234_new_n1572_; 
wire _abc_41234_new_n1573_; 
wire _abc_41234_new_n1574_; 
wire _abc_41234_new_n1575_; 
wire _abc_41234_new_n1576_; 
wire _abc_41234_new_n1577_; 
wire _abc_41234_new_n1578_; 
wire _abc_41234_new_n1579_; 
wire _abc_41234_new_n1580_; 
wire _abc_41234_new_n1581_; 
wire _abc_41234_new_n1582_; 
wire _abc_41234_new_n1583_; 
wire _abc_41234_new_n1584_; 
wire _abc_41234_new_n1585_; 
wire _abc_41234_new_n1586_; 
wire _abc_41234_new_n1587_; 
wire _abc_41234_new_n1588_; 
wire _abc_41234_new_n1589_; 
wire _abc_41234_new_n1590_; 
wire _abc_41234_new_n1591_; 
wire _abc_41234_new_n1592_; 
wire _abc_41234_new_n1593_; 
wire _abc_41234_new_n1594_; 
wire _abc_41234_new_n1595_; 
wire _abc_41234_new_n1596_; 
wire _abc_41234_new_n1597_; 
wire _abc_41234_new_n1598_; 
wire _abc_41234_new_n1599_; 
wire _abc_41234_new_n1600_; 
wire _abc_41234_new_n1601_; 
wire _abc_41234_new_n1602_; 
wire _abc_41234_new_n1603_; 
wire _abc_41234_new_n1605_; 
wire _abc_41234_new_n1606_; 
wire _abc_41234_new_n1607_; 
wire _abc_41234_new_n1608_; 
wire _abc_41234_new_n1609_; 
wire _abc_41234_new_n1610_; 
wire _abc_41234_new_n1611_; 
wire _abc_41234_new_n1612_; 
wire _abc_41234_new_n1613_; 
wire _abc_41234_new_n1614_; 
wire _abc_41234_new_n1615_; 
wire _abc_41234_new_n1616_; 
wire _abc_41234_new_n1617_; 
wire _abc_41234_new_n1618_; 
wire _abc_41234_new_n1619_; 
wire _abc_41234_new_n1620_; 
wire _abc_41234_new_n1621_; 
wire _abc_41234_new_n1622_; 
wire _abc_41234_new_n1623_; 
wire _abc_41234_new_n1624_; 
wire _abc_41234_new_n1625_; 
wire _abc_41234_new_n1626_; 
wire _abc_41234_new_n1627_; 
wire _abc_41234_new_n1628_; 
wire _abc_41234_new_n1629_; 
wire _abc_41234_new_n1630_; 
wire _abc_41234_new_n1631_; 
wire _abc_41234_new_n1632_; 
wire _abc_41234_new_n1633_; 
wire _abc_41234_new_n1634_; 
wire _abc_41234_new_n1635_; 
wire _abc_41234_new_n1636_; 
wire _abc_41234_new_n1637_; 
wire _abc_41234_new_n1638_; 
wire _abc_41234_new_n1639_; 
wire _abc_41234_new_n1639__bF_buf0; 
wire _abc_41234_new_n1639__bF_buf1; 
wire _abc_41234_new_n1639__bF_buf2; 
wire _abc_41234_new_n1639__bF_buf3; 
wire _abc_41234_new_n1640_; 
wire _abc_41234_new_n1641_; 
wire _abc_41234_new_n1642_; 
wire _abc_41234_new_n1643_; 
wire _abc_41234_new_n1643__bF_buf0; 
wire _abc_41234_new_n1643__bF_buf1; 
wire _abc_41234_new_n1643__bF_buf2; 
wire _abc_41234_new_n1643__bF_buf3; 
wire _abc_41234_new_n1643__bF_buf4; 
wire _abc_41234_new_n1643__bF_buf5; 
wire _abc_41234_new_n1644_; 
wire _abc_41234_new_n1645_; 
wire _abc_41234_new_n1646_; 
wire _abc_41234_new_n1647_; 
wire _abc_41234_new_n1648_; 
wire _abc_41234_new_n1649_; 
wire _abc_41234_new_n1650_; 
wire _abc_41234_new_n1651_; 
wire _abc_41234_new_n1652_; 
wire _abc_41234_new_n1653_; 
wire _abc_41234_new_n1654_; 
wire _abc_41234_new_n1655_; 
wire _abc_41234_new_n1656_; 
wire _abc_41234_new_n1657_; 
wire _abc_41234_new_n1658_; 
wire _abc_41234_new_n1659_; 
wire _abc_41234_new_n1660_; 
wire _abc_41234_new_n1661_; 
wire _abc_41234_new_n1662_; 
wire _abc_41234_new_n1663_; 
wire _abc_41234_new_n1664_; 
wire _abc_41234_new_n1666_; 
wire _abc_41234_new_n1667_; 
wire _abc_41234_new_n1668_; 
wire _abc_41234_new_n1669_; 
wire _abc_41234_new_n1670_; 
wire _abc_41234_new_n1671_; 
wire _abc_41234_new_n1672_; 
wire _abc_41234_new_n1673_; 
wire _abc_41234_new_n1674_; 
wire _abc_41234_new_n1675_; 
wire _abc_41234_new_n1676_; 
wire _abc_41234_new_n1677_; 
wire _abc_41234_new_n1678_; 
wire _abc_41234_new_n1679_; 
wire _abc_41234_new_n1680_; 
wire _abc_41234_new_n1681_; 
wire _abc_41234_new_n1682_; 
wire _abc_41234_new_n1683_; 
wire _abc_41234_new_n1684_; 
wire _abc_41234_new_n1685_; 
wire _abc_41234_new_n1686_; 
wire _abc_41234_new_n1687_; 
wire _abc_41234_new_n1688_; 
wire _abc_41234_new_n1689_; 
wire _abc_41234_new_n1690_; 
wire _abc_41234_new_n1691_; 
wire _abc_41234_new_n1692_; 
wire _abc_41234_new_n1693_; 
wire _abc_41234_new_n1694_; 
wire _abc_41234_new_n1695_; 
wire _abc_41234_new_n1697_; 
wire _abc_41234_new_n1698_; 
wire _abc_41234_new_n1699_; 
wire _abc_41234_new_n1700_; 
wire _abc_41234_new_n1701_; 
wire _abc_41234_new_n1702_; 
wire _abc_41234_new_n1703_; 
wire _abc_41234_new_n1704_; 
wire _abc_41234_new_n1705_; 
wire _abc_41234_new_n1706_; 
wire _abc_41234_new_n1707_; 
wire _abc_41234_new_n1708_; 
wire _abc_41234_new_n1709_; 
wire _abc_41234_new_n1710_; 
wire _abc_41234_new_n1711_; 
wire _abc_41234_new_n1712_; 
wire _abc_41234_new_n1713_; 
wire _abc_41234_new_n1714_; 
wire _abc_41234_new_n1715_; 
wire _abc_41234_new_n1716_; 
wire _abc_41234_new_n1717_; 
wire _abc_41234_new_n1718_; 
wire _abc_41234_new_n1719_; 
wire _abc_41234_new_n1720_; 
wire _abc_41234_new_n1721_; 
wire _abc_41234_new_n1722_; 
wire _abc_41234_new_n1724_; 
wire _abc_41234_new_n1725_; 
wire _abc_41234_new_n1726_; 
wire _abc_41234_new_n1727_; 
wire _abc_41234_new_n1728_; 
wire _abc_41234_new_n1729_; 
wire _abc_41234_new_n1730_; 
wire _abc_41234_new_n1731_; 
wire _abc_41234_new_n1732_; 
wire _abc_41234_new_n1733_; 
wire _abc_41234_new_n1734_; 
wire _abc_41234_new_n1735_; 
wire _abc_41234_new_n1736_; 
wire _abc_41234_new_n1737_; 
wire _abc_41234_new_n1738_; 
wire _abc_41234_new_n1739_; 
wire _abc_41234_new_n1740_; 
wire _abc_41234_new_n1741_; 
wire _abc_41234_new_n1742_; 
wire _abc_41234_new_n1743_; 
wire _abc_41234_new_n1744_; 
wire _abc_41234_new_n1746_; 
wire _abc_41234_new_n1747_; 
wire _abc_41234_new_n1748_; 
wire _abc_41234_new_n1749_; 
wire _abc_41234_new_n1750_; 
wire _abc_41234_new_n1751_; 
wire _abc_41234_new_n1752_; 
wire _abc_41234_new_n1753_; 
wire _abc_41234_new_n1754_; 
wire _abc_41234_new_n1755_; 
wire _abc_41234_new_n1756_; 
wire _abc_41234_new_n1757_; 
wire _abc_41234_new_n1758_; 
wire _abc_41234_new_n1759_; 
wire _abc_41234_new_n1760_; 
wire _abc_41234_new_n1761_; 
wire _abc_41234_new_n1762_; 
wire _abc_41234_new_n1763_; 
wire _abc_41234_new_n1764_; 
wire _abc_41234_new_n1765_; 
wire _abc_41234_new_n1766_; 
wire _abc_41234_new_n1767_; 
wire _abc_41234_new_n1768_; 
wire _abc_41234_new_n1769_; 
wire _abc_41234_new_n1771_; 
wire _abc_41234_new_n1772_; 
wire _abc_41234_new_n1773_; 
wire _abc_41234_new_n1774_; 
wire _abc_41234_new_n1775_; 
wire _abc_41234_new_n1776_; 
wire _abc_41234_new_n1777_; 
wire _abc_41234_new_n1778_; 
wire _abc_41234_new_n1779_; 
wire _abc_41234_new_n1780_; 
wire _abc_41234_new_n1781_; 
wire _abc_41234_new_n1782_; 
wire _abc_41234_new_n1783_; 
wire _abc_41234_new_n1784_; 
wire _abc_41234_new_n1785_; 
wire _abc_41234_new_n1786_; 
wire _abc_41234_new_n1787_; 
wire _abc_41234_new_n1788_; 
wire _abc_41234_new_n1789_; 
wire _abc_41234_new_n1790_; 
wire _abc_41234_new_n1791_; 
wire _abc_41234_new_n1793_; 
wire _abc_41234_new_n1794_; 
wire _abc_41234_new_n1795_; 
wire _abc_41234_new_n1796_; 
wire _abc_41234_new_n1797_; 
wire _abc_41234_new_n1798_; 
wire _abc_41234_new_n1799_; 
wire _abc_41234_new_n1800_; 
wire _abc_41234_new_n1801_; 
wire _abc_41234_new_n1802_; 
wire _abc_41234_new_n1803_; 
wire _abc_41234_new_n1804_; 
wire _abc_41234_new_n1805_; 
wire _abc_41234_new_n1806_; 
wire _abc_41234_new_n1807_; 
wire _abc_41234_new_n1808_; 
wire _abc_41234_new_n1809_; 
wire _abc_41234_new_n1810_; 
wire _abc_41234_new_n1811_; 
wire _abc_41234_new_n1812_; 
wire _abc_41234_new_n1813_; 
wire _abc_41234_new_n1814_; 
wire _abc_41234_new_n1815_; 
wire _abc_41234_new_n1816_; 
wire _abc_41234_new_n1817_; 
wire _abc_41234_new_n1818_; 
wire _abc_41234_new_n1819_; 
wire _abc_41234_new_n1821_; 
wire _abc_41234_new_n1822_; 
wire _abc_41234_new_n1823_; 
wire _abc_41234_new_n1824_; 
wire _abc_41234_new_n1825_; 
wire _abc_41234_new_n1826_; 
wire _abc_41234_new_n1827_; 
wire _abc_41234_new_n1828_; 
wire _abc_41234_new_n1829_; 
wire _abc_41234_new_n1830_; 
wire _abc_41234_new_n1831_; 
wire _abc_41234_new_n1832_; 
wire _abc_41234_new_n1833_; 
wire _abc_41234_new_n1834_; 
wire _abc_41234_new_n1835_; 
wire _abc_41234_new_n1836_; 
wire _abc_41234_new_n1837_; 
wire _abc_41234_new_n1838_; 
wire _abc_41234_new_n1839_; 
wire _abc_41234_new_n1840_; 
wire _abc_41234_new_n1841_; 
wire _abc_41234_new_n1842_; 
wire _abc_41234_new_n1843_; 
wire _abc_41234_new_n1844_; 
wire _abc_41234_new_n1846_; 
wire _abc_41234_new_n1847_; 
wire _abc_41234_new_n1848_; 
wire _abc_41234_new_n1849_; 
wire _abc_41234_new_n1850_; 
wire _abc_41234_new_n1851_; 
wire _abc_41234_new_n1852_; 
wire _abc_41234_new_n1853_; 
wire _abc_41234_new_n1854_; 
wire _abc_41234_new_n1855_; 
wire _abc_41234_new_n1856_; 
wire _abc_41234_new_n1857_; 
wire _abc_41234_new_n1858_; 
wire _abc_41234_new_n1859_; 
wire _abc_41234_new_n1860_; 
wire _abc_41234_new_n1861_; 
wire _abc_41234_new_n1862_; 
wire _abc_41234_new_n1863_; 
wire _abc_41234_new_n1864_; 
wire _abc_41234_new_n1865_; 
wire _abc_41234_new_n1866_; 
wire _abc_41234_new_n1868_; 
wire _abc_41234_new_n1869_; 
wire _abc_41234_new_n1870_; 
wire _abc_41234_new_n1871_; 
wire _abc_41234_new_n1872_; 
wire _abc_41234_new_n1873_; 
wire _abc_41234_new_n1874_; 
wire _abc_41234_new_n1875_; 
wire _abc_41234_new_n1876_; 
wire _abc_41234_new_n1877_; 
wire _abc_41234_new_n1878_; 
wire _abc_41234_new_n1879_; 
wire _abc_41234_new_n1880_; 
wire _abc_41234_new_n1881_; 
wire _abc_41234_new_n1882_; 
wire _abc_41234_new_n1884_; 
wire _abc_41234_new_n1885_; 
wire _abc_41234_new_n1886_; 
wire _abc_41234_new_n1887_; 
wire _abc_41234_new_n1888_; 
wire _abc_41234_new_n1889_; 
wire _abc_41234_new_n1890_; 
wire _abc_41234_new_n1891_; 
wire _abc_41234_new_n1892_; 
wire _abc_41234_new_n1893_; 
wire _abc_41234_new_n1894_; 
wire _abc_41234_new_n1895_; 
wire _abc_41234_new_n1897_; 
wire _abc_41234_new_n1898_; 
wire _abc_41234_new_n1899_; 
wire _abc_41234_new_n1900_; 
wire _abc_41234_new_n1901_; 
wire _abc_41234_new_n1902_; 
wire _abc_41234_new_n1903_; 
wire _abc_41234_new_n1904_; 
wire _abc_41234_new_n1905_; 
wire _abc_41234_new_n1906_; 
wire _abc_41234_new_n1908_; 
wire _abc_41234_new_n1909_; 
wire _abc_41234_new_n1910_; 
wire _abc_41234_new_n1911_; 
wire _abc_41234_new_n1912_; 
wire _abc_41234_new_n1913_; 
wire _abc_41234_new_n1914_; 
wire _abc_41234_new_n1915_; 
wire _abc_41234_new_n1916_; 
wire _abc_41234_new_n1917_; 
wire _abc_41234_new_n1918_; 
wire _abc_41234_new_n1919_; 
wire _abc_41234_new_n1920_; 
wire _abc_41234_new_n1922_; 
wire _abc_41234_new_n1923_; 
wire _abc_41234_new_n1924_; 
wire _abc_41234_new_n1925_; 
wire _abc_41234_new_n1926_; 
wire _abc_41234_new_n1927_; 
wire _abc_41234_new_n1928_; 
wire _abc_41234_new_n1929_; 
wire _abc_41234_new_n1930_; 
wire _abc_41234_new_n1931_; 
wire _abc_41234_new_n1932_; 
wire _abc_41234_new_n1933_; 
wire _abc_41234_new_n1934_; 
wire _abc_41234_new_n1936_; 
wire _abc_41234_new_n1937_; 
wire _abc_41234_new_n1938_; 
wire _abc_41234_new_n1939_; 
wire _abc_41234_new_n1940_; 
wire _abc_41234_new_n1941_; 
wire _abc_41234_new_n1942_; 
wire _abc_41234_new_n1943_; 
wire _abc_41234_new_n1944_; 
wire _abc_41234_new_n1945_; 
wire _abc_41234_new_n1946_; 
wire _abc_41234_new_n1947_; 
wire _abc_41234_new_n1949_; 
wire _abc_41234_new_n1950_; 
wire _abc_41234_new_n1951_; 
wire _abc_41234_new_n1952_; 
wire _abc_41234_new_n1953_; 
wire _abc_41234_new_n1954_; 
wire _abc_41234_new_n1955_; 
wire _abc_41234_new_n1956_; 
wire _abc_41234_new_n1957_; 
wire _abc_41234_new_n1958_; 
wire _abc_41234_new_n1959_; 
wire _abc_41234_new_n1960_; 
wire _abc_41234_new_n1961_; 
wire _abc_41234_new_n1962_; 
wire _abc_41234_new_n1963_; 
wire _abc_41234_new_n1964_; 
wire _abc_41234_new_n1966_; 
wire _abc_41234_new_n1967_; 
wire _abc_41234_new_n1968_; 
wire _abc_41234_new_n1969_; 
wire _abc_41234_new_n1970_; 
wire _abc_41234_new_n1971_; 
wire _abc_41234_new_n1973_; 
wire _abc_41234_new_n1974_; 
wire _abc_41234_new_n1975_; 
wire _abc_41234_new_n1976_; 
wire _abc_41234_new_n1977_; 
wire _abc_41234_new_n1978_; 
wire _abc_41234_new_n1979_; 
wire _abc_41234_new_n1980_; 
wire _abc_41234_new_n1982_; 
wire _abc_41234_new_n1983_; 
wire _abc_41234_new_n1984_; 
wire _abc_41234_new_n1985_; 
wire _abc_41234_new_n1986_; 
wire _abc_41234_new_n1987_; 
wire _abc_41234_new_n1988_; 
wire _abc_41234_new_n1989_; 
wire _abc_41234_new_n1991_; 
wire _abc_41234_new_n1992_; 
wire _abc_41234_new_n1993_; 
wire _abc_41234_new_n1994_; 
wire _abc_41234_new_n1995_; 
wire _abc_41234_new_n1996_; 
wire _abc_41234_new_n1997_; 
wire _abc_41234_new_n1998_; 
wire _abc_41234_new_n1999_; 
wire _abc_41234_new_n2001_; 
wire _abc_41234_new_n2002_; 
wire _abc_41234_new_n2003_; 
wire _abc_41234_new_n2004_; 
wire _abc_41234_new_n2005_; 
wire _abc_41234_new_n2006_; 
wire _abc_41234_new_n2008_; 
wire _abc_41234_new_n2009_; 
wire _abc_41234_new_n2010_; 
wire _abc_41234_new_n2011_; 
wire _abc_41234_new_n2012_; 
wire _abc_41234_new_n2013_; 
wire _abc_41234_new_n2014_; 
wire _abc_41234_new_n2015_; 
wire _abc_41234_new_n2017_; 
wire _abc_41234_new_n2018_; 
wire _abc_41234_new_n2019_; 
wire _abc_41234_new_n2020_; 
wire _abc_41234_new_n2021_; 
wire _abc_41234_new_n2022_; 
wire _abc_41234_new_n2023_; 
wire _abc_41234_new_n2024_; 
wire _abc_41234_new_n2026_; 
wire _abc_41234_new_n2027_; 
wire _abc_41234_new_n2028_; 
wire _abc_41234_new_n2029_; 
wire _abc_41234_new_n2030_; 
wire _abc_41234_new_n2031_; 
wire _abc_41234_new_n2032_; 
wire _abc_41234_new_n2033_; 
wire _abc_41234_new_n2035_; 
wire _abc_41234_new_n2036_; 
wire _abc_41234_new_n2038_; 
wire _abc_41234_new_n2040_; 
wire _abc_41234_new_n2042_; 
wire _abc_41234_new_n2044_; 
wire _abc_41234_new_n2046_; 
wire _abc_41234_new_n2048_; 
wire _abc_41234_new_n2049_; 
wire _abc_41234_new_n2051_; 
wire _abc_41234_new_n2053_; 
wire _abc_41234_new_n2054_; 
wire _abc_41234_new_n2055_; 
wire _abc_41234_new_n2056_; 
wire _abc_41234_new_n2057_; 
wire _abc_41234_new_n2058_; 
wire _abc_41234_new_n2059_; 
wire _abc_41234_new_n2060_; 
wire _abc_41234_new_n2061_; 
wire _abc_41234_new_n2062_; 
wire _abc_41234_new_n2063_; 
wire _abc_41234_new_n2064_; 
wire _abc_41234_new_n2065_; 
wire _abc_41234_new_n2066_; 
wire _abc_41234_new_n2068_; 
wire _abc_41234_new_n2069_; 
wire _abc_41234_new_n2070_; 
wire _abc_41234_new_n2071_; 
wire _abc_41234_new_n2072_; 
wire _abc_41234_new_n2073_; 
wire _abc_41234_new_n2074_; 
wire _abc_41234_new_n2075_; 
wire _abc_41234_new_n2076_; 
wire _abc_41234_new_n2077_; 
wire _abc_41234_new_n2078_; 
wire _abc_41234_new_n2080_; 
wire _abc_41234_new_n2081_; 
wire _abc_41234_new_n2082_; 
wire _abc_41234_new_n2083_; 
wire _abc_41234_new_n2084_; 
wire _abc_41234_new_n2085_; 
wire _abc_41234_new_n2086_; 
wire _abc_41234_new_n2087_; 
wire _abc_41234_new_n2088_; 
wire _abc_41234_new_n2089_; 
wire _abc_41234_new_n2090_; 
wire _abc_41234_new_n2092_; 
wire _abc_41234_new_n2093_; 
wire _abc_41234_new_n2094_; 
wire _abc_41234_new_n2095_; 
wire _abc_41234_new_n2096_; 
wire _abc_41234_new_n2097_; 
wire _abc_41234_new_n2098_; 
wire _abc_41234_new_n2099_; 
wire _abc_41234_new_n2100_; 
wire _abc_41234_new_n2101_; 
wire _abc_41234_new_n2102_; 
wire _abc_41234_new_n2103_; 
wire _abc_41234_new_n2104_; 
wire _abc_41234_new_n2106_; 
wire _abc_41234_new_n2107_; 
wire _abc_41234_new_n2108_; 
wire _abc_41234_new_n2109_; 
wire _abc_41234_new_n2110_; 
wire _abc_41234_new_n2111_; 
wire _abc_41234_new_n2112_; 
wire _abc_41234_new_n2113_; 
wire _abc_41234_new_n2114_; 
wire _abc_41234_new_n2115_; 
wire _abc_41234_new_n2116_; 
wire _abc_41234_new_n2118_; 
wire _abc_41234_new_n2119_; 
wire _abc_41234_new_n2120_; 
wire _abc_41234_new_n2121_; 
wire _abc_41234_new_n2122_; 
wire _abc_41234_new_n2123_; 
wire _abc_41234_new_n2124_; 
wire _abc_41234_new_n2125_; 
wire _abc_41234_new_n2126_; 
wire _abc_41234_new_n2127_; 
wire _abc_41234_new_n2128_; 
wire _abc_41234_new_n2130_; 
wire _abc_41234_new_n2131_; 
wire _abc_41234_new_n2132_; 
wire _abc_41234_new_n2133_; 
wire _abc_41234_new_n2134_; 
wire _abc_41234_new_n2135_; 
wire _abc_41234_new_n2136_; 
wire _abc_41234_new_n2137_; 
wire _abc_41234_new_n2138_; 
wire _abc_41234_new_n2139_; 
wire _abc_41234_new_n2140_; 
wire _abc_41234_new_n2141_; 
wire _abc_41234_new_n2142_; 
wire _abc_41234_new_n2143_; 
wire _abc_41234_new_n2144_; 
wire _abc_41234_new_n2145_; 
wire _abc_41234_new_n2146_; 
wire _abc_41234_new_n2147_; 
wire _abc_41234_new_n2148_; 
wire _abc_41234_new_n2149_; 
wire _abc_41234_new_n2150_; 
wire _abc_41234_new_n2151_; 
wire _abc_41234_new_n2152_; 
wire _abc_41234_new_n2153_; 
wire _abc_41234_new_n2154_; 
wire _abc_41234_new_n2155_; 
wire _abc_41234_new_n2156_; 
wire _abc_41234_new_n2157_; 
wire _abc_41234_new_n2159_; 
wire _abc_41234_new_n2160_; 
wire _abc_41234_new_n2161_; 
wire _abc_41234_new_n2162_; 
wire _abc_41234_new_n2163_; 
wire _abc_41234_new_n2164_; 
wire _abc_41234_new_n2165_; 
wire _abc_41234_new_n2166_; 
wire _abc_41234_new_n2167_; 
wire _abc_41234_new_n2168_; 
wire _abc_41234_new_n2169_; 
wire _abc_41234_new_n2170_; 
wire _abc_41234_new_n2171_; 
wire _abc_41234_new_n2172_; 
wire _abc_41234_new_n2174_; 
wire _abc_41234_new_n2175_; 
wire _abc_41234_new_n2176_; 
wire _abc_41234_new_n2177_; 
wire _abc_41234_new_n2178_; 
wire _abc_41234_new_n2179_; 
wire _abc_41234_new_n2180_; 
wire _abc_41234_new_n2181_; 
wire _abc_41234_new_n2182_; 
wire _abc_41234_new_n2184_; 
wire _abc_41234_new_n2185_; 
wire _abc_41234_new_n2185__bF_buf0; 
wire _abc_41234_new_n2185__bF_buf1; 
wire _abc_41234_new_n2185__bF_buf2; 
wire _abc_41234_new_n2185__bF_buf3; 
wire _abc_41234_new_n2185__bF_buf4; 
wire _abc_41234_new_n2185__bF_buf5; 
wire _abc_41234_new_n2186_; 
wire _abc_41234_new_n2187_; 
wire _abc_41234_new_n2188_; 
wire _abc_41234_new_n2189_; 
wire _abc_41234_new_n2189__bF_buf0; 
wire _abc_41234_new_n2189__bF_buf1; 
wire _abc_41234_new_n2189__bF_buf2; 
wire _abc_41234_new_n2189__bF_buf3; 
wire _abc_41234_new_n2189__bF_buf4; 
wire _abc_41234_new_n2189__bF_buf5; 
wire _abc_41234_new_n2190_; 
wire _abc_41234_new_n2190__bF_buf0; 
wire _abc_41234_new_n2190__bF_buf1; 
wire _abc_41234_new_n2190__bF_buf2; 
wire _abc_41234_new_n2190__bF_buf3; 
wire _abc_41234_new_n2191_; 
wire _abc_41234_new_n2192_; 
wire _abc_41234_new_n2193_; 
wire _abc_41234_new_n2195_; 
wire _abc_41234_new_n2196_; 
wire _abc_41234_new_n2197_; 
wire _abc_41234_new_n2198_; 
wire _abc_41234_new_n2199_; 
wire _abc_41234_new_n2201_; 
wire _abc_41234_new_n2202_; 
wire _abc_41234_new_n2203_; 
wire _abc_41234_new_n2205_; 
wire _abc_41234_new_n2206_; 
wire _abc_41234_new_n2207_; 
wire _abc_41234_new_n2207__bF_buf0; 
wire _abc_41234_new_n2207__bF_buf1; 
wire _abc_41234_new_n2207__bF_buf2; 
wire _abc_41234_new_n2207__bF_buf3; 
wire _abc_41234_new_n2208_; 
wire _abc_41234_new_n2209_; 
wire _abc_41234_new_n2210_; 
wire _abc_41234_new_n2211_; 
wire _abc_41234_new_n2212_; 
wire _abc_41234_new_n2213_; 
wire _abc_41234_new_n2214_; 
wire _abc_41234_new_n2215_; 
wire _abc_41234_new_n2216_; 
wire _abc_41234_new_n2217_; 
wire _abc_41234_new_n2218_; 
wire _abc_41234_new_n2220_; 
wire _abc_41234_new_n2221_; 
wire _abc_41234_new_n2222_; 
wire _abc_41234_new_n2223_; 
wire _abc_41234_new_n2224_; 
wire _abc_41234_new_n2225_; 
wire _abc_41234_new_n2227_; 
wire _abc_41234_new_n2228_; 
wire _abc_41234_new_n2230_; 
wire _abc_41234_new_n2231_; 
wire _abc_41234_new_n2233_; 
wire _abc_41234_new_n2234_; 
wire _abc_41234_new_n2236_; 
wire _abc_41234_new_n2237_; 
wire _abc_41234_new_n2239_; 
wire _abc_41234_new_n2240_; 
wire _abc_41234_new_n2242_; 
wire _abc_41234_new_n2243_; 
wire _abc_41234_new_n2245_; 
wire _abc_41234_new_n2246_; 
wire _abc_41234_new_n2247_; 
wire _abc_41234_new_n2248_; 
wire _abc_41234_new_n2249_; 
wire _abc_41234_new_n2250_; 
wire _abc_41234_new_n2251_; 
wire _abc_41234_new_n2252_; 
wire _abc_41234_new_n2253_; 
wire _abc_41234_new_n2254_; 
wire _abc_41234_new_n2255_; 
wire _abc_41234_new_n2256_; 
wire _abc_41234_new_n2257_; 
wire _abc_41234_new_n2258_; 
wire _abc_41234_new_n2259_; 
wire _abc_41234_new_n2260_; 
wire _abc_41234_new_n2261_; 
wire _abc_41234_new_n2262_; 
wire _abc_41234_new_n2263_; 
wire _abc_41234_new_n2264_; 
wire _abc_41234_new_n2265_; 
wire _abc_41234_new_n2266_; 
wire _abc_41234_new_n2267_; 
wire _abc_41234_new_n2269_; 
wire _abc_41234_new_n2270_; 
wire _abc_41234_new_n2271_; 
wire _abc_41234_new_n2272_; 
wire _abc_41234_new_n2273_; 
wire _abc_41234_new_n2274_; 
wire _abc_41234_new_n2275_; 
wire _abc_41234_new_n2276_; 
wire _abc_41234_new_n2277_; 
wire _abc_41234_new_n2278_; 
wire _abc_41234_new_n2279_; 
wire _abc_41234_new_n2281_; 
wire _abc_41234_new_n2282_; 
wire _abc_41234_new_n2283_; 
wire _abc_41234_new_n2284_; 
wire _abc_41234_new_n2285_; 
wire _abc_41234_new_n2286_; 
wire _abc_41234_new_n2287_; 
wire _abc_41234_new_n2288_; 
wire _abc_41234_new_n2289_; 
wire _abc_41234_new_n2290_; 
wire _abc_41234_new_n2291_; 
wire _abc_41234_new_n2293_; 
wire _abc_41234_new_n2294_; 
wire _abc_41234_new_n2295_; 
wire _abc_41234_new_n2296_; 
wire _abc_41234_new_n2297_; 
wire _abc_41234_new_n2298_; 
wire _abc_41234_new_n2299_; 
wire _abc_41234_new_n2300_; 
wire _abc_41234_new_n2301_; 
wire _abc_41234_new_n2302_; 
wire _abc_41234_new_n2303_; 
wire _abc_41234_new_n2305_; 
wire _abc_41234_new_n2306_; 
wire _abc_41234_new_n2307_; 
wire _abc_41234_new_n2308_; 
wire _abc_41234_new_n2309_; 
wire _abc_41234_new_n2310_; 
wire _abc_41234_new_n2311_; 
wire _abc_41234_new_n2312_; 
wire _abc_41234_new_n2313_; 
wire _abc_41234_new_n2314_; 
wire _abc_41234_new_n2315_; 
wire _abc_41234_new_n2317_; 
wire _abc_41234_new_n2318_; 
wire _abc_41234_new_n2319_; 
wire _abc_41234_new_n2320_; 
wire _abc_41234_new_n2321_; 
wire _abc_41234_new_n2322_; 
wire _abc_41234_new_n2323_; 
wire _abc_41234_new_n2324_; 
wire _abc_41234_new_n2325_; 
wire _abc_41234_new_n2326_; 
wire _abc_41234_new_n2327_; 
wire _abc_41234_new_n2328_; 
wire _abc_41234_new_n2330_; 
wire _abc_41234_new_n2331_; 
wire _abc_41234_new_n2332_; 
wire _abc_41234_new_n2333_; 
wire _abc_41234_new_n2334_; 
wire _abc_41234_new_n2335_; 
wire _abc_41234_new_n2336_; 
wire _abc_41234_new_n2337_; 
wire _abc_41234_new_n2338_; 
wire _abc_41234_new_n2339_; 
wire _abc_41234_new_n2340_; 
wire _abc_41234_new_n2342_; 
wire _abc_41234_new_n2343_; 
wire _abc_41234_new_n2344_; 
wire _abc_41234_new_n2345_; 
wire _abc_41234_new_n2346_; 
wire _abc_41234_new_n2347_; 
wire _abc_41234_new_n2348_; 
wire _abc_41234_new_n2349_; 
wire _abc_41234_new_n2350_; 
wire _abc_41234_new_n2351_; 
wire _abc_41234_new_n2353_; 
wire _abc_41234_new_n2354_; 
wire _abc_41234_new_n2355_; 
wire _abc_41234_new_n2356_; 
wire _abc_41234_new_n2357_; 
wire _abc_41234_new_n2358_; 
wire _abc_41234_new_n2359_; 
wire _abc_41234_new_n2361_; 
wire _abc_41234_new_n2362_; 
wire _abc_41234_new_n2363_; 
wire _abc_41234_new_n2364_; 
wire _abc_41234_new_n2365_; 
wire _abc_41234_new_n2366_; 
wire _abc_41234_new_n2367_; 
wire _abc_41234_new_n2368_; 
wire _abc_41234_new_n2370_; 
wire _abc_41234_new_n2371_; 
wire _abc_41234_new_n2372_; 
wire _abc_41234_new_n2373_; 
wire _abc_41234_new_n2374_; 
wire _abc_41234_new_n2376_; 
wire _abc_41234_new_n2377_; 
wire _abc_41234_new_n2378_; 
wire _abc_41234_new_n2379_; 
wire _abc_41234_new_n2380_; 
wire _abc_41234_new_n2381_; 
wire _abc_41234_new_n2382_; 
wire _abc_41234_new_n2384_; 
wire _abc_41234_new_n2385_; 
wire _abc_41234_new_n2386_; 
wire _abc_41234_new_n2387_; 
wire _abc_41234_new_n2388_; 
wire _abc_41234_new_n2389_; 
wire _abc_41234_new_n2390_; 
wire _abc_41234_new_n2391_; 
wire _abc_41234_new_n2393_; 
wire _abc_41234_new_n2394_; 
wire _abc_41234_new_n2395_; 
wire _abc_41234_new_n2396_; 
wire _abc_41234_new_n2397_; 
wire _abc_41234_new_n2398_; 
wire _abc_41234_new_n2399_; 
wire _abc_41234_new_n2400_; 
wire _abc_41234_new_n2401_; 
wire _abc_41234_new_n2402_; 
wire _abc_41234_new_n2403_; 
wire _abc_41234_new_n2404_; 
wire _abc_41234_new_n2405_; 
wire _abc_41234_new_n2406_; 
wire _abc_41234_new_n2407_; 
wire _abc_41234_new_n2408_; 
wire _abc_41234_new_n2409_; 
wire _abc_41234_new_n2410_; 
wire _abc_41234_new_n2411_; 
wire _abc_41234_new_n2412_; 
wire _abc_41234_new_n2413_; 
wire _abc_41234_new_n2414_; 
wire _abc_41234_new_n2415_; 
wire _abc_41234_new_n2415__bF_buf0; 
wire _abc_41234_new_n2415__bF_buf1; 
wire _abc_41234_new_n2415__bF_buf2; 
wire _abc_41234_new_n2415__bF_buf3; 
wire _abc_41234_new_n2415__bF_buf4; 
wire _abc_41234_new_n2416_; 
wire _abc_41234_new_n2417_; 
wire _abc_41234_new_n2418_; 
wire _abc_41234_new_n2419_; 
wire _abc_41234_new_n2420_; 
wire _abc_41234_new_n2421_; 
wire _abc_41234_new_n2422_; 
wire _abc_41234_new_n2423_; 
wire _abc_41234_new_n2424_; 
wire _abc_41234_new_n2425_; 
wire _abc_41234_new_n2427_; 
wire _abc_41234_new_n2428_; 
wire _abc_41234_new_n2429_; 
wire _abc_41234_new_n2430_; 
wire _abc_41234_new_n2432_; 
wire _abc_41234_new_n2433_; 
wire _abc_41234_new_n2435_; 
wire _abc_41234_new_n2437_; 
wire _abc_41234_new_n2438_; 
wire _abc_41234_new_n2441_; 
wire _abc_41234_new_n2443_; 
wire _abc_41234_new_n2444_; 
wire _abc_41234_new_n2446_; 
wire _abc_41234_new_n2448_; 
wire _abc_41234_new_n2449_; 
wire _abc_41234_new_n2450_; 
wire _abc_41234_new_n2451_; 
wire _abc_41234_new_n2452_; 
wire _abc_41234_new_n2453_; 
wire _abc_41234_new_n2455_; 
wire _abc_41234_new_n2456_; 
wire _abc_41234_new_n2457_; 
wire _abc_41234_new_n2458_; 
wire _abc_41234_new_n2459_; 
wire _abc_41234_new_n2460_; 
wire _abc_41234_new_n2461_; 
wire _abc_41234_new_n2462_; 
wire _abc_41234_new_n2463_; 
wire _abc_41234_new_n2464_; 
wire _abc_41234_new_n2465_; 
wire _abc_41234_new_n2466_; 
wire _abc_41234_new_n2467_; 
wire _abc_41234_new_n2468_; 
wire _abc_41234_new_n2469_; 
wire _abc_41234_new_n2470_; 
wire _abc_41234_new_n2471_; 
wire _abc_41234_new_n2472_; 
wire _abc_41234_new_n2473_; 
wire _abc_41234_new_n2474_; 
wire _abc_41234_new_n2475_; 
wire _abc_41234_new_n2476_; 
wire _abc_41234_new_n2477_; 
wire _abc_41234_new_n2478_; 
wire _abc_41234_new_n2479_; 
wire _abc_41234_new_n2480_; 
wire _abc_41234_new_n2481_; 
wire _abc_41234_new_n2482_; 
wire _abc_41234_new_n2483_; 
wire _abc_41234_new_n2484_; 
wire _abc_41234_new_n2485_; 
wire _abc_41234_new_n2486_; 
wire _abc_41234_new_n2487_; 
wire _abc_41234_new_n2488_; 
wire _abc_41234_new_n2489_; 
wire _abc_41234_new_n2490_; 
wire _abc_41234_new_n2491_; 
wire _abc_41234_new_n2492_; 
wire _abc_41234_new_n2493_; 
wire _abc_41234_new_n2494_; 
wire _abc_41234_new_n2495_; 
wire _abc_41234_new_n2496_; 
wire _abc_41234_new_n2497_; 
wire _abc_41234_new_n2498_; 
wire _abc_41234_new_n2499_; 
wire _abc_41234_new_n2500_; 
wire _abc_41234_new_n2501_; 
wire _abc_41234_new_n2502_; 
wire _abc_41234_new_n2503_; 
wire _abc_41234_new_n2504_; 
wire _abc_41234_new_n2505_; 
wire _abc_41234_new_n2506_; 
wire _abc_41234_new_n2507_; 
wire _abc_41234_new_n2508_; 
wire _abc_41234_new_n2509_; 
wire _abc_41234_new_n2510_; 
wire _abc_41234_new_n2511_; 
wire _abc_41234_new_n2512_; 
wire _abc_41234_new_n2513_; 
wire _abc_41234_new_n2514_; 
wire _abc_41234_new_n2515_; 
wire _abc_41234_new_n2516_; 
wire _abc_41234_new_n2517_; 
wire _abc_41234_new_n2518_; 
wire _abc_41234_new_n2519_; 
wire _abc_41234_new_n2520_; 
wire _abc_41234_new_n2521_; 
wire _abc_41234_new_n2522_; 
wire _abc_41234_new_n2523_; 
wire _abc_41234_new_n2524_; 
wire _abc_41234_new_n2525_; 
wire _abc_41234_new_n2526_; 
wire _abc_41234_new_n2527_; 
wire _abc_41234_new_n2528_; 
wire _abc_41234_new_n2529_; 
wire _abc_41234_new_n2530_; 
wire _abc_41234_new_n2531_; 
wire _abc_41234_new_n2532_; 
wire _abc_41234_new_n2533_; 
wire _abc_41234_new_n2534_; 
wire _abc_41234_new_n2535_; 
wire _abc_41234_new_n2536_; 
wire _abc_41234_new_n2538_; 
wire _abc_41234_new_n2539_; 
wire _abc_41234_new_n2540_; 
wire _abc_41234_new_n2541_; 
wire _abc_41234_new_n2542_; 
wire _abc_41234_new_n2543_; 
wire _abc_41234_new_n2544_; 
wire _abc_41234_new_n2545_; 
wire _abc_41234_new_n2546_; 
wire _abc_41234_new_n2547_; 
wire _abc_41234_new_n2548_; 
wire _abc_41234_new_n2549_; 
wire _abc_41234_new_n2550_; 
wire _abc_41234_new_n2551_; 
wire _abc_41234_new_n2552_; 
wire _abc_41234_new_n2553_; 
wire _abc_41234_new_n2554_; 
wire _abc_41234_new_n2555_; 
wire _abc_41234_new_n2556_; 
wire _abc_41234_new_n2557_; 
wire _abc_41234_new_n2558_; 
wire _abc_41234_new_n2559_; 
wire _abc_41234_new_n2560_; 
wire _abc_41234_new_n2561_; 
wire _abc_41234_new_n2563_; 
wire _abc_41234_new_n2564_; 
wire _abc_41234_new_n2565_; 
wire _abc_41234_new_n2566_; 
wire _abc_41234_new_n2567_; 
wire _abc_41234_new_n2568_; 
wire _abc_41234_new_n2569_; 
wire _abc_41234_new_n2570_; 
wire _abc_41234_new_n2571_; 
wire _abc_41234_new_n2572_; 
wire _abc_41234_new_n2573_; 
wire _abc_41234_new_n2574_; 
wire _abc_41234_new_n2575_; 
wire _abc_41234_new_n2576_; 
wire _abc_41234_new_n2577_; 
wire _abc_41234_new_n2578_; 
wire _abc_41234_new_n2579_; 
wire _abc_41234_new_n2580_; 
wire _abc_41234_new_n2581_; 
wire _abc_41234_new_n2582_; 
wire _abc_41234_new_n2583_; 
wire _abc_41234_new_n2584_; 
wire _abc_41234_new_n2585_; 
wire _abc_41234_new_n2586_; 
wire _abc_41234_new_n2588_; 
wire _abc_41234_new_n2589_; 
wire _abc_41234_new_n2590_; 
wire _abc_41234_new_n2591_; 
wire _abc_41234_new_n2592_; 
wire _abc_41234_new_n2593_; 
wire _abc_41234_new_n2594_; 
wire _abc_41234_new_n2595_; 
wire _abc_41234_new_n2596_; 
wire _abc_41234_new_n2597_; 
wire _abc_41234_new_n2598_; 
wire _abc_41234_new_n2599_; 
wire _abc_41234_new_n2600_; 
wire _abc_41234_new_n2601_; 
wire _abc_41234_new_n2602_; 
wire _abc_41234_new_n2603_; 
wire _abc_41234_new_n2604_; 
wire _abc_41234_new_n2605_; 
wire _abc_41234_new_n2606_; 
wire _abc_41234_new_n2607_; 
wire _abc_41234_new_n2608_; 
wire _abc_41234_new_n2609_; 
wire _abc_41234_new_n2611_; 
wire _abc_41234_new_n2612_; 
wire _abc_41234_new_n2613_; 
wire _abc_41234_new_n2614_; 
wire _abc_41234_new_n2615_; 
wire _abc_41234_new_n2616_; 
wire _abc_41234_new_n2617_; 
wire _abc_41234_new_n2618_; 
wire _abc_41234_new_n2619_; 
wire _abc_41234_new_n2620_; 
wire _abc_41234_new_n2621_; 
wire _abc_41234_new_n2622_; 
wire _abc_41234_new_n2623_; 
wire _abc_41234_new_n2624_; 
wire _abc_41234_new_n2625_; 
wire _abc_41234_new_n2626_; 
wire _abc_41234_new_n2627_; 
wire _abc_41234_new_n2629_; 
wire _abc_41234_new_n2630_; 
wire _abc_41234_new_n2631_; 
wire _abc_41234_new_n2632_; 
wire _abc_41234_new_n2633_; 
wire _abc_41234_new_n2634_; 
wire _abc_41234_new_n2635_; 
wire _abc_41234_new_n2636_; 
wire _abc_41234_new_n2637_; 
wire _abc_41234_new_n2638_; 
wire _abc_41234_new_n2639_; 
wire _abc_41234_new_n2640_; 
wire _abc_41234_new_n2641_; 
wire _abc_41234_new_n2642_; 
wire _abc_41234_new_n2644_; 
wire _abc_41234_new_n2645_; 
wire _abc_41234_new_n2647_; 
wire _abc_41234_new_n2649_; 
wire _abc_41234_new_n2651_; 
wire _abc_41234_new_n2654_; 
wire _abc_41234_new_n2656_; 
wire _abc_41234_new_n2658_; 
wire _abc_41234_new_n2670_; 
wire _abc_41234_new_n2671_; 
wire _abc_41234_new_n2672_; 
wire _abc_41234_new_n2673_; 
wire _abc_41234_new_n2674_; 
wire _abc_41234_new_n2675_; 
wire _abc_41234_new_n2676_; 
wire _abc_41234_new_n2677_; 
wire _abc_41234_new_n2678_; 
wire _abc_41234_new_n2679_; 
wire _abc_41234_new_n2680_; 
wire _abc_41234_new_n2681_; 
wire _abc_41234_new_n2682_; 
wire _abc_41234_new_n2683_; 
wire _abc_41234_new_n2684_; 
wire _abc_41234_new_n2685_; 
wire _abc_41234_new_n2686_; 
wire _abc_41234_new_n2687_; 
wire _abc_41234_new_n2688_; 
wire _abc_41234_new_n2689_; 
wire _abc_41234_new_n2690_; 
wire _abc_41234_new_n2691_; 
wire _abc_41234_new_n2692_; 
wire _abc_41234_new_n2693_; 
wire _abc_41234_new_n2694_; 
wire _abc_41234_new_n2695_; 
wire _abc_41234_new_n2696_; 
wire _abc_41234_new_n2696__bF_buf0; 
wire _abc_41234_new_n2696__bF_buf1; 
wire _abc_41234_new_n2696__bF_buf2; 
wire _abc_41234_new_n2696__bF_buf3; 
wire _abc_41234_new_n2696__bF_buf4; 
wire _abc_41234_new_n2697_; 
wire _abc_41234_new_n2698_; 
wire _abc_41234_new_n2699_; 
wire _abc_41234_new_n2701_; 
wire _abc_41234_new_n2702_; 
wire _abc_41234_new_n2703_; 
wire _abc_41234_new_n2704_; 
wire _abc_41234_new_n2705_; 
wire _abc_41234_new_n2706_; 
wire _abc_41234_new_n2707_; 
wire _abc_41234_new_n2708_; 
wire _abc_41234_new_n2709_; 
wire _abc_41234_new_n2710_; 
wire _abc_41234_new_n2711_; 
wire _abc_41234_new_n2712_; 
wire _abc_41234_new_n2713_; 
wire _abc_41234_new_n2714_; 
wire _abc_41234_new_n2715_; 
wire _abc_41234_new_n2716_; 
wire _abc_41234_new_n2717_; 
wire _abc_41234_new_n2718_; 
wire _abc_41234_new_n2719_; 
wire _abc_41234_new_n2720_; 
wire _abc_41234_new_n2721_; 
wire _abc_41234_new_n2722_; 
wire _abc_41234_new_n2723_; 
wire _abc_41234_new_n2724_; 
wire _abc_41234_new_n2725_; 
wire _abc_41234_new_n2726_; 
wire _abc_41234_new_n2727_; 
wire _abc_41234_new_n2728_; 
wire _abc_41234_new_n2729_; 
wire _abc_41234_new_n2731_; 
wire _abc_41234_new_n2732_; 
wire _abc_41234_new_n2733_; 
wire _abc_41234_new_n2734_; 
wire _abc_41234_new_n2735_; 
wire _abc_41234_new_n2736_; 
wire _abc_41234_new_n2737_; 
wire _abc_41234_new_n2738_; 
wire _abc_41234_new_n2739_; 
wire _abc_41234_new_n2740_; 
wire _abc_41234_new_n2741_; 
wire _abc_41234_new_n2742_; 
wire _abc_41234_new_n2743_; 
wire _abc_41234_new_n2744_; 
wire _abc_41234_new_n2745_; 
wire _abc_41234_new_n2746_; 
wire _abc_41234_new_n2747_; 
wire _abc_41234_new_n2748_; 
wire _abc_41234_new_n2749_; 
wire _abc_41234_new_n2750_; 
wire _abc_41234_new_n2751_; 
wire _abc_41234_new_n2752_; 
wire _abc_41234_new_n2753_; 
wire _abc_41234_new_n2754_; 
wire _abc_41234_new_n2755_; 
wire _abc_41234_new_n2756_; 
wire _abc_41234_new_n2757_; 
wire _abc_41234_new_n2758_; 
wire _abc_41234_new_n2759_; 
wire _abc_41234_new_n2760_; 
wire _abc_41234_new_n2761_; 
wire _abc_41234_new_n2762_; 
wire _abc_41234_new_n2764_; 
wire _abc_41234_new_n2765_; 
wire _abc_41234_new_n2766_; 
wire _abc_41234_new_n2767_; 
wire _abc_41234_new_n2768_; 
wire _abc_41234_new_n2769_; 
wire _abc_41234_new_n2770_; 
wire _abc_41234_new_n2771_; 
wire _abc_41234_new_n2772_; 
wire _abc_41234_new_n2773_; 
wire _abc_41234_new_n2774_; 
wire _abc_41234_new_n2775_; 
wire _abc_41234_new_n2776_; 
wire _abc_41234_new_n2777_; 
wire _abc_41234_new_n2778_; 
wire _abc_41234_new_n2779_; 
wire _abc_41234_new_n2780_; 
wire _abc_41234_new_n2781_; 
wire _abc_41234_new_n2782_; 
wire _abc_41234_new_n2783_; 
wire _abc_41234_new_n2784_; 
wire _abc_41234_new_n2785_; 
wire _abc_41234_new_n2786_; 
wire _abc_41234_new_n2787_; 
wire _abc_41234_new_n2788_; 
wire _abc_41234_new_n2789_; 
wire _abc_41234_new_n2790_; 
wire _abc_41234_new_n2792_; 
wire _abc_41234_new_n2793_; 
wire _abc_41234_new_n2794_; 
wire _abc_41234_new_n2795_; 
wire _abc_41234_new_n2796_; 
wire _abc_41234_new_n2797_; 
wire _abc_41234_new_n2798_; 
wire _abc_41234_new_n2799_; 
wire _abc_41234_new_n2800_; 
wire _abc_41234_new_n2801_; 
wire _abc_41234_new_n2802_; 
wire _abc_41234_new_n2803_; 
wire _abc_41234_new_n2804_; 
wire _abc_41234_new_n2805_; 
wire _abc_41234_new_n2806_; 
wire _abc_41234_new_n2807_; 
wire _abc_41234_new_n2808_; 
wire _abc_41234_new_n2809_; 
wire _abc_41234_new_n2810_; 
wire _abc_41234_new_n2811_; 
wire _abc_41234_new_n2812_; 
wire _abc_41234_new_n2813_; 
wire _abc_41234_new_n2814_; 
wire _abc_41234_new_n2815_; 
wire _abc_41234_new_n2816_; 
wire _abc_41234_new_n2817_; 
wire _abc_41234_new_n2818_; 
wire _abc_41234_new_n2819_; 
wire _abc_41234_new_n2820_; 
wire _abc_41234_new_n2821_; 
wire _abc_41234_new_n2822_; 
wire _abc_41234_new_n2824_; 
wire _abc_41234_new_n2825_; 
wire _abc_41234_new_n2826_; 
wire _abc_41234_new_n2827_; 
wire _abc_41234_new_n2828_; 
wire _abc_41234_new_n2829_; 
wire _abc_41234_new_n2830_; 
wire _abc_41234_new_n2831_; 
wire _abc_41234_new_n2832_; 
wire _abc_41234_new_n2833_; 
wire _abc_41234_new_n2834_; 
wire _abc_41234_new_n2835_; 
wire _abc_41234_new_n2836_; 
wire _abc_41234_new_n2837_; 
wire _abc_41234_new_n2838_; 
wire _abc_41234_new_n2839_; 
wire _abc_41234_new_n2840_; 
wire _abc_41234_new_n2841_; 
wire _abc_41234_new_n2842_; 
wire _abc_41234_new_n2843_; 
wire _abc_41234_new_n2844_; 
wire _abc_41234_new_n2845_; 
wire _abc_41234_new_n2846_; 
wire _abc_41234_new_n2847_; 
wire _abc_41234_new_n2848_; 
wire _abc_41234_new_n2849_; 
wire _abc_41234_new_n2851_; 
wire _abc_41234_new_n2852_; 
wire _abc_41234_new_n2853_; 
wire _abc_41234_new_n2854_; 
wire _abc_41234_new_n2855_; 
wire _abc_41234_new_n2856_; 
wire _abc_41234_new_n2857_; 
wire _abc_41234_new_n2858_; 
wire _abc_41234_new_n2859_; 
wire _abc_41234_new_n2860_; 
wire _abc_41234_new_n2861_; 
wire _abc_41234_new_n2862_; 
wire _abc_41234_new_n2863_; 
wire _abc_41234_new_n2864_; 
wire _abc_41234_new_n2865_; 
wire _abc_41234_new_n2866_; 
wire _abc_41234_new_n2867_; 
wire _abc_41234_new_n2868_; 
wire _abc_41234_new_n2869_; 
wire _abc_41234_new_n2870_; 
wire _abc_41234_new_n2871_; 
wire _abc_41234_new_n2872_; 
wire _abc_41234_new_n2873_; 
wire _abc_41234_new_n2874_; 
wire _abc_41234_new_n2875_; 
wire _abc_41234_new_n2876_; 
wire _abc_41234_new_n2877_; 
wire _abc_41234_new_n2878_; 
wire _abc_41234_new_n2879_; 
wire _abc_41234_new_n2881_; 
wire _abc_41234_new_n2882_; 
wire _abc_41234_new_n2883_; 
wire _abc_41234_new_n2884_; 
wire _abc_41234_new_n2885_; 
wire _abc_41234_new_n2886_; 
wire _abc_41234_new_n2887_; 
wire _abc_41234_new_n2888_; 
wire _abc_41234_new_n2889_; 
wire _abc_41234_new_n2890_; 
wire _abc_41234_new_n2891_; 
wire _abc_41234_new_n2892_; 
wire _abc_41234_new_n2893_; 
wire _abc_41234_new_n2894_; 
wire _abc_41234_new_n2895_; 
wire _abc_41234_new_n2896_; 
wire _abc_41234_new_n2897_; 
wire _abc_41234_new_n2898_; 
wire _abc_41234_new_n2899_; 
wire _abc_41234_new_n2900_; 
wire _abc_41234_new_n2901_; 
wire _abc_41234_new_n2902_; 
wire _abc_41234_new_n2903_; 
wire _abc_41234_new_n2904_; 
wire _abc_41234_new_n2905_; 
wire _abc_41234_new_n2906_; 
wire _abc_41234_new_n2907_; 
wire _abc_41234_new_n2908_; 
wire _abc_41234_new_n2910_; 
wire _abc_41234_new_n2911_; 
wire _abc_41234_new_n2912_; 
wire _abc_41234_new_n2913_; 
wire _abc_41234_new_n2914_; 
wire _abc_41234_new_n2915_; 
wire _abc_41234_new_n2916_; 
wire _abc_41234_new_n2917_; 
wire _abc_41234_new_n2918_; 
wire _abc_41234_new_n2919_; 
wire _abc_41234_new_n2919__bF_buf0; 
wire _abc_41234_new_n2919__bF_buf1; 
wire _abc_41234_new_n2919__bF_buf2; 
wire _abc_41234_new_n2919__bF_buf3; 
wire _abc_41234_new_n2920_; 
wire _abc_41234_new_n2921_; 
wire _abc_41234_new_n2922_; 
wire _abc_41234_new_n2923_; 
wire _abc_41234_new_n2924_; 
wire _abc_41234_new_n2925_; 
wire _abc_41234_new_n2926_; 
wire _abc_41234_new_n2927_; 
wire _abc_41234_new_n2928_; 
wire _abc_41234_new_n2929_; 
wire _abc_41234_new_n2930_; 
wire _abc_41234_new_n2931_; 
wire _abc_41234_new_n2932_; 
wire _abc_41234_new_n2933_; 
wire _abc_41234_new_n2934_; 
wire _abc_41234_new_n2935_; 
wire _abc_41234_new_n2936_; 
wire _abc_41234_new_n2937_; 
wire _abc_41234_new_n2938_; 
wire _abc_41234_new_n2939_; 
wire _abc_41234_new_n2940_; 
wire _abc_41234_new_n2941_; 
wire _abc_41234_new_n2942_; 
wire _abc_41234_new_n2942__bF_buf0; 
wire _abc_41234_new_n2942__bF_buf1; 
wire _abc_41234_new_n2942__bF_buf2; 
wire _abc_41234_new_n2942__bF_buf3; 
wire _abc_41234_new_n2943_; 
wire _abc_41234_new_n2944_; 
wire _abc_41234_new_n2945_; 
wire _abc_41234_new_n2946_; 
wire _abc_41234_new_n2947_; 
wire _abc_41234_new_n2947__bF_buf0; 
wire _abc_41234_new_n2947__bF_buf1; 
wire _abc_41234_new_n2947__bF_buf2; 
wire _abc_41234_new_n2947__bF_buf3; 
wire _abc_41234_new_n2948_; 
wire _abc_41234_new_n2949_; 
wire _abc_41234_new_n2950_; 
wire _abc_41234_new_n2951_; 
wire _abc_41234_new_n2951__bF_buf0; 
wire _abc_41234_new_n2951__bF_buf1; 
wire _abc_41234_new_n2951__bF_buf2; 
wire _abc_41234_new_n2951__bF_buf3; 
wire _abc_41234_new_n2952_; 
wire _abc_41234_new_n2953_; 
wire _abc_41234_new_n2954_; 
wire _abc_41234_new_n2955_; 
wire _abc_41234_new_n2956_; 
wire _abc_41234_new_n2957_; 
wire _abc_41234_new_n2958_; 
wire _abc_41234_new_n2959_; 
wire _abc_41234_new_n2959__bF_buf0; 
wire _abc_41234_new_n2959__bF_buf1; 
wire _abc_41234_new_n2959__bF_buf2; 
wire _abc_41234_new_n2959__bF_buf3; 
wire _abc_41234_new_n2960_; 
wire _abc_41234_new_n2961_; 
wire _abc_41234_new_n2963_; 
wire _abc_41234_new_n2964_; 
wire _abc_41234_new_n2965_; 
wire _abc_41234_new_n2966_; 
wire _abc_41234_new_n2967_; 
wire _abc_41234_new_n2968_; 
wire _abc_41234_new_n2969_; 
wire _abc_41234_new_n2970_; 
wire _abc_41234_new_n2971_; 
wire _abc_41234_new_n2972_; 
wire _abc_41234_new_n2973_; 
wire _abc_41234_new_n2974_; 
wire _abc_41234_new_n2975_; 
wire _abc_41234_new_n2976_; 
wire _abc_41234_new_n2977_; 
wire _abc_41234_new_n2978_; 
wire _abc_41234_new_n2979_; 
wire _abc_41234_new_n2980_; 
wire _abc_41234_new_n2981_; 
wire _abc_41234_new_n2982_; 
wire _abc_41234_new_n2983_; 
wire _abc_41234_new_n2984_; 
wire _abc_41234_new_n2985_; 
wire _abc_41234_new_n2986_; 
wire _abc_41234_new_n2987_; 
wire _abc_41234_new_n2988_; 
wire _abc_41234_new_n2989_; 
wire _abc_41234_new_n2990_; 
wire _abc_41234_new_n2991_; 
wire _abc_41234_new_n2993_; 
wire _abc_41234_new_n2994_; 
wire _abc_41234_new_n2995_; 
wire _abc_41234_new_n2996_; 
wire _abc_41234_new_n2997_; 
wire _abc_41234_new_n2998_; 
wire _abc_41234_new_n2999_; 
wire _abc_41234_new_n3000_; 
wire _abc_41234_new_n3001_; 
wire _abc_41234_new_n3002_; 
wire _abc_41234_new_n3003_; 
wire _abc_41234_new_n3004_; 
wire _abc_41234_new_n3005_; 
wire _abc_41234_new_n3006_; 
wire _abc_41234_new_n3007_; 
wire _abc_41234_new_n3008_; 
wire _abc_41234_new_n3009_; 
wire _abc_41234_new_n3010_; 
wire _abc_41234_new_n3011_; 
wire _abc_41234_new_n3012_; 
wire _abc_41234_new_n3013_; 
wire _abc_41234_new_n3014_; 
wire _abc_41234_new_n3015_; 
wire _abc_41234_new_n3016_; 
wire _abc_41234_new_n3017_; 
wire _abc_41234_new_n3018_; 
wire _abc_41234_new_n3019_; 
wire _abc_41234_new_n3020_; 
wire _abc_41234_new_n3021_; 
wire _abc_41234_new_n3023_; 
wire _abc_41234_new_n3024_; 
wire _abc_41234_new_n3025_; 
wire _abc_41234_new_n3026_; 
wire _abc_41234_new_n3027_; 
wire _abc_41234_new_n3028_; 
wire _abc_41234_new_n3029_; 
wire _abc_41234_new_n3030_; 
wire _abc_41234_new_n3031_; 
wire _abc_41234_new_n3032_; 
wire _abc_41234_new_n3033_; 
wire _abc_41234_new_n3034_; 
wire _abc_41234_new_n3035_; 
wire _abc_41234_new_n3036_; 
wire _abc_41234_new_n3037_; 
wire _abc_41234_new_n3038_; 
wire _abc_41234_new_n3039_; 
wire _abc_41234_new_n3040_; 
wire _abc_41234_new_n3041_; 
wire _abc_41234_new_n3042_; 
wire _abc_41234_new_n3043_; 
wire _abc_41234_new_n3044_; 
wire _abc_41234_new_n3045_; 
wire _abc_41234_new_n3046_; 
wire _abc_41234_new_n3047_; 
wire _abc_41234_new_n3049_; 
wire _abc_41234_new_n3050_; 
wire _abc_41234_new_n3051_; 
wire _abc_41234_new_n3052_; 
wire _abc_41234_new_n3053_; 
wire _abc_41234_new_n3054_; 
wire _abc_41234_new_n3055_; 
wire _abc_41234_new_n3056_; 
wire _abc_41234_new_n3057_; 
wire _abc_41234_new_n3058_; 
wire _abc_41234_new_n3059_; 
wire _abc_41234_new_n3060_; 
wire _abc_41234_new_n3061_; 
wire _abc_41234_new_n3062_; 
wire _abc_41234_new_n3063_; 
wire _abc_41234_new_n3064_; 
wire _abc_41234_new_n3065_; 
wire _abc_41234_new_n3066_; 
wire _abc_41234_new_n3067_; 
wire _abc_41234_new_n3068_; 
wire _abc_41234_new_n3069_; 
wire _abc_41234_new_n3070_; 
wire _abc_41234_new_n3071_; 
wire _abc_41234_new_n3072_; 
wire _abc_41234_new_n3074_; 
wire _abc_41234_new_n3075_; 
wire _abc_41234_new_n3076_; 
wire _abc_41234_new_n3077_; 
wire _abc_41234_new_n3078_; 
wire _abc_41234_new_n3079_; 
wire _abc_41234_new_n3080_; 
wire _abc_41234_new_n3081_; 
wire _abc_41234_new_n3082_; 
wire _abc_41234_new_n3083_; 
wire _abc_41234_new_n3084_; 
wire _abc_41234_new_n3085_; 
wire _abc_41234_new_n3086_; 
wire _abc_41234_new_n3087_; 
wire _abc_41234_new_n3088_; 
wire _abc_41234_new_n3089_; 
wire _abc_41234_new_n3090_; 
wire _abc_41234_new_n3091_; 
wire _abc_41234_new_n3092_; 
wire _abc_41234_new_n3093_; 
wire _abc_41234_new_n3094_; 
wire _abc_41234_new_n3095_; 
wire _abc_41234_new_n3096_; 
wire _abc_41234_new_n3097_; 
wire _abc_41234_new_n3098_; 
wire _abc_41234_new_n3099_; 
wire _abc_41234_new_n3101_; 
wire _abc_41234_new_n3102_; 
wire _abc_41234_new_n3103_; 
wire _abc_41234_new_n3104_; 
wire _abc_41234_new_n3105_; 
wire _abc_41234_new_n3106_; 
wire _abc_41234_new_n3107_; 
wire _abc_41234_new_n3108_; 
wire _abc_41234_new_n3109_; 
wire _abc_41234_new_n3110_; 
wire _abc_41234_new_n3111_; 
wire _abc_41234_new_n3112_; 
wire _abc_41234_new_n3113_; 
wire _abc_41234_new_n3114_; 
wire _abc_41234_new_n3115_; 
wire _abc_41234_new_n3116_; 
wire _abc_41234_new_n3117_; 
wire _abc_41234_new_n3118_; 
wire _abc_41234_new_n3119_; 
wire _abc_41234_new_n3120_; 
wire _abc_41234_new_n3121_; 
wire _abc_41234_new_n3122_; 
wire _abc_41234_new_n3123_; 
wire _abc_41234_new_n3125_; 
wire _abc_41234_new_n3126_; 
wire _abc_41234_new_n3127_; 
wire _abc_41234_new_n3128_; 
wire _abc_41234_new_n3129_; 
wire _abc_41234_new_n3130_; 
wire _abc_41234_new_n3131_; 
wire _abc_41234_new_n3132_; 
wire _abc_41234_new_n3133_; 
wire _abc_41234_new_n3134_; 
wire _abc_41234_new_n3135_; 
wire _abc_41234_new_n3136_; 
wire _abc_41234_new_n3137_; 
wire _abc_41234_new_n3138_; 
wire _abc_41234_new_n3139_; 
wire _abc_41234_new_n3140_; 
wire _abc_41234_new_n3141_; 
wire _abc_41234_new_n3142_; 
wire _abc_41234_new_n3143_; 
wire _abc_41234_new_n3144_; 
wire _abc_41234_new_n3145_; 
wire _abc_41234_new_n3146_; 
wire _abc_41234_new_n3147_; 
wire _abc_41234_new_n3148_; 
wire _abc_41234_new_n3149_; 
wire _abc_41234_new_n3151_; 
wire _abc_41234_new_n3152_; 
wire _abc_41234_new_n3153_; 
wire _abc_41234_new_n3154_; 
wire _abc_41234_new_n3155_; 
wire _abc_41234_new_n3156_; 
wire _abc_41234_new_n3157_; 
wire _abc_41234_new_n3158_; 
wire _abc_41234_new_n3159_; 
wire _abc_41234_new_n3160_; 
wire _abc_41234_new_n3161_; 
wire _abc_41234_new_n3162_; 
wire _abc_41234_new_n3163_; 
wire _abc_41234_new_n3164_; 
wire _abc_41234_new_n3165_; 
wire _abc_41234_new_n3166_; 
wire _abc_41234_new_n3167_; 
wire _abc_41234_new_n3168_; 
wire _abc_41234_new_n3169_; 
wire _abc_41234_new_n3170_; 
wire _abc_41234_new_n3171_; 
wire _abc_41234_new_n3172_; 
wire _abc_41234_new_n3173_; 
wire _abc_41234_new_n3175_; 
wire _abc_41234_new_n3176_; 
wire _abc_41234_new_n3177_; 
wire _abc_41234_new_n3178_; 
wire _abc_41234_new_n3179_; 
wire _abc_41234_new_n3180_; 
wire _abc_41234_new_n3181_; 
wire _abc_41234_new_n3182_; 
wire _abc_41234_new_n3183_; 
wire _abc_41234_new_n3184_; 
wire _abc_41234_new_n3185_; 
wire _abc_41234_new_n3186_; 
wire _abc_41234_new_n3187_; 
wire _abc_41234_new_n3188_; 
wire _abc_41234_new_n3189_; 
wire _abc_41234_new_n3190_; 
wire _abc_41234_new_n3191_; 
wire _abc_41234_new_n3192_; 
wire _abc_41234_new_n3193_; 
wire _abc_41234_new_n3194_; 
wire _abc_41234_new_n3195_; 
wire _abc_41234_new_n3196_; 
wire _abc_41234_new_n3197_; 
wire _abc_41234_new_n3198_; 
wire _abc_41234_new_n3200_; 
wire _abc_41234_new_n3201_; 
wire _abc_41234_new_n3202_; 
wire _abc_41234_new_n3203_; 
wire _abc_41234_new_n3204_; 
wire _abc_41234_new_n3205_; 
wire _abc_41234_new_n3206_; 
wire _abc_41234_new_n3207_; 
wire _abc_41234_new_n3208_; 
wire _abc_41234_new_n3209_; 
wire _abc_41234_new_n3210_; 
wire _abc_41234_new_n3211_; 
wire _abc_41234_new_n3212_; 
wire _abc_41234_new_n3213_; 
wire _abc_41234_new_n3214_; 
wire _abc_41234_new_n3215_; 
wire _abc_41234_new_n3216_; 
wire _abc_41234_new_n3217_; 
wire _abc_41234_new_n3218_; 
wire _abc_41234_new_n3219_; 
wire _abc_41234_new_n3220_; 
wire _abc_41234_new_n3221_; 
wire _abc_41234_new_n3222_; 
wire _abc_41234_new_n3223_; 
wire _abc_41234_new_n3225_; 
wire _abc_41234_new_n3226_; 
wire _abc_41234_new_n3227_; 
wire _abc_41234_new_n3228_; 
wire _abc_41234_new_n3229_; 
wire _abc_41234_new_n3230_; 
wire _abc_41234_new_n3231_; 
wire _abc_41234_new_n3232_; 
wire _abc_41234_new_n3233_; 
wire _abc_41234_new_n3234_; 
wire _abc_41234_new_n3235_; 
wire _abc_41234_new_n3236_; 
wire _abc_41234_new_n3237_; 
wire _abc_41234_new_n3238_; 
wire _abc_41234_new_n3239_; 
wire _abc_41234_new_n3240_; 
wire _abc_41234_new_n3241_; 
wire _abc_41234_new_n3242_; 
wire _abc_41234_new_n3243_; 
wire _abc_41234_new_n3244_; 
wire _abc_41234_new_n3245_; 
wire _abc_41234_new_n3246_; 
wire _abc_41234_new_n3248_; 
wire _abc_41234_new_n3249_; 
wire _abc_41234_new_n3250_; 
wire _abc_41234_new_n3251_; 
wire _abc_41234_new_n3252_; 
wire _abc_41234_new_n3253_; 
wire _abc_41234_new_n3254_; 
wire _abc_41234_new_n3255_; 
wire _abc_41234_new_n3256_; 
wire _abc_41234_new_n3257_; 
wire _abc_41234_new_n3258_; 
wire _abc_41234_new_n3259_; 
wire _abc_41234_new_n3260_; 
wire _abc_41234_new_n3261_; 
wire _abc_41234_new_n3262_; 
wire _abc_41234_new_n3263_; 
wire _abc_41234_new_n3264_; 
wire _abc_41234_new_n3265_; 
wire _abc_41234_new_n3266_; 
wire _abc_41234_new_n3267_; 
wire _abc_41234_new_n3268_; 
wire _abc_41234_new_n3269_; 
wire _abc_41234_new_n3270_; 
wire _abc_41234_new_n3272_; 
wire _abc_41234_new_n3273_; 
wire _abc_41234_new_n3274_; 
wire _abc_41234_new_n3275_; 
wire _abc_41234_new_n3276_; 
wire _abc_41234_new_n3277_; 
wire _abc_41234_new_n3278_; 
wire _abc_41234_new_n3279_; 
wire _abc_41234_new_n3280_; 
wire _abc_41234_new_n3281_; 
wire _abc_41234_new_n3282_; 
wire _abc_41234_new_n3283_; 
wire _abc_41234_new_n3284_; 
wire _abc_41234_new_n3285_; 
wire _abc_41234_new_n3286_; 
wire _abc_41234_new_n3287_; 
wire _abc_41234_new_n3288_; 
wire _abc_41234_new_n3289_; 
wire _abc_41234_new_n3290_; 
wire _abc_41234_new_n3291_; 
wire _abc_41234_new_n3292_; 
wire _abc_41234_new_n3294_; 
wire _abc_41234_new_n3295_; 
wire _abc_41234_new_n3296_; 
wire _abc_41234_new_n3297_; 
wire _abc_41234_new_n3298_; 
wire _abc_41234_new_n3299_; 
wire _abc_41234_new_n3300_; 
wire _abc_41234_new_n3301_; 
wire _abc_41234_new_n3302_; 
wire _abc_41234_new_n3303_; 
wire _abc_41234_new_n3304_; 
wire _abc_41234_new_n3305_; 
wire _abc_41234_new_n3306_; 
wire _abc_41234_new_n3307_; 
wire _abc_41234_new_n3308_; 
wire _abc_41234_new_n3309_; 
wire _abc_41234_new_n3310_; 
wire _abc_41234_new_n3311_; 
wire _abc_41234_new_n3312_; 
wire _abc_41234_new_n3313_; 
wire _abc_41234_new_n3314_; 
wire _abc_41234_new_n3316_; 
wire _abc_41234_new_n3317_; 
wire _abc_41234_new_n3318_; 
wire _abc_41234_new_n3319_; 
wire _abc_41234_new_n3320_; 
wire _abc_41234_new_n3321_; 
wire _abc_41234_new_n3322_; 
wire _abc_41234_new_n3323_; 
wire _abc_41234_new_n3324_; 
wire _abc_41234_new_n3325_; 
wire _abc_41234_new_n3326_; 
wire _abc_41234_new_n3327_; 
wire _abc_41234_new_n3328_; 
wire _abc_41234_new_n3329_; 
wire _abc_41234_new_n3330_; 
wire _abc_41234_new_n3331_; 
wire _abc_41234_new_n3332_; 
wire _abc_41234_new_n3333_; 
wire _abc_41234_new_n3334_; 
wire _abc_41234_new_n3335_; 
wire _abc_41234_new_n3337_; 
wire _abc_41234_new_n3338_; 
wire _abc_41234_new_n3339_; 
wire _abc_41234_new_n3340_; 
wire _abc_41234_new_n3341_; 
wire _abc_41234_new_n3342_; 
wire _abc_41234_new_n3343_; 
wire _abc_41234_new_n3344_; 
wire _abc_41234_new_n3345_; 
wire _abc_41234_new_n3346_; 
wire _abc_41234_new_n3347_; 
wire _abc_41234_new_n3348_; 
wire _abc_41234_new_n3349_; 
wire _abc_41234_new_n3350_; 
wire _abc_41234_new_n3351_; 
wire _abc_41234_new_n3352_; 
wire _abc_41234_new_n3353_; 
wire _abc_41234_new_n3354_; 
wire _abc_41234_new_n3355_; 
wire _abc_41234_new_n3356_; 
wire _abc_41234_new_n3358_; 
wire _abc_41234_new_n3359_; 
wire _abc_41234_new_n3360_; 
wire _abc_41234_new_n3361_; 
wire _abc_41234_new_n3362_; 
wire _abc_41234_new_n3363_; 
wire _abc_41234_new_n3364_; 
wire _abc_41234_new_n3365_; 
wire _abc_41234_new_n3366_; 
wire _abc_41234_new_n3367_; 
wire _abc_41234_new_n3368_; 
wire _abc_41234_new_n3369_; 
wire _abc_41234_new_n3370_; 
wire _abc_41234_new_n3371_; 
wire _abc_41234_new_n3372_; 
wire _abc_41234_new_n3373_; 
wire _abc_41234_new_n3374_; 
wire _abc_41234_new_n3375_; 
wire _abc_41234_new_n3376_; 
wire _abc_41234_new_n3377_; 
wire _abc_41234_new_n3378_; 
wire _abc_41234_new_n3379_; 
wire _abc_41234_new_n3381_; 
wire _abc_41234_new_n3382_; 
wire _abc_41234_new_n3383_; 
wire _abc_41234_new_n3384_; 
wire _abc_41234_new_n3385_; 
wire _abc_41234_new_n3386_; 
wire _abc_41234_new_n3387_; 
wire _abc_41234_new_n3388_; 
wire _abc_41234_new_n3389_; 
wire _abc_41234_new_n3390_; 
wire _abc_41234_new_n3391_; 
wire _abc_41234_new_n3392_; 
wire _abc_41234_new_n3393_; 
wire _abc_41234_new_n3394_; 
wire _abc_41234_new_n3395_; 
wire _abc_41234_new_n3396_; 
wire _abc_41234_new_n3397_; 
wire _abc_41234_new_n3398_; 
wire _abc_41234_new_n3399_; 
wire _abc_41234_new_n3400_; 
wire _abc_41234_new_n3401_; 
wire _abc_41234_new_n3403_; 
wire _abc_41234_new_n3404_; 
wire _abc_41234_new_n3405_; 
wire _abc_41234_new_n3406_; 
wire _abc_41234_new_n3407_; 
wire _abc_41234_new_n3408_; 
wire _abc_41234_new_n3409_; 
wire _abc_41234_new_n3410_; 
wire _abc_41234_new_n3411_; 
wire _abc_41234_new_n3412_; 
wire _abc_41234_new_n3413_; 
wire _abc_41234_new_n3414_; 
wire _abc_41234_new_n3415_; 
wire _abc_41234_new_n3416_; 
wire _abc_41234_new_n3417_; 
wire _abc_41234_new_n3418_; 
wire _abc_41234_new_n3419_; 
wire _abc_41234_new_n3420_; 
wire _abc_41234_new_n3422_; 
wire _abc_41234_new_n3423_; 
wire _abc_41234_new_n3424_; 
wire _abc_41234_new_n3425_; 
wire _abc_41234_new_n3426_; 
wire _abc_41234_new_n3427_; 
wire _abc_41234_new_n3428_; 
wire _abc_41234_new_n3429_; 
wire _abc_41234_new_n3430_; 
wire _abc_41234_new_n3431_; 
wire _abc_41234_new_n3432_; 
wire _abc_41234_new_n3433_; 
wire _abc_41234_new_n3434_; 
wire _abc_41234_new_n3435_; 
wire _abc_41234_new_n3436_; 
wire _abc_41234_new_n3437_; 
wire _abc_41234_new_n3438_; 
wire _abc_41234_new_n3439_; 
wire _abc_41234_new_n3440_; 
wire _abc_41234_new_n3441_; 
wire _abc_41234_new_n3442_; 
wire _abc_41234_new_n3443_; 
wire _abc_41234_new_n3445_; 
wire _abc_41234_new_n3446_; 
wire _abc_41234_new_n3447_; 
wire _abc_41234_new_n3448_; 
wire _abc_41234_new_n3449_; 
wire _abc_41234_new_n3450_; 
wire _abc_41234_new_n3451_; 
wire _abc_41234_new_n3452_; 
wire _abc_41234_new_n3453_; 
wire _abc_41234_new_n3454_; 
wire _abc_41234_new_n3455_; 
wire _abc_41234_new_n3456_; 
wire _abc_41234_new_n3457_; 
wire _abc_41234_new_n3458_; 
wire _abc_41234_new_n3459_; 
wire _abc_41234_new_n3460_; 
wire _abc_41234_new_n3461_; 
wire _abc_41234_new_n3462_; 
wire _abc_41234_new_n3463_; 
wire _abc_41234_new_n3464_; 
wire _abc_41234_new_n3466_; 
wire _abc_41234_new_n3467_; 
wire _abc_41234_new_n3468_; 
wire _abc_41234_new_n3469_; 
wire _abc_41234_new_n3470_; 
wire _abc_41234_new_n3471_; 
wire _abc_41234_new_n3472_; 
wire _abc_41234_new_n3473_; 
wire _abc_41234_new_n3474_; 
wire _abc_41234_new_n3475_; 
wire _abc_41234_new_n3476_; 
wire _abc_41234_new_n3477_; 
wire _abc_41234_new_n3478_; 
wire _abc_41234_new_n3479_; 
wire _abc_41234_new_n3480_; 
wire _abc_41234_new_n3481_; 
wire _abc_41234_new_n3482_; 
wire _abc_41234_new_n3483_; 
wire _abc_41234_new_n3484_; 
wire _abc_41234_new_n3485_; 
wire _abc_41234_new_n3487_; 
wire _abc_41234_new_n3488_; 
wire _abc_41234_new_n3489_; 
wire _abc_41234_new_n3490_; 
wire _abc_41234_new_n3491_; 
wire _abc_41234_new_n3492_; 
wire _abc_41234_new_n3493_; 
wire _abc_41234_new_n3494_; 
wire _abc_41234_new_n3495_; 
wire _abc_41234_new_n3496_; 
wire _abc_41234_new_n3497_; 
wire _abc_41234_new_n3498_; 
wire _abc_41234_new_n3499_; 
wire _abc_41234_new_n3500_; 
wire _abc_41234_new_n3501_; 
wire _abc_41234_new_n3502_; 
wire _abc_41234_new_n3503_; 
wire _abc_41234_new_n3504_; 
wire _abc_41234_new_n3505_; 
wire _abc_41234_new_n3507_; 
wire _abc_41234_new_n3508_; 
wire _abc_41234_new_n3509_; 
wire _abc_41234_new_n3510_; 
wire _abc_41234_new_n3511_; 
wire _abc_41234_new_n3512_; 
wire _abc_41234_new_n3513_; 
wire _abc_41234_new_n3514_; 
wire _abc_41234_new_n3515_; 
wire _abc_41234_new_n3516_; 
wire _abc_41234_new_n3517_; 
wire _abc_41234_new_n3518_; 
wire _abc_41234_new_n3519_; 
wire _abc_41234_new_n3520_; 
wire _abc_41234_new_n3521_; 
wire _abc_41234_new_n3522_; 
wire _abc_41234_new_n3523_; 
wire _abc_41234_new_n3524_; 
wire _abc_41234_new_n3526_; 
wire _abc_41234_new_n3527_; 
wire _abc_41234_new_n3528_; 
wire _abc_41234_new_n3529_; 
wire _abc_41234_new_n3530_; 
wire _abc_41234_new_n3531_; 
wire _abc_41234_new_n3532_; 
wire _abc_41234_new_n3533_; 
wire _abc_41234_new_n3534_; 
wire _abc_41234_new_n3535_; 
wire _abc_41234_new_n3536_; 
wire _abc_41234_new_n3537_; 
wire _abc_41234_new_n3538_; 
wire _abc_41234_new_n3539_; 
wire _abc_41234_new_n3540_; 
wire _abc_41234_new_n3541_; 
wire _abc_41234_new_n3542_; 
wire _abc_41234_new_n3543_; 
wire _abc_41234_new_n3544_; 
wire _abc_41234_new_n3545_; 
wire _abc_41234_new_n3547_; 
wire _abc_41234_new_n3548_; 
wire _abc_41234_new_n3549_; 
wire _abc_41234_new_n3550_; 
wire _abc_41234_new_n3551_; 
wire _abc_41234_new_n3552_; 
wire _abc_41234_new_n3553_; 
wire _abc_41234_new_n3554_; 
wire _abc_41234_new_n3555_; 
wire _abc_41234_new_n3556_; 
wire _abc_41234_new_n3557_; 
wire _abc_41234_new_n3558_; 
wire _abc_41234_new_n3559_; 
wire _abc_41234_new_n3560_; 
wire _abc_41234_new_n3561_; 
wire _abc_41234_new_n3562_; 
wire _abc_41234_new_n3563_; 
wire _abc_41234_new_n3564_; 
wire _abc_41234_new_n3565_; 
wire _abc_41234_new_n3566_; 
wire _abc_41234_new_n3567_; 
wire _abc_41234_new_n3569_; 
wire _abc_41234_new_n3570_; 
wire _abc_41234_new_n3571_; 
wire _abc_41234_new_n3572_; 
wire _abc_41234_new_n3573_; 
wire _abc_41234_new_n3574_; 
wire _abc_41234_new_n3575_; 
wire _abc_41234_new_n3576_; 
wire _abc_41234_new_n3577_; 
wire _abc_41234_new_n3578_; 
wire _abc_41234_new_n3579_; 
wire _abc_41234_new_n3580_; 
wire _abc_41234_new_n3581_; 
wire _abc_41234_new_n3582_; 
wire _abc_41234_new_n3583_; 
wire _abc_41234_new_n3584_; 
wire _abc_41234_new_n3585_; 
wire _abc_41234_new_n3586_; 
wire _abc_41234_new_n3587_; 
wire _abc_41234_new_n3588_; 
wire _abc_41234_new_n3589_; 
wire _abc_41234_new_n3591_; 
wire _abc_41234_new_n3592_; 
wire _abc_41234_new_n3593_; 
wire _abc_41234_new_n3594_; 
wire _abc_41234_new_n3595_; 
wire _abc_41234_new_n3596_; 
wire _abc_41234_new_n3597_; 
wire _abc_41234_new_n3598_; 
wire _abc_41234_new_n3599_; 
wire _abc_41234_new_n3600_; 
wire _abc_41234_new_n3601_; 
wire _abc_41234_new_n3602_; 
wire _abc_41234_new_n3603_; 
wire _abc_41234_new_n3604_; 
wire _abc_41234_new_n3605_; 
wire _abc_41234_new_n3606_; 
wire _abc_41234_new_n3607_; 
wire _abc_41234_new_n3608_; 
wire _abc_41234_new_n3609_; 
wire _abc_41234_new_n3610_; 
wire _abc_41234_new_n3611_; 
wire _abc_41234_new_n3612_; 
wire _abc_41234_new_n3614_; 
wire _abc_41234_new_n3615_; 
wire _abc_41234_new_n3616_; 
wire _abc_41234_new_n3617_; 
wire _abc_41234_new_n3618_; 
wire _abc_41234_new_n3619_; 
wire _abc_41234_new_n3620_; 
wire _abc_41234_new_n3621_; 
wire _abc_41234_new_n3622_; 
wire _abc_41234_new_n3623_; 
wire _abc_41234_new_n3624_; 
wire _abc_41234_new_n3625_; 
wire _abc_41234_new_n3626_; 
wire _abc_41234_new_n3627_; 
wire _abc_41234_new_n3628_; 
wire _abc_41234_new_n3629_; 
wire _abc_41234_new_n3630_; 
wire _abc_41234_new_n3631_; 
wire _abc_41234_new_n3632_; 
wire _abc_41234_new_n3633_; 
wire _abc_41234_new_n3634_; 
wire _abc_41234_new_n3635_; 
wire _abc_41234_new_n3637_; 
wire _abc_41234_new_n3638_; 
wire _abc_41234_new_n3639_; 
wire _abc_41234_new_n3640_; 
wire _abc_41234_new_n3641_; 
wire _abc_41234_new_n3642_; 
wire _abc_41234_new_n3643_; 
wire _abc_41234_new_n3644_; 
wire _abc_41234_new_n3645_; 
wire _abc_41234_new_n3646_; 
wire _abc_41234_new_n3647_; 
wire _abc_41234_new_n3648_; 
wire _abc_41234_new_n3649_; 
wire _abc_41234_new_n3650_; 
wire _abc_41234_new_n3651_; 
wire _abc_41234_new_n3652_; 
wire _abc_41234_new_n3653_; 
wire _abc_41234_new_n3654_; 
wire _abc_41234_new_n3656_; 
wire _abc_41234_new_n3657_; 
wire _abc_41234_new_n3658_; 
wire _abc_41234_new_n3659_; 
wire _abc_41234_new_n3660_; 
wire _abc_41234_new_n3661_; 
wire _abc_41234_new_n3662_; 
wire _abc_41234_new_n3663_; 
wire _abc_41234_new_n3664_; 
wire _abc_41234_new_n3665_; 
wire _abc_41234_new_n3666_; 
wire _abc_41234_new_n3667_; 
wire _abc_41234_new_n3668_; 
wire _abc_41234_new_n3669_; 
wire _abc_41234_new_n3670_; 
wire _abc_41234_new_n3671_; 
wire _abc_41234_new_n3672_; 
wire _abc_41234_new_n3673_; 
wire _abc_41234_new_n3674_; 
wire _abc_41234_new_n3676_; 
wire _abc_41234_new_n3677_; 
wire _abc_41234_new_n3678_; 
wire _abc_41234_new_n3680_; 
wire _abc_41234_new_n3682_; 
wire _abc_41234_new_n3684_; 
wire _abc_41234_new_n3686_; 
wire _abc_41234_new_n3688_; 
wire _abc_41234_new_n3690_; 
wire _abc_41234_new_n3692_; 
wire _abc_41234_new_n3694_; 
wire _abc_41234_new_n3695_; 
wire _abc_41234_new_n3696_; 
wire _abc_41234_new_n3697_; 
wire _abc_41234_new_n3698_; 
wire _abc_41234_new_n3699_; 
wire _abc_41234_new_n3700_; 
wire _abc_41234_new_n3702_; 
wire _abc_41234_new_n3703_; 
wire _abc_41234_new_n3704_; 
wire _abc_41234_new_n3705_; 
wire _abc_41234_new_n3706_; 
wire _abc_41234_new_n3708_; 
wire _abc_41234_new_n3709_; 
wire _abc_41234_new_n3710_; 
wire _abc_41234_new_n3711_; 
wire _abc_41234_new_n3712_; 
wire _abc_41234_new_n3714_; 
wire _abc_41234_new_n3715_; 
wire _abc_41234_new_n3716_; 
wire _abc_41234_new_n3717_; 
wire _abc_41234_new_n3718_; 
wire _abc_41234_new_n3719_; 
wire _abc_41234_new_n3720_; 
wire _abc_41234_new_n3721_; 
wire _abc_41234_new_n3722_; 
wire _abc_41234_new_n3723_; 
wire _abc_41234_new_n3724_; 
wire _abc_41234_new_n3725_; 
wire _abc_41234_new_n3726_; 
wire _abc_41234_new_n3727_; 
wire _abc_41234_new_n3728_; 
wire _abc_41234_new_n3730_; 
wire _abc_41234_new_n3731_; 
wire _abc_41234_new_n3732_; 
wire _abc_41234_new_n3733_; 
wire _abc_41234_new_n3734_; 
wire _abc_41234_new_n3735_; 
wire _abc_41234_new_n3736_; 
wire _abc_41234_new_n3737_; 
wire _abc_41234_new_n3738_; 
wire _abc_41234_new_n3739_; 
wire _abc_41234_new_n3740_; 
wire _abc_41234_new_n3741_; 
wire _abc_41234_new_n3742_; 
wire _abc_41234_new_n3743_; 
wire _abc_41234_new_n3744_; 
wire _abc_41234_new_n3745_; 
wire _abc_41234_new_n3746_; 
wire _abc_41234_new_n3747_; 
wire _abc_41234_new_n3748_; 
wire _abc_41234_new_n3749_; 
wire _abc_41234_new_n3750_; 
wire _abc_41234_new_n3751_; 
wire _abc_41234_new_n3752_; 
wire _abc_41234_new_n3753_; 
wire _abc_41234_new_n3754_; 
wire _abc_41234_new_n3756_; 
wire _abc_41234_new_n3757_; 
wire _abc_41234_new_n3758_; 
wire _abc_41234_new_n3759_; 
wire _abc_41234_new_n3760_; 
wire _abc_41234_new_n3761_; 
wire _abc_41234_new_n3762_; 
wire _abc_41234_new_n3763_; 
wire _abc_41234_new_n3764_; 
wire _abc_41234_new_n3765_; 
wire _abc_41234_new_n3766_; 
wire _abc_41234_new_n3767_; 
wire _abc_41234_new_n3768_; 
wire _abc_41234_new_n3769_; 
wire _abc_41234_new_n3770_; 
wire _abc_41234_new_n3771_; 
wire _abc_41234_new_n3772_; 
wire _abc_41234_new_n3773_; 
wire _abc_41234_new_n3774_; 
wire _abc_41234_new_n3775_; 
wire _abc_41234_new_n3776_; 
wire _abc_41234_new_n3777_; 
wire _abc_41234_new_n3778_; 
wire _abc_41234_new_n3780_; 
wire _abc_41234_new_n3781_; 
wire _abc_41234_new_n3782_; 
wire _abc_41234_new_n3783_; 
wire _abc_41234_new_n3784_; 
wire _abc_41234_new_n3785_; 
wire _abc_41234_new_n3786_; 
wire _abc_41234_new_n3787_; 
wire _abc_41234_new_n3788_; 
wire _abc_41234_new_n3789_; 
wire _abc_41234_new_n3790_; 
wire _abc_41234_new_n3791_; 
wire _abc_41234_new_n3792_; 
wire _abc_41234_new_n3793_; 
wire _abc_41234_new_n3794_; 
wire _abc_41234_new_n3795_; 
wire _abc_41234_new_n3796_; 
wire _abc_41234_new_n3797_; 
wire _abc_41234_new_n3798_; 
wire _abc_41234_new_n3799_; 
wire _abc_41234_new_n3800_; 
wire _abc_41234_new_n3801_; 
wire _abc_41234_new_n3803_; 
wire _abc_41234_new_n3804_; 
wire _abc_41234_new_n3805_; 
wire _abc_41234_new_n3806_; 
wire _abc_41234_new_n3807_; 
wire _abc_41234_new_n3808_; 
wire _abc_41234_new_n3809_; 
wire _abc_41234_new_n3810_; 
wire _abc_41234_new_n3811_; 
wire _abc_41234_new_n3812_; 
wire _abc_41234_new_n3813_; 
wire _abc_41234_new_n3814_; 
wire _abc_41234_new_n3815_; 
wire _abc_41234_new_n3816_; 
wire _abc_41234_new_n3817_; 
wire _abc_41234_new_n3818_; 
wire _abc_41234_new_n3819_; 
wire _abc_41234_new_n3820_; 
wire _abc_41234_new_n3821_; 
wire _abc_41234_new_n3822_; 
wire _abc_41234_new_n3823_; 
wire _abc_41234_new_n3824_; 
wire _abc_41234_new_n3825_; 
wire _abc_41234_new_n3827_; 
wire _abc_41234_new_n3828_; 
wire _abc_41234_new_n3829_; 
wire _abc_41234_new_n3830_; 
wire _abc_41234_new_n3831_; 
wire _abc_41234_new_n3832_; 
wire _abc_41234_new_n3833_; 
wire _abc_41234_new_n3834_; 
wire _abc_41234_new_n3835_; 
wire _abc_41234_new_n3836_; 
wire _abc_41234_new_n3837_; 
wire _abc_41234_new_n3838_; 
wire _abc_41234_new_n3839_; 
wire _abc_41234_new_n3840_; 
wire _abc_41234_new_n3841_; 
wire _abc_41234_new_n3842_; 
wire _abc_41234_new_n3843_; 
wire _abc_41234_new_n3844_; 
wire _abc_41234_new_n3845_; 
wire _abc_41234_new_n3846_; 
wire _abc_41234_new_n3847_; 
wire _abc_41234_new_n3848_; 
wire _abc_41234_new_n3849_; 
wire _abc_41234_new_n3850_; 
wire _abc_41234_new_n3852_; 
wire _abc_41234_new_n3853_; 
wire _abc_41234_new_n3854_; 
wire _abc_41234_new_n3855_; 
wire _abc_41234_new_n3856_; 
wire _abc_41234_new_n3857_; 
wire _abc_41234_new_n3858_; 
wire _abc_41234_new_n3859_; 
wire _abc_41234_new_n3860_; 
wire _abc_41234_new_n3861_; 
wire _abc_41234_new_n3862_; 
wire _abc_41234_new_n3863_; 
wire _abc_41234_new_n3864_; 
wire _abc_41234_new_n3865_; 
wire _abc_41234_new_n3866_; 
wire _abc_41234_new_n3867_; 
wire _abc_41234_new_n3868_; 
wire _abc_41234_new_n3869_; 
wire _abc_41234_new_n3870_; 
wire _abc_41234_new_n3871_; 
wire _abc_41234_new_n3872_; 
wire _abc_41234_new_n3873_; 
wire _abc_41234_new_n3874_; 
wire _abc_41234_new_n3875_; 
wire _abc_41234_new_n3876_; 
wire _abc_41234_new_n3877_; 
wire _abc_41234_new_n3878_; 
wire _abc_41234_new_n3879_; 
wire _abc_41234_new_n3881_; 
wire _abc_41234_new_n3882_; 
wire _abc_41234_new_n3883_; 
wire _abc_41234_new_n3884_; 
wire _abc_41234_new_n3885_; 
wire _abc_41234_new_n3886_; 
wire _abc_41234_new_n3887_; 
wire _abc_41234_new_n3888_; 
wire _abc_41234_new_n3889_; 
wire _abc_41234_new_n3890_; 
wire _abc_41234_new_n3891_; 
wire _abc_41234_new_n3892_; 
wire _abc_41234_new_n3893_; 
wire _abc_41234_new_n3894_; 
wire _abc_41234_new_n3895_; 
wire _abc_41234_new_n3896_; 
wire _abc_41234_new_n3897_; 
wire _abc_41234_new_n3898_; 
wire _abc_41234_new_n3899_; 
wire _abc_41234_new_n3900_; 
wire _abc_41234_new_n3901_; 
wire _abc_41234_new_n3902_; 
wire _abc_41234_new_n3903_; 
wire _abc_41234_new_n3904_; 
wire _abc_41234_new_n3905_; 
wire _abc_41234_new_n3906_; 
wire _abc_41234_new_n3907_; 
wire _abc_41234_new_n3908_; 
wire _abc_41234_new_n3910_; 
wire _abc_41234_new_n3911_; 
wire _abc_41234_new_n3912_; 
wire _abc_41234_new_n3913_; 
wire _abc_41234_new_n3914_; 
wire _abc_41234_new_n3914__bF_buf0; 
wire _abc_41234_new_n3914__bF_buf1; 
wire _abc_41234_new_n3914__bF_buf2; 
wire _abc_41234_new_n3914__bF_buf3; 
wire _abc_41234_new_n3915_; 
wire _abc_41234_new_n3916_; 
wire _abc_41234_new_n3917_; 
wire _abc_41234_new_n3918_; 
wire _abc_41234_new_n3919_; 
wire _abc_41234_new_n3920_; 
wire _abc_41234_new_n3921_; 
wire _abc_41234_new_n3922_; 
wire _abc_41234_new_n3923_; 
wire _abc_41234_new_n3924_; 
wire _abc_41234_new_n3925_; 
wire _abc_41234_new_n3927_; 
wire _abc_41234_new_n3928_; 
wire _abc_41234_new_n3929_; 
wire _abc_41234_new_n3930_; 
wire _abc_41234_new_n3931_; 
wire _abc_41234_new_n3932_; 
wire _abc_41234_new_n3933_; 
wire _abc_41234_new_n3934_; 
wire _abc_41234_new_n3935_; 
wire _abc_41234_new_n3936_; 
wire _abc_41234_new_n3937_; 
wire _abc_41234_new_n3938_; 
wire _abc_41234_new_n3939_; 
wire _abc_41234_new_n3940_; 
wire _abc_41234_new_n3941_; 
wire _abc_41234_new_n3942_; 
wire _abc_41234_new_n3944_; 
wire _abc_41234_new_n3945_; 
wire _abc_41234_new_n3946_; 
wire _abc_41234_new_n3947_; 
wire _abc_41234_new_n3948_; 
wire _abc_41234_new_n3949_; 
wire _abc_41234_new_n3950_; 
wire _abc_41234_new_n3951_; 
wire _abc_41234_new_n3952_; 
wire _abc_41234_new_n3953_; 
wire _abc_41234_new_n3954_; 
wire _abc_41234_new_n3955_; 
wire _abc_41234_new_n3956_; 
wire _abc_41234_new_n3957_; 
wire _abc_41234_new_n3958_; 
wire _abc_41234_new_n3959_; 
wire _abc_41234_new_n3960_; 
wire _abc_41234_new_n3961_; 
wire _abc_41234_new_n3962_; 
wire _abc_41234_new_n3963_; 
wire _abc_41234_new_n3964_; 
wire _abc_41234_new_n3965_; 
wire _abc_41234_new_n3966_; 
wire _abc_41234_new_n3967_; 
wire _abc_41234_new_n3969_; 
wire _abc_41234_new_n3970_; 
wire _abc_41234_new_n3971_; 
wire _abc_41234_new_n3972_; 
wire _abc_41234_new_n3973_; 
wire _abc_41234_new_n3974_; 
wire _abc_41234_new_n3975_; 
wire _abc_41234_new_n3976_; 
wire _abc_41234_new_n3977_; 
wire _abc_41234_new_n3978_; 
wire _abc_41234_new_n3979_; 
wire _abc_41234_new_n3980_; 
wire _abc_41234_new_n3981_; 
wire _abc_41234_new_n3982_; 
wire _abc_41234_new_n3983_; 
wire _abc_41234_new_n3984_; 
wire _abc_41234_new_n3985_; 
wire _abc_41234_new_n3986_; 
wire _abc_41234_new_n3987_; 
wire _abc_41234_new_n3988_; 
wire _abc_41234_new_n3990_; 
wire _abc_41234_new_n3991_; 
wire _abc_41234_new_n3992_; 
wire _abc_41234_new_n3993_; 
wire _abc_41234_new_n3994_; 
wire _abc_41234_new_n3995_; 
wire _abc_41234_new_n3996_; 
wire _abc_41234_new_n3997_; 
wire _abc_41234_new_n3998_; 
wire _abc_41234_new_n3999_; 
wire _abc_41234_new_n4000_; 
wire _abc_41234_new_n4001_; 
wire _abc_41234_new_n4002_; 
wire _abc_41234_new_n4003_; 
wire _abc_41234_new_n4004_; 
wire _abc_41234_new_n4005_; 
wire _abc_41234_new_n4006_; 
wire _abc_41234_new_n4007_; 
wire _abc_41234_new_n4009_; 
wire _abc_41234_new_n4010_; 
wire _abc_41234_new_n4011_; 
wire _abc_41234_new_n4012_; 
wire _abc_41234_new_n4013_; 
wire _abc_41234_new_n4014_; 
wire _abc_41234_new_n4015_; 
wire _abc_41234_new_n4016_; 
wire _abc_41234_new_n4017_; 
wire _abc_41234_new_n4018_; 
wire _abc_41234_new_n4019_; 
wire _abc_41234_new_n4020_; 
wire _abc_41234_new_n4021_; 
wire _abc_41234_new_n4022_; 
wire _abc_41234_new_n4023_; 
wire _abc_41234_new_n4024_; 
wire _abc_41234_new_n4025_; 
wire _abc_41234_new_n4026_; 
wire _abc_41234_new_n4027_; 
wire _abc_41234_new_n4028_; 
wire _abc_41234_new_n4029_; 
wire _abc_41234_new_n4030_; 
wire _abc_41234_new_n4031_; 
wire _abc_41234_new_n4032_; 
wire _abc_41234_new_n4033_; 
wire _abc_41234_new_n4034_; 
wire _abc_41234_new_n4036_; 
wire _abc_41234_new_n4037_; 
wire _abc_41234_new_n4038_; 
wire _abc_41234_new_n4039_; 
wire _abc_41234_new_n4040_; 
wire _abc_41234_new_n4041_; 
wire _abc_41234_new_n4042_; 
wire _abc_41234_new_n4043_; 
wire _abc_41234_new_n4044_; 
wire _abc_41234_new_n4045_; 
wire _abc_41234_new_n4046_; 
wire _abc_41234_new_n4047_; 
wire _abc_41234_new_n4048_; 
wire _abc_41234_new_n4049_; 
wire _abc_41234_new_n4050_; 
wire _abc_41234_new_n4051_; 
wire _abc_41234_new_n4052_; 
wire _abc_41234_new_n4053_; 
wire _abc_41234_new_n4054_; 
wire _abc_41234_new_n4055_; 
wire _abc_41234_new_n4056_; 
wire _abc_41234_new_n4057_; 
wire _abc_41234_new_n4059_; 
wire _abc_41234_new_n4060_; 
wire _abc_41234_new_n4061_; 
wire _abc_41234_new_n4062_; 
wire _abc_41234_new_n4063_; 
wire _abc_41234_new_n4064_; 
wire _abc_41234_new_n4065_; 
wire _abc_41234_new_n4066_; 
wire _abc_41234_new_n4067_; 
wire _abc_41234_new_n4068_; 
wire _abc_41234_new_n4069_; 
wire _abc_41234_new_n4070_; 
wire _abc_41234_new_n4071_; 
wire _abc_41234_new_n4072_; 
wire _abc_41234_new_n4073_; 
wire _abc_41234_new_n4074_; 
wire _abc_41234_new_n4075_; 
wire _abc_41234_new_n4076_; 
wire _abc_41234_new_n4077_; 
wire _abc_41234_new_n4079_; 
wire _abc_41234_new_n4080_; 
wire _abc_41234_new_n4081_; 
wire _abc_41234_new_n4082_; 
wire _abc_41234_new_n4083_; 
wire _abc_41234_new_n4084_; 
wire _abc_41234_new_n4085_; 
wire _abc_41234_new_n4086_; 
wire _abc_41234_new_n4087_; 
wire _abc_41234_new_n4088_; 
wire _abc_41234_new_n4089_; 
wire _abc_41234_new_n4090_; 
wire _abc_41234_new_n4091_; 
wire _abc_41234_new_n4092_; 
wire _abc_41234_new_n4093_; 
wire _abc_41234_new_n4094_; 
wire _abc_41234_new_n4095_; 
wire _abc_41234_new_n4096_; 
wire _abc_41234_new_n4097_; 
wire _abc_41234_new_n4098_; 
wire _abc_41234_new_n4099_; 
wire _abc_41234_new_n4101_; 
wire _abc_41234_new_n4102_; 
wire _abc_41234_new_n4103_; 
wire _abc_41234_new_n4104_; 
wire _abc_41234_new_n4105_; 
wire _abc_41234_new_n4106_; 
wire _abc_41234_new_n4107_; 
wire _abc_41234_new_n4108_; 
wire _abc_41234_new_n4109_; 
wire _abc_41234_new_n4110_; 
wire _abc_41234_new_n4111_; 
wire _abc_41234_new_n4112_; 
wire _abc_41234_new_n4113_; 
wire _abc_41234_new_n4114_; 
wire _abc_41234_new_n4115_; 
wire _abc_41234_new_n4116_; 
wire _abc_41234_new_n4117_; 
wire _abc_41234_new_n4118_; 
wire _abc_41234_new_n4119_; 
wire _abc_41234_new_n4120_; 
wire _abc_41234_new_n4121_; 
wire _abc_41234_new_n4123_; 
wire _abc_41234_new_n4124_; 
wire _abc_41234_new_n4125_; 
wire _abc_41234_new_n4126_; 
wire _abc_41234_new_n4127_; 
wire _abc_41234_new_n4128_; 
wire _abc_41234_new_n4129_; 
wire _abc_41234_new_n4130_; 
wire _abc_41234_new_n4131_; 
wire _abc_41234_new_n4132_; 
wire _abc_41234_new_n4133_; 
wire _abc_41234_new_n4134_; 
wire _abc_41234_new_n4135_; 
wire _abc_41234_new_n4136_; 
wire _abc_41234_new_n4137_; 
wire _abc_41234_new_n4138_; 
wire _abc_41234_new_n4139_; 
wire _abc_41234_new_n4140_; 
wire _abc_41234_new_n4141_; 
wire _abc_41234_new_n4142_; 
wire _abc_41234_new_n4143_; 
wire _abc_41234_new_n4144_; 
wire _abc_41234_new_n4146_; 
wire _abc_41234_new_n4147_; 
wire _abc_41234_new_n4148_; 
wire _abc_41234_new_n4149_; 
wire _abc_41234_new_n4150_; 
wire _abc_41234_new_n4151_; 
wire _abc_41234_new_n4152_; 
wire _abc_41234_new_n4153_; 
wire _abc_41234_new_n4154_; 
wire _abc_41234_new_n4155_; 
wire _abc_41234_new_n4156_; 
wire _abc_41234_new_n4157_; 
wire _abc_41234_new_n4158_; 
wire _abc_41234_new_n4159_; 
wire _abc_41234_new_n4160_; 
wire _abc_41234_new_n4161_; 
wire _abc_41234_new_n4162_; 
wire _abc_41234_new_n4163_; 
wire _abc_41234_new_n4164_; 
wire _abc_41234_new_n4165_; 
wire _abc_41234_new_n4166_; 
wire _abc_41234_new_n4167_; 
wire _abc_41234_new_n4169_; 
wire _abc_41234_new_n4170_; 
wire _abc_41234_new_n4171_; 
wire _abc_41234_new_n4172_; 
wire _abc_41234_new_n4173_; 
wire _abc_41234_new_n4174_; 
wire _abc_41234_new_n4175_; 
wire _abc_41234_new_n4176_; 
wire _abc_41234_new_n4177_; 
wire _abc_41234_new_n4178_; 
wire _abc_41234_new_n4179_; 
wire _abc_41234_new_n4180_; 
wire _abc_41234_new_n4181_; 
wire _abc_41234_new_n4182_; 
wire _abc_41234_new_n4183_; 
wire _abc_41234_new_n4184_; 
wire _abc_41234_new_n4185_; 
wire _abc_41234_new_n4186_; 
wire _abc_41234_new_n4187_; 
wire _abc_41234_new_n4189_; 
wire _abc_41234_new_n4190_; 
wire _abc_41234_new_n4191_; 
wire _abc_41234_new_n4192_; 
wire _abc_41234_new_n4193_; 
wire _abc_41234_new_n4194_; 
wire _abc_41234_new_n4195_; 
wire _abc_41234_new_n4196_; 
wire _abc_41234_new_n4197_; 
wire _abc_41234_new_n4198_; 
wire _abc_41234_new_n4199_; 
wire _abc_41234_new_n4200_; 
wire _abc_41234_new_n4201_; 
wire _abc_41234_new_n4202_; 
wire _abc_41234_new_n4203_; 
wire _abc_41234_new_n4204_; 
wire _abc_41234_new_n4205_; 
wire _abc_41234_new_n4206_; 
wire _abc_41234_new_n4207_; 
wire _abc_41234_new_n4208_; 
wire _abc_41234_new_n4210_; 
wire _abc_41234_new_n4211_; 
wire _abc_41234_new_n4212_; 
wire _abc_41234_new_n4213_; 
wire _abc_41234_new_n4214_; 
wire _abc_41234_new_n4215_; 
wire _abc_41234_new_n4216_; 
wire _abc_41234_new_n4217_; 
wire _abc_41234_new_n4218_; 
wire _abc_41234_new_n4219_; 
wire _abc_41234_new_n4220_; 
wire _abc_41234_new_n4221_; 
wire _abc_41234_new_n4222_; 
wire _abc_41234_new_n4223_; 
wire _abc_41234_new_n4224_; 
wire _abc_41234_new_n4225_; 
wire _abc_41234_new_n4226_; 
wire _abc_41234_new_n4227_; 
wire _abc_41234_new_n4228_; 
wire _abc_41234_new_n4229_; 
wire _abc_41234_new_n4230_; 
wire _abc_41234_new_n4231_; 
wire _abc_41234_new_n4232_; 
wire _abc_41234_new_n4234_; 
wire _abc_41234_new_n4235_; 
wire _abc_41234_new_n4236_; 
wire _abc_41234_new_n4237_; 
wire _abc_41234_new_n4238_; 
wire _abc_41234_new_n4239_; 
wire _abc_41234_new_n4240_; 
wire _abc_41234_new_n4241_; 
wire _abc_41234_new_n4242_; 
wire _abc_41234_new_n4243_; 
wire _abc_41234_new_n4244_; 
wire _abc_41234_new_n4245_; 
wire _abc_41234_new_n4246_; 
wire _abc_41234_new_n4247_; 
wire _abc_41234_new_n4248_; 
wire _abc_41234_new_n4249_; 
wire _abc_41234_new_n4250_; 
wire _abc_41234_new_n4251_; 
wire _abc_41234_new_n4252_; 
wire _abc_41234_new_n4253_; 
wire _abc_41234_new_n4254_; 
wire _abc_41234_new_n4255_; 
wire _abc_41234_new_n4257_; 
wire _abc_41234_new_n4258_; 
wire _abc_41234_new_n4260_; 
wire _abc_41234_new_n4262_; 
wire _abc_41234_new_n4264_; 
wire _abc_41234_new_n4266_; 
wire _abc_41234_new_n4268_; 
wire _abc_41234_new_n4270_; 
wire _abc_41234_new_n4272_; 
wire _abc_41234_new_n4274_; 
wire _abc_41234_new_n4274__bF_buf0; 
wire _abc_41234_new_n4274__bF_buf1; 
wire _abc_41234_new_n4274__bF_buf2; 
wire _abc_41234_new_n4274__bF_buf3; 
wire _abc_41234_new_n4275_; 
wire _abc_41234_new_n4276_; 
wire _abc_41234_new_n4277_; 
wire _abc_41234_new_n4278_; 
wire _abc_41234_new_n4279_; 
wire _abc_41234_new_n4280_; 
wire _abc_41234_new_n4281_; 
wire _abc_41234_new_n4282_; 
wire _abc_41234_new_n4283_; 
wire _abc_41234_new_n4284_; 
wire _abc_41234_new_n4285_; 
wire _abc_41234_new_n4286_; 
wire _abc_41234_new_n4287_; 
wire _abc_41234_new_n4288_; 
wire _abc_41234_new_n4289_; 
wire _abc_41234_new_n4290_; 
wire _abc_41234_new_n4291_; 
wire _abc_41234_new_n4292_; 
wire _abc_41234_new_n4293_; 
wire _abc_41234_new_n4294_; 
wire _abc_41234_new_n4295_; 
wire _abc_41234_new_n4296_; 
wire _abc_41234_new_n4297_; 
wire _abc_41234_new_n4297__bF_buf0; 
wire _abc_41234_new_n4297__bF_buf1; 
wire _abc_41234_new_n4297__bF_buf2; 
wire _abc_41234_new_n4297__bF_buf3; 
wire _abc_41234_new_n4298_; 
wire _abc_41234_new_n4299_; 
wire _abc_41234_new_n4300_; 
wire _abc_41234_new_n4301_; 
wire _abc_41234_new_n4302_; 
wire _abc_41234_new_n4303_; 
wire _abc_41234_new_n4304_; 
wire _abc_41234_new_n4305_; 
wire _abc_41234_new_n4306_; 
wire _abc_41234_new_n4307_; 
wire _abc_41234_new_n4308_; 
wire _abc_41234_new_n4309_; 
wire _abc_41234_new_n4310_; 
wire _abc_41234_new_n4311_; 
wire _abc_41234_new_n4312_; 
wire _abc_41234_new_n4313_; 
wire _abc_41234_new_n4314_; 
wire _abc_41234_new_n4315_; 
wire _abc_41234_new_n4316_; 
wire _abc_41234_new_n4317_; 
wire _abc_41234_new_n4318_; 
wire _abc_41234_new_n4320_; 
wire _abc_41234_new_n4321_; 
wire _abc_41234_new_n4322_; 
wire _abc_41234_new_n4323_; 
wire _abc_41234_new_n4324_; 
wire _abc_41234_new_n4325_; 
wire _abc_41234_new_n4326_; 
wire _abc_41234_new_n4327_; 
wire _abc_41234_new_n4328_; 
wire _abc_41234_new_n4329_; 
wire _abc_41234_new_n4330_; 
wire _abc_41234_new_n4331_; 
wire _abc_41234_new_n4332_; 
wire _abc_41234_new_n4333_; 
wire _abc_41234_new_n4334_; 
wire _abc_41234_new_n4335_; 
wire _abc_41234_new_n4336_; 
wire _abc_41234_new_n4338_; 
wire _abc_41234_new_n4339_; 
wire _abc_41234_new_n4340_; 
wire _abc_41234_new_n4341_; 
wire _abc_41234_new_n4342_; 
wire _abc_41234_new_n4343_; 
wire _abc_41234_new_n4344_; 
wire _abc_41234_new_n4345_; 
wire _abc_41234_new_n4346_; 
wire _abc_41234_new_n4347_; 
wire _abc_41234_new_n4348_; 
wire _abc_41234_new_n4349_; 
wire _abc_41234_new_n4350_; 
wire _abc_41234_new_n4351_; 
wire _abc_41234_new_n4353_; 
wire _abc_41234_new_n4354_; 
wire _abc_41234_new_n4355_; 
wire _abc_41234_new_n4356_; 
wire _abc_41234_new_n4357_; 
wire _abc_41234_new_n4358_; 
wire _abc_41234_new_n4359_; 
wire _abc_41234_new_n4360_; 
wire _abc_41234_new_n4361_; 
wire _abc_41234_new_n4362_; 
wire _abc_41234_new_n4363_; 
wire _abc_41234_new_n4364_; 
wire _abc_41234_new_n4365_; 
wire _abc_41234_new_n4366_; 
wire _abc_41234_new_n4367_; 
wire _abc_41234_new_n4368_; 
wire _abc_41234_new_n4369_; 
wire _abc_41234_new_n4371_; 
wire _abc_41234_new_n4372_; 
wire _abc_41234_new_n4373_; 
wire _abc_41234_new_n4374_; 
wire _abc_41234_new_n4375_; 
wire _abc_41234_new_n4376_; 
wire _abc_41234_new_n4377_; 
wire _abc_41234_new_n4378_; 
wire _abc_41234_new_n4379_; 
wire _abc_41234_new_n4380_; 
wire _abc_41234_new_n4381_; 
wire _abc_41234_new_n4382_; 
wire _abc_41234_new_n4383_; 
wire _abc_41234_new_n4384_; 
wire _abc_41234_new_n4385_; 
wire _abc_41234_new_n4386_; 
wire _abc_41234_new_n4388_; 
wire _abc_41234_new_n4389_; 
wire _abc_41234_new_n4390_; 
wire _abc_41234_new_n4391_; 
wire _abc_41234_new_n4392_; 
wire _abc_41234_new_n4393_; 
wire _abc_41234_new_n4394_; 
wire _abc_41234_new_n4395_; 
wire _abc_41234_new_n4396_; 
wire _abc_41234_new_n4397_; 
wire _abc_41234_new_n4398_; 
wire _abc_41234_new_n4399_; 
wire _abc_41234_new_n4400_; 
wire _abc_41234_new_n4401_; 
wire _abc_41234_new_n4402_; 
wire _abc_41234_new_n4403_; 
wire _abc_41234_new_n4404_; 
wire _abc_41234_new_n4405_; 
wire _abc_41234_new_n4407_; 
wire _abc_41234_new_n4408_; 
wire _abc_41234_new_n4409_; 
wire _abc_41234_new_n4410_; 
wire _abc_41234_new_n4411_; 
wire _abc_41234_new_n4412_; 
wire _abc_41234_new_n4413_; 
wire _abc_41234_new_n4414_; 
wire _abc_41234_new_n4415_; 
wire _abc_41234_new_n4416_; 
wire _abc_41234_new_n4417_; 
wire _abc_41234_new_n4418_; 
wire _abc_41234_new_n4419_; 
wire _abc_41234_new_n4420_; 
wire _abc_41234_new_n4421_; 
wire _abc_41234_new_n4422_; 
wire _abc_41234_new_n4423_; 
wire _abc_41234_new_n4424_; 
wire _abc_41234_new_n4426_; 
wire _abc_41234_new_n4427_; 
wire _abc_41234_new_n4428_; 
wire _abc_41234_new_n4429_; 
wire _abc_41234_new_n4430_; 
wire _abc_41234_new_n4431_; 
wire _abc_41234_new_n4432_; 
wire _abc_41234_new_n4433_; 
wire _abc_41234_new_n4434_; 
wire _abc_41234_new_n4435_; 
wire _abc_41234_new_n4436_; 
wire _abc_41234_new_n4437_; 
wire _abc_41234_new_n4438_; 
wire _abc_41234_new_n4439_; 
wire _abc_41234_new_n4440_; 
wire _abc_41234_new_n4441_; 
wire _abc_41234_new_n4442_; 
wire _abc_41234_new_n4443_; 
wire _abc_41234_new_n4445_; 
wire _abc_41234_new_n4446_; 
wire _abc_41234_new_n4447_; 
wire _abc_41234_new_n4448_; 
wire _abc_41234_new_n4449_; 
wire _abc_41234_new_n4450_; 
wire _abc_41234_new_n4451_; 
wire _abc_41234_new_n4452_; 
wire _abc_41234_new_n4453_; 
wire _abc_41234_new_n4454_; 
wire _abc_41234_new_n4455_; 
wire _abc_41234_new_n4456_; 
wire _abc_41234_new_n4457_; 
wire _abc_41234_new_n4458_; 
wire _abc_41234_new_n4459_; 
wire _abc_41234_new_n4460_; 
wire _abc_41234_new_n4461_; 
wire _abc_41234_new_n4463_; 
wire _abc_41234_new_n4464_; 
wire _abc_41234_new_n4465_; 
wire _abc_41234_new_n4466_; 
wire _abc_41234_new_n4467_; 
wire _abc_41234_new_n4468_; 
wire _abc_41234_new_n4469_; 
wire _abc_41234_new_n4470_; 
wire _abc_41234_new_n4471_; 
wire _abc_41234_new_n4472_; 
wire _abc_41234_new_n4473_; 
wire _abc_41234_new_n4474_; 
wire _abc_41234_new_n4475_; 
wire _abc_41234_new_n4476_; 
wire _abc_41234_new_n4477_; 
wire _abc_41234_new_n4478_; 
wire _abc_41234_new_n4480_; 
wire _abc_41234_new_n4481_; 
wire _abc_41234_new_n4482_; 
wire _abc_41234_new_n4483_; 
wire _abc_41234_new_n4484_; 
wire _abc_41234_new_n4485_; 
wire _abc_41234_new_n4486_; 
wire _abc_41234_new_n4487_; 
wire _abc_41234_new_n4488_; 
wire _abc_41234_new_n4489_; 
wire _abc_41234_new_n4490_; 
wire _abc_41234_new_n4491_; 
wire _abc_41234_new_n4492_; 
wire _abc_41234_new_n4493_; 
wire _abc_41234_new_n4494_; 
wire _abc_41234_new_n4495_; 
wire _abc_41234_new_n4496_; 
wire _abc_41234_new_n4497_; 
wire _abc_41234_new_n4499_; 
wire _abc_41234_new_n4500_; 
wire _abc_41234_new_n4501_; 
wire _abc_41234_new_n4502_; 
wire _abc_41234_new_n4503_; 
wire _abc_41234_new_n4504_; 
wire _abc_41234_new_n4505_; 
wire _abc_41234_new_n4506_; 
wire _abc_41234_new_n4507_; 
wire _abc_41234_new_n4508_; 
wire _abc_41234_new_n4509_; 
wire _abc_41234_new_n4510_; 
wire _abc_41234_new_n4511_; 
wire _abc_41234_new_n4512_; 
wire _abc_41234_new_n4513_; 
wire _abc_41234_new_n4514_; 
wire _abc_41234_new_n4515_; 
wire _abc_41234_new_n4517_; 
wire _abc_41234_new_n4518_; 
wire _abc_41234_new_n4519_; 
wire _abc_41234_new_n4520_; 
wire _abc_41234_new_n4521_; 
wire _abc_41234_new_n4522_; 
wire _abc_41234_new_n4523_; 
wire _abc_41234_new_n4524_; 
wire _abc_41234_new_n4525_; 
wire _abc_41234_new_n4526_; 
wire _abc_41234_new_n4527_; 
wire _abc_41234_new_n4528_; 
wire _abc_41234_new_n4529_; 
wire _abc_41234_new_n4530_; 
wire _abc_41234_new_n4531_; 
wire _abc_41234_new_n4532_; 
wire _abc_41234_new_n4533_; 
wire _abc_41234_new_n4534_; 
wire _abc_41234_new_n4535_; 
wire _abc_41234_new_n4537_; 
wire _abc_41234_new_n4538_; 
wire _abc_41234_new_n4539_; 
wire _abc_41234_new_n4540_; 
wire _abc_41234_new_n4541_; 
wire _abc_41234_new_n4542_; 
wire _abc_41234_new_n4543_; 
wire _abc_41234_new_n4544_; 
wire _abc_41234_new_n4545_; 
wire _abc_41234_new_n4546_; 
wire _abc_41234_new_n4547_; 
wire _abc_41234_new_n4548_; 
wire _abc_41234_new_n4549_; 
wire _abc_41234_new_n4550_; 
wire _abc_41234_new_n4551_; 
wire _abc_41234_new_n4552_; 
wire _abc_41234_new_n4553_; 
wire _abc_41234_new_n4555_; 
wire _abc_41234_new_n4556_; 
wire _abc_41234_new_n4557_; 
wire _abc_41234_new_n4558_; 
wire _abc_41234_new_n4559_; 
wire _abc_41234_new_n4560_; 
wire _abc_41234_new_n4561_; 
wire _abc_41234_new_n4562_; 
wire _abc_41234_new_n4563_; 
wire _abc_41234_new_n4564_; 
wire _abc_41234_new_n4565_; 
wire _abc_41234_new_n4566_; 
wire _abc_41234_new_n4567_; 
wire _abc_41234_new_n4568_; 
wire _abc_41234_new_n4569_; 
wire _abc_41234_new_n4570_; 
wire _abc_41234_new_n4571_; 
wire _abc_41234_new_n4572_; 
wire _abc_41234_new_n4573_; 
wire _abc_41234_new_n4574_; 
wire _abc_41234_new_n4576_; 
wire _abc_41234_new_n4577_; 
wire _abc_41234_new_n4578_; 
wire _abc_41234_new_n4579_; 
wire _abc_41234_new_n4580_; 
wire _abc_41234_new_n4581_; 
wire _abc_41234_new_n4582_; 
wire _abc_41234_new_n4583_; 
wire _abc_41234_new_n4584_; 
wire _abc_41234_new_n4585_; 
wire _abc_41234_new_n4586_; 
wire _abc_41234_new_n4587_; 
wire _abc_41234_new_n4588_; 
wire _abc_41234_new_n4589_; 
wire _abc_41234_new_n4590_; 
wire _abc_41234_new_n4591_; 
wire _abc_41234_new_n4592_; 
wire _abc_41234_new_n4593_; 
wire _abc_41234_new_n4594_; 
wire _abc_41234_new_n4595_; 
wire _abc_41234_new_n4596_; 
wire _abc_41234_new_n4597_; 
wire _abc_41234_new_n4599_; 
wire _abc_41234_new_n4600_; 
wire _abc_41234_new_n4601_; 
wire _abc_41234_new_n4602_; 
wire _abc_41234_new_n4604_; 
wire _abc_41234_new_n4605_; 
wire _abc_41234_new_n4606_; 
wire _abc_41234_new_n4607_; 
wire _abc_41234_new_n4608_; 
wire _abc_41234_new_n4609_; 
wire _abc_41234_new_n4611_; 
wire _abc_41234_new_n4612_; 
wire _abc_41234_new_n4613_; 
wire _abc_41234_new_n4614_; 
wire _abc_41234_new_n4615_; 
wire _abc_41234_new_n4616_; 
wire _abc_41234_new_n4617_; 
wire _abc_41234_new_n4618_; 
wire _abc_41234_new_n4620_; 
wire _abc_41234_new_n4621_; 
wire _abc_41234_new_n4622_; 
wire _abc_41234_new_n4623_; 
wire _abc_41234_new_n4625_; 
wire _abc_41234_new_n4626_; 
wire _abc_41234_new_n4627_; 
wire _abc_41234_new_n4628_; 
wire _abc_41234_new_n4630_; 
wire _abc_41234_new_n4631_; 
wire _abc_41234_new_n4632_; 
wire _abc_41234_new_n4633_; 
wire _abc_41234_new_n4635_; 
wire _abc_41234_new_n4636_; 
wire _abc_41234_new_n4637_; 
wire _abc_41234_new_n4638_; 
wire _abc_41234_new_n4640_; 
wire _abc_41234_new_n4641_; 
wire _abc_41234_new_n4642_; 
wire _abc_41234_new_n4643_; 
wire _abc_41234_new_n4645_; 
wire _abc_41234_new_n4646_; 
wire _abc_41234_new_n4647_; 
wire _abc_41234_new_n4648_; 
wire _abc_41234_new_n4650_; 
wire _abc_41234_new_n4651_; 
wire _abc_41234_new_n4652_; 
wire _abc_41234_new_n4653_; 
wire _abc_41234_new_n4655_; 
wire _abc_41234_new_n4656_; 
wire _abc_41234_new_n4657_; 
wire _abc_41234_new_n4659_; 
wire _abc_41234_new_n4660_; 
wire _abc_41234_new_n4661_; 
wire _abc_41234_new_n4662_; 
wire _abc_41234_new_n4663_; 
wire _abc_41234_new_n4664_; 
wire _abc_41234_new_n4666_; 
wire _abc_41234_new_n4667_; 
wire _abc_41234_new_n4668_; 
wire _abc_41234_new_n4669_; 
wire _abc_41234_new_n4671_; 
wire _abc_41234_new_n4672_; 
wire _abc_41234_new_n4673_; 
wire _abc_41234_new_n4674_; 
wire _abc_41234_new_n4676_; 
wire _abc_41234_new_n4677_; 
wire _abc_41234_new_n4678_; 
wire _abc_41234_new_n4680_; 
wire _abc_41234_new_n4681_; 
wire _abc_41234_new_n4682_; 
wire _abc_41234_new_n4684_; 
wire _abc_41234_new_n4685_; 
wire _abc_41234_new_n4686_; 
wire _abc_41234_new_n4687_; 
wire _abc_41234_new_n4689_; 
wire _abc_41234_new_n4690_; 
wire _abc_41234_new_n4691_; 
wire _abc_41234_new_n4693_; 
wire _abc_41234_new_n4695_; 
wire _abc_41234_new_n4696_; 
wire _abc_41234_new_n4697_; 
wire _abc_41234_new_n4698_; 
wire _abc_41234_new_n4699_; 
wire _abc_41234_new_n4700_; 
wire _abc_41234_new_n4701_; 
wire _abc_41234_new_n4703_; 
wire _abc_41234_new_n4704_; 
wire _abc_41234_new_n4705_; 
wire _abc_41234_new_n4706_; 
wire _abc_41234_new_n4708_; 
wire _abc_41234_new_n4709_; 
wire _abc_41234_new_n4710_; 
wire _abc_41234_new_n4711_; 
wire _abc_41234_new_n4712_; 
wire _abc_41234_new_n4713_; 
wire _abc_41234_new_n4714_; 
wire _abc_41234_new_n4715_; 
wire _abc_41234_new_n4716_; 
wire _abc_41234_new_n4717_; 
wire _abc_41234_new_n4718_; 
wire _abc_41234_new_n4719_; 
wire _abc_41234_new_n4720_; 
wire _abc_41234_new_n4721_; 
wire _abc_41234_new_n4722_; 
wire _abc_41234_new_n4723_; 
wire _abc_41234_new_n4724_; 
wire _abc_41234_new_n4725_; 
wire _abc_41234_new_n4726_; 
wire _abc_41234_new_n4727_; 
wire _abc_41234_new_n4728_; 
wire _abc_41234_new_n4729_; 
wire _abc_41234_new_n4730_; 
wire _abc_41234_new_n4731_; 
wire _abc_41234_new_n4732_; 
wire _abc_41234_new_n4733_; 
wire _abc_41234_new_n4734_; 
wire _abc_41234_new_n4735_; 
wire _abc_41234_new_n4736_; 
wire _abc_41234_new_n4737_; 
wire _abc_41234_new_n4738_; 
wire _abc_41234_new_n4739_; 
wire _abc_41234_new_n4740_; 
wire _abc_41234_new_n4741_; 
wire _abc_41234_new_n4742_; 
wire _abc_41234_new_n4743_; 
wire _abc_41234_new_n4744_; 
wire _abc_41234_new_n4745_; 
wire _abc_41234_new_n4746_; 
wire _abc_41234_new_n4747_; 
wire _abc_41234_new_n4748_; 
wire _abc_41234_new_n4749_; 
wire _abc_41234_new_n4750_; 
wire _abc_41234_new_n4751_; 
wire _abc_41234_new_n4752_; 
wire _abc_41234_new_n4753_; 
wire _abc_41234_new_n4754_; 
wire _abc_41234_new_n4755_; 
wire _abc_41234_new_n4756_; 
wire _abc_41234_new_n4757_; 
wire _abc_41234_new_n4758_; 
wire _abc_41234_new_n4759_; 
wire _abc_41234_new_n4760_; 
wire _abc_41234_new_n4761_; 
wire _abc_41234_new_n4762_; 
wire _abc_41234_new_n4763_; 
wire _abc_41234_new_n4764_; 
wire _abc_41234_new_n4765_; 
wire _abc_41234_new_n4766_; 
wire _abc_41234_new_n4767_; 
wire _abc_41234_new_n4768_; 
wire _abc_41234_new_n4769_; 
wire _abc_41234_new_n4770_; 
wire _abc_41234_new_n4771_; 
wire _abc_41234_new_n4772_; 
wire _abc_41234_new_n4773_; 
wire _abc_41234_new_n4774_; 
wire _abc_41234_new_n4775_; 
wire _abc_41234_new_n4776_; 
wire _abc_41234_new_n4777_; 
wire _abc_41234_new_n4778_; 
wire _abc_41234_new_n4779_; 
wire _abc_41234_new_n4780_; 
wire _abc_41234_new_n4781_; 
wire _abc_41234_new_n4782_; 
wire _abc_41234_new_n4783_; 
wire _abc_41234_new_n4784_; 
wire _abc_41234_new_n4785_; 
wire _abc_41234_new_n4786_; 
wire _abc_41234_new_n4787_; 
wire _abc_41234_new_n4788_; 
wire _abc_41234_new_n4789_; 
wire _abc_41234_new_n4790_; 
wire _abc_41234_new_n4791_; 
wire _abc_41234_new_n4792_; 
wire _abc_41234_new_n4793_; 
wire _abc_41234_new_n4794_; 
wire _abc_41234_new_n4795_; 
wire _abc_41234_new_n4796_; 
wire _abc_41234_new_n4797_; 
wire _abc_41234_new_n4798_; 
wire _abc_41234_new_n4799_; 
wire _abc_41234_new_n4800_; 
wire _abc_41234_new_n4801_; 
wire _abc_41234_new_n4802_; 
wire _abc_41234_new_n4803_; 
wire _abc_41234_new_n4804_; 
wire _abc_41234_new_n4805_; 
wire _abc_41234_new_n4806_; 
wire _abc_41234_new_n4807_; 
wire _abc_41234_new_n4808_; 
wire _abc_41234_new_n4809_; 
wire _abc_41234_new_n4810_; 
wire _abc_41234_new_n4811_; 
wire _abc_41234_new_n4812_; 
wire _abc_41234_new_n4813_; 
wire _abc_41234_new_n4814_; 
wire _abc_41234_new_n4815_; 
wire _abc_41234_new_n4816_; 
wire _abc_41234_new_n4817_; 
wire _abc_41234_new_n4818_; 
wire _abc_41234_new_n4820_; 
wire _abc_41234_new_n4821_; 
wire _abc_41234_new_n4822_; 
wire _abc_41234_new_n4823_; 
wire _abc_41234_new_n4824_; 
wire _abc_41234_new_n4825_; 
wire _abc_41234_new_n4826_; 
wire _abc_41234_new_n4827_; 
wire _abc_41234_new_n4828_; 
wire _abc_41234_new_n4829_; 
wire _abc_41234_new_n4830_; 
wire _abc_41234_new_n4831_; 
wire _abc_41234_new_n4832_; 
wire _abc_41234_new_n4833_; 
wire _abc_41234_new_n4834_; 
wire _abc_41234_new_n4835_; 
wire _abc_41234_new_n4836_; 
wire _abc_41234_new_n4837_; 
wire _abc_41234_new_n4838_; 
wire _abc_41234_new_n4840_; 
wire _abc_41234_new_n4841_; 
wire _abc_41234_new_n4842_; 
wire _abc_41234_new_n4843_; 
wire _abc_41234_new_n4844_; 
wire _abc_41234_new_n4845_; 
wire _abc_41234_new_n4846_; 
wire _abc_41234_new_n4847_; 
wire _abc_41234_new_n4848_; 
wire _abc_41234_new_n4849_; 
wire _abc_41234_new_n4850_; 
wire _abc_41234_new_n4851_; 
wire _abc_41234_new_n4852_; 
wire _abc_41234_new_n4853_; 
wire _abc_41234_new_n4854_; 
wire _abc_41234_new_n4855_; 
wire _abc_41234_new_n4856_; 
wire _abc_41234_new_n4858_; 
wire _abc_41234_new_n4859_; 
wire _abc_41234_new_n4860_; 
wire _abc_41234_new_n4861_; 
wire _abc_41234_new_n4862_; 
wire _abc_41234_new_n4863_; 
wire _abc_41234_new_n4864_; 
wire _abc_41234_new_n4865_; 
wire _abc_41234_new_n4866_; 
wire _abc_41234_new_n4867_; 
wire _abc_41234_new_n4869_; 
wire _abc_41234_new_n4870_; 
wire _abc_41234_new_n4871_; 
wire _abc_41234_new_n4872_; 
wire _abc_41234_new_n4873_; 
wire _abc_41234_new_n4874_; 
wire _abc_41234_new_n4875_; 
wire _abc_41234_new_n4876_; 
wire _abc_41234_new_n4877_; 
wire _abc_41234_new_n4878_; 
wire _abc_41234_new_n4879_; 
wire _abc_41234_new_n4880_; 
wire _abc_41234_new_n4882_; 
wire _abc_41234_new_n4883_; 
wire _abc_41234_new_n4884_; 
wire _abc_41234_new_n4885_; 
wire _abc_41234_new_n4886_; 
wire _abc_41234_new_n4887_; 
wire _abc_41234_new_n4889_; 
wire _abc_41234_new_n4890_; 
wire _abc_41234_new_n4891_; 
wire _abc_41234_new_n4892_; 
wire _abc_41234_new_n501_; 
wire _abc_41234_new_n502_; 
wire _abc_41234_new_n503_; 
wire _abc_41234_new_n504_; 
wire _abc_41234_new_n505_; 
wire _abc_41234_new_n506_; 
wire _abc_41234_new_n507_; 
wire _abc_41234_new_n508_; 
wire _abc_41234_new_n509_; 
wire _abc_41234_new_n510_; 
wire _abc_41234_new_n511_; 
wire _abc_41234_new_n512_; 
wire _abc_41234_new_n513_; 
wire _abc_41234_new_n514_; 
wire _abc_41234_new_n515_; 
wire _abc_41234_new_n515__bF_buf0; 
wire _abc_41234_new_n515__bF_buf1; 
wire _abc_41234_new_n515__bF_buf2; 
wire _abc_41234_new_n515__bF_buf3; 
wire _abc_41234_new_n515__bF_buf4; 
wire _abc_41234_new_n515__bF_buf5; 
wire _abc_41234_new_n515__bF_buf6; 
wire _abc_41234_new_n516_; 
wire _abc_41234_new_n516__bF_buf0; 
wire _abc_41234_new_n516__bF_buf1; 
wire _abc_41234_new_n516__bF_buf2; 
wire _abc_41234_new_n516__bF_buf3; 
wire _abc_41234_new_n516__bF_buf4; 
wire _abc_41234_new_n516__bF_buf5; 
wire _abc_41234_new_n517_; 
wire _abc_41234_new_n518_; 
wire _abc_41234_new_n519_; 
wire _abc_41234_new_n520_; 
wire _abc_41234_new_n521_; 
wire _abc_41234_new_n522_; 
wire _abc_41234_new_n523_; 
wire _abc_41234_new_n523__bF_buf0; 
wire _abc_41234_new_n523__bF_buf1; 
wire _abc_41234_new_n523__bF_buf2; 
wire _abc_41234_new_n523__bF_buf3; 
wire _abc_41234_new_n523__bF_buf4; 
wire _abc_41234_new_n524_; 
wire _abc_41234_new_n525_; 
wire _abc_41234_new_n525__bF_buf0; 
wire _abc_41234_new_n525__bF_buf1; 
wire _abc_41234_new_n525__bF_buf2; 
wire _abc_41234_new_n525__bF_buf3; 
wire _abc_41234_new_n526_; 
wire _abc_41234_new_n526__bF_buf0; 
wire _abc_41234_new_n526__bF_buf1; 
wire _abc_41234_new_n526__bF_buf2; 
wire _abc_41234_new_n526__bF_buf3; 
wire _abc_41234_new_n527_; 
wire _abc_41234_new_n528_; 
wire _abc_41234_new_n529_; 
wire _abc_41234_new_n530_; 
wire _abc_41234_new_n531_; 
wire _abc_41234_new_n532_; 
wire _abc_41234_new_n533_; 
wire _abc_41234_new_n534_; 
wire _abc_41234_new_n534__bF_buf0; 
wire _abc_41234_new_n534__bF_buf1; 
wire _abc_41234_new_n534__bF_buf2; 
wire _abc_41234_new_n534__bF_buf3; 
wire _abc_41234_new_n534__bF_buf4; 
wire _abc_41234_new_n534__bF_buf5; 
wire _abc_41234_new_n535_; 
wire _abc_41234_new_n536_; 
wire _abc_41234_new_n536__bF_buf0; 
wire _abc_41234_new_n536__bF_buf1; 
wire _abc_41234_new_n536__bF_buf2; 
wire _abc_41234_new_n536__bF_buf3; 
wire _abc_41234_new_n536__bF_buf4; 
wire _abc_41234_new_n536__bF_buf5; 
wire _abc_41234_new_n537_; 
wire _abc_41234_new_n537__bF_buf0; 
wire _abc_41234_new_n537__bF_buf1; 
wire _abc_41234_new_n537__bF_buf2; 
wire _abc_41234_new_n537__bF_buf3; 
wire _abc_41234_new_n538_; 
wire _abc_41234_new_n539_; 
wire _abc_41234_new_n540_; 
wire _abc_41234_new_n541_; 
wire _abc_41234_new_n542_; 
wire _abc_41234_new_n543_; 
wire _abc_41234_new_n544_; 
wire _abc_41234_new_n544__bF_buf0; 
wire _abc_41234_new_n544__bF_buf1; 
wire _abc_41234_new_n544__bF_buf2; 
wire _abc_41234_new_n544__bF_buf3; 
wire _abc_41234_new_n545_; 
wire _abc_41234_new_n546_; 
wire _abc_41234_new_n546__bF_buf0; 
wire _abc_41234_new_n546__bF_buf1; 
wire _abc_41234_new_n546__bF_buf2; 
wire _abc_41234_new_n546__bF_buf3; 
wire _abc_41234_new_n546__bF_buf4; 
wire _abc_41234_new_n546__bF_buf5; 
wire _abc_41234_new_n547_; 
wire _abc_41234_new_n548_; 
wire _abc_41234_new_n549_; 
wire _abc_41234_new_n550_; 
wire _abc_41234_new_n551_; 
wire _abc_41234_new_n552_; 
wire _abc_41234_new_n553_; 
wire _abc_41234_new_n554_; 
wire _abc_41234_new_n555_; 
wire _abc_41234_new_n556_; 
wire _abc_41234_new_n557_; 
wire _abc_41234_new_n558_; 
wire _abc_41234_new_n559_; 
wire _abc_41234_new_n560_; 
wire _abc_41234_new_n561_; 
wire _abc_41234_new_n562_; 
wire _abc_41234_new_n563_; 
wire _abc_41234_new_n564_; 
wire _abc_41234_new_n565_; 
wire _abc_41234_new_n566_; 
wire _abc_41234_new_n567_; 
wire _abc_41234_new_n568_; 
wire _abc_41234_new_n569_; 
wire _abc_41234_new_n570_; 
wire _abc_41234_new_n571_; 
wire _abc_41234_new_n572_; 
wire _abc_41234_new_n573_; 
wire _abc_41234_new_n574_; 
wire _abc_41234_new_n575_; 
wire _abc_41234_new_n576_; 
wire _abc_41234_new_n577_; 
wire _abc_41234_new_n578_; 
wire _abc_41234_new_n579_; 
wire _abc_41234_new_n580_; 
wire _abc_41234_new_n581_; 
wire _abc_41234_new_n582_; 
wire _abc_41234_new_n583_; 
wire _abc_41234_new_n584_; 
wire _abc_41234_new_n585_; 
wire _abc_41234_new_n586_; 
wire _abc_41234_new_n587_; 
wire _abc_41234_new_n588_; 
wire _abc_41234_new_n589_; 
wire _abc_41234_new_n590_; 
wire _abc_41234_new_n591_; 
wire _abc_41234_new_n592_; 
wire _abc_41234_new_n593_; 
wire _abc_41234_new_n594_; 
wire _abc_41234_new_n595_; 
wire _abc_41234_new_n596_; 
wire _abc_41234_new_n597_; 
wire _abc_41234_new_n598_; 
wire _abc_41234_new_n599_; 
wire _abc_41234_new_n600_; 
wire _abc_41234_new_n601_; 
wire _abc_41234_new_n602_; 
wire _abc_41234_new_n603_; 
wire _abc_41234_new_n604_; 
wire _abc_41234_new_n605_; 
wire _abc_41234_new_n606_; 
wire _abc_41234_new_n607_; 
wire _abc_41234_new_n608_; 
wire _abc_41234_new_n609_; 
wire _abc_41234_new_n610_; 
wire _abc_41234_new_n611_; 
wire _abc_41234_new_n612_; 
wire _abc_41234_new_n613_; 
wire _abc_41234_new_n614_; 
wire _abc_41234_new_n615_; 
wire _abc_41234_new_n616_; 
wire _abc_41234_new_n617_; 
wire _abc_41234_new_n618_; 
wire _abc_41234_new_n619_; 
wire _abc_41234_new_n620_; 
wire _abc_41234_new_n620__bF_buf0; 
wire _abc_41234_new_n620__bF_buf1; 
wire _abc_41234_new_n620__bF_buf2; 
wire _abc_41234_new_n620__bF_buf3; 
wire _abc_41234_new_n620__bF_buf4; 
wire _abc_41234_new_n620__bF_buf5; 
wire _abc_41234_new_n621_; 
wire _abc_41234_new_n622_; 
wire _abc_41234_new_n623_; 
wire _abc_41234_new_n624_; 
wire _abc_41234_new_n625_; 
wire _abc_41234_new_n626_; 
wire _abc_41234_new_n627_; 
wire _abc_41234_new_n628_; 
wire _abc_41234_new_n629_; 
wire _abc_41234_new_n630_; 
wire _abc_41234_new_n631_; 
wire _abc_41234_new_n632_; 
wire _abc_41234_new_n633_; 
wire _abc_41234_new_n634_; 
wire _abc_41234_new_n635_; 
wire _abc_41234_new_n636_; 
wire _abc_41234_new_n637_; 
wire _abc_41234_new_n638_; 
wire _abc_41234_new_n639_; 
wire _abc_41234_new_n640_; 
wire _abc_41234_new_n641_; 
wire _abc_41234_new_n642_; 
wire _abc_41234_new_n643_; 
wire _abc_41234_new_n644_; 
wire _abc_41234_new_n645_; 
wire _abc_41234_new_n646_; 
wire _abc_41234_new_n647_; 
wire _abc_41234_new_n648_; 
wire _abc_41234_new_n649_; 
wire _abc_41234_new_n650_; 
wire _abc_41234_new_n651_; 
wire _abc_41234_new_n652_; 
wire _abc_41234_new_n653_; 
wire _abc_41234_new_n654_; 
wire _abc_41234_new_n655_; 
wire _abc_41234_new_n656_; 
wire _abc_41234_new_n657_; 
wire _abc_41234_new_n658_; 
wire _abc_41234_new_n659_; 
wire _abc_41234_new_n660_; 
wire _abc_41234_new_n660__bF_buf0; 
wire _abc_41234_new_n660__bF_buf1; 
wire _abc_41234_new_n660__bF_buf2; 
wire _abc_41234_new_n660__bF_buf3; 
wire _abc_41234_new_n660__bF_buf4; 
wire _abc_41234_new_n660__bF_buf5; 
wire _abc_41234_new_n660__bF_buf6; 
wire _abc_41234_new_n660__bF_buf7; 
wire _abc_41234_new_n661_; 
wire _abc_41234_new_n662_; 
wire _abc_41234_new_n663_; 
wire _abc_41234_new_n664_; 
wire _abc_41234_new_n665_; 
wire _abc_41234_new_n665__bF_buf0; 
wire _abc_41234_new_n665__bF_buf1; 
wire _abc_41234_new_n665__bF_buf2; 
wire _abc_41234_new_n665__bF_buf3; 
wire _abc_41234_new_n666_; 
wire _abc_41234_new_n667_; 
wire _abc_41234_new_n668_; 
wire _abc_41234_new_n668__bF_buf0; 
wire _abc_41234_new_n668__bF_buf1; 
wire _abc_41234_new_n668__bF_buf2; 
wire _abc_41234_new_n668__bF_buf3; 
wire _abc_41234_new_n668__bF_buf4; 
wire _abc_41234_new_n668__bF_buf5; 
wire _abc_41234_new_n669_; 
wire _abc_41234_new_n669__bF_buf0; 
wire _abc_41234_new_n669__bF_buf1; 
wire _abc_41234_new_n669__bF_buf2; 
wire _abc_41234_new_n669__bF_buf3; 
wire _abc_41234_new_n670_; 
wire _abc_41234_new_n671_; 
wire _abc_41234_new_n672_; 
wire _abc_41234_new_n673_; 
wire _abc_41234_new_n674_; 
wire _abc_41234_new_n675_; 
wire _abc_41234_new_n676_; 
wire _abc_41234_new_n677_; 
wire _abc_41234_new_n678_; 
wire _abc_41234_new_n679_; 
wire _abc_41234_new_n680_; 
wire _abc_41234_new_n681_; 
wire _abc_41234_new_n682_; 
wire _abc_41234_new_n683_; 
wire _abc_41234_new_n684_; 
wire _abc_41234_new_n685_; 
wire _abc_41234_new_n686_; 
wire _abc_41234_new_n687_; 
wire _abc_41234_new_n688_; 
wire _abc_41234_new_n689_; 
wire _abc_41234_new_n690_; 
wire _abc_41234_new_n691_; 
wire _abc_41234_new_n692_; 
wire _abc_41234_new_n693_; 
wire _abc_41234_new_n694_; 
wire _abc_41234_new_n695_; 
wire _abc_41234_new_n696_; 
wire _abc_41234_new_n697_; 
wire _abc_41234_new_n698_; 
wire _abc_41234_new_n699_; 
wire _abc_41234_new_n700_; 
wire _abc_41234_new_n701_; 
wire _abc_41234_new_n702_; 
wire _abc_41234_new_n703_; 
wire _abc_41234_new_n704_; 
wire _abc_41234_new_n705_; 
wire _abc_41234_new_n706_; 
wire _abc_41234_new_n707_; 
wire _abc_41234_new_n708_; 
wire _abc_41234_new_n709_; 
wire _abc_41234_new_n710_; 
wire _abc_41234_new_n711_; 
wire _abc_41234_new_n712_; 
wire _abc_41234_new_n713_; 
wire _abc_41234_new_n714_; 
wire _abc_41234_new_n715_; 
wire _abc_41234_new_n716_; 
wire _abc_41234_new_n718_; 
wire _abc_41234_new_n719_; 
wire _abc_41234_new_n720_; 
wire _abc_41234_new_n721_; 
wire _abc_41234_new_n722_; 
wire _abc_41234_new_n722__bF_buf0; 
wire _abc_41234_new_n722__bF_buf1; 
wire _abc_41234_new_n722__bF_buf2; 
wire _abc_41234_new_n722__bF_buf3; 
wire _abc_41234_new_n723_; 
wire _abc_41234_new_n724_; 
wire _abc_41234_new_n725_; 
wire _abc_41234_new_n726_; 
wire _abc_41234_new_n727_; 
wire _abc_41234_new_n728_; 
wire _abc_41234_new_n729_; 
wire _abc_41234_new_n730_; 
wire _abc_41234_new_n731_; 
wire _abc_41234_new_n732_; 
wire _abc_41234_new_n733_; 
wire _abc_41234_new_n734_; 
wire _abc_41234_new_n735_; 
wire _abc_41234_new_n736_; 
wire _abc_41234_new_n737_; 
wire _abc_41234_new_n738_; 
wire _abc_41234_new_n739_; 
wire _abc_41234_new_n740_; 
wire _abc_41234_new_n741_; 
wire _abc_41234_new_n742_; 
wire _abc_41234_new_n743_; 
wire _abc_41234_new_n744_; 
wire _abc_41234_new_n745_; 
wire _abc_41234_new_n746_; 
wire _abc_41234_new_n747_; 
wire _abc_41234_new_n748_; 
wire _abc_41234_new_n749_; 
wire _abc_41234_new_n750_; 
wire _abc_41234_new_n751_; 
wire _abc_41234_new_n752_; 
wire _abc_41234_new_n753_; 
wire _abc_41234_new_n754_; 
wire _abc_41234_new_n755_; 
wire _abc_41234_new_n756_; 
wire _abc_41234_new_n757_; 
wire _abc_41234_new_n758_; 
wire _abc_41234_new_n759_; 
wire _abc_41234_new_n760_; 
wire _abc_41234_new_n761_; 
wire _abc_41234_new_n762_; 
wire _abc_41234_new_n763_; 
wire _abc_41234_new_n765_; 
wire _abc_41234_new_n766_; 
wire _abc_41234_new_n767_; 
wire _abc_41234_new_n768_; 
wire _abc_41234_new_n769_; 
wire _abc_41234_new_n770_; 
wire _abc_41234_new_n771_; 
wire _abc_41234_new_n772_; 
wire _abc_41234_new_n773_; 
wire _abc_41234_new_n774_; 
wire _abc_41234_new_n775_; 
wire _abc_41234_new_n776_; 
wire _abc_41234_new_n777_; 
wire _abc_41234_new_n778_; 
wire _abc_41234_new_n779_; 
wire _abc_41234_new_n780_; 
wire _abc_41234_new_n781_; 
wire _abc_41234_new_n782_; 
wire _abc_41234_new_n783_; 
wire _abc_41234_new_n784_; 
wire _abc_41234_new_n785_; 
wire _abc_41234_new_n786_; 
wire _abc_41234_new_n787_; 
wire _abc_41234_new_n788_; 
wire _abc_41234_new_n789_; 
wire _abc_41234_new_n790_; 
wire _abc_41234_new_n791_; 
wire _abc_41234_new_n792_; 
wire _abc_41234_new_n793_; 
wire _abc_41234_new_n794_; 
wire _abc_41234_new_n795_; 
wire _abc_41234_new_n796_; 
wire _abc_41234_new_n797_; 
wire _abc_41234_new_n798_; 
wire _abc_41234_new_n799_; 
wire _abc_41234_new_n800_; 
wire _abc_41234_new_n801_; 
wire _abc_41234_new_n802_; 
wire _abc_41234_new_n803_; 
wire _abc_41234_new_n805_; 
wire _abc_41234_new_n806_; 
wire _abc_41234_new_n807_; 
wire _abc_41234_new_n808_; 
wire _abc_41234_new_n809_; 
wire _abc_41234_new_n810_; 
wire _abc_41234_new_n811_; 
wire _abc_41234_new_n812_; 
wire _abc_41234_new_n813_; 
wire _abc_41234_new_n814_; 
wire _abc_41234_new_n815_; 
wire _abc_41234_new_n816_; 
wire _abc_41234_new_n817_; 
wire _abc_41234_new_n818_; 
wire _abc_41234_new_n819_; 
wire _abc_41234_new_n820_; 
wire _abc_41234_new_n821_; 
wire _abc_41234_new_n822_; 
wire _abc_41234_new_n823_; 
wire _abc_41234_new_n824_; 
wire _abc_41234_new_n825_; 
wire _abc_41234_new_n826_; 
wire _abc_41234_new_n827_; 
wire _abc_41234_new_n828_; 
wire _abc_41234_new_n829_; 
wire _abc_41234_new_n830_; 
wire _abc_41234_new_n831_; 
wire _abc_41234_new_n832_; 
wire _abc_41234_new_n833_; 
wire _abc_41234_new_n834_; 
wire _abc_41234_new_n835_; 
wire _abc_41234_new_n836_; 
wire _abc_41234_new_n837_; 
wire _abc_41234_new_n838_; 
wire _abc_41234_new_n839_; 
wire _abc_41234_new_n840_; 
wire _abc_41234_new_n841_; 
wire _abc_41234_new_n842_; 
wire _abc_41234_new_n843_; 
wire _abc_41234_new_n844_; 
wire _abc_41234_new_n845_; 
wire _abc_41234_new_n847_; 
wire _abc_41234_new_n848_; 
wire _abc_41234_new_n849_; 
wire _abc_41234_new_n850_; 
wire _abc_41234_new_n851_; 
wire _abc_41234_new_n852_; 
wire _abc_41234_new_n853_; 
wire _abc_41234_new_n854_; 
wire _abc_41234_new_n855_; 
wire _abc_41234_new_n856_; 
wire _abc_41234_new_n857_; 
wire _abc_41234_new_n858_; 
wire _abc_41234_new_n859_; 
wire _abc_41234_new_n860_; 
wire _abc_41234_new_n861_; 
wire _abc_41234_new_n862_; 
wire _abc_41234_new_n863_; 
wire _abc_41234_new_n864_; 
wire _abc_41234_new_n865_; 
wire _abc_41234_new_n866_; 
wire _abc_41234_new_n867_; 
wire _abc_41234_new_n868_; 
wire _abc_41234_new_n869_; 
wire _abc_41234_new_n870_; 
wire _abc_41234_new_n871_; 
wire _abc_41234_new_n872_; 
wire _abc_41234_new_n873_; 
wire _abc_41234_new_n874_; 
wire _abc_41234_new_n875_; 
wire _abc_41234_new_n876_; 
wire _abc_41234_new_n877_; 
wire _abc_41234_new_n878_; 
wire _abc_41234_new_n879_; 
wire _abc_41234_new_n880_; 
wire _abc_41234_new_n881_; 
wire _abc_41234_new_n882_; 
wire _abc_41234_new_n883_; 
wire _abc_41234_new_n884_; 
wire _abc_41234_new_n885_; 
wire _abc_41234_new_n886_; 
wire _abc_41234_new_n887_; 
wire _abc_41234_new_n888_; 
wire _abc_41234_new_n889_; 
wire _abc_41234_new_n890_; 
wire _abc_41234_new_n891_; 
wire _abc_41234_new_n892_; 
wire _abc_41234_new_n893_; 
wire _abc_41234_new_n895_; 
wire _abc_41234_new_n896_; 
wire _abc_41234_new_n897_; 
wire _abc_41234_new_n898_; 
wire _abc_41234_new_n899_; 
wire _abc_41234_new_n900_; 
wire _abc_41234_new_n901_; 
wire _abc_41234_new_n902_; 
wire _abc_41234_new_n903_; 
wire _abc_41234_new_n904_; 
wire _abc_41234_new_n905_; 
wire _abc_41234_new_n906_; 
wire _abc_41234_new_n907_; 
wire _abc_41234_new_n908_; 
wire _abc_41234_new_n909_; 
wire _abc_41234_new_n910_; 
wire _abc_41234_new_n911_; 
wire _abc_41234_new_n912_; 
wire _abc_41234_new_n913_; 
wire _abc_41234_new_n914_; 
wire _abc_41234_new_n915_; 
wire _abc_41234_new_n916_; 
wire _abc_41234_new_n917_; 
wire _abc_41234_new_n918_; 
wire _abc_41234_new_n919_; 
wire _abc_41234_new_n920_; 
wire _abc_41234_new_n921_; 
wire _abc_41234_new_n922_; 
wire _abc_41234_new_n923_; 
wire _abc_41234_new_n924_; 
wire _abc_41234_new_n925_; 
wire _abc_41234_new_n926_; 
wire _abc_41234_new_n927_; 
wire _abc_41234_new_n928_; 
wire _abc_41234_new_n929_; 
wire _abc_41234_new_n930_; 
wire _abc_41234_new_n931_; 
wire _abc_41234_new_n932_; 
wire _abc_41234_new_n933_; 
wire _abc_41234_new_n934_; 
wire _abc_41234_new_n935_; 
wire _abc_41234_new_n936_; 
wire _abc_41234_new_n937_; 
wire _abc_41234_new_n938_; 
wire _abc_41234_new_n940_; 
wire _abc_41234_new_n941_; 
wire _abc_41234_new_n942_; 
wire _abc_41234_new_n943_; 
wire _abc_41234_new_n944_; 
wire _abc_41234_new_n945_; 
wire _abc_41234_new_n946_; 
wire _abc_41234_new_n947_; 
wire _abc_41234_new_n948_; 
wire _abc_41234_new_n949_; 
wire _abc_41234_new_n950_; 
wire _abc_41234_new_n951_; 
wire _abc_41234_new_n952_; 
wire _abc_41234_new_n953_; 
wire _abc_41234_new_n954_; 
wire _abc_41234_new_n955_; 
wire _abc_41234_new_n956_; 
wire _abc_41234_new_n957_; 
wire _abc_41234_new_n958_; 
wire _abc_41234_new_n959_; 
wire _abc_41234_new_n960_; 
wire _abc_41234_new_n961_; 
wire _abc_41234_new_n962_; 
wire _abc_41234_new_n963_; 
wire _abc_41234_new_n964_; 
wire _abc_41234_new_n965_; 
wire _abc_41234_new_n966_; 
wire _abc_41234_new_n967_; 
wire _abc_41234_new_n968_; 
wire _abc_41234_new_n969_; 
wire _abc_41234_new_n970_; 
wire _abc_41234_new_n971_; 
wire _abc_41234_new_n972_; 
wire _abc_41234_new_n973_; 
wire _abc_41234_new_n974_; 
wire _abc_41234_new_n975_; 
wire _abc_41234_new_n976_; 
wire _abc_41234_new_n977_; 
wire _abc_41234_new_n978_; 
wire _abc_41234_new_n979_; 
wire _abc_41234_new_n980_; 
wire _abc_41234_new_n981_; 
wire _abc_41234_new_n983_; 
wire _abc_41234_new_n984_; 
wire _abc_41234_new_n985_; 
wire _abc_41234_new_n986_; 
wire _abc_41234_new_n987_; 
wire _abc_41234_new_n988_; 
wire _abc_41234_new_n989_; 
wire _abc_41234_new_n990_; 
wire _abc_41234_new_n991_; 
wire _abc_41234_new_n992_; 
wire _abc_41234_new_n993_; 
wire _abc_41234_new_n994_; 
wire _abc_41234_new_n995_; 
wire _abc_41234_new_n996_; 
wire _abc_41234_new_n997_; 
wire _abc_41234_new_n998_; 
wire _abc_41234_new_n999_; 
wire _auto_iopadmap_cc_368_execute_45628_0_; 
wire _auto_iopadmap_cc_368_execute_45628_10_; 
wire _auto_iopadmap_cc_368_execute_45628_11_; 
wire _auto_iopadmap_cc_368_execute_45628_12_; 
wire _auto_iopadmap_cc_368_execute_45628_13_; 
wire _auto_iopadmap_cc_368_execute_45628_14_; 
wire _auto_iopadmap_cc_368_execute_45628_15_; 
wire _auto_iopadmap_cc_368_execute_45628_1_; 
wire _auto_iopadmap_cc_368_execute_45628_2_; 
wire _auto_iopadmap_cc_368_execute_45628_3_; 
wire _auto_iopadmap_cc_368_execute_45628_4_; 
wire _auto_iopadmap_cc_368_execute_45628_5_; 
wire _auto_iopadmap_cc_368_execute_45628_6_; 
wire _auto_iopadmap_cc_368_execute_45628_7_; 
wire _auto_iopadmap_cc_368_execute_45628_8_; 
wire _auto_iopadmap_cc_368_execute_45628_9_; 
wire _auto_iopadmap_cc_368_execute_45645; 
wire _auto_iopadmap_cc_368_execute_45647; 
wire _auto_iopadmap_cc_368_execute_45649; 
wire _auto_iopadmap_cc_368_execute_45651; 
wire _auto_iopadmap_cc_368_execute_45653; 
output \addr[0] ;
output \addr[10] ;
output \addr[11] ;
output \addr[12] ;
output \addr[13] ;
output \addr[14] ;
output \addr[15] ;
output \addr[1] ;
output \addr[2] ;
output \addr[3] ;
output \addr[4] ;
output \addr[5] ;
output \addr[6] ;
output \addr[7] ;
output \addr[8] ;
output \addr[9] ;
wire alu__abc_40887_new_n100_; 
wire alu__abc_40887_new_n101_; 
wire alu__abc_40887_new_n102_; 
wire alu__abc_40887_new_n103_; 
wire alu__abc_40887_new_n104_; 
wire alu__abc_40887_new_n105_; 
wire alu__abc_40887_new_n106_; 
wire alu__abc_40887_new_n107_; 
wire alu__abc_40887_new_n108_; 
wire alu__abc_40887_new_n109_; 
wire alu__abc_40887_new_n110_; 
wire alu__abc_40887_new_n111_; 
wire alu__abc_40887_new_n112_; 
wire alu__abc_40887_new_n113_; 
wire alu__abc_40887_new_n114_; 
wire alu__abc_40887_new_n115_; 
wire alu__abc_40887_new_n116_; 
wire alu__abc_40887_new_n117_; 
wire alu__abc_40887_new_n118_; 
wire alu__abc_40887_new_n119_; 
wire alu__abc_40887_new_n120_; 
wire alu__abc_40887_new_n121_; 
wire alu__abc_40887_new_n122_; 
wire alu__abc_40887_new_n123_; 
wire alu__abc_40887_new_n124_; 
wire alu__abc_40887_new_n125_; 
wire alu__abc_40887_new_n126_; 
wire alu__abc_40887_new_n127_; 
wire alu__abc_40887_new_n128_; 
wire alu__abc_40887_new_n129_; 
wire alu__abc_40887_new_n130_; 
wire alu__abc_40887_new_n131_; 
wire alu__abc_40887_new_n132_; 
wire alu__abc_40887_new_n133_; 
wire alu__abc_40887_new_n134_; 
wire alu__abc_40887_new_n135_; 
wire alu__abc_40887_new_n136_; 
wire alu__abc_40887_new_n137_; 
wire alu__abc_40887_new_n138_; 
wire alu__abc_40887_new_n139_; 
wire alu__abc_40887_new_n140_; 
wire alu__abc_40887_new_n141_; 
wire alu__abc_40887_new_n142_; 
wire alu__abc_40887_new_n143_; 
wire alu__abc_40887_new_n144_; 
wire alu__abc_40887_new_n145_; 
wire alu__abc_40887_new_n146_; 
wire alu__abc_40887_new_n147_; 
wire alu__abc_40887_new_n148_; 
wire alu__abc_40887_new_n149_; 
wire alu__abc_40887_new_n150_; 
wire alu__abc_40887_new_n151_; 
wire alu__abc_40887_new_n152_; 
wire alu__abc_40887_new_n153_; 
wire alu__abc_40887_new_n154_; 
wire alu__abc_40887_new_n155_; 
wire alu__abc_40887_new_n156_; 
wire alu__abc_40887_new_n157_; 
wire alu__abc_40887_new_n158_; 
wire alu__abc_40887_new_n159_; 
wire alu__abc_40887_new_n160_; 
wire alu__abc_40887_new_n161_; 
wire alu__abc_40887_new_n162_; 
wire alu__abc_40887_new_n163_; 
wire alu__abc_40887_new_n164_; 
wire alu__abc_40887_new_n165_; 
wire alu__abc_40887_new_n166_; 
wire alu__abc_40887_new_n167_; 
wire alu__abc_40887_new_n168_; 
wire alu__abc_40887_new_n169_; 
wire alu__abc_40887_new_n170_; 
wire alu__abc_40887_new_n171_; 
wire alu__abc_40887_new_n172_; 
wire alu__abc_40887_new_n173_; 
wire alu__abc_40887_new_n174_; 
wire alu__abc_40887_new_n175_; 
wire alu__abc_40887_new_n176_; 
wire alu__abc_40887_new_n177_; 
wire alu__abc_40887_new_n178_; 
wire alu__abc_40887_new_n179_; 
wire alu__abc_40887_new_n180_; 
wire alu__abc_40887_new_n181_; 
wire alu__abc_40887_new_n182_; 
wire alu__abc_40887_new_n183_; 
wire alu__abc_40887_new_n184_; 
wire alu__abc_40887_new_n185_; 
wire alu__abc_40887_new_n186_; 
wire alu__abc_40887_new_n187_; 
wire alu__abc_40887_new_n188_; 
wire alu__abc_40887_new_n189_; 
wire alu__abc_40887_new_n190_; 
wire alu__abc_40887_new_n191_; 
wire alu__abc_40887_new_n192_; 
wire alu__abc_40887_new_n193_; 
wire alu__abc_40887_new_n194_; 
wire alu__abc_40887_new_n195_; 
wire alu__abc_40887_new_n196_; 
wire alu__abc_40887_new_n197_; 
wire alu__abc_40887_new_n198_; 
wire alu__abc_40887_new_n199_; 
wire alu__abc_40887_new_n200_; 
wire alu__abc_40887_new_n201_; 
wire alu__abc_40887_new_n202_; 
wire alu__abc_40887_new_n203_; 
wire alu__abc_40887_new_n204_; 
wire alu__abc_40887_new_n205_; 
wire alu__abc_40887_new_n206_; 
wire alu__abc_40887_new_n207_; 
wire alu__abc_40887_new_n208_; 
wire alu__abc_40887_new_n209_; 
wire alu__abc_40887_new_n210_; 
wire alu__abc_40887_new_n211_; 
wire alu__abc_40887_new_n212_; 
wire alu__abc_40887_new_n213_; 
wire alu__abc_40887_new_n214_; 
wire alu__abc_40887_new_n215_; 
wire alu__abc_40887_new_n217_; 
wire alu__abc_40887_new_n218_; 
wire alu__abc_40887_new_n219_; 
wire alu__abc_40887_new_n220_; 
wire alu__abc_40887_new_n221_; 
wire alu__abc_40887_new_n222_; 
wire alu__abc_40887_new_n223_; 
wire alu__abc_40887_new_n224_; 
wire alu__abc_40887_new_n225_; 
wire alu__abc_40887_new_n226_; 
wire alu__abc_40887_new_n227_; 
wire alu__abc_40887_new_n228_; 
wire alu__abc_40887_new_n229_; 
wire alu__abc_40887_new_n230_; 
wire alu__abc_40887_new_n231_; 
wire alu__abc_40887_new_n232_; 
wire alu__abc_40887_new_n233_; 
wire alu__abc_40887_new_n234_; 
wire alu__abc_40887_new_n235_; 
wire alu__abc_40887_new_n236_; 
wire alu__abc_40887_new_n237_; 
wire alu__abc_40887_new_n238_; 
wire alu__abc_40887_new_n239_; 
wire alu__abc_40887_new_n240_; 
wire alu__abc_40887_new_n241_; 
wire alu__abc_40887_new_n242_; 
wire alu__abc_40887_new_n243_; 
wire alu__abc_40887_new_n244_; 
wire alu__abc_40887_new_n245_; 
wire alu__abc_40887_new_n246_; 
wire alu__abc_40887_new_n247_; 
wire alu__abc_40887_new_n248_; 
wire alu__abc_40887_new_n249_; 
wire alu__abc_40887_new_n250_; 
wire alu__abc_40887_new_n251_; 
wire alu__abc_40887_new_n252_; 
wire alu__abc_40887_new_n253_; 
wire alu__abc_40887_new_n254_; 
wire alu__abc_40887_new_n255_; 
wire alu__abc_40887_new_n256_; 
wire alu__abc_40887_new_n257_; 
wire alu__abc_40887_new_n258_; 
wire alu__abc_40887_new_n259_; 
wire alu__abc_40887_new_n260_; 
wire alu__abc_40887_new_n261_; 
wire alu__abc_40887_new_n262_; 
wire alu__abc_40887_new_n263_; 
wire alu__abc_40887_new_n264_; 
wire alu__abc_40887_new_n265_; 
wire alu__abc_40887_new_n266_; 
wire alu__abc_40887_new_n267_; 
wire alu__abc_40887_new_n268_; 
wire alu__abc_40887_new_n269_; 
wire alu__abc_40887_new_n270_; 
wire alu__abc_40887_new_n271_; 
wire alu__abc_40887_new_n272_; 
wire alu__abc_40887_new_n273_; 
wire alu__abc_40887_new_n274_; 
wire alu__abc_40887_new_n275_; 
wire alu__abc_40887_new_n276_; 
wire alu__abc_40887_new_n277_; 
wire alu__abc_40887_new_n278_; 
wire alu__abc_40887_new_n279_; 
wire alu__abc_40887_new_n280_; 
wire alu__abc_40887_new_n281_; 
wire alu__abc_40887_new_n282_; 
wire alu__abc_40887_new_n283_; 
wire alu__abc_40887_new_n284_; 
wire alu__abc_40887_new_n285_; 
wire alu__abc_40887_new_n286_; 
wire alu__abc_40887_new_n287_; 
wire alu__abc_40887_new_n288_; 
wire alu__abc_40887_new_n289_; 
wire alu__abc_40887_new_n290_; 
wire alu__abc_40887_new_n291_; 
wire alu__abc_40887_new_n292_; 
wire alu__abc_40887_new_n293_; 
wire alu__abc_40887_new_n294_; 
wire alu__abc_40887_new_n295_; 
wire alu__abc_40887_new_n296_; 
wire alu__abc_40887_new_n297_; 
wire alu__abc_40887_new_n298_; 
wire alu__abc_40887_new_n299_; 
wire alu__abc_40887_new_n300_; 
wire alu__abc_40887_new_n301_; 
wire alu__abc_40887_new_n302_; 
wire alu__abc_40887_new_n303_; 
wire alu__abc_40887_new_n304_; 
wire alu__abc_40887_new_n305_; 
wire alu__abc_40887_new_n306_; 
wire alu__abc_40887_new_n307_; 
wire alu__abc_40887_new_n308_; 
wire alu__abc_40887_new_n309_; 
wire alu__abc_40887_new_n310_; 
wire alu__abc_40887_new_n311_; 
wire alu__abc_40887_new_n312_; 
wire alu__abc_40887_new_n313_; 
wire alu__abc_40887_new_n314_; 
wire alu__abc_40887_new_n315_; 
wire alu__abc_40887_new_n316_; 
wire alu__abc_40887_new_n317_; 
wire alu__abc_40887_new_n318_; 
wire alu__abc_40887_new_n319_; 
wire alu__abc_40887_new_n320_; 
wire alu__abc_40887_new_n321_; 
wire alu__abc_40887_new_n322_; 
wire alu__abc_40887_new_n323_; 
wire alu__abc_40887_new_n324_; 
wire alu__abc_40887_new_n325_; 
wire alu__abc_40887_new_n326_; 
wire alu__abc_40887_new_n327_; 
wire alu__abc_40887_new_n328_; 
wire alu__abc_40887_new_n329_; 
wire alu__abc_40887_new_n330_; 
wire alu__abc_40887_new_n331_; 
wire alu__abc_40887_new_n332_; 
wire alu__abc_40887_new_n333_; 
wire alu__abc_40887_new_n334_; 
wire alu__abc_40887_new_n335_; 
wire alu__abc_40887_new_n336_; 
wire alu__abc_40887_new_n337_; 
wire alu__abc_40887_new_n338_; 
wire alu__abc_40887_new_n339_; 
wire alu__abc_40887_new_n33_; 
wire alu__abc_40887_new_n340_; 
wire alu__abc_40887_new_n341_; 
wire alu__abc_40887_new_n342_; 
wire alu__abc_40887_new_n343_; 
wire alu__abc_40887_new_n344_; 
wire alu__abc_40887_new_n345_; 
wire alu__abc_40887_new_n346_; 
wire alu__abc_40887_new_n347_; 
wire alu__abc_40887_new_n348_; 
wire alu__abc_40887_new_n34_; 
wire alu__abc_40887_new_n350_; 
wire alu__abc_40887_new_n351_; 
wire alu__abc_40887_new_n352_; 
wire alu__abc_40887_new_n354_; 
wire alu__abc_40887_new_n356_; 
wire alu__abc_40887_new_n358_; 
wire alu__abc_40887_new_n35_; 
wire alu__abc_40887_new_n360_; 
wire alu__abc_40887_new_n362_; 
wire alu__abc_40887_new_n365_; 
wire alu__abc_40887_new_n367_; 
wire alu__abc_40887_new_n368_; 
wire alu__abc_40887_new_n36_; 
wire alu__abc_40887_new_n370_; 
wire alu__abc_40887_new_n371_; 
wire alu__abc_40887_new_n372_; 
wire alu__abc_40887_new_n373_; 
wire alu__abc_40887_new_n374_; 
wire alu__abc_40887_new_n375_; 
wire alu__abc_40887_new_n376_; 
wire alu__abc_40887_new_n377_; 
wire alu__abc_40887_new_n37_; 
wire alu__abc_40887_new_n38_; 
wire alu__abc_40887_new_n39_; 
wire alu__abc_40887_new_n40_; 
wire alu__abc_40887_new_n41_; 
wire alu__abc_40887_new_n42_; 
wire alu__abc_40887_new_n43_; 
wire alu__abc_40887_new_n44_; 
wire alu__abc_40887_new_n45_; 
wire alu__abc_40887_new_n46_; 
wire alu__abc_40887_new_n47_; 
wire alu__abc_40887_new_n48_; 
wire alu__abc_40887_new_n49_; 
wire alu__abc_40887_new_n50_; 
wire alu__abc_40887_new_n51_; 
wire alu__abc_40887_new_n52_; 
wire alu__abc_40887_new_n53_; 
wire alu__abc_40887_new_n54_; 
wire alu__abc_40887_new_n55_; 
wire alu__abc_40887_new_n56_; 
wire alu__abc_40887_new_n57_; 
wire alu__abc_40887_new_n58_; 
wire alu__abc_40887_new_n59_; 
wire alu__abc_40887_new_n60_; 
wire alu__abc_40887_new_n61_; 
wire alu__abc_40887_new_n62_; 
wire alu__abc_40887_new_n63_; 
wire alu__abc_40887_new_n64_; 
wire alu__abc_40887_new_n65_; 
wire alu__abc_40887_new_n66_; 
wire alu__abc_40887_new_n67_; 
wire alu__abc_40887_new_n68_; 
wire alu__abc_40887_new_n69_; 
wire alu__abc_40887_new_n70_; 
wire alu__abc_40887_new_n71_; 
wire alu__abc_40887_new_n72_; 
wire alu__abc_40887_new_n73_; 
wire alu__abc_40887_new_n74_; 
wire alu__abc_40887_new_n75_; 
wire alu__abc_40887_new_n76_; 
wire alu__abc_40887_new_n77_; 
wire alu__abc_40887_new_n78_; 
wire alu__abc_40887_new_n79_; 
wire alu__abc_40887_new_n80_; 
wire alu__abc_40887_new_n81_; 
wire alu__abc_40887_new_n82_; 
wire alu__abc_40887_new_n83_; 
wire alu__abc_40887_new_n84_; 
wire alu__abc_40887_new_n85_; 
wire alu__abc_40887_new_n86_; 
wire alu__abc_40887_new_n87_; 
wire alu__abc_40887_new_n88_; 
wire alu__abc_40887_new_n89_; 
wire alu__abc_40887_new_n90_; 
wire alu__abc_40887_new_n91_; 
wire alu__abc_40887_new_n92_; 
wire alu__abc_40887_new_n93_; 
wire alu__abc_40887_new_n94_; 
wire alu__abc_40887_new_n95_; 
wire alu__abc_40887_new_n96_; 
wire alu__abc_40887_new_n97_; 
wire alu__abc_40887_new_n98_; 
wire alu__abc_40887_new_n99_; 
wire alu_cin; 
wire alu_cout; 
wire alu_opra_0_; 
wire alu_opra_1_; 
wire alu_opra_2_; 
wire alu_opra_3_; 
wire alu_opra_4_; 
wire alu_opra_5_; 
wire alu_opra_6_; 
wire alu_opra_7_; 
wire alu_oprb_0_; 
wire alu_oprb_1_; 
wire alu_oprb_2_; 
wire alu_oprb_3_; 
wire alu_oprb_4_; 
wire alu_oprb_5_; 
wire alu_oprb_6_; 
wire alu_oprb_7_; 
wire alu_parity; 
wire alu_res_0_; 
wire alu_res_1_; 
wire alu_res_2_; 
wire alu_res_3_; 
wire alu_res_4_; 
wire alu_res_5_; 
wire alu_res_6_; 
wire alu_res_7_; 
wire alu_sel_0_; 
wire alu_sel_1_; 
wire alu_sel_2_; 
wire alu_sout; 
wire alu_zout; 
wire auxcar; 
wire carry; 
input clock;
wire clock_bF_buf0; 
wire clock_bF_buf1; 
wire clock_bF_buf10; 
wire clock_bF_buf11; 
wire clock_bF_buf12; 
wire clock_bF_buf13; 
wire clock_bF_buf13_bF_buf0; 
wire clock_bF_buf13_bF_buf1; 
wire clock_bF_buf13_bF_buf2; 
wire clock_bF_buf13_bF_buf3; 
wire clock_bF_buf14; 
wire clock_bF_buf14_bF_buf0; 
wire clock_bF_buf14_bF_buf1; 
wire clock_bF_buf14_bF_buf2; 
wire clock_bF_buf14_bF_buf3; 
wire clock_bF_buf2; 
wire clock_bF_buf3; 
wire clock_bF_buf4; 
wire clock_bF_buf5; 
wire clock_bF_buf6; 
wire clock_bF_buf7; 
wire clock_bF_buf8; 
wire clock_bF_buf9; 
input \data[0] ;
input \data[1] ;
input \data[2] ;
input \data[3] ;
input \data[4] ;
input \data[5] ;
input \data[6] ;
input \data[7] ;
wire ei; 
wire eienb; 
output inta;
wire intcyc; 
wire intcyc_bF_buf0; 
wire intcyc_bF_buf1; 
wire intcyc_bF_buf2; 
wire intcyc_bF_buf3; 
input intr;
wire opcode_0_; 
wire opcode_1_; 
wire opcode_2_; 
wire opcode_3_; 
wire opcode_3_bF_buf0_; 
wire opcode_3_bF_buf1_; 
wire opcode_3_bF_buf2_; 
wire opcode_3_bF_buf3_; 
wire opcode_4_; 
wire opcode_4_bF_buf0_; 
wire opcode_4_bF_buf1_; 
wire opcode_4_bF_buf2_; 
wire opcode_4_bF_buf3_; 
wire opcode_4_bF_buf4_; 
wire opcode_4_bF_buf5_; 
wire opcode_4_bF_buf6_; 
wire opcode_5_; 
wire opcode_5_bF_buf0_; 
wire opcode_5_bF_buf1_; 
wire opcode_5_bF_buf2_; 
wire opcode_5_bF_buf3_; 
wire opcode_5_bF_buf4_; 
wire opcode_6_; 
wire opcode_7_; 
wire parity; 
wire pc_0_; 
wire pc_10_; 
wire pc_11_; 
wire pc_12_; 
wire pc_13_; 
wire pc_14_; 
wire pc_15_; 
wire pc_1_; 
wire pc_2_; 
wire pc_3_; 
wire pc_4_; 
wire pc_5_; 
wire pc_6_; 
wire pc_7_; 
wire pc_8_; 
wire pc_9_; 
wire popdes_0_; 
wire popdes_1_; 
wire raddrhold_0_; 
wire raddrhold_10_; 
wire raddrhold_11_; 
wire raddrhold_12_; 
wire raddrhold_13_; 
wire raddrhold_14_; 
wire raddrhold_15_; 
wire raddrhold_1_; 
wire raddrhold_2_; 
wire raddrhold_3_; 
wire raddrhold_4_; 
wire raddrhold_5_; 
wire raddrhold_6_; 
wire raddrhold_7_; 
wire raddrhold_8_; 
wire raddrhold_9_; 
wire rdatahold2_0_; 
wire rdatahold2_1_; 
wire rdatahold2_2_; 
wire rdatahold2_3_; 
wire rdatahold2_4_; 
wire rdatahold2_5_; 
wire rdatahold2_6_; 
wire rdatahold2_7_; 
wire rdatahold_0_; 
wire rdatahold_1_; 
wire rdatahold_2_; 
wire rdatahold_3_; 
wire rdatahold_4_; 
wire rdatahold_5_; 
wire rdatahold_6_; 
wire rdatahold_7_; 
output readio;
output readmem;
wire regd_0_; 
wire regd_1_; 
wire regd_2_; 
wire regfil_0__0_; 
wire regfil_0__1_; 
wire regfil_0__2_; 
wire regfil_0__3_; 
wire regfil_0__4_; 
wire regfil_0__5_; 
wire regfil_0__6_; 
wire regfil_0__7_; 
wire regfil_1__0_; 
wire regfil_1__1_; 
wire regfil_1__2_; 
wire regfil_1__3_; 
wire regfil_1__4_; 
wire regfil_1__5_; 
wire regfil_1__6_; 
wire regfil_1__7_; 
wire regfil_2__0_; 
wire regfil_2__1_; 
wire regfil_2__2_; 
wire regfil_2__3_; 
wire regfil_2__4_; 
wire regfil_2__5_; 
wire regfil_2__6_; 
wire regfil_2__7_; 
wire regfil_3__0_; 
wire regfil_3__1_; 
wire regfil_3__2_; 
wire regfil_3__3_; 
wire regfil_3__4_; 
wire regfil_3__5_; 
wire regfil_3__6_; 
wire regfil_3__7_; 
wire regfil_4__0_; 
wire regfil_4__1_; 
wire regfil_4__1_bF_buf0_; 
wire regfil_4__1_bF_buf1_; 
wire regfil_4__1_bF_buf2_; 
wire regfil_4__1_bF_buf3_; 
wire regfil_4__2_; 
wire regfil_4__2_bF_buf0_; 
wire regfil_4__2_bF_buf1_; 
wire regfil_4__2_bF_buf2_; 
wire regfil_4__2_bF_buf3_; 
wire regfil_4__3_; 
wire regfil_4__4_; 
wire regfil_4__5_; 
wire regfil_4__6_; 
wire regfil_4__7_; 
wire regfil_5__0_; 
wire regfil_5__1_; 
wire regfil_5__2_; 
wire regfil_5__3_; 
wire regfil_5__3_bF_buf0_; 
wire regfil_5__3_bF_buf1_; 
wire regfil_5__3_bF_buf2_; 
wire regfil_5__3_bF_buf3_; 
wire regfil_5__4_; 
wire regfil_5__5_; 
wire regfil_5__6_; 
wire regfil_5__6_bF_buf0_; 
wire regfil_5__6_bF_buf1_; 
wire regfil_5__6_bF_buf2_; 
wire regfil_5__6_bF_buf3_; 
wire regfil_5__7_; 
wire regfil_6__0_; 
wire regfil_6__1_; 
wire regfil_6__2_; 
wire regfil_6__3_; 
wire regfil_6__4_; 
wire regfil_6__5_; 
wire regfil_6__6_; 
wire regfil_6__7_; 
wire regfil_7__0_; 
wire regfil_7__1_; 
wire regfil_7__2_; 
wire regfil_7__3_; 
wire regfil_7__4_; 
wire regfil_7__5_; 
wire regfil_7__6_; 
wire regfil_7__7_; 
input reset;
wire reset_bF_buf0; 
wire reset_bF_buf1; 
wire reset_bF_buf2; 
wire reset_bF_buf3; 
wire reset_bF_buf4; 
wire reset_bF_buf5; 
wire reset_bF_buf6; 
wire reset_bF_buf7; 
wire reset_bF_buf8; 
wire reset_bF_buf9; 
wire sign; 
wire sp_0_; 
wire sp_0_bF_buf0_; 
wire sp_0_bF_buf1_; 
wire sp_0_bF_buf2_; 
wire sp_0_bF_buf3_; 
wire sp_10_; 
wire sp_11_; 
wire sp_12_; 
wire sp_13_; 
wire sp_14_; 
wire sp_15_; 
wire sp_1_; 
wire sp_2_; 
wire sp_3_; 
wire sp_4_; 
wire sp_5_; 
wire sp_6_; 
wire sp_7_; 
wire sp_8_; 
wire sp_9_; 
wire state_0_; 
wire state_1_; 
wire state_2_; 
wire state_3_; 
wire state_4_; 
wire state_5_; 
wire statesel_0_; 
wire statesel_1_; 
wire statesel_2_; 
wire statesel_3_; 
wire statesel_4_; 
wire statesel_5_; 
wire waddrhold_0_; 
wire waddrhold_10_; 
wire waddrhold_11_; 
wire waddrhold_12_; 
wire waddrhold_13_; 
wire waddrhold_14_; 
wire waddrhold_15_; 
wire waddrhold_1_; 
wire waddrhold_2_; 
wire waddrhold_3_; 
wire waddrhold_4_; 
wire waddrhold_5_; 
wire waddrhold_6_; 
wire waddrhold_7_; 
wire waddrhold_8_; 
wire waddrhold_9_; 
input waitr;
wire wdatahold2_0_; 
wire wdatahold2_1_; 
wire wdatahold2_2_; 
wire wdatahold2_3_; 
wire wdatahold2_4_; 
wire wdatahold2_5_; 
wire wdatahold2_6_; 
wire wdatahold2_7_; 
wire wdatahold_0_; 
wire wdatahold_1_; 
wire wdatahold_2_; 
wire wdatahold_3_; 
wire wdatahold_4_; 
wire wdatahold_5_; 
wire wdatahold_6_; 
wire wdatahold_7_; 
output writeio;
output writemem;
wire zero; 
AND2X2 AND2X2_1 ( .A(_abc_41234_new_n789_), .B(_abc_41234_new_n765_), .Y(_abc_41234_new_n790_));
AND2X2 AND2X2_10 ( .A(_abc_41234_new_n1153_), .B(_abc_41234_new_n1149_), .Y(_abc_41234_new_n1154_));
AND2X2 AND2X2_100 ( .A(alu_oprb_2_), .B(alu_opra_2_), .Y(alu__abc_40887_new_n47_));
AND2X2 AND2X2_101 ( .A(alu_oprb_3_), .B(alu_opra_3_), .Y(alu__abc_40887_new_n50_));
AND2X2 AND2X2_102 ( .A(alu__abc_40887_new_n57_), .B(alu__abc_40887_new_n56_), .Y(alu__abc_40887_new_n58_));
AND2X2 AND2X2_103 ( .A(alu__abc_40887_new_n53_), .B(alu__abc_40887_new_n55_), .Y(alu__abc_40887_new_n78_));
AND2X2 AND2X2_104 ( .A(alu__abc_40887_new_n46_), .B(alu__abc_40887_new_n49_), .Y(alu__abc_40887_new_n82_));
AND2X2 AND2X2_105 ( .A(alu__abc_40887_new_n98_), .B(alu__abc_40887_new_n75_), .Y(alu__abc_40887_new_n99_));
AND2X2 AND2X2_106 ( .A(alu__abc_40887_new_n117_), .B(alu__abc_40887_new_n115_), .Y(alu__abc_40887_new_n118_));
AND2X2 AND2X2_107 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_40887_new_n127_));
AND2X2 AND2X2_108 ( .A(alu__abc_40887_new_n161_), .B(alu__abc_40887_new_n164_), .Y(alu__abc_40887_new_n287_));
AND2X2 AND2X2_109 ( .A(alu__abc_40887_new_n263_), .B(alu__abc_40887_new_n265_), .Y(alu__abc_40887_new_n292_));
AND2X2 AND2X2_11 ( .A(regfil_1__3_), .B(regfil_5__3_bF_buf3_), .Y(_abc_41234_new_n1161_));
AND2X2 AND2X2_110 ( .A(alu_sout), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n345_));
AND2X2 AND2X2_111 ( .A(alu__abc_40887_new_n352_), .B(alu__abc_40887_new_n344_), .Y(alu_zout));
AND2X2 AND2X2_12 ( .A(regfil_1__2_), .B(regfil_5__2_), .Y(_abc_41234_new_n1164_));
AND2X2 AND2X2_13 ( .A(regfil_1__7_), .B(regfil_5__7_), .Y(_abc_41234_new_n1171_));
AND2X2 AND2X2_14 ( .A(regfil_1__6_), .B(regfil_5__6_bF_buf2_), .Y(_abc_41234_new_n1174_));
AND2X2 AND2X2_15 ( .A(regfil_1__4_), .B(regfil_5__4_), .Y(_abc_41234_new_n1178_));
AND2X2 AND2X2_16 ( .A(regfil_1__5_), .B(regfil_5__5_), .Y(_abc_41234_new_n1181_));
AND2X2 AND2X2_17 ( .A(_abc_41234_new_n1241_), .B(_abc_41234_new_n1242_), .Y(_abc_41234_new_n1243_));
AND2X2 AND2X2_18 ( .A(_abc_41234_new_n1282_), .B(_abc_41234_new_n1263_), .Y(_abc_41234_new_n1283_));
AND2X2 AND2X2_19 ( .A(_abc_41234_new_n1374_), .B(_abc_41234_new_n1378_), .Y(_abc_41234_new_n1379_));
AND2X2 AND2X2_2 ( .A(_abc_41234_new_n920_), .B(_abc_41234_new_n631_), .Y(_abc_41234_new_n921_));
AND2X2 AND2X2_20 ( .A(_abc_41234_new_n1406_), .B(_abc_41234_new_n1410_), .Y(_abc_41234_new_n1411_));
AND2X2 AND2X2_21 ( .A(_abc_41234_new_n1433_), .B(_abc_41234_new_n1427_), .Y(_abc_41234_new_n1434_));
AND2X2 AND2X2_22 ( .A(_abc_41234_new_n1438_), .B(_abc_41234_new_n1263_), .Y(_abc_41234_new_n1439_));
AND2X2 AND2X2_23 ( .A(_abc_41234_new_n1461_), .B(_abc_41234_new_n1409_), .Y(_abc_41234_new_n1465_));
AND2X2 AND2X2_24 ( .A(_abc_41234_new_n1464_), .B(_abc_41234_new_n1466_), .Y(_abc_41234_new_n1467_));
AND2X2 AND2X2_25 ( .A(_abc_41234_new_n1513_), .B(_abc_41234_new_n1514_), .Y(_abc_41234_new_n1515_));
AND2X2 AND2X2_26 ( .A(_abc_41234_new_n1533_), .B(_abc_41234_new_n1538_), .Y(_abc_41234_new_n1540_));
AND2X2 AND2X2_27 ( .A(_abc_41234_new_n1621_), .B(_abc_41234_new_n1623_), .Y(_abc_41234_new_n1624_));
AND2X2 AND2X2_28 ( .A(_abc_41234_new_n1678_), .B(_abc_41234_new_n1679_), .Y(_abc_41234_new_n1680_));
AND2X2 AND2X2_29 ( .A(_abc_41234_new_n1715_), .B(_abc_41234_new_n1714_), .Y(_abc_41234_new_n1716_));
AND2X2 AND2X2_3 ( .A(_abc_41234_new_n942_), .B(_abc_41234_new_n941_), .Y(_abc_41234_new_n943_));
AND2X2 AND2X2_30 ( .A(_abc_41234_new_n1751_), .B(_abc_41234_new_n1749_), .Y(_abc_41234_new_n1752_));
AND2X2 AND2X2_31 ( .A(_abc_41234_new_n1779_), .B(_abc_41234_new_n1778_), .Y(_abc_41234_new_n1780_));
AND2X2 AND2X2_32 ( .A(_abc_41234_new_n1781_), .B(_abc_41234_new_n1785_), .Y(_abc_41234_new_n1786_));
AND2X2 AND2X2_33 ( .A(_abc_41234_new_n1797_), .B(_abc_41234_new_n1799_), .Y(_abc_41234_new_n1800_));
AND2X2 AND2X2_34 ( .A(_abc_41234_new_n1834_), .B(_abc_41234_new_n1838_), .Y(_abc_41234_new_n1839_));
AND2X2 AND2X2_35 ( .A(_abc_41234_new_n594_), .B(_abc_41234_new_n1879_), .Y(_abc_41234_new_n1880_));
AND2X2 AND2X2_36 ( .A(_abc_41234_new_n1888_), .B(_abc_41234_new_n1889_), .Y(_abc_41234_new_n1890_));
AND2X2 AND2X2_37 ( .A(_abc_41234_new_n535_), .B(_abc_41234_new_n1954_), .Y(_abc_41234_new_n1955_));
AND2X2 AND2X2_38 ( .A(_abc_41234_new_n1940_), .B(_abc_41234_new_n992_), .Y(_abc_41234_new_n1956_));
AND2X2 AND2X2_39 ( .A(_abc_41234_new_n572_), .B(_abc_41234_new_n1986_), .Y(_abc_41234_new_n1987_));
AND2X2 AND2X2_4 ( .A(_abc_41234_new_n978_), .B(_abc_41234_new_n979_), .Y(_abc_41234_new_n980_));
AND2X2 AND2X2_40 ( .A(_abc_41234_new_n1995_), .B(_abc_41234_new_n1996_), .Y(_abc_41234_new_n1997_));
AND2X2 AND2X2_41 ( .A(_abc_41234_new_n2009_), .B(_abc_41234_new_n2010_), .Y(_abc_41234_new_n2011_));
AND2X2 AND2X2_42 ( .A(_abc_41234_new_n2063_), .B(_abc_41234_new_n2059_), .Y(_abc_41234_new_n2064_));
AND2X2 AND2X2_43 ( .A(_abc_41234_new_n2073_), .B(_abc_41234_new_n2072_), .Y(_abc_41234_new_n2074_));
AND2X2 AND2X2_44 ( .A(_abc_41234_new_n2087_), .B(_abc_41234_new_n2084_), .Y(_abc_41234_new_n2088_));
AND2X2 AND2X2_45 ( .A(_abc_41234_new_n2100_), .B(_abc_41234_new_n1049__bF_buf0), .Y(_abc_41234_new_n2101_));
AND2X2 AND2X2_46 ( .A(_abc_41234_new_n2140_), .B(_abc_41234_new_n2141_), .Y(_abc_41234_new_n2142_));
AND2X2 AND2X2_47 ( .A(_abc_41234_new_n1953_), .B(_abc_41234_new_n2142_), .Y(_abc_41234_new_n2143_));
AND2X2 AND2X2_48 ( .A(_abc_41234_new_n2163_), .B(regfil_2__7_), .Y(_abc_41234_new_n2164_));
AND2X2 AND2X2_49 ( .A(_abc_41234_new_n507_), .B(_abc_41234_new_n692_), .Y(_abc_41234_new_n2261_));
AND2X2 AND2X2_5 ( .A(_abc_41234_new_n975_), .B(_abc_41234_new_n980_), .Y(_abc_41234_new_n981_));
AND2X2 AND2X2_50 ( .A(_abc_41234_new_n2417_), .B(_abc_41234_new_n2424_), .Y(_abc_41234_new_n2425_));
AND2X2 AND2X2_51 ( .A(_abc_41234_new_n2523_), .B(_abc_41234_new_n2517_), .Y(_abc_41234_new_n2524_));
AND2X2 AND2X2_52 ( .A(_abc_41234_new_n2546_), .B(_abc_41234_new_n2467_), .Y(_abc_41234_new_n2547_));
AND2X2 AND2X2_53 ( .A(_abc_41234_new_n2709_), .B(_abc_41234_new_n2715_), .Y(_abc_41234_new_n2716_));
AND2X2 AND2X2_54 ( .A(_abc_41234_new_n2726_), .B(_abc_41234_new_n2728_), .Y(_abc_41234_new_n2729_));
AND2X2 AND2X2_55 ( .A(_abc_41234_new_n2733_), .B(_abc_41234_new_n2734_), .Y(_abc_41234_new_n2735_));
AND2X2 AND2X2_56 ( .A(_abc_41234_new_n2759_), .B(_abc_41234_new_n2761_), .Y(_abc_41234_new_n2762_));
AND2X2 AND2X2_57 ( .A(_abc_41234_new_n2772_), .B(_abc_41234_new_n1649_), .Y(_abc_41234_new_n2773_));
AND2X2 AND2X2_58 ( .A(_abc_41234_new_n1616_), .B(_abc_41234_new_n2775_), .Y(_abc_41234_new_n2776_));
AND2X2 AND2X2_59 ( .A(_abc_41234_new_n2815_), .B(_abc_41234_new_n2808_), .Y(_abc_41234_new_n2816_));
AND2X2 AND2X2_6 ( .A(_abc_41234_new_n1014_), .B(_abc_41234_new_n689_), .Y(_abc_41234_new_n1015_));
AND2X2 AND2X2_60 ( .A(_abc_41234_new_n2975_), .B(_abc_41234_new_n2982_), .Y(_abc_41234_new_n2983_));
AND2X2 AND2X2_61 ( .A(_abc_41234_new_n3112_), .B(_abc_41234_new_n3117_), .Y(_abc_41234_new_n3118_));
AND2X2 AND2X2_62 ( .A(_abc_41234_new_n3136_), .B(_abc_41234_new_n3141_), .Y(_abc_41234_new_n3142_));
AND2X2 AND2X2_63 ( .A(_abc_41234_new_n3161_), .B(_abc_41234_new_n3166_), .Y(_abc_41234_new_n3167_));
AND2X2 AND2X2_64 ( .A(_abc_41234_new_n3309_), .B(raddrhold_14_), .Y(_abc_41234_new_n3311_));
AND2X2 AND2X2_65 ( .A(_abc_41234_new_n3374_), .B(_abc_41234_new_n3375_), .Y(_abc_41234_new_n3376_));
AND2X2 AND2X2_66 ( .A(_abc_41234_new_n3397_), .B(_abc_41234_new_n3396_), .Y(_abc_41234_new_n3398_));
AND2X2 AND2X2_67 ( .A(_abc_41234_new_n3632_), .B(waddrhold_13_), .Y(_abc_41234_new_n3633_));
AND2X2 AND2X2_68 ( .A(_abc_41234_new_n3731_), .B(_abc_41234_new_n3753_), .Y(_abc_41234_new_n3754_));
AND2X2 AND2X2_69 ( .A(_abc_41234_new_n1325_), .B(_abc_41234_new_n3788_), .Y(_abc_41234_new_n3789_));
AND2X2 AND2X2_7 ( .A(regfil_5__3_bF_buf1_), .B(regfil_3__3_), .Y(_abc_41234_new_n1112_));
AND2X2 AND2X2_70 ( .A(_abc_41234_new_n1229_), .B(_abc_41234_new_n903_), .Y(_abc_41234_new_n3846_));
AND2X2 AND2X2_71 ( .A(_abc_41234_new_n3866_), .B(_abc_41234_new_n3864_), .Y(_abc_41234_new_n3867_));
AND2X2 AND2X2_72 ( .A(_abc_41234_new_n1214_), .B(_abc_41234_new_n3885_), .Y(_abc_41234_new_n3886_));
AND2X2 AND2X2_73 ( .A(_abc_41234_new_n3944_), .B(_abc_41234_new_n3946_), .Y(_abc_41234_new_n3947_));
AND2X2 AND2X2_74 ( .A(_abc_41234_new_n3969_), .B(_abc_41234_new_n3970_), .Y(_abc_41234_new_n3971_));
AND2X2 AND2X2_75 ( .A(_abc_41234_new_n3984_), .B(_abc_41234_new_n3987_), .Y(_abc_41234_new_n3988_));
AND2X2 AND2X2_76 ( .A(_abc_41234_new_n4014_), .B(_abc_41234_new_n4015_), .Y(_abc_41234_new_n4016_));
AND2X2 AND2X2_77 ( .A(_abc_41234_new_n4016_), .B(_abc_41234_new_n2462_), .Y(_abc_41234_new_n4017_));
AND2X2 AND2X2_78 ( .A(_abc_41234_new_n4080_), .B(_abc_41234_new_n4081_), .Y(_abc_41234_new_n4082_));
AND2X2 AND2X2_79 ( .A(_abc_41234_new_n4085_), .B(_abc_41234_new_n4083_), .Y(_abc_41234_new_n4086_));
AND2X2 AND2X2_8 ( .A(regfil_5__7_), .B(regfil_3__7_), .Y(_abc_41234_new_n1125_));
AND2X2 AND2X2_80 ( .A(_abc_41234_new_n4088_), .B(_abc_41234_new_n3936_), .Y(_abc_41234_new_n4089_));
AND2X2 AND2X2_81 ( .A(_abc_41234_new_n4102_), .B(_abc_41234_new_n4113_), .Y(_abc_41234_new_n4114_));
AND2X2 AND2X2_82 ( .A(_abc_41234_new_n4116_), .B(_abc_41234_new_n4117_), .Y(_abc_41234_new_n4118_));
AND2X2 AND2X2_83 ( .A(_abc_41234_new_n4132_), .B(_abc_41234_new_n4131_), .Y(_abc_41234_new_n4133_));
AND2X2 AND2X2_84 ( .A(_abc_41234_new_n4162_), .B(_abc_41234_new_n4166_), .Y(_abc_41234_new_n4167_));
AND2X2 AND2X2_85 ( .A(_abc_41234_new_n4189_), .B(_abc_41234_new_n4197_), .Y(_abc_41234_new_n4198_));
AND2X2 AND2X2_86 ( .A(_abc_41234_new_n4286_), .B(_abc_41234_new_n1640_), .Y(_abc_41234_new_n4287_));
AND2X2 AND2X2_87 ( .A(_abc_41234_new_n2471_), .B(_abc_41234_new_n4288_), .Y(_abc_41234_new_n4289_));
AND2X2 AND2X2_88 ( .A(_abc_41234_new_n4287_), .B(_abc_41234_new_n4289_), .Y(_abc_41234_new_n4290_));
AND2X2 AND2X2_89 ( .A(_abc_41234_new_n4408_), .B(_abc_41234_new_n4409_), .Y(_abc_41234_new_n4410_));
AND2X2 AND2X2_9 ( .A(regfil_5__6_bF_buf0_), .B(regfil_3__6_), .Y(_abc_41234_new_n1128_));
AND2X2 AND2X2_90 ( .A(_abc_41234_new_n1680_), .B(_abc_41234_new_n1606_), .Y(_abc_41234_new_n4463_));
AND2X2 AND2X2_91 ( .A(_abc_41234_new_n4481_), .B(_abc_41234_new_n4482_), .Y(_abc_41234_new_n4483_));
AND2X2 AND2X2_92 ( .A(_abc_41234_new_n1728_), .B(_abc_41234_new_n4309_), .Y(_abc_41234_new_n4509_));
AND2X2 AND2X2_93 ( .A(_abc_41234_new_n1752_), .B(_abc_41234_new_n4309_), .Y(_abc_41234_new_n4525_));
AND2X2 AND2X2_94 ( .A(_abc_41234_new_n1774_), .B(_abc_41234_new_n4309_), .Y(_abc_41234_new_n4545_));
AND2X2 AND2X2_95 ( .A(_abc_41234_new_n1800_), .B(_abc_41234_new_n4309_), .Y(_abc_41234_new_n4566_));
AND2X2 AND2X2_96 ( .A(_abc_41234_new_n4852_), .B(_abc_41234_new_n4851_), .Y(_abc_41234_new_n4853_));
AND2X2 AND2X2_97 ( .A(_abc_41234_new_n4864_), .B(_abc_41234_new_n4861_), .Y(_abc_41234_new_n4865_));
AND2X2 AND2X2_98 ( .A(_abc_41234_new_n4885_), .B(_abc_41234_new_n4886_), .Y(_abc_41234_new_n4887_));
AND2X2 AND2X2_99 ( .A(_abc_41234_new_n4891_), .B(_abc_41234_new_n516__bF_buf0), .Y(_abc_41234_new_n4892_));
AOI21X1 AOI21X1_1 ( .A(_abc_41234_new_n559_), .B(_abc_41234_new_n562_), .C(_abc_41234_new_n533_), .Y(_abc_41234_new_n563_));
AOI21X1 AOI21X1_10 ( .A(_abc_41234_new_n743_), .B(_abc_41234_new_n766_), .C(_abc_41234_new_n805_), .Y(_abc_41234_new_n808_));
AOI21X1 AOI21X1_100 ( .A(_abc_41234_new_n1644_), .B(_abc_41234_new_n1821_), .C(_abc_41234_new_n1047__bF_buf3), .Y(_abc_41234_new_n1843_));
AOI21X1 AOI21X1_101 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n1848_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n1860_));
AOI21X1 AOI21X1_102 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n730_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n1868_));
AOI21X1 AOI21X1_103 ( .A(_abc_41234_new_n1875_), .B(_abc_41234_new_n1872_), .C(_abc_41234_new_n1066__bF_buf0), .Y(_abc_41234_new_n1876_));
AOI21X1 AOI21X1_104 ( .A(_abc_41234_new_n1066__bF_buf3), .B(_abc_41234_new_n719_), .C(_abc_41234_new_n1880_), .Y(_abc_41234_new_n1881_));
AOI21X1 AOI21X1_105 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n768_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n1884_));
AOI21X1 AOI21X1_106 ( .A(regfil_5__2_), .B(_abc_41234_new_n1066__bF_buf2), .C(_abc_41234_new_n1894_), .Y(_abc_41234_new_n1895_));
AOI21X1 AOI21X1_107 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n814_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n1897_));
AOI21X1 AOI21X1_108 ( .A(regfil_5__3_bF_buf2_), .B(_abc_41234_new_n1066__bF_buf1), .C(_abc_41234_new_n1905_), .Y(_abc_41234_new_n1906_));
AOI21X1 AOI21X1_109 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n858_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n1908_));
AOI21X1 AOI21X1_11 ( .A(_abc_41234_new_n784_), .B(regfil_0__3_), .C(_abc_41234_new_n584_), .Y(_abc_41234_new_n810_));
AOI21X1 AOI21X1_110 ( .A(regfil_5__4_), .B(_abc_41234_new_n1066__bF_buf0), .C(_abc_41234_new_n1919_), .Y(_abc_41234_new_n1920_));
AOI21X1 AOI21X1_111 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n899_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n1922_));
AOI21X1 AOI21X1_112 ( .A(regfil_5__5_), .B(_abc_41234_new_n1066__bF_buf3), .C(_abc_41234_new_n1933_), .Y(_abc_41234_new_n1934_));
AOI21X1 AOI21X1_113 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n1936_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n1937_));
AOI21X1 AOI21X1_114 ( .A(regfil_5__6_bF_buf2_), .B(_abc_41234_new_n1066__bF_buf2), .C(_abc_41234_new_n1946_), .Y(_abc_41234_new_n1947_));
AOI21X1 AOI21X1_115 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n992_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n1949_));
AOI21X1 AOI21X1_116 ( .A(_abc_41234_new_n1066__bF_buf1), .B(_abc_41234_new_n996_), .C(_abc_41234_new_n1853_), .Y(_abc_41234_new_n1952_));
AOI21X1 AOI21X1_117 ( .A(_abc_41234_new_n1967_), .B(_abc_41234_new_n569_), .C(_abc_41234_new_n648_), .Y(_abc_41234_new_n1968_));
AOI21X1 AOI21X1_118 ( .A(_abc_41234_new_n1967_), .B(_abc_41234_new_n570_), .C(_abc_41234_new_n648_), .Y(_abc_41234_new_n1973_));
AOI21X1 AOI21X1_119 ( .A(_abc_41234_new_n1967_), .B(_abc_41234_new_n634_), .C(_abc_41234_new_n648_), .Y(_abc_41234_new_n1982_));
AOI21X1 AOI21X1_12 ( .A(rdatahold_3_), .B(_abc_41234_new_n633_), .C(_abc_41234_new_n827_), .Y(_abc_41234_new_n828_));
AOI21X1 AOI21X1_120 ( .A(_abc_41234_new_n1967_), .B(_abc_41234_new_n568_), .C(_abc_41234_new_n648_), .Y(_abc_41234_new_n1991_));
AOI21X1 AOI21X1_121 ( .A(rdatahold2_4_), .B(_abc_41234_new_n596_), .C(_abc_41234_new_n2005_), .Y(_abc_41234_new_n2006_));
AOI21X1 AOI21X1_122 ( .A(rdatahold2_5_), .B(_abc_41234_new_n596_), .C(_abc_41234_new_n2014_), .Y(_abc_41234_new_n2015_));
AOI21X1 AOI21X1_123 ( .A(rdatahold2_6_), .B(_abc_41234_new_n596_), .C(_abc_41234_new_n2023_), .Y(_abc_41234_new_n2024_));
AOI21X1 AOI21X1_124 ( .A(_abc_41234_new_n2019_), .B(regfil_1__6_), .C(regfil_1__7_), .Y(_abc_41234_new_n2030_));
AOI21X1 AOI21X1_125 ( .A(rdatahold2_7_), .B(_abc_41234_new_n596_), .C(_abc_41234_new_n2032_), .Y(_abc_41234_new_n2033_));
AOI21X1 AOI21X1_126 ( .A(_abc_41234_new_n1056_), .B(_abc_41234_new_n2035_), .C(_abc_41234_new_n2036_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_0_));
AOI21X1 AOI21X1_127 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n1143_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n2054_));
AOI21X1 AOI21X1_128 ( .A(rdatahold_0_), .B(_abc_41234_new_n1855_), .C(_abc_41234_new_n2065_), .Y(_abc_41234_new_n2066_));
AOI21X1 AOI21X1_129 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n731_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n2068_));
AOI21X1 AOI21X1_13 ( .A(_abc_41234_new_n836_), .B(_abc_41234_new_n837_), .C(_abc_41234_new_n559_), .Y(_abc_41234_new_n838_));
AOI21X1 AOI21X1_130 ( .A(regfil_4__1_bF_buf0_), .B(_abc_41234_new_n1066__bF_buf3), .C(_abc_41234_new_n2077_), .Y(_abc_41234_new_n2078_));
AOI21X1 AOI21X1_131 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n769_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n2080_));
AOI21X1 AOI21X1_132 ( .A(_abc_41234_new_n1956_), .B(_abc_41234_new_n2071_), .C(_abc_41234_new_n769_), .Y(_abc_41234_new_n2083_));
AOI21X1 AOI21X1_133 ( .A(rdatahold_2_), .B(_abc_41234_new_n1855_), .C(_abc_41234_new_n2089_), .Y(_abc_41234_new_n2090_));
AOI21X1 AOI21X1_134 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n815_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n2092_));
AOI21X1 AOI21X1_135 ( .A(_abc_41234_new_n1066__bF_buf2), .B(_abc_41234_new_n819_), .C(_abc_41234_new_n1880_), .Y(_abc_41234_new_n2103_));
AOI21X1 AOI21X1_136 ( .A(_abc_41234_new_n2112_), .B(_abc_41234_new_n1873_), .C(_abc_41234_new_n1066__bF_buf1), .Y(_abc_41234_new_n2113_));
AOI21X1 AOI21X1_137 ( .A(_abc_41234_new_n1066__bF_buf0), .B(_abc_41234_new_n849_), .C(_abc_41234_new_n1880_), .Y(_abc_41234_new_n2115_));
AOI21X1 AOI21X1_138 ( .A(_abc_41234_new_n2124_), .B(_abc_41234_new_n1873_), .C(_abc_41234_new_n1066__bF_buf3), .Y(_abc_41234_new_n2125_));
AOI21X1 AOI21X1_139 ( .A(_abc_41234_new_n1066__bF_buf2), .B(_abc_41234_new_n904_), .C(_abc_41234_new_n1880_), .Y(_abc_41234_new_n2127_));
AOI21X1 AOI21X1_14 ( .A(_abc_41234_new_n533_), .B(regfil_7__4_), .C(_abc_41234_new_n513_), .Y(_abc_41234_new_n841_));
AOI21X1 AOI21X1_140 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n1535_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n2130_));
AOI21X1 AOI21X1_141 ( .A(_abc_41234_new_n2145_), .B(_abc_41234_new_n2148_), .C(_abc_41234_new_n2139_), .Y(_abc_41234_new_n2149_));
AOI21X1 AOI21X1_142 ( .A(_abc_41234_new_n2098_), .B(_abc_41234_new_n2121_), .C(regfil_2__6_), .Y(_abc_41234_new_n2151_));
AOI21X1 AOI21X1_143 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n993_), .C(_abc_41234_new_n1859_), .Y(_abc_41234_new_n2159_));
AOI21X1 AOI21X1_144 ( .A(_abc_41234_new_n1066__bF_buf1), .B(_abc_41234_new_n997_), .C(_abc_41234_new_n1853_), .Y(_abc_41234_new_n2162_));
AOI21X1 AOI21X1_145 ( .A(_abc_41234_new_n2205_), .B(_abc_41234_new_n2189__bF_buf2), .C(_abc_41234_new_n2210_), .Y(_abc_41234_new_n2211_));
AOI21X1 AOI21X1_146 ( .A(_abc_41234_new_n524_), .B(_abc_41234_new_n2221_), .C(_abc_41234_new_n2216_), .Y(_abc_41234_new_n2222_));
AOI21X1 AOI21X1_147 ( .A(_abc_41234_new_n2245_), .B(regfil_7__0_), .C(_abc_41234_new_n536__bF_buf0), .Y(_abc_41234_new_n2246_));
AOI21X1 AOI21X1_148 ( .A(_abc_41234_new_n2245_), .B(regfil_7__1_), .C(_abc_41234_new_n536__bF_buf4), .Y(_abc_41234_new_n2269_));
AOI21X1 AOI21X1_149 ( .A(_abc_41234_new_n2245_), .B(regfil_7__2_), .C(_abc_41234_new_n536__bF_buf2), .Y(_abc_41234_new_n2281_));
AOI21X1 AOI21X1_15 ( .A(_abc_41234_new_n842_), .B(_abc_41234_new_n833_), .C(_abc_41234_new_n844_), .Y(_abc_41234_new_n845_));
AOI21X1 AOI21X1_150 ( .A(_abc_41234_new_n2245_), .B(regfil_7__3_), .C(_abc_41234_new_n536__bF_buf0), .Y(_abc_41234_new_n2293_));
AOI21X1 AOI21X1_151 ( .A(_abc_41234_new_n2245_), .B(regfil_7__4_), .C(_abc_41234_new_n536__bF_buf4), .Y(_abc_41234_new_n2305_));
AOI21X1 AOI21X1_152 ( .A(regfil_7__5_), .B(_abc_41234_new_n2201_), .C(_abc_41234_new_n2326_), .Y(_abc_41234_new_n2327_));
AOI21X1 AOI21X1_153 ( .A(regfil_7__6_), .B(_abc_41234_new_n2201_), .C(_abc_41234_new_n2338_), .Y(_abc_41234_new_n2339_));
AOI21X1 AOI21X1_154 ( .A(_abc_41234_new_n2213_), .B(_abc_41234_new_n2357_), .C(_abc_41234_new_n2359_), .Y(_0intcyc_0_0_));
AOI21X1 AOI21X1_155 ( .A(_abc_41234_new_n509_), .B(_abc_41234_new_n2378_), .C(_abc_41234_new_n2381_), .Y(_abc_41234_new_n2382_));
AOI21X1 AOI21X1_156 ( .A(_abc_41234_new_n2386_), .B(_abc_41234_new_n660__bF_buf2), .C(_abc_41234_new_n2389_), .Y(_abc_41234_new_n2390_));
AOI21X1 AOI21X1_157 ( .A(_abc_41234_new_n1591_), .B(_abc_41234_new_n1536_), .C(_abc_41234_new_n1590_), .Y(_abc_41234_new_n2401_));
AOI21X1 AOI21X1_158 ( .A(regfil_7__7_), .B(_abc_41234_new_n1634_), .C(_abc_41234_new_n2405_), .Y(_abc_41234_new_n2406_));
AOI21X1 AOI21X1_159 ( .A(_abc_41234_new_n2403_), .B(_abc_41234_new_n1307_), .C(_abc_41234_new_n2407_), .Y(_abc_41234_new_n2408_));
AOI21X1 AOI21X1_16 ( .A(_abc_41234_new_n806_), .B(regfil_0__4_), .C(_abc_41234_new_n600_), .Y(_abc_41234_new_n876_));
AOI21X1 AOI21X1_160 ( .A(_abc_41234_new_n1013_), .B(_abc_41234_new_n534__bF_buf0), .C(_abc_41234_new_n2415__bF_buf4), .Y(_abc_41234_new_n2416_));
AOI21X1 AOI21X1_161 ( .A(_abc_41234_new_n509_), .B(_abc_41234_new_n2423_), .C(_abc_41234_new_n2420_), .Y(_abc_41234_new_n2424_));
AOI21X1 AOI21X1_162 ( .A(_abc_41234_new_n2415__bF_buf3), .B(_abc_41234_new_n2448_), .C(_abc_41234_new_n2453_), .Y(_0eienb_0_0_));
AOI21X1 AOI21X1_163 ( .A(_abc_41234_new_n536__bF_buf2), .B(_abc_41234_new_n2462_), .C(_abc_41234_new_n2490_), .Y(_abc_41234_new_n2491_));
AOI21X1 AOI21X1_164 ( .A(_abc_41234_new_n515__bF_buf5), .B(_abc_41234_new_n2500_), .C(_abc_41234_new_n2507_), .Y(_abc_41234_new_n2508_));
AOI21X1 AOI21X1_165 ( .A(_abc_41234_new_n2485_), .B(_abc_41234_new_n1046__bF_buf7), .C(_abc_41234_new_n2509_), .Y(_abc_41234_new_n2510_));
AOI21X1 AOI21X1_166 ( .A(_abc_41234_new_n2538_), .B(statesel_1_), .C(_abc_41234_new_n2539_), .Y(_abc_41234_new_n2540_));
AOI21X1 AOI21X1_167 ( .A(_abc_41234_new_n668__bF_buf3), .B(_abc_41234_new_n665__bF_buf1), .C(statesel_1_), .Y(_abc_41234_new_n2550_));
AOI21X1 AOI21X1_168 ( .A(_abc_41234_new_n2548_), .B(_abc_41234_new_n515__bF_buf4), .C(_abc_41234_new_n2552_), .Y(_abc_41234_new_n2553_));
AOI21X1 AOI21X1_169 ( .A(_abc_41234_new_n530_), .B(_abc_41234_new_n2563_), .C(_abc_41234_new_n665__bF_buf3), .Y(_abc_41234_new_n2564_));
AOI21X1 AOI21X1_17 ( .A(_abc_41234_new_n875_), .B(_abc_41234_new_n876_), .C(_abc_41234_new_n647_), .Y(_abc_41234_new_n877_));
AOI21X1 AOI21X1_170 ( .A(_abc_41234_new_n2538_), .B(statesel_2_), .C(_abc_41234_new_n2565_), .Y(_abc_41234_new_n2566_));
AOI21X1 AOI21X1_171 ( .A(opcode_5_bF_buf4_), .B(_abc_41234_new_n2466_), .C(_abc_41234_new_n2569_), .Y(_abc_41234_new_n2570_));
AOI21X1 AOI21X1_172 ( .A(_abc_41234_new_n2568_), .B(_abc_41234_new_n2570_), .C(_abc_41234_new_n2572_), .Y(_abc_41234_new_n2573_));
AOI21X1 AOI21X1_173 ( .A(statesel_2_), .B(_abc_41234_new_n2567_), .C(_abc_41234_new_n2573_), .Y(_abc_41234_new_n2574_));
AOI21X1 AOI21X1_174 ( .A(_abc_41234_new_n2582_), .B(_abc_41234_new_n2581_), .C(reset_bF_buf7), .Y(_abc_41234_new_n2585_));
AOI21X1 AOI21X1_175 ( .A(_abc_41234_new_n2538_), .B(statesel_3_), .C(_abc_41234_new_n2589_), .Y(_abc_41234_new_n2590_));
AOI21X1 AOI21X1_176 ( .A(_abc_41234_new_n2593_), .B(_abc_41234_new_n2592_), .C(_abc_41234_new_n2594_), .Y(_abc_41234_new_n2595_));
AOI21X1 AOI21X1_177 ( .A(_abc_41234_new_n2596_), .B(_abc_41234_new_n2597_), .C(_abc_41234_new_n2595_), .Y(_abc_41234_new_n2598_));
AOI21X1 AOI21X1_178 ( .A(_abc_41234_new_n2599_), .B(_abc_41234_new_n660__bF_buf6), .C(_abc_41234_new_n2608_), .Y(_abc_41234_new_n2609_));
AOI21X1 AOI21X1_179 ( .A(_abc_41234_new_n2538_), .B(statesel_4_), .C(_abc_41234_new_n2461_), .Y(_abc_41234_new_n2612_));
AOI21X1 AOI21X1_18 ( .A(_abc_41234_new_n851_), .B(_abc_41234_new_n541_), .C(_abc_41234_new_n883_), .Y(_abc_41234_new_n884_));
AOI21X1 AOI21X1_180 ( .A(_abc_41234_new_n2614_), .B(statesel_4_), .C(_abc_41234_new_n2617_), .Y(_abc_41234_new_n2618_));
AOI21X1 AOI21X1_181 ( .A(_abc_41234_new_n2619_), .B(_abc_41234_new_n660__bF_buf5), .C(_abc_41234_new_n2626_), .Y(_abc_41234_new_n2627_));
AOI21X1 AOI21X1_182 ( .A(_abc_41234_new_n2614_), .B(statesel_5_), .C(_abc_41234_new_n2630_), .Y(_abc_41234_new_n2631_));
AOI21X1 AOI21X1_183 ( .A(_abc_41234_new_n1610_), .B(_abc_41234_new_n2670_), .C(_abc_41234_new_n534__bF_buf5), .Y(_abc_41234_new_n2679_));
AOI21X1 AOI21X1_184 ( .A(_abc_41234_new_n536__bF_buf5), .B(_abc_41234_new_n2685_), .C(_abc_41234_new_n2677_), .Y(_abc_41234_new_n2686_));
AOI21X1 AOI21X1_185 ( .A(_abc_41234_new_n2691_), .B(_abc_41234_new_n1046__bF_buf5), .C(_abc_41234_new_n2683_), .Y(_abc_41234_new_n2692_));
AOI21X1 AOI21X1_186 ( .A(_abc_41234_new_n2693_), .B(_abc_41234_new_n660__bF_buf3), .C(_abc_41234_new_n2698_), .Y(_abc_41234_new_n2699_));
AOI21X1 AOI21X1_187 ( .A(_abc_41234_new_n661_), .B(_abc_41234_new_n2720_), .C(_abc_41234_new_n2722_), .Y(_abc_41234_new_n2723_));
AOI21X1 AOI21X1_188 ( .A(_abc_41234_new_n2701_), .B(_abc_41234_new_n2189__bF_buf3), .C(_abc_41234_new_n2415__bF_buf2), .Y(_abc_41234_new_n2725_));
AOI21X1 AOI21X1_189 ( .A(_abc_41234_new_n1637_), .B(_abc_41234_new_n2735_), .C(_abc_41234_new_n2744_), .Y(_abc_41234_new_n2745_));
AOI21X1 AOI21X1_19 ( .A(regfil_7__5_), .B(_abc_41234_new_n533_), .C(_abc_41234_new_n887_), .Y(_abc_41234_new_n888_));
AOI21X1 AOI21X1_190 ( .A(_abc_41234_new_n2739_), .B(_abc_41234_new_n1729_), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n2746_));
AOI21X1 AOI21X1_191 ( .A(_abc_41234_new_n1644_), .B(wdatahold_2_), .C(_abc_41234_new_n2748_), .Y(_abc_41234_new_n2749_));
AOI21X1 AOI21X1_192 ( .A(_abc_41234_new_n2749_), .B(_abc_41234_new_n2745_), .C(_abc_41234_new_n1047__bF_buf1), .Y(_abc_41234_new_n2750_));
AOI21X1 AOI21X1_193 ( .A(_abc_41234_new_n1610_), .B(_abc_41234_new_n2731_), .C(_abc_41234_new_n534__bF_buf4), .Y(_abc_41234_new_n2754_));
AOI21X1 AOI21X1_194 ( .A(alu_res_2_), .B(_abc_41234_new_n2695_), .C(_abc_41234_new_n2760_), .Y(_abc_41234_new_n2761_));
AOI21X1 AOI21X1_195 ( .A(_abc_41234_new_n2504_), .B(_abc_41234_new_n2764_), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n2768_));
AOI21X1 AOI21X1_196 ( .A(_abc_41234_new_n536__bF_buf1), .B(_abc_41234_new_n2779_), .C(_abc_41234_new_n2765_), .Y(_abc_41234_new_n2780_));
AOI21X1 AOI21X1_197 ( .A(_abc_41234_new_n1630_), .B(_abc_41234_new_n2778_), .C(_abc_41234_new_n2783_), .Y(_abc_41234_new_n2784_));
AOI21X1 AOI21X1_198 ( .A(_abc_41234_new_n2785_), .B(_abc_41234_new_n1046__bF_buf3), .C(_abc_41234_new_n2770_), .Y(_abc_41234_new_n2786_));
AOI21X1 AOI21X1_199 ( .A(_abc_41234_new_n2787_), .B(_abc_41234_new_n660__bF_buf1), .C(_abc_41234_new_n2789_), .Y(_abc_41234_new_n2790_));
AOI21X1 AOI21X1_2 ( .A(_abc_41234_new_n679_), .B(_abc_41234_new_n680_), .C(_abc_41234_new_n711_), .Y(_abc_41234_new_n712_));
AOI21X1 AOI21X1_20 ( .A(_abc_41234_new_n847_), .B(_abc_41234_new_n513_), .C(_abc_41234_new_n888_), .Y(_abc_41234_new_n889_));
AOI21X1 AOI21X1_200 ( .A(_abc_41234_new_n2504_), .B(_abc_41234_new_n2792_), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n2798_));
AOI21X1 AOI21X1_201 ( .A(_abc_41234_new_n2806_), .B(intcyc_bF_buf1), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n2807_));
AOI21X1 AOI21X1_202 ( .A(_abc_41234_new_n536__bF_buf0), .B(_abc_41234_new_n2811_), .C(_abc_41234_new_n2810_), .Y(_abc_41234_new_n2812_));
AOI21X1 AOI21X1_203 ( .A(_abc_41234_new_n2805_), .B(_abc_41234_new_n1627_), .C(_abc_41234_new_n2814_), .Y(_abc_41234_new_n2815_));
AOI21X1 AOI21X1_204 ( .A(_abc_41234_new_n2817_), .B(_abc_41234_new_n1046__bF_buf2), .C(_abc_41234_new_n2800_), .Y(_abc_41234_new_n2818_));
AOI21X1 AOI21X1_205 ( .A(_abc_41234_new_n2793_), .B(_abc_41234_new_n2818_), .C(_abc_41234_new_n2415__bF_buf1), .Y(_abc_41234_new_n2819_));
AOI21X1 AOI21X1_206 ( .A(_abc_41234_new_n2504_), .B(_abc_41234_new_n2824_), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n2828_));
AOI21X1 AOI21X1_207 ( .A(_abc_41234_new_n536__bF_buf5), .B(_abc_41234_new_n2839_), .C(_abc_41234_new_n2825_), .Y(_abc_41234_new_n2840_));
AOI21X1 AOI21X1_208 ( .A(_abc_41234_new_n2837_), .B(_abc_41234_new_n2838_), .C(_abc_41234_new_n2842_), .Y(_abc_41234_new_n2843_));
AOI21X1 AOI21X1_209 ( .A(_abc_41234_new_n2844_), .B(_abc_41234_new_n1046__bF_buf1), .C(_abc_41234_new_n2830_), .Y(_abc_41234_new_n2845_));
AOI21X1 AOI21X1_21 ( .A(_abc_41234_new_n921_), .B(_abc_41234_new_n919_), .C(_abc_41234_new_n647_), .Y(_abc_41234_new_n922_));
AOI21X1 AOI21X1_210 ( .A(_abc_41234_new_n2846_), .B(_abc_41234_new_n660__bF_buf0), .C(_abc_41234_new_n2848_), .Y(_abc_41234_new_n2849_));
AOI21X1 AOI21X1_211 ( .A(_abc_41234_new_n2858_), .B(_abc_41234_new_n2859_), .C(_abc_41234_new_n2868_), .Y(_abc_41234_new_n2869_));
AOI21X1 AOI21X1_212 ( .A(_abc_41234_new_n1610_), .B(_abc_41234_new_n2851_), .C(_abc_41234_new_n534__bF_buf0), .Y(_abc_41234_new_n2872_));
AOI21X1 AOI21X1_213 ( .A(_abc_41234_new_n2870_), .B(_abc_41234_new_n1046__bF_buf0), .C(_abc_41234_new_n2874_), .Y(_abc_41234_new_n2875_));
AOI21X1 AOI21X1_214 ( .A(_abc_41234_new_n2876_), .B(_abc_41234_new_n660__bF_buf7), .C(_abc_41234_new_n2878_), .Y(_abc_41234_new_n2879_));
AOI21X1 AOI21X1_215 ( .A(_abc_41234_new_n2884_), .B(_abc_41234_new_n1729_), .C(_abc_41234_new_n2885_), .Y(_abc_41234_new_n2886_));
AOI21X1 AOI21X1_216 ( .A(wdatahold_7_), .B(_abc_41234_new_n2189__bF_buf1), .C(_abc_41234_new_n2903_), .Y(_abc_41234_new_n2904_));
AOI21X1 AOI21X1_217 ( .A(_abc_41234_new_n2905_), .B(_abc_41234_new_n660__bF_buf6), .C(_abc_41234_new_n2907_), .Y(_abc_41234_new_n2908_));
AOI21X1 AOI21X1_218 ( .A(_abc_41234_new_n2189__bF_buf0), .B(_abc_41234_new_n2930_), .C(_abc_41234_new_n2955_), .Y(_abc_41234_new_n2956_));
AOI21X1 AOI21X1_219 ( .A(_abc_41234_new_n2957_), .B(_abc_41234_new_n660__bF_buf5), .C(_abc_41234_new_n2960_), .Y(_abc_41234_new_n2961_));
AOI21X1 AOI21X1_22 ( .A(_abc_41234_new_n533_), .B(regfil_7__6_), .C(_abc_41234_new_n513_), .Y(_abc_41234_new_n928_));
AOI21X1 AOI21X1_220 ( .A(_abc_41234_new_n668__bF_buf3), .B(_abc_41234_new_n2965_), .C(_abc_41234_new_n2207__bF_buf2), .Y(_abc_41234_new_n2966_));
AOI21X1 AOI21X1_221 ( .A(_abc_41234_new_n2977_), .B(_abc_41234_new_n2980_), .C(_abc_41234_new_n2981_), .Y(_abc_41234_new_n2982_));
AOI21X1 AOI21X1_222 ( .A(_abc_41234_new_n2994_), .B(raddrhold_2_), .C(_abc_41234_new_n3001_), .Y(_abc_41234_new_n3002_));
AOI21X1 AOI21X1_223 ( .A(_abc_41234_new_n2951__bF_buf1), .B(_abc_41234_new_n3003_), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n3007_));
AOI21X1 AOI21X1_224 ( .A(rdatahold2_2_), .B(_abc_41234_new_n2513_), .C(_abc_41234_new_n3015_), .Y(_abc_41234_new_n3016_));
AOI21X1 AOI21X1_225 ( .A(_abc_41234_new_n3028_), .B(raddrhold_3_), .C(_abc_41234_new_n3033_), .Y(_abc_41234_new_n3034_));
AOI21X1 AOI21X1_226 ( .A(_abc_41234_new_n2951__bF_buf3), .B(_abc_41234_new_n3023_), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n3038_));
AOI21X1 AOI21X1_227 ( .A(raddrhold_4_), .B(_abc_41234_new_n3024_), .C(_abc_41234_new_n3050_), .Y(_abc_41234_new_n3051_));
AOI21X1 AOI21X1_228 ( .A(_abc_41234_new_n3053_), .B(raddrhold_4_), .C(_abc_41234_new_n3058_), .Y(_abc_41234_new_n3059_));
AOI21X1 AOI21X1_229 ( .A(_abc_41234_new_n2951__bF_buf1), .B(_abc_41234_new_n3049_), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n3063_));
AOI21X1 AOI21X1_23 ( .A(_abc_41234_new_n933_), .B(_abc_41234_new_n932_), .C(_abc_41234_new_n559_), .Y(_abc_41234_new_n934_));
AOI21X1 AOI21X1_230 ( .A(_abc_41234_new_n3077_), .B(_abc_41234_new_n3074_), .C(_abc_41234_new_n2959__bF_buf2), .Y(_abc_41234_new_n3078_));
AOI21X1 AOI21X1_231 ( .A(_abc_41234_new_n3080_), .B(raddrhold_5_), .C(_abc_41234_new_n3085_), .Y(_abc_41234_new_n3086_));
AOI21X1 AOI21X1_232 ( .A(_abc_41234_new_n2951__bF_buf3), .B(_abc_41234_new_n3074_), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n3090_));
AOI21X1 AOI21X1_233 ( .A(_abc_41234_new_n3076_), .B(_abc_41234_new_n3078_), .C(_abc_41234_new_n3098_), .Y(_abc_41234_new_n3099_));
AOI21X1 AOI21X1_234 ( .A(_abc_41234_new_n668__bF_buf2), .B(_abc_41234_new_n3101_), .C(_abc_41234_new_n2207__bF_buf1), .Y(_abc_41234_new_n3102_));
AOI21X1 AOI21X1_235 ( .A(_abc_41234_new_n2977_), .B(_abc_41234_new_n3115_), .C(_abc_41234_new_n3116_), .Y(_abc_41234_new_n3117_));
AOI21X1 AOI21X1_236 ( .A(_abc_41234_new_n3076_), .B(_abc_41234_new_n3101_), .C(_abc_41234_new_n2959__bF_buf1), .Y(_abc_41234_new_n3120_));
AOI21X1 AOI21X1_237 ( .A(_abc_41234_new_n3119_), .B(_abc_41234_new_n660__bF_buf7), .C(_abc_41234_new_n3122_), .Y(_abc_41234_new_n3123_));
AOI21X1 AOI21X1_238 ( .A(_abc_41234_new_n2977_), .B(_abc_41234_new_n3138_), .C(_abc_41234_new_n3140_), .Y(_abc_41234_new_n3141_));
AOI21X1 AOI21X1_239 ( .A(_abc_41234_new_n3143_), .B(_abc_41234_new_n660__bF_buf6), .C(_abc_41234_new_n3148_), .Y(_abc_41234_new_n3149_));
AOI21X1 AOI21X1_24 ( .A(_abc_41234_new_n935_), .B(_abc_41234_new_n927_), .C(_abc_41234_new_n937_), .Y(_abc_41234_new_n938_));
AOI21X1 AOI21X1_240 ( .A(_abc_41234_new_n2977_), .B(_abc_41234_new_n3163_), .C(_abc_41234_new_n3165_), .Y(_abc_41234_new_n3166_));
AOI21X1 AOI21X1_241 ( .A(_abc_41234_new_n3168_), .B(_abc_41234_new_n660__bF_buf5), .C(_abc_41234_new_n3172_), .Y(_abc_41234_new_n3173_));
AOI21X1 AOI21X1_242 ( .A(_abc_41234_new_n2951__bF_buf1), .B(_abc_41234_new_n3175_), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n3188_));
AOI21X1 AOI21X1_243 ( .A(_abc_41234_new_n3176_), .B(_abc_41234_new_n3178_), .C(_abc_41234_new_n3197_), .Y(_abc_41234_new_n3198_));
AOI21X1 AOI21X1_244 ( .A(_abc_41234_new_n2920_), .B(_abc_41234_new_n3200_), .C(_abc_41234_new_n534__bF_buf1), .Y(_abc_41234_new_n3211_));
AOI21X1 AOI21X1_245 ( .A(raddrhold_10_), .B(_abc_41234_new_n2951__bF_buf3), .C(_abc_41234_new_n3214_), .Y(_abc_41234_new_n3215_));
AOI21X1 AOI21X1_246 ( .A(_abc_41234_new_n3211_), .B(_abc_41234_new_n3210_), .C(_abc_41234_new_n3216_), .Y(_abc_41234_new_n3217_));
AOI21X1 AOI21X1_247 ( .A(_abc_41234_new_n3218_), .B(_abc_41234_new_n660__bF_buf3), .C(_abc_41234_new_n3222_), .Y(_abc_41234_new_n3223_));
AOI21X1 AOI21X1_248 ( .A(_abc_41234_new_n3177_), .B(raddrhold_10_), .C(raddrhold_11_), .Y(_abc_41234_new_n3243_));
AOI21X1 AOI21X1_249 ( .A(_abc_41234_new_n3242_), .B(_abc_41234_new_n660__bF_buf2), .C(_abc_41234_new_n3245_), .Y(_abc_41234_new_n3246_));
AOI21X1 AOI21X1_25 ( .A(_abc_41234_new_n919_), .B(regfil_0__6_), .C(_abc_41234_new_n600_), .Y(_abc_41234_new_n960_));
AOI21X1 AOI21X1_250 ( .A(_abc_41234_new_n668__bF_buf1), .B(_abc_41234_new_n3248_), .C(_abc_41234_new_n2207__bF_buf0), .Y(_abc_41234_new_n3251_));
AOI21X1 AOI21X1_251 ( .A(_abc_41234_new_n3262_), .B(_abc_41234_new_n660__bF_buf1), .C(_abc_41234_new_n3269_), .Y(_abc_41234_new_n3270_));
AOI21X1 AOI21X1_252 ( .A(_abc_41234_new_n3282_), .B(raddrhold_13_), .C(_abc_41234_new_n3286_), .Y(_abc_41234_new_n3287_));
AOI21X1 AOI21X1_253 ( .A(_abc_41234_new_n3288_), .B(_abc_41234_new_n660__bF_buf0), .C(_abc_41234_new_n3291_), .Y(_abc_41234_new_n3292_));
AOI21X1 AOI21X1_254 ( .A(_abc_41234_new_n2920_), .B(_abc_41234_new_n3294_), .C(_abc_41234_new_n534__bF_buf3), .Y(_abc_41234_new_n3300_));
AOI21X1 AOI21X1_255 ( .A(_abc_41234_new_n3308_), .B(_abc_41234_new_n660__bF_buf7), .C(_abc_41234_new_n3313_), .Y(_abc_41234_new_n3314_));
AOI21X1 AOI21X1_256 ( .A(_abc_41234_new_n1831_), .B(_abc_41234_new_n1832_), .C(_abc_41234_new_n2918_), .Y(_abc_41234_new_n3317_));
AOI21X1 AOI21X1_257 ( .A(_abc_41234_new_n2920_), .B(_abc_41234_new_n3316_), .C(_abc_41234_new_n534__bF_buf2), .Y(_abc_41234_new_n3323_));
AOI21X1 AOI21X1_258 ( .A(_abc_41234_new_n1831_), .B(_abc_41234_new_n1832_), .C(_abc_41234_new_n2944_), .Y(_abc_41234_new_n3325_));
AOI21X1 AOI21X1_259 ( .A(_abc_41234_new_n3331_), .B(_abc_41234_new_n660__bF_buf6), .C(_abc_41234_new_n3334_), .Y(_abc_41234_new_n3335_));
AOI21X1 AOI21X1_26 ( .A(_abc_41234_new_n960_), .B(_abc_41234_new_n959_), .C(_abc_41234_new_n647_), .Y(_abc_41234_new_n961_));
AOI21X1 AOI21X1_260 ( .A(_abc_41234_new_n3337_), .B(_abc_41234_new_n668__bF_buf3), .C(_abc_41234_new_n2922_), .Y(_abc_41234_new_n3345_));
AOI21X1 AOI21X1_261 ( .A(_abc_41234_new_n3345_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf3), .Y(_abc_41234_new_n3348_));
AOI21X1 AOI21X1_262 ( .A(waddrhold_0_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3349_), .Y(_abc_41234_new_n3350_));
AOI21X1 AOI21X1_263 ( .A(_abc_41234_new_n3337_), .B(_abc_41234_new_n2189__bF_buf2), .C(_abc_41234_new_n2415__bF_buf4), .Y(_abc_41234_new_n3352_));
AOI21X1 AOI21X1_264 ( .A(_abc_41234_new_n3351_), .B(_abc_41234_new_n3352_), .C(_abc_41234_new_n3355_), .Y(_abc_41234_new_n3356_));
AOI21X1 AOI21X1_265 ( .A(_abc_41234_new_n2497_), .B(_abc_41234_new_n3365_), .C(_abc_41234_new_n3369_), .Y(_abc_41234_new_n3370_));
AOI21X1 AOI21X1_266 ( .A(_abc_41234_new_n3358_), .B(_abc_41234_new_n2189__bF_buf1), .C(_abc_41234_new_n2415__bF_buf3), .Y(_abc_41234_new_n3372_));
AOI21X1 AOI21X1_267 ( .A(_abc_41234_new_n3371_), .B(_abc_41234_new_n3372_), .C(_abc_41234_new_n3378_), .Y(_abc_41234_new_n3379_));
AOI21X1 AOI21X1_268 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3385_), .C(_abc_41234_new_n3386_), .Y(_abc_41234_new_n3387_));
AOI21X1 AOI21X1_269 ( .A(_abc_41234_new_n3381_), .B(_abc_41234_new_n668__bF_buf1), .C(_abc_41234_new_n2993_), .Y(_abc_41234_new_n3390_));
AOI21X1 AOI21X1_27 ( .A(_abc_41234_new_n703_), .B(_abc_41234_new_n1015_), .C(_abc_41234_new_n1018_), .Y(_abc_41234_new_n1019_));
AOI21X1 AOI21X1_270 ( .A(_abc_41234_new_n3390_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf0), .Y(_abc_41234_new_n3391_));
AOI21X1 AOI21X1_271 ( .A(waddrhold_2_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3392_), .Y(_abc_41234_new_n3393_));
AOI21X1 AOI21X1_272 ( .A(_abc_41234_new_n3381_), .B(_abc_41234_new_n2189__bF_buf5), .C(_abc_41234_new_n2415__bF_buf2), .Y(_abc_41234_new_n3395_));
AOI21X1 AOI21X1_273 ( .A(_abc_41234_new_n3394_), .B(_abc_41234_new_n3395_), .C(_abc_41234_new_n3400_), .Y(_abc_41234_new_n3401_));
AOI21X1 AOI21X1_274 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3404_), .C(_abc_41234_new_n3405_), .Y(_abc_41234_new_n3406_));
AOI21X1 AOI21X1_275 ( .A(_abc_41234_new_n3403_), .B(_abc_41234_new_n668__bF_buf0), .C(_abc_41234_new_n3027_), .Y(_abc_41234_new_n3409_));
AOI21X1 AOI21X1_276 ( .A(_abc_41234_new_n3409_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf4), .Y(_abc_41234_new_n3410_));
AOI21X1 AOI21X1_277 ( .A(waddrhold_3_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3411_), .Y(_abc_41234_new_n3412_));
AOI21X1 AOI21X1_278 ( .A(_abc_41234_new_n3403_), .B(_abc_41234_new_n2189__bF_buf3), .C(_abc_41234_new_n2415__bF_buf1), .Y(_abc_41234_new_n3414_));
AOI21X1 AOI21X1_279 ( .A(_abc_41234_new_n3403_), .B(_abc_41234_new_n3397_), .C(_abc_41234_new_n2671_), .Y(_abc_41234_new_n3417_));
AOI21X1 AOI21X1_28 ( .A(_abc_41234_new_n1027_), .B(_abc_41234_new_n1028_), .C(_abc_41234_new_n1021_), .Y(_abc_41234_new_n1029_));
AOI21X1 AOI21X1_280 ( .A(_abc_41234_new_n3413_), .B(_abc_41234_new_n3414_), .C(_abc_41234_new_n3419_), .Y(_abc_41234_new_n3420_));
AOI21X1 AOI21X1_281 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3427_), .C(_abc_41234_new_n3428_), .Y(_abc_41234_new_n3429_));
AOI21X1 AOI21X1_282 ( .A(_abc_41234_new_n3422_), .B(_abc_41234_new_n668__bF_buf5), .C(_abc_41234_new_n3052_), .Y(_abc_41234_new_n3432_));
AOI21X1 AOI21X1_283 ( .A(_abc_41234_new_n3432_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf2), .Y(_abc_41234_new_n3433_));
AOI21X1 AOI21X1_284 ( .A(waddrhold_4_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3434_), .Y(_abc_41234_new_n3435_));
AOI21X1 AOI21X1_285 ( .A(_abc_41234_new_n3422_), .B(_abc_41234_new_n2189__bF_buf1), .C(_abc_41234_new_n2415__bF_buf0), .Y(_abc_41234_new_n3437_));
AOI21X1 AOI21X1_286 ( .A(_abc_41234_new_n3436_), .B(_abc_41234_new_n3437_), .C(_abc_41234_new_n3442_), .Y(_abc_41234_new_n3443_));
AOI21X1 AOI21X1_287 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3449_), .C(_abc_41234_new_n3450_), .Y(_abc_41234_new_n3451_));
AOI21X1 AOI21X1_288 ( .A(_abc_41234_new_n3445_), .B(_abc_41234_new_n668__bF_buf4), .C(_abc_41234_new_n3079_), .Y(_abc_41234_new_n3454_));
AOI21X1 AOI21X1_289 ( .A(_abc_41234_new_n3454_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf0), .Y(_abc_41234_new_n3455_));
AOI21X1 AOI21X1_29 ( .A(_abc_41234_new_n1077_), .B(_abc_41234_new_n1076_), .C(_abc_41234_new_n1072_), .Y(_abc_41234_new_n1078_));
AOI21X1 AOI21X1_290 ( .A(waddrhold_5_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3456_), .Y(_abc_41234_new_n3457_));
AOI21X1 AOI21X1_291 ( .A(_abc_41234_new_n3445_), .B(_abc_41234_new_n2189__bF_buf5), .C(_abc_41234_new_n2415__bF_buf4), .Y(_abc_41234_new_n3459_));
AOI21X1 AOI21X1_292 ( .A(_abc_41234_new_n3458_), .B(_abc_41234_new_n3459_), .C(_abc_41234_new_n3463_), .Y(_abc_41234_new_n3464_));
AOI21X1 AOI21X1_293 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3469_), .C(_abc_41234_new_n3470_), .Y(_abc_41234_new_n3471_));
AOI21X1 AOI21X1_294 ( .A(_abc_41234_new_n3474_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf4), .Y(_abc_41234_new_n3475_));
AOI21X1 AOI21X1_295 ( .A(waddrhold_6_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3476_), .Y(_abc_41234_new_n3477_));
AOI21X1 AOI21X1_296 ( .A(_abc_41234_new_n3466_), .B(_abc_41234_new_n2189__bF_buf3), .C(_abc_41234_new_n2415__bF_buf3), .Y(_abc_41234_new_n3479_));
AOI21X1 AOI21X1_297 ( .A(_abc_41234_new_n3478_), .B(_abc_41234_new_n3479_), .C(_abc_41234_new_n3484_), .Y(_abc_41234_new_n3485_));
AOI21X1 AOI21X1_298 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3490_), .C(_abc_41234_new_n3491_), .Y(_abc_41234_new_n3492_));
AOI21X1 AOI21X1_299 ( .A(_abc_41234_new_n3487_), .B(_abc_41234_new_n668__bF_buf2), .C(_abc_41234_new_n3127_), .Y(_abc_41234_new_n3495_));
AOI21X1 AOI21X1_3 ( .A(alu_res_0_), .B(_abc_41234_new_n707_), .C(_abc_41234_new_n715_), .Y(_abc_41234_new_n716_));
AOI21X1 AOI21X1_30 ( .A(_abc_41234_new_n1083_), .B(_abc_41234_new_n1086_), .C(_abc_41234_new_n1081_), .Y(_abc_41234_new_n1100_));
AOI21X1 AOI21X1_300 ( .A(_abc_41234_new_n3495_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf2), .Y(_abc_41234_new_n3496_));
AOI21X1 AOI21X1_301 ( .A(waddrhold_7_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3497_), .Y(_abc_41234_new_n3498_));
AOI21X1 AOI21X1_302 ( .A(_abc_41234_new_n3487_), .B(_abc_41234_new_n2189__bF_buf1), .C(_abc_41234_new_n2415__bF_buf2), .Y(_abc_41234_new_n3500_));
AOI21X1 AOI21X1_303 ( .A(_abc_41234_new_n3499_), .B(_abc_41234_new_n3500_), .C(_abc_41234_new_n3504_), .Y(_abc_41234_new_n3505_));
AOI21X1 AOI21X1_304 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3508_), .C(_abc_41234_new_n3509_), .Y(_abc_41234_new_n3510_));
AOI21X1 AOI21X1_305 ( .A(_abc_41234_new_n3507_), .B(_abc_41234_new_n668__bF_buf1), .C(_abc_41234_new_n3152_), .Y(_abc_41234_new_n3513_));
AOI21X1 AOI21X1_306 ( .A(_abc_41234_new_n3513_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf0), .Y(_abc_41234_new_n3514_));
AOI21X1 AOI21X1_307 ( .A(waddrhold_8_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3515_), .Y(_abc_41234_new_n3516_));
AOI21X1 AOI21X1_308 ( .A(_abc_41234_new_n3507_), .B(_abc_41234_new_n2189__bF_buf5), .C(_abc_41234_new_n2415__bF_buf1), .Y(_abc_41234_new_n3518_));
AOI21X1 AOI21X1_309 ( .A(_abc_41234_new_n3517_), .B(_abc_41234_new_n3518_), .C(_abc_41234_new_n3523_), .Y(_abc_41234_new_n3524_));
AOI21X1 AOI21X1_31 ( .A(_abc_41234_new_n1097_), .B(_abc_41234_new_n1091_), .C(_abc_41234_new_n1095_), .Y(_abc_41234_new_n1101_));
AOI21X1 AOI21X1_310 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3530_), .C(_abc_41234_new_n3531_), .Y(_abc_41234_new_n3532_));
AOI21X1 AOI21X1_311 ( .A(_abc_41234_new_n3526_), .B(_abc_41234_new_n668__bF_buf0), .C(_abc_41234_new_n3179_), .Y(_abc_41234_new_n3535_));
AOI21X1 AOI21X1_312 ( .A(_abc_41234_new_n3535_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf4), .Y(_abc_41234_new_n3536_));
AOI21X1 AOI21X1_313 ( .A(waddrhold_9_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3537_), .Y(_abc_41234_new_n3538_));
AOI21X1 AOI21X1_314 ( .A(_abc_41234_new_n3526_), .B(_abc_41234_new_n2189__bF_buf3), .C(_abc_41234_new_n2415__bF_buf0), .Y(_abc_41234_new_n3540_));
AOI21X1 AOI21X1_315 ( .A(_abc_41234_new_n3539_), .B(_abc_41234_new_n3540_), .C(_abc_41234_new_n3544_), .Y(_abc_41234_new_n3545_));
AOI21X1 AOI21X1_316 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3551_), .C(_abc_41234_new_n3552_), .Y(_abc_41234_new_n3553_));
AOI21X1 AOI21X1_317 ( .A(_abc_41234_new_n3547_), .B(_abc_41234_new_n668__bF_buf5), .C(_abc_41234_new_n3205_), .Y(_abc_41234_new_n3556_));
AOI21X1 AOI21X1_318 ( .A(_abc_41234_new_n3556_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf2), .Y(_abc_41234_new_n3557_));
AOI21X1 AOI21X1_319 ( .A(waddrhold_10_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3558_), .Y(_abc_41234_new_n3559_));
AOI21X1 AOI21X1_32 ( .A(_abc_41234_new_n1099_), .B(_abc_41234_new_n1079_), .C(_abc_41234_new_n1102_), .Y(_abc_41234_new_n1103_));
AOI21X1 AOI21X1_320 ( .A(_abc_41234_new_n3547_), .B(_abc_41234_new_n2189__bF_buf1), .C(_abc_41234_new_n2415__bF_buf4), .Y(_abc_41234_new_n3561_));
AOI21X1 AOI21X1_321 ( .A(_abc_41234_new_n3560_), .B(_abc_41234_new_n3561_), .C(_abc_41234_new_n3566_), .Y(_abc_41234_new_n3567_));
AOI21X1 AOI21X1_322 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3573_), .C(_abc_41234_new_n3574_), .Y(_abc_41234_new_n3575_));
AOI21X1 AOI21X1_323 ( .A(_abc_41234_new_n3569_), .B(_abc_41234_new_n668__bF_buf4), .C(_abc_41234_new_n3226_), .Y(_abc_41234_new_n3578_));
AOI21X1 AOI21X1_324 ( .A(_abc_41234_new_n3578_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf0), .Y(_abc_41234_new_n3579_));
AOI21X1 AOI21X1_325 ( .A(waddrhold_11_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3580_), .Y(_abc_41234_new_n3581_));
AOI21X1 AOI21X1_326 ( .A(_abc_41234_new_n3569_), .B(_abc_41234_new_n2189__bF_buf5), .C(_abc_41234_new_n2415__bF_buf3), .Y(_abc_41234_new_n3583_));
AOI21X1 AOI21X1_327 ( .A(_abc_41234_new_n3582_), .B(_abc_41234_new_n3583_), .C(_abc_41234_new_n3588_), .Y(_abc_41234_new_n3589_));
AOI21X1 AOI21X1_328 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3595_), .C(_abc_41234_new_n3596_), .Y(_abc_41234_new_n3597_));
AOI21X1 AOI21X1_329 ( .A(_abc_41234_new_n2497_), .B(_abc_41234_new_n3600_), .C(_abc_41234_new_n2189__bF_buf4), .Y(_abc_41234_new_n3601_));
AOI21X1 AOI21X1_33 ( .A(_abc_41234_new_n1103_), .B(_abc_41234_new_n1104_), .C(_abc_41234_new_n1109_), .Y(_abc_41234_new_n1110_));
AOI21X1 AOI21X1_330 ( .A(waddrhold_12_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3602_), .Y(_abc_41234_new_n3603_));
AOI21X1 AOI21X1_331 ( .A(_abc_41234_new_n3605_), .B(_abc_41234_new_n2189__bF_buf3), .C(_abc_41234_new_n2415__bF_buf2), .Y(_abc_41234_new_n3606_));
AOI21X1 AOI21X1_332 ( .A(_abc_41234_new_n3604_), .B(_abc_41234_new_n3606_), .C(_abc_41234_new_n3591_), .Y(_abc_41234_new_n3607_));
AOI21X1 AOI21X1_333 ( .A(_abc_41234_new_n3585_), .B(_abc_41234_new_n3605_), .C(_abc_41234_new_n3610_), .Y(_abc_41234_new_n3611_));
AOI21X1 AOI21X1_334 ( .A(_abc_41234_new_n3359_), .B(_abc_41234_new_n3619_), .C(_abc_41234_new_n3620_), .Y(_abc_41234_new_n3621_));
AOI21X1 AOI21X1_335 ( .A(_abc_41234_new_n3624_), .B(_abc_41234_new_n668__bF_buf3), .C(_abc_41234_new_n3275_), .Y(_abc_41234_new_n3625_));
AOI21X1 AOI21X1_336 ( .A(_abc_41234_new_n3625_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf2), .Y(_abc_41234_new_n3626_));
AOI21X1 AOI21X1_337 ( .A(waddrhold_13_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3627_), .Y(_abc_41234_new_n3628_));
AOI21X1 AOI21X1_338 ( .A(_abc_41234_new_n3624_), .B(_abc_41234_new_n2189__bF_buf1), .C(_abc_41234_new_n2415__bF_buf1), .Y(_abc_41234_new_n3630_));
AOI21X1 AOI21X1_339 ( .A(_abc_41234_new_n3629_), .B(_abc_41234_new_n3630_), .C(_abc_41234_new_n3614_), .Y(_abc_41234_new_n3631_));
AOI21X1 AOI21X1_34 ( .A(_abc_41234_new_n1115_), .B(_abc_41234_new_n1114_), .C(_abc_41234_new_n1112_), .Y(_abc_41234_new_n1116_));
AOI21X1 AOI21X1_340 ( .A(_abc_41234_new_n3592_), .B(_abc_41234_new_n3617_), .C(_abc_41234_new_n1524_), .Y(_abc_41234_new_n3639_));
AOI21X1 AOI21X1_341 ( .A(waddrhold_14_), .B(_abc_41234_new_n1644_), .C(_abc_41234_new_n3641_), .Y(_abc_41234_new_n3642_));
AOI21X1 AOI21X1_342 ( .A(_abc_41234_new_n3644_), .B(_abc_41234_new_n668__bF_buf2), .C(_abc_41234_new_n3295_), .Y(_abc_41234_new_n3645_));
AOI21X1 AOI21X1_343 ( .A(_abc_41234_new_n3645_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf0), .Y(_abc_41234_new_n3646_));
AOI21X1 AOI21X1_344 ( .A(waddrhold_14_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3647_), .Y(_abc_41234_new_n3648_));
AOI21X1 AOI21X1_345 ( .A(_abc_41234_new_n3644_), .B(_abc_41234_new_n2189__bF_buf5), .C(_abc_41234_new_n2415__bF_buf0), .Y(_abc_41234_new_n3650_));
AOI21X1 AOI21X1_346 ( .A(_abc_41234_new_n3649_), .B(_abc_41234_new_n3650_), .C(_abc_41234_new_n3637_), .Y(_abc_41234_new_n3651_));
AOI21X1 AOI21X1_347 ( .A(_abc_41234_new_n1644_), .B(_abc_41234_new_n3661_), .C(_abc_41234_new_n1047__bF_buf0), .Y(_abc_41234_new_n3662_));
AOI21X1 AOI21X1_348 ( .A(_abc_41234_new_n3661_), .B(_abc_41234_new_n668__bF_buf1), .C(_abc_41234_new_n3318_), .Y(_abc_41234_new_n3665_));
AOI21X1 AOI21X1_349 ( .A(_abc_41234_new_n3665_), .B(_abc_41234_new_n3347_), .C(_abc_41234_new_n2189__bF_buf4), .Y(_abc_41234_new_n3666_));
AOI21X1 AOI21X1_35 ( .A(_abc_41234_new_n1127_), .B(_abc_41234_new_n1128_), .C(_abc_41234_new_n1125_), .Y(_abc_41234_new_n1139_));
AOI21X1 AOI21X1_350 ( .A(waddrhold_15_), .B(_abc_41234_new_n3343_), .C(_abc_41234_new_n3667_), .Y(_abc_41234_new_n3668_));
AOI21X1 AOI21X1_351 ( .A(_abc_41234_new_n3663_), .B(_abc_41234_new_n3668_), .C(_abc_41234_new_n3669_), .Y(_abc_41234_new_n3670_));
AOI21X1 AOI21X1_352 ( .A(_abc_41234_new_n3653_), .B(_abc_41234_new_n3661_), .C(_abc_41234_new_n3610_), .Y(_abc_41234_new_n3672_));
AOI21X1 AOI21X1_353 ( .A(_abc_41234_new_n2466_), .B(_abc_41234_new_n544__bF_buf0), .C(_abc_41234_new_n3697_), .Y(_abc_41234_new_n3698_));
AOI21X1 AOI21X1_354 ( .A(_abc_41234_new_n665__bF_buf1), .B(_abc_41234_new_n536__bF_buf2), .C(_abc_41234_new_n663_), .Y(_abc_41234_new_n3710_));
AOI21X1 AOI21X1_355 ( .A(_abc_41234_new_n1066__bF_buf3), .B(_abc_41234_new_n1848_), .C(_abc_41234_new_n1035_), .Y(_abc_41234_new_n3718_));
AOI21X1 AOI21X1_356 ( .A(_abc_41234_new_n1043_), .B(_abc_41234_new_n1221_), .C(_abc_41234_new_n1066__bF_buf2), .Y(_abc_41234_new_n3726_));
AOI21X1 AOI21X1_357 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n719_), .C(_abc_41234_new_n1344_), .Y(_abc_41234_new_n3730_));
AOI21X1 AOI21X1_358 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n1207_), .C(_abc_41234_new_n3759_), .Y(_abc_41234_new_n3760_));
AOI21X1 AOI21X1_359 ( .A(_abc_41234_new_n818_), .B(_abc_41234_new_n3714_), .C(_abc_41234_new_n3780_), .Y(_abc_41234_new_n3781_));
AOI21X1 AOI21X1_36 ( .A(_abc_41234_new_n1135_), .B(_abc_41234_new_n1124_), .C(_abc_41234_new_n1140_), .Y(_abc_41234_new_n1141_));
AOI21X1 AOI21X1_360 ( .A(_abc_41234_new_n1218_), .B(_abc_41234_new_n3782_), .C(_abc_41234_new_n1066__bF_buf0), .Y(_abc_41234_new_n3783_));
AOI21X1 AOI21X1_361 ( .A(_abc_41234_new_n1163_), .B(_abc_41234_new_n3787_), .C(_abc_41234_new_n1309_), .Y(_abc_41234_new_n3790_));
AOI21X1 AOI21X1_362 ( .A(_abc_41234_new_n848_), .B(_abc_41234_new_n3714_), .C(_abc_41234_new_n3803_), .Y(_abc_41234_new_n3804_));
AOI21X1 AOI21X1_363 ( .A(_abc_41234_new_n3821_), .B(_abc_41234_new_n1108_), .C(_abc_41234_new_n1206_), .Y(_abc_41234_new_n3822_));
AOI21X1 AOI21X1_364 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n903_), .C(_abc_41234_new_n1344_), .Y(_abc_41234_new_n3827_));
AOI21X1 AOI21X1_365 ( .A(_abc_41234_new_n1079_), .B(_abc_41234_new_n1093_), .C(_abc_41234_new_n1091_), .Y(_abc_41234_new_n3832_));
AOI21X1 AOI21X1_366 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n1084_), .C(_abc_41234_new_n1344_), .Y(_abc_41234_new_n3852_));
AOI21X1 AOI21X1_367 ( .A(_abc_41234_new_n1167_), .B(_abc_41234_new_n1169_), .C(_abc_41234_new_n1184_), .Y(_abc_41234_new_n3865_));
AOI21X1 AOI21X1_368 ( .A(_abc_41234_new_n3873_), .B(_abc_41234_new_n1108_), .C(_abc_41234_new_n1206_), .Y(_abc_41234_new_n3874_));
AOI21X1 AOI21X1_369 ( .A(_abc_41234_new_n3903_), .B(_abc_41234_new_n3901_), .C(_abc_41234_new_n1109_), .Y(_abc_41234_new_n3904_));
AOI21X1 AOI21X1_37 ( .A(_abc_41234_new_n1141_), .B(_abc_41234_new_n1147_), .C(_abc_41234_new_n1152_), .Y(_abc_41234_new_n1153_));
AOI21X1 AOI21X1_370 ( .A(_abc_41234_new_n3907_), .B(_abc_41234_new_n3890_), .C(_abc_41234_new_n3887_), .Y(_abc_41234_new_n3908_));
AOI21X1 AOI21X1_371 ( .A(_abc_41234_new_n3910_), .B(_abc_41234_new_n3912_), .C(reset_bF_buf4), .Y(_abc_41234_new_n3913_));
AOI21X1 AOI21X1_372 ( .A(_abc_41234_new_n2947__bF_buf3), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n3918_), .Y(_abc_41234_new_n3919_));
AOI21X1 AOI21X1_373 ( .A(_abc_41234_new_n1106_), .B(regfil_5__0_), .C(_abc_41234_new_n1047__bF_buf4), .Y(_abc_41234_new_n3921_));
AOI21X1 AOI21X1_374 ( .A(_abc_41234_new_n3920_), .B(_abc_41234_new_n3922_), .C(_abc_41234_new_n3924_), .Y(_abc_41234_new_n3925_));
AOI21X1 AOI21X1_375 ( .A(_abc_41234_new_n2482_), .B(_abc_41234_new_n2973_), .C(_abc_41234_new_n3928_), .Y(_abc_41234_new_n3929_));
AOI21X1 AOI21X1_376 ( .A(_abc_41234_new_n3936_), .B(_abc_41234_new_n3934_), .C(_abc_41234_new_n3937_), .Y(_abc_41234_new_n3938_));
AOI21X1 AOI21X1_377 ( .A(_abc_41234_new_n3938_), .B(_abc_41234_new_n3933_), .C(_abc_41234_new_n3939_), .Y(_abc_41234_new_n3940_));
AOI21X1 AOI21X1_378 ( .A(_abc_41234_new_n3930_), .B(_abc_41234_new_n3940_), .C(_abc_41234_new_n3941_), .Y(_abc_41234_new_n3942_));
AOI21X1 AOI21X1_379 ( .A(_abc_41234_new_n1106_), .B(regfil_5__2_), .C(_abc_41234_new_n3945_), .Y(_abc_41234_new_n3946_));
AOI21X1 AOI21X1_38 ( .A(_abc_41234_new_n1168_), .B(_abc_41234_new_n1164_), .C(_abc_41234_new_n1161_), .Y(_abc_41234_new_n1169_));
AOI21X1 AOI21X1_380 ( .A(_abc_41234_new_n2452_), .B(_abc_41234_new_n3955_), .C(_abc_41234_new_n534__bF_buf4), .Y(_abc_41234_new_n3956_));
AOI21X1 AOI21X1_381 ( .A(_abc_41234_new_n3952_), .B(_abc_41234_new_n3956_), .C(_abc_41234_new_n3957_), .Y(_abc_41234_new_n3958_));
AOI21X1 AOI21X1_382 ( .A(_abc_41234_new_n3948_), .B(_abc_41234_new_n3958_), .C(_abc_41234_new_n3966_), .Y(_abc_41234_new_n3967_));
AOI21X1 AOI21X1_383 ( .A(_abc_41234_new_n2463_), .B(_abc_41234_new_n3404_), .C(_abc_41234_new_n3973_), .Y(_abc_41234_new_n3974_));
AOI21X1 AOI21X1_384 ( .A(_abc_41234_new_n3916_), .B(sp_3_), .C(_abc_41234_new_n534__bF_buf3), .Y(_abc_41234_new_n3976_));
AOI21X1 AOI21X1_385 ( .A(_abc_41234_new_n3981_), .B(_abc_41234_new_n3976_), .C(_abc_41234_new_n3982_), .Y(_abc_41234_new_n3983_));
AOI21X1 AOI21X1_386 ( .A(_abc_41234_new_n3960_), .B(_abc_41234_new_n3971_), .C(_abc_41234_new_n3986_), .Y(_abc_41234_new_n3987_));
AOI21X1 AOI21X1_387 ( .A(_abc_41234_new_n2463_), .B(_abc_41234_new_n3427_), .C(_abc_41234_new_n3992_), .Y(_abc_41234_new_n3993_));
AOI21X1 AOI21X1_388 ( .A(_abc_41234_new_n4000_), .B(_abc_41234_new_n2452_), .C(_abc_41234_new_n534__bF_buf2), .Y(_abc_41234_new_n4001_));
AOI21X1 AOI21X1_389 ( .A(_abc_41234_new_n3998_), .B(_abc_41234_new_n4001_), .C(_abc_41234_new_n4002_), .Y(_abc_41234_new_n4003_));
AOI21X1 AOI21X1_39 ( .A(_abc_41234_new_n1186_), .B(_abc_41234_new_n1187_), .C(_abc_41234_new_n1182_), .Y(_abc_41234_new_n1188_));
AOI21X1 AOI21X1_390 ( .A(_abc_41234_new_n3427_), .B(_abc_41234_new_n3963_), .C(_abc_41234_new_n4004_), .Y(_abc_41234_new_n4005_));
AOI21X1 AOI21X1_391 ( .A(_abc_41234_new_n3994_), .B(_abc_41234_new_n4003_), .C(_abc_41234_new_n4006_), .Y(_abc_41234_new_n4007_));
AOI21X1 AOI21X1_392 ( .A(_abc_41234_new_n4023_), .B(_abc_41234_new_n1094_), .C(_abc_41234_new_n2451_), .Y(_abc_41234_new_n4024_));
AOI21X1 AOI21X1_393 ( .A(sp_5_), .B(_abc_41234_new_n4012_), .C(_abc_41234_new_n4028_), .Y(_abc_41234_new_n4029_));
AOI21X1 AOI21X1_394 ( .A(_abc_41234_new_n3447_), .B(_abc_41234_new_n2947__bF_buf0), .C(_abc_41234_new_n1085_), .Y(_abc_41234_new_n4037_));
AOI21X1 AOI21X1_395 ( .A(_abc_41234_new_n4053_), .B(_abc_41234_new_n4054_), .C(_abc_41234_new_n4049_), .Y(_abc_41234_new_n4055_));
AOI21X1 AOI21X1_396 ( .A(_abc_41234_new_n1106_), .B(regfil_5__7_), .C(_abc_41234_new_n1047__bF_buf1), .Y(_abc_41234_new_n4062_));
AOI21X1 AOI21X1_397 ( .A(_abc_41234_new_n2463_), .B(_abc_41234_new_n3490_), .C(_abc_41234_new_n4063_), .Y(_abc_41234_new_n4064_));
AOI21X1 AOI21X1_398 ( .A(_abc_41234_new_n4041_), .B(_abc_41234_new_n1080_), .C(_abc_41234_new_n3935_), .Y(_abc_41234_new_n4066_));
AOI21X1 AOI21X1_399 ( .A(sp_7_), .B(_abc_41234_new_n4068_), .C(_abc_41234_new_n4071_), .Y(_abc_41234_new_n4072_));
AOI21X1 AOI21X1_4 ( .A(regfil_0__1_), .B(_abc_41234_new_n642_), .C(_abc_41234_new_n600_), .Y(_abc_41234_new_n745_));
AOI21X1 AOI21X1_40 ( .A(_abc_41234_new_n1173_), .B(_abc_41234_new_n1174_), .C(_abc_41234_new_n1171_), .Y(_abc_41234_new_n1190_));
AOI21X1 AOI21X1_400 ( .A(_abc_41234_new_n4072_), .B(_abc_41234_new_n4067_), .C(_abc_41234_new_n4073_), .Y(_abc_41234_new_n4074_));
AOI21X1 AOI21X1_401 ( .A(_abc_41234_new_n4074_), .B(_abc_41234_new_n4065_), .C(_abc_41234_new_n4076_), .Y(_abc_41234_new_n4077_));
AOI21X1 AOI21X1_402 ( .A(_abc_41234_new_n2463_), .B(_abc_41234_new_n3508_), .C(_abc_41234_new_n4084_), .Y(_abc_41234_new_n4085_));
AOI21X1 AOI21X1_403 ( .A(sp_8_), .B(_abc_41234_new_n4091_), .C(_abc_41234_new_n4093_), .Y(_abc_41234_new_n4094_));
AOI21X1 AOI21X1_404 ( .A(_abc_41234_new_n4094_), .B(_abc_41234_new_n4090_), .C(_abc_41234_new_n4095_), .Y(_abc_41234_new_n4096_));
AOI21X1 AOI21X1_405 ( .A(_abc_41234_new_n4096_), .B(_abc_41234_new_n4087_), .C(_abc_41234_new_n4098_), .Y(_abc_41234_new_n4099_));
AOI21X1 AOI21X1_406 ( .A(_abc_41234_new_n4108_), .B(_abc_41234_new_n4106_), .C(_abc_41234_new_n534__bF_buf1), .Y(_abc_41234_new_n4109_));
AOI21X1 AOI21X1_407 ( .A(_abc_41234_new_n1251_), .B(_abc_41234_new_n1606_), .C(_abc_41234_new_n2415__bF_buf1), .Y(_abc_41234_new_n4117_));
AOI21X1 AOI21X1_408 ( .A(_abc_41234_new_n4118_), .B(_abc_41234_new_n4110_), .C(_abc_41234_new_n4120_), .Y(_abc_41234_new_n4121_));
AOI21X1 AOI21X1_409 ( .A(_abc_41234_new_n4069_), .B(_abc_41234_new_n3528_), .C(_abc_41234_new_n1358_), .Y(_abc_41234_new_n4124_));
AOI21X1 AOI21X1_41 ( .A(_abc_41234_new_n1185_), .B(_abc_41234_new_n1170_), .C(_abc_41234_new_n1191_), .Y(_abc_41234_new_n1192_));
AOI21X1 AOI21X1_410 ( .A(_abc_41234_new_n4138_), .B(_abc_41234_new_n4130_), .C(_abc_41234_new_n2415__bF_buf0), .Y(_abc_41234_new_n4139_));
AOI21X1 AOI21X1_411 ( .A(_abc_41234_new_n4112_), .B(sp_11_), .C(_abc_41234_new_n4151_), .Y(_abc_41234_new_n4152_));
AOI21X1 AOI21X1_412 ( .A(_abc_41234_new_n4155_), .B(_abc_41234_new_n2452_), .C(_abc_41234_new_n4156_), .Y(_abc_41234_new_n4157_));
AOI21X1 AOI21X1_413 ( .A(_abc_41234_new_n1362_), .B(_abc_41234_new_n1606_), .C(_abc_41234_new_n2415__bF_buf4), .Y(_abc_41234_new_n4161_));
AOI21X1 AOI21X1_414 ( .A(_abc_41234_new_n3592_), .B(_abc_41234_new_n2947__bF_buf1), .C(_abc_41234_new_n1408_), .Y(_abc_41234_new_n4171_));
AOI21X1 AOI21X1_415 ( .A(_abc_41234_new_n4183_), .B(_abc_41234_new_n4178_), .C(_abc_41234_new_n2415__bF_buf3), .Y(_abc_41234_new_n4184_));
AOI21X1 AOI21X1_416 ( .A(_abc_41234_new_n4193_), .B(_abc_41234_new_n2452_), .C(_abc_41234_new_n4194_), .Y(_abc_41234_new_n4195_));
AOI21X1 AOI21X1_417 ( .A(_abc_41234_new_n1106_), .B(regfil_4__5_), .C(_abc_41234_new_n1047__bF_buf0), .Y(_abc_41234_new_n4201_));
AOI21X1 AOI21X1_418 ( .A(_abc_41234_new_n4198_), .B(_abc_41234_new_n2462_), .C(_abc_41234_new_n4202_), .Y(_abc_41234_new_n4203_));
AOI21X1 AOI21X1_419 ( .A(_abc_41234_new_n4205_), .B(_abc_41234_new_n4196_), .C(_abc_41234_new_n4207_), .Y(_abc_41234_new_n4208_));
AOI21X1 AOI21X1_42 ( .A(_abc_41234_new_n1155_), .B(_abc_41234_new_n996_), .C(_abc_41234_new_n1108_), .Y(_abc_41234_new_n1203_));
AOI21X1 AOI21X1_420 ( .A(_abc_41234_new_n4215_), .B(_abc_41234_new_n2452_), .C(_abc_41234_new_n4216_), .Y(_abc_41234_new_n4217_));
AOI21X1 AOI21X1_421 ( .A(_abc_41234_new_n1106_), .B(regfil_4__6_), .C(_abc_41234_new_n1047__bF_buf4), .Y(_abc_41234_new_n4223_));
AOI21X1 AOI21X1_422 ( .A(_abc_41234_new_n4220_), .B(_abc_41234_new_n4225_), .C(_abc_41234_new_n4226_), .Y(_abc_41234_new_n4227_));
AOI21X1 AOI21X1_423 ( .A(_abc_41234_new_n4227_), .B(_abc_41234_new_n4218_), .C(_abc_41234_new_n4231_), .Y(_abc_41234_new_n4232_));
AOI21X1 AOI21X1_424 ( .A(_abc_41234_new_n3916_), .B(sp_15_), .C(_abc_41234_new_n534__bF_buf0), .Y(_abc_41234_new_n4240_));
AOI21X1 AOI21X1_425 ( .A(_abc_41234_new_n1106_), .B(regfil_4__7_), .C(_abc_41234_new_n1047__bF_buf3), .Y(_abc_41234_new_n4246_));
AOI21X1 AOI21X1_426 ( .A(_abc_41234_new_n4245_), .B(_abc_41234_new_n2463_), .C(_abc_41234_new_n4247_), .Y(_abc_41234_new_n4248_));
AOI21X1 AOI21X1_427 ( .A(_abc_41234_new_n4248_), .B(_abc_41234_new_n4244_), .C(_abc_41234_new_n4249_), .Y(_abc_41234_new_n4250_));
AOI21X1 AOI21X1_428 ( .A(_abc_41234_new_n4241_), .B(_abc_41234_new_n4250_), .C(_abc_41234_new_n4254_), .Y(_abc_41234_new_n4255_));
AOI21X1 AOI21X1_429 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n2563_), .C(_abc_41234_new_n1634_), .Y(_abc_41234_new_n4281_));
AOI21X1 AOI21X1_43 ( .A(_abc_41234_new_n1214_), .B(regfil_4__0_), .C(_abc_41234_new_n1219_), .Y(_abc_41234_new_n1220_));
AOI21X1 AOI21X1_430 ( .A(_abc_41234_new_n4318_), .B(_abc_41234_new_n4276_), .C(reset_bF_buf1), .Y(_0pc_15_0__0_));
AOI21X1 AOI21X1_431 ( .A(_abc_41234_new_n1646_), .B(_abc_41234_new_n4297__bF_buf1), .C(_abc_41234_new_n4324_), .Y(_abc_41234_new_n4325_));
AOI21X1 AOI21X1_432 ( .A(_abc_41234_new_n1646_), .B(_abc_41234_new_n4301_), .C(_abc_41234_new_n4330_), .Y(_abc_41234_new_n4331_));
AOI21X1 AOI21X1_433 ( .A(_abc_41234_new_n4335_), .B(_abc_41234_new_n4336_), .C(reset_bF_buf0), .Y(_0pc_15_0__1_));
AOI21X1 AOI21X1_434 ( .A(_abc_41234_new_n665__bF_buf3), .B(_abc_41234_new_n4338_), .C(_abc_41234_new_n4297__bF_buf0), .Y(_abc_41234_new_n4339_));
AOI21X1 AOI21X1_435 ( .A(_abc_41234_new_n4295_), .B(_abc_41234_new_n2735_), .C(_abc_41234_new_n4340_), .Y(_abc_41234_new_n4341_));
AOI21X1 AOI21X1_436 ( .A(_abc_41234_new_n4301_), .B(_abc_41234_new_n4338_), .C(_abc_41234_new_n4345_), .Y(_abc_41234_new_n4346_));
AOI21X1 AOI21X1_437 ( .A(_abc_41234_new_n4350_), .B(_abc_41234_new_n4351_), .C(reset_bF_buf9), .Y(_0pc_15_0__2_));
AOI21X1 AOI21X1_438 ( .A(_abc_41234_new_n1303_), .B(regfil_5__3_bF_buf2_), .C(_abc_41234_new_n528_), .Y(_abc_41234_new_n4362_));
AOI21X1 AOI21X1_439 ( .A(_abc_41234_new_n2776_), .B(_abc_41234_new_n4309_), .C(_abc_41234_new_n4363_), .Y(_abc_41234_new_n4364_));
AOI21X1 AOI21X1_44 ( .A(_abc_41234_new_n1205_), .B(_abc_41234_new_n1233_), .C(_abc_41234_new_n1066__bF_buf3), .Y(_abc_41234_new_n1234_));
AOI21X1 AOI21X1_440 ( .A(_abc_41234_new_n4368_), .B(_abc_41234_new_n4369_), .C(reset_bF_buf8), .Y(_0pc_15_0__3_));
AOI21X1 AOI21X1_441 ( .A(_abc_41234_new_n2806_), .B(_abc_41234_new_n4297__bF_buf0), .C(_abc_41234_new_n4374_), .Y(_abc_41234_new_n4375_));
AOI21X1 AOI21X1_442 ( .A(_abc_41234_new_n2805_), .B(_abc_41234_new_n4309_), .C(_abc_41234_new_n4378_), .Y(_abc_41234_new_n4379_));
AOI21X1 AOI21X1_443 ( .A(_abc_41234_new_n2801_), .B(_abc_41234_new_n4308_), .C(_abc_41234_new_n4380_), .Y(_abc_41234_new_n4381_));
AOI21X1 AOI21X1_444 ( .A(_abc_41234_new_n4382_), .B(_abc_41234_new_n4054_), .C(_abc_41234_new_n4385_), .Y(_abc_41234_new_n4386_));
AOI21X1 AOI21X1_445 ( .A(_abc_41234_new_n4377_), .B(_abc_41234_new_n4386_), .C(reset_bF_buf7), .Y(_0pc_15_0__4_));
AOI21X1 AOI21X1_446 ( .A(_abc_41234_new_n4389_), .B(_abc_41234_new_n4393_), .C(_abc_41234_new_n4394_), .Y(_abc_41234_new_n4395_));
AOI21X1 AOI21X1_447 ( .A(regfil_5__5_), .B(_abc_41234_new_n1303_), .C(_abc_41234_new_n4397_), .Y(_abc_41234_new_n4398_));
AOI21X1 AOI21X1_448 ( .A(opcode_5_bF_buf1_), .B(_abc_41234_new_n1637_), .C(_abc_41234_new_n4399_), .Y(_abc_41234_new_n4400_));
AOI21X1 AOI21X1_449 ( .A(_abc_41234_new_n4404_), .B(_abc_41234_new_n4405_), .C(reset_bF_buf6), .Y(_0pc_15_0__5_));
AOI21X1 AOI21X1_45 ( .A(_abc_41234_new_n1149_), .B(_abc_41234_new_n1267_), .C(_abc_41234_new_n1269_), .Y(_abc_41234_new_n1270_));
AOI21X1 AOI21X1_450 ( .A(_abc_41234_new_n4295_), .B(_abc_41234_new_n2854_), .C(_abc_41234_new_n4412_), .Y(_abc_41234_new_n4413_));
AOI21X1 AOI21X1_451 ( .A(_abc_41234_new_n4308_), .B(_abc_41234_new_n2854_), .C(_abc_41234_new_n4418_), .Y(_abc_41234_new_n4419_));
AOI21X1 AOI21X1_452 ( .A(_abc_41234_new_n4423_), .B(_abc_41234_new_n4424_), .C(reset_bF_buf5), .Y(_0pc_15_0__6_));
AOI21X1 AOI21X1_453 ( .A(_abc_41234_new_n4407_), .B(pc_6_), .C(pc_7_), .Y(_abc_41234_new_n4428_));
AOI21X1 AOI21X1_454 ( .A(_abc_41234_new_n4301_), .B(_abc_41234_new_n4429_), .C(_abc_41234_new_n4432_), .Y(_abc_41234_new_n4433_));
AOI21X1 AOI21X1_455 ( .A(_abc_41234_new_n4429_), .B(_abc_41234_new_n665__bF_buf1), .C(_abc_41234_new_n4297__bF_buf2), .Y(_abc_41234_new_n4437_));
AOI21X1 AOI21X1_456 ( .A(_abc_41234_new_n4295_), .B(_abc_41234_new_n4436_), .C(_abc_41234_new_n4438_), .Y(_abc_41234_new_n4439_));
AOI21X1 AOI21X1_457 ( .A(_abc_41234_new_n4442_), .B(_abc_41234_new_n4443_), .C(reset_bF_buf4), .Y(_0pc_15_0__7_));
AOI21X1 AOI21X1_458 ( .A(_abc_41234_new_n1622_), .B(_abc_41234_new_n4297__bF_buf0), .C(_abc_41234_new_n4451_), .Y(_abc_41234_new_n4452_));
AOI21X1 AOI21X1_459 ( .A(_abc_41234_new_n4460_), .B(_abc_41234_new_n4461_), .C(reset_bF_buf3), .Y(_0pc_15_0__8_));
AOI21X1 AOI21X1_46 ( .A(_abc_41234_new_n1195_), .B(_abc_41234_new_n1273_), .C(_abc_41234_new_n1199_), .Y(_abc_41234_new_n1278_));
AOI21X1 AOI21X1_460 ( .A(_abc_41234_new_n4308_), .B(_abc_41234_new_n1680_), .C(_abc_41234_new_n4468_), .Y(_abc_41234_new_n4469_));
AOI21X1 AOI21X1_461 ( .A(_abc_41234_new_n4477_), .B(_abc_41234_new_n4478_), .C(reset_bF_buf2), .Y(_0pc_15_0__9_));
AOI21X1 AOI21X1_462 ( .A(_abc_41234_new_n4295_), .B(_abc_41234_new_n1716_), .C(_abc_41234_new_n4485_), .Y(_abc_41234_new_n4486_));
AOI21X1 AOI21X1_463 ( .A(_abc_41234_new_n4486_), .B(_abc_41234_new_n4484_), .C(_abc_41234_new_n4487_), .Y(_abc_41234_new_n4488_));
AOI21X1 AOI21X1_464 ( .A(_abc_41234_new_n4496_), .B(_abc_41234_new_n4497_), .C(reset_bF_buf1), .Y(_0pc_15_0__10_));
AOI21X1 AOI21X1_465 ( .A(_abc_41234_new_n4514_), .B(_abc_41234_new_n4515_), .C(reset_bF_buf0), .Y(_0pc_15_0__11_));
AOI21X1 AOI21X1_466 ( .A(_abc_41234_new_n4534_), .B(_abc_41234_new_n4535_), .C(reset_bF_buf9), .Y(_0pc_15_0__12_));
AOI21X1 AOI21X1_467 ( .A(_abc_41234_new_n4297__bF_buf0), .B(_abc_41234_new_n1775_), .C(_abc_41234_new_n534__bF_buf3), .Y(_abc_41234_new_n4542_));
AOI21X1 AOI21X1_468 ( .A(_abc_41234_new_n4552_), .B(_abc_41234_new_n4553_), .C(reset_bF_buf8), .Y(_0pc_15_0__13_));
AOI21X1 AOI21X1_469 ( .A(_abc_41234_new_n4297__bF_buf2), .B(_abc_41234_new_n1798_), .C(_abc_41234_new_n534__bF_buf2), .Y(_abc_41234_new_n4563_));
AOI21X1 AOI21X1_47 ( .A(_abc_41234_new_n1155_), .B(_abc_41234_new_n1144_), .C(_abc_41234_new_n1108_), .Y(_abc_41234_new_n1281_));
AOI21X1 AOI21X1_470 ( .A(_abc_41234_new_n4312_), .B(pc_14_), .C(_abc_41234_new_n1576_), .Y(_abc_41234_new_n4569_));
AOI21X1 AOI21X1_471 ( .A(_abc_41234_new_n4573_), .B(_abc_41234_new_n4574_), .C(reset_bF_buf7), .Y(_0pc_15_0__14_));
AOI21X1 AOI21X1_472 ( .A(_abc_41234_new_n1826_), .B(_abc_41234_new_n1825_), .C(_abc_41234_new_n4329_), .Y(_abc_41234_new_n4588_));
AOI21X1 AOI21X1_473 ( .A(_abc_41234_new_n4596_), .B(_abc_41234_new_n4597_), .C(reset_bF_buf6), .Y(_0pc_15_0__15_));
AOI21X1 AOI21X1_474 ( .A(waitr), .B(_abc_41234_new_n4604_), .C(_abc_41234_new_n4606_), .Y(_abc_41234_new_n4607_));
AOI21X1 AOI21X1_475 ( .A(_abc_41234_new_n4607_), .B(_abc_41234_new_n4604_), .C(_abc_41234_new_n4609_), .Y(_0readmem_0_0_));
AOI21X1 AOI21X1_476 ( .A(rdatahold_0_), .B(_abc_41234_new_n4613_), .C(_abc_41234_new_n4617_), .Y(_abc_41234_new_n4618_));
AOI21X1 AOI21X1_477 ( .A(rdatahold_1_), .B(_abc_41234_new_n4613_), .C(_abc_41234_new_n4622_), .Y(_abc_41234_new_n4623_));
AOI21X1 AOI21X1_478 ( .A(rdatahold_2_), .B(_abc_41234_new_n4613_), .C(_abc_41234_new_n4627_), .Y(_abc_41234_new_n4628_));
AOI21X1 AOI21X1_479 ( .A(rdatahold_3_), .B(_abc_41234_new_n4613_), .C(_abc_41234_new_n4632_), .Y(_abc_41234_new_n4633_));
AOI21X1 AOI21X1_48 ( .A(_abc_41234_new_n1284_), .B(_abc_41234_new_n1249_), .C(_abc_41234_new_n1244_), .Y(_abc_41234_new_n1285_));
AOI21X1 AOI21X1_480 ( .A(rdatahold_4_), .B(_abc_41234_new_n4613_), .C(_abc_41234_new_n4637_), .Y(_abc_41234_new_n4638_));
AOI21X1 AOI21X1_481 ( .A(rdatahold_5_), .B(_abc_41234_new_n4613_), .C(_abc_41234_new_n4642_), .Y(_abc_41234_new_n4643_));
AOI21X1 AOI21X1_482 ( .A(rdatahold_6_), .B(_abc_41234_new_n4613_), .C(_abc_41234_new_n4647_), .Y(_abc_41234_new_n4648_));
AOI21X1 AOI21X1_483 ( .A(rdatahold_7_), .B(_abc_41234_new_n4613_), .C(_abc_41234_new_n4652_), .Y(_abc_41234_new_n4653_));
AOI21X1 AOI21X1_484 ( .A(raddrhold_8_), .B(_abc_41234_new_n2911_), .C(_abc_41234_new_n4656_), .Y(_abc_41234_new_n4657_));
AOI21X1 AOI21X1_485 ( .A(waddrhold_9_), .B(_abc_41234_new_n3609_), .C(_abc_41234_new_n4663_), .Y(_abc_41234_new_n4664_));
AOI21X1 AOI21X1_486 ( .A(waddrhold_10_), .B(_abc_41234_new_n3609_), .C(_abc_41234_new_n4668_), .Y(_abc_41234_new_n4669_));
AOI21X1 AOI21X1_487 ( .A(waddrhold_11_), .B(_abc_41234_new_n3609_), .C(_abc_41234_new_n4673_), .Y(_abc_41234_new_n4674_));
AOI21X1 AOI21X1_488 ( .A(raddrhold_12_), .B(_abc_41234_new_n2911_), .C(_abc_41234_new_n4677_), .Y(_abc_41234_new_n4678_));
AOI21X1 AOI21X1_489 ( .A(raddrhold_13_), .B(_abc_41234_new_n2911_), .C(_abc_41234_new_n4681_), .Y(_abc_41234_new_n4682_));
AOI21X1 AOI21X1_49 ( .A(_abc_41234_new_n1241_), .B(regfil_4__2_bF_buf1_), .C(_abc_41234_new_n1219_), .Y(_abc_41234_new_n1291_));
AOI21X1 AOI21X1_490 ( .A(waddrhold_14_), .B(_abc_41234_new_n3609_), .C(_abc_41234_new_n4686_), .Y(_abc_41234_new_n4687_));
AOI21X1 AOI21X1_491 ( .A(raddrhold_15_), .B(_abc_41234_new_n2911_), .C(_abc_41234_new_n4690_), .Y(_abc_41234_new_n4691_));
AOI21X1 AOI21X1_492 ( .A(_abc_41234_new_n4693_), .B(_abc_41234_new_n4612_), .C(reset_bF_buf0), .Y(_0readio_0_0_));
AOI21X1 AOI21X1_493 ( .A(_abc_41234_new_n4696_), .B(_abc_41234_new_n4607_), .C(_abc_41234_new_n4701_), .Y(_0inta_0_0_));
AOI21X1 AOI21X1_494 ( .A(_abc_41234_new_n2376_), .B(opcode_5_bF_buf4_), .C(_abc_41234_new_n2255_), .Y(_abc_41234_new_n4743_));
AOI21X1 AOI21X1_495 ( .A(_abc_41234_new_n555_), .B(zero), .C(_abc_41234_new_n4745_), .Y(_abc_41234_new_n4746_));
AOI21X1 AOI21X1_496 ( .A(_abc_41234_new_n669__bF_buf2), .B(_abc_41234_new_n2376_), .C(_abc_41234_new_n4746_), .Y(_abc_41234_new_n4747_));
AOI21X1 AOI21X1_497 ( .A(_abc_41234_new_n4747_), .B(_abc_41234_new_n4744_), .C(_abc_41234_new_n4740_), .Y(_abc_41234_new_n4748_));
AOI21X1 AOI21X1_498 ( .A(_abc_41234_new_n516__bF_buf1), .B(_abc_41234_new_n2630_), .C(_abc_41234_new_n4754_), .Y(_abc_41234_new_n4755_));
AOI21X1 AOI21X1_499 ( .A(_abc_41234_new_n692_), .B(_abc_41234_new_n2213_), .C(_abc_41234_new_n4758_), .Y(_abc_41234_new_n4759_));
AOI21X1 AOI21X1_5 ( .A(_abc_41234_new_n745_), .B(_abc_41234_new_n744_), .C(_abc_41234_new_n647_), .Y(_abc_41234_new_n746_));
AOI21X1 AOI21X1_50 ( .A(_abc_41234_new_n1257_), .B(_abc_41234_new_n1256_), .C(_abc_41234_new_n1252_), .Y(_abc_41234_new_n1296_));
AOI21X1 AOI21X1_500 ( .A(_abc_41234_new_n2535_), .B(_abc_41234_new_n4811_), .C(_abc_41234_new_n551_), .Y(_abc_41234_new_n4883_));
AOI21X1 AOI21X1_501 ( .A(_abc_41234_new_n2355_), .B(ei), .C(eienb), .Y(_abc_41234_new_n4889_));
AOI21X1 AOI21X1_502 ( .A(alu__abc_40887_new_n54_), .B(alu__abc_40887_new_n47_), .C(alu__abc_40887_new_n50_), .Y(alu__abc_40887_new_n55_));
AOI21X1 AOI21X1_503 ( .A(alu__abc_40887_new_n53_), .B(alu__abc_40887_new_n55_), .C(alu__abc_40887_new_n63_), .Y(alu__abc_40887_new_n64_));
AOI21X1 AOI21X1_504 ( .A(alu__abc_40887_new_n66_), .B(alu__abc_40887_new_n38_), .C(alu__abc_40887_new_n37_), .Y(alu__abc_40887_new_n67_));
AOI21X1 AOI21X1_505 ( .A(alu__abc_40887_new_n75_), .B(alu__abc_40887_new_n77_), .C(alu__abc_40887_new_n80_), .Y(alu__abc_40887_new_n81_));
AOI21X1 AOI21X1_506 ( .A(alu__abc_40887_new_n85_), .B(alu__abc_40887_new_n88_), .C(alu__abc_40887_new_n95_), .Y(alu__abc_40887_new_n96_));
AOI21X1 AOI21X1_507 ( .A(alu__abc_40887_new_n130_), .B(alu__abc_40887_new_n126_), .C(alu__abc_40887_new_n131_), .Y(alu__abc_40887_new_n132_));
AOI21X1 AOI21X1_508 ( .A(alu__abc_40887_new_n84_), .B(alu__abc_40887_new_n146_), .C(alu__abc_40887_new_n120_), .Y(alu__abc_40887_new_n147_));
AOI21X1 AOI21X1_509 ( .A(alu__abc_40887_new_n153_), .B(alu__abc_40887_new_n147_), .C(alu__abc_40887_new_n133_), .Y(alu__abc_40887_new_n154_));
AOI21X1 AOI21X1_51 ( .A(_abc_41234_new_n1340_), .B(_abc_41234_new_n1292_), .C(_abc_41234_new_n1066__bF_buf2), .Y(_abc_41234_new_n1341_));
AOI21X1 AOI21X1_510 ( .A(alu__abc_40887_new_n130_), .B(alu__abc_40887_new_n126_), .C(alu__abc_40887_new_n49_), .Y(alu__abc_40887_new_n160_));
AOI21X1 AOI21X1_511 ( .A(alu__abc_40887_new_n91_), .B(alu__abc_40887_new_n45_), .C(alu__abc_40887_new_n167_), .Y(alu__abc_40887_new_n168_));
AOI21X1 AOI21X1_512 ( .A(alu__abc_40887_new_n171_), .B(alu__abc_40887_new_n130_), .C(alu__abc_40887_new_n169_), .Y(alu__abc_40887_new_n172_));
AOI21X1 AOI21X1_513 ( .A(alu__abc_40887_new_n161_), .B(alu__abc_40887_new_n164_), .C(alu__abc_40887_new_n173_), .Y(alu__abc_40887_new_n174_));
AOI21X1 AOI21X1_514 ( .A(alu__abc_40887_new_n176_), .B(alu__abc_40887_new_n152_), .C(alu__abc_40887_new_n124_), .Y(alu__abc_40887_new_n177_));
AOI21X1 AOI21X1_515 ( .A(alu__abc_40887_new_n145_), .B(alu__abc_40887_new_n157_), .C(alu__abc_40887_new_n185_), .Y(alu__abc_40887_new_n186_));
AOI21X1 AOI21X1_516 ( .A(alu__abc_40887_new_n175_), .B(alu__abc_40887_new_n179_), .C(alu__abc_40887_new_n188_), .Y(alu__abc_40887_new_n189_));
AOI21X1 AOI21X1_517 ( .A(alu__abc_40887_new_n163_), .B(alu__abc_40887_new_n165_), .C(alu__abc_40887_new_n193_), .Y(alu__abc_40887_new_n194_));
AOI21X1 AOI21X1_518 ( .A(alu__abc_40887_new_n196_), .B(alu__abc_40887_new_n159_), .C(alu__abc_40887_new_n187_), .Y(alu__abc_40887_new_n197_));
AOI21X1 AOI21X1_519 ( .A(alu__abc_40887_new_n207_), .B(alu__abc_40887_new_n209_), .C(alu__abc_40887_new_n212_), .Y(alu__abc_40887_new_n213_));
AOI21X1 AOI21X1_52 ( .A(_abc_41234_new_n1061_), .B(_abc_41234_new_n819_), .C(_abc_41234_new_n1344_), .Y(_abc_41234_new_n1345_));
AOI21X1 AOI21X1_520 ( .A(alu__abc_40887_new_n108_), .B(alu__abc_40887_new_n201_), .C(alu__abc_40887_new_n214_), .Y(alu__abc_40887_new_n215_));
AOI21X1 AOI21X1_521 ( .A(alu__abc_40887_new_n42_), .B(alu__abc_40887_new_n227_), .C(alu__abc_40887_new_n228_), .Y(alu__abc_40887_new_n229_));
AOI21X1 AOI21X1_522 ( .A(alu__abc_40887_new_n170_), .B(alu__abc_40887_new_n227_), .C(alu__abc_40887_new_n245_), .Y(alu__abc_40887_new_n246_));
AOI21X1 AOI21X1_523 ( .A(alu__abc_40887_new_n240_), .B(alu__abc_40887_new_n242_), .C(alu__abc_40887_new_n247_), .Y(alu__abc_40887_new_n248_));
AOI21X1 AOI21X1_524 ( .A(alu__abc_40887_new_n250_), .B(alu__abc_40887_new_n243_), .C(alu__abc_40887_new_n239_), .Y(alu__abc_40887_new_n251_));
AOI21X1 AOI21X1_525 ( .A(alu__abc_40887_new_n167_), .B(alu__abc_40887_new_n239_), .C(alu__abc_40887_new_n252_), .Y(alu__abc_40887_new_n253_));
AOI21X1 AOI21X1_526 ( .A(alu__abc_40887_new_n227_), .B(alu__abc_40887_new_n52_), .C(alu__abc_40887_new_n264_), .Y(alu__abc_40887_new_n265_));
AOI21X1 AOI21X1_527 ( .A(alu__abc_40887_new_n261_), .B(alu__abc_40887_new_n262_), .C(alu__abc_40887_new_n268_), .Y(alu__abc_40887_new_n269_));
AOI21X1 AOI21X1_528 ( .A(alu__abc_40887_new_n272_), .B(alu__abc_40887_new_n173_), .C(alu__abc_40887_new_n270_), .Y(alu__abc_40887_new_n273_));
AOI21X1 AOI21X1_529 ( .A(alu__abc_40887_new_n151_), .B(alu__abc_40887_new_n209_), .C(alu__abc_40887_new_n281_), .Y(alu__abc_40887_new_n282_));
AOI21X1 AOI21X1_53 ( .A(_abc_41234_new_n1370_), .B(_abc_41234_new_n1371_), .C(_abc_41234_new_n1152_), .Y(_abc_41234_new_n1372_));
AOI21X1 AOI21X1_530 ( .A(alu__abc_40887_new_n288_), .B(alu__abc_40887_new_n286_), .C(alu__abc_40887_new_n270_), .Y(alu__abc_40887_new_n289_));
AOI21X1 AOI21X1_531 ( .A(alu__abc_40887_new_n271_), .B(alu__abc_40887_new_n205_), .C(alu__abc_40887_new_n296_), .Y(alu__abc_40887_new_n297_));
AOI21X1 AOI21X1_532 ( .A(alu__abc_40887_new_n269_), .B(alu__abc_40887_new_n260_), .C(alu__abc_40887_new_n284_), .Y(alu__abc_40887_new_n303_));
AOI21X1 AOI21X1_533 ( .A(alu__abc_40887_new_n189_), .B(alu__abc_40887_new_n205_), .C(alu__abc_40887_new_n316_), .Y(alu__abc_40887_new_n317_));
AOI21X1 AOI21X1_534 ( .A(alu__abc_40887_new_n290_), .B(alu__abc_40887_new_n306_), .C(alu__abc_40887_new_n241_), .Y(alu__abc_40887_new_n320_));
AOI21X1 AOI21X1_535 ( .A(alu__abc_40887_new_n99_), .B(alu__abc_40887_new_n201_), .C(alu__abc_40887_new_n329_), .Y(alu__abc_40887_new_n330_));
AOI21X1 AOI21X1_536 ( .A(alu__abc_40887_new_n340_), .B(alu__abc_40887_new_n341_), .C(alu__abc_40887_new_n339_), .Y(alu__abc_40887_new_n346_));
AOI21X1 AOI21X1_537 ( .A(alu__abc_40887_new_n332_), .B(alu__abc_40887_new_n335_), .C(alu__abc_40887_new_n305_), .Y(alu__abc_40887_new_n347_));
AOI21X1 AOI21X1_54 ( .A(_abc_41234_new_n1329_), .B(_abc_41234_new_n1333_), .C(_abc_41234_new_n1332_), .Y(_abc_41234_new_n1374_));
AOI21X1 AOI21X1_55 ( .A(_abc_41234_new_n1383_), .B(_abc_41234_new_n1352_), .C(_abc_41234_new_n1066__bF_buf1), .Y(_abc_41234_new_n1384_));
AOI21X1 AOI21X1_56 ( .A(_abc_41234_new_n1061_), .B(_abc_41234_new_n849_), .C(_abc_41234_new_n1344_), .Y(_abc_41234_new_n1388_));
AOI21X1 AOI21X1_57 ( .A(_abc_41234_new_n1413_), .B(_abc_41234_new_n1313_), .C(_abc_41234_new_n1416_), .Y(_abc_41234_new_n1417_));
AOI21X1 AOI21X1_58 ( .A(_abc_41234_new_n1418_), .B(_abc_41234_new_n1421_), .C(_abc_41234_new_n1422_), .Y(_abc_41234_new_n1423_));
AOI21X1 AOI21X1_59 ( .A(_abc_41234_new_n1430_), .B(_abc_41234_new_n1327_), .C(_abc_41234_new_n1428_), .Y(_abc_41234_new_n1431_));
AOI21X1 AOI21X1_6 ( .A(alu_res_1_), .B(_abc_41234_new_n707_), .C(_abc_41234_new_n760_), .Y(_abc_41234_new_n761_));
AOI21X1 AOI21X1_60 ( .A(_abc_41234_new_n1155_), .B(_abc_41234_new_n819_), .C(_abc_41234_new_n1108_), .Y(_abc_41234_new_n1437_));
AOI21X1 AOI21X1_61 ( .A(_abc_41234_new_n1440_), .B(_abc_41234_new_n1399_), .C(_abc_41234_new_n1395_), .Y(_abc_41234_new_n1441_));
AOI21X1 AOI21X1_62 ( .A(_abc_41234_new_n1061_), .B(_abc_41234_new_n904_), .C(_abc_41234_new_n1344_), .Y(_abc_41234_new_n1445_));
AOI21X1 AOI21X1_63 ( .A(_abc_41234_new_n1426_), .B(_abc_41234_new_n1476_), .C(_abc_41234_new_n1199_), .Y(_abc_41234_new_n1480_));
AOI21X1 AOI21X1_64 ( .A(_abc_41234_new_n1418_), .B(_abc_41234_new_n1421_), .C(_abc_41234_new_n1485_), .Y(_abc_41234_new_n1486_));
AOI21X1 AOI21X1_65 ( .A(_abc_41234_new_n1487_), .B(_abc_41234_new_n1488_), .C(_abc_41234_new_n1489_), .Y(_abc_41234_new_n1490_));
AOI21X1 AOI21X1_66 ( .A(_abc_41234_new_n1116_), .B(_abc_41234_new_n1123_), .C(_abc_41234_new_n1491_), .Y(_abc_41234_new_n1492_));
AOI21X1 AOI21X1_67 ( .A(_abc_41234_new_n1495_), .B(_abc_41234_new_n1417_), .C(_abc_41234_new_n1497_), .Y(_abc_41234_new_n1498_));
AOI21X1 AOI21X1_68 ( .A(_abc_41234_new_n535_), .B(_abc_41234_new_n1470_), .C(_abc_41234_new_n1502_), .Y(_abc_41234_new_n1503_));
AOI21X1 AOI21X1_69 ( .A(_abc_41234_new_n1504_), .B(_abc_41234_new_n1455_), .C(_abc_41234_new_n1451_), .Y(_abc_41234_new_n1505_));
AOI21X1 AOI21X1_7 ( .A(_abc_41234_new_n744_), .B(regfil_0__2_), .C(_abc_41234_new_n600_), .Y(_abc_41234_new_n787_));
AOI21X1 AOI21X1_70 ( .A(_abc_41234_new_n1061_), .B(_abc_41234_new_n1509_), .C(_abc_41234_new_n1344_), .Y(_abc_41234_new_n1510_));
AOI21X1 AOI21X1_71 ( .A(_abc_41234_new_n1517_), .B(regfil_4__6_), .C(_abc_41234_new_n1218_), .Y(_abc_41234_new_n1518_));
AOI21X1 AOI21X1_72 ( .A(_abc_41234_new_n1406_), .B(_abc_41234_new_n1463_), .C(_abc_41234_new_n1521_), .Y(_abc_41234_new_n1522_));
AOI21X1 AOI21X1_73 ( .A(_abc_41234_new_n1418_), .B(_abc_41234_new_n1531_), .C(_abc_41234_new_n1532_), .Y(_abc_41234_new_n1533_));
AOI21X1 AOI21X1_74 ( .A(_abc_41234_new_n1433_), .B(_abc_41234_new_n1478_), .C(_abc_41234_new_n1542_), .Y(_abc_41234_new_n1549_));
AOI21X1 AOI21X1_75 ( .A(_abc_41234_new_n1155_), .B(_abc_41234_new_n904_), .C(_abc_41234_new_n1108_), .Y(_abc_41234_new_n1553_));
AOI21X1 AOI21X1_76 ( .A(_abc_41234_new_n1520_), .B(_abc_41234_new_n1555_), .C(_abc_41234_new_n1516_), .Y(_abc_41234_new_n1556_));
AOI21X1 AOI21X1_77 ( .A(_abc_41234_new_n1448_), .B(_abc_41234_new_n1509_), .C(regfil_4__7_), .Y(_abc_41234_new_n1563_));
AOI21X1 AOI21X1_78 ( .A(_abc_41234_new_n1546_), .B(_abc_41234_new_n1581_), .C(_abc_41234_new_n1199_), .Y(_abc_41234_new_n1585_));
AOI21X1 AOI21X1_79 ( .A(_abc_41234_new_n1588_), .B(_abc_41234_new_n1587_), .C(_abc_41234_new_n1592_), .Y(_abc_41234_new_n1593_));
AOI21X1 AOI21X1_8 ( .A(_abc_41234_new_n787_), .B(_abc_41234_new_n786_), .C(_abc_41234_new_n647_), .Y(_abc_41234_new_n788_));
AOI21X1 AOI21X1_80 ( .A(_abc_41234_new_n535_), .B(_abc_41234_new_n1576_), .C(_abc_41234_new_n1596_), .Y(_abc_41234_new_n1597_));
AOI21X1 AOI21X1_81 ( .A(_abc_41234_new_n1599_), .B(_abc_41234_new_n997_), .C(_abc_41234_new_n1263_), .Y(_abc_41234_new_n1600_));
AOI21X1 AOI21X1_82 ( .A(_abc_41234_new_n1622_), .B(intcyc_bF_buf3), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n1632_));
AOI21X1 AOI21X1_83 ( .A(_abc_41234_new_n1632_), .B(intcyc_bF_buf2), .C(_abc_41234_new_n1659_), .Y(_abc_41234_new_n1660_));
AOI21X1 AOI21X1_84 ( .A(intcyc_bF_buf1), .B(_abc_41234_new_n1670_), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n1675_));
AOI21X1 AOI21X1_85 ( .A(_abc_41234_new_n1682_), .B(_abc_41234_new_n1640_), .C(_abc_41234_new_n544__bF_buf3), .Y(_abc_41234_new_n1683_));
AOI21X1 AOI21X1_86 ( .A(regfil_4__1_bF_buf1_), .B(_abc_41234_new_n1683_), .C(_abc_41234_new_n1690_), .Y(_abc_41234_new_n1691_));
AOI21X1 AOI21X1_87 ( .A(intcyc_bF_buf3), .B(_abc_41234_new_n1705_), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n1711_));
AOI21X1 AOI21X1_88 ( .A(_abc_41234_new_n1644_), .B(_abc_41234_new_n1697_), .C(_abc_41234_new_n1047__bF_buf3), .Y(_abc_41234_new_n1721_));
AOI21X1 AOI21X1_89 ( .A(_abc_41234_new_n1734_), .B(_abc_41234_new_n1637_), .C(_abc_41234_new_n1740_), .Y(_abc_41234_new_n1741_));
AOI21X1 AOI21X1_9 ( .A(_abc_41234_new_n533_), .B(regfil_7__3_), .C(_abc_41234_new_n513_), .Y(_abc_41234_new_n799_));
AOI21X1 AOI21X1_90 ( .A(_abc_41234_new_n1644_), .B(_abc_41234_new_n1724_), .C(_abc_41234_new_n1047__bF_buf2), .Y(_abc_41234_new_n1743_));
AOI21X1 AOI21X1_91 ( .A(intcyc_bF_buf3), .B(_abc_41234_new_n1750_), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n1758_));
AOI21X1 AOI21X1_92 ( .A(_abc_41234_new_n1644_), .B(_abc_41234_new_n1746_), .C(_abc_41234_new_n1047__bF_buf1), .Y(_abc_41234_new_n1768_));
AOI21X1 AOI21X1_93 ( .A(intcyc_bF_buf1), .B(_abc_41234_new_n1775_), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n1776_));
AOI21X1 AOI21X1_94 ( .A(_abc_41234_new_n1780_), .B(_abc_41234_new_n1637_), .C(_abc_41234_new_n1787_), .Y(_abc_41234_new_n1788_));
AOI21X1 AOI21X1_95 ( .A(_abc_41234_new_n1644_), .B(_abc_41234_new_n1771_), .C(_abc_41234_new_n1047__bF_buf0), .Y(_abc_41234_new_n1790_));
AOI21X1 AOI21X1_96 ( .A(intcyc_bF_buf3), .B(_abc_41234_new_n1798_), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n1807_));
AOI21X1 AOI21X1_97 ( .A(_abc_41234_new_n1644_), .B(_abc_41234_new_n1793_), .C(_abc_41234_new_n1047__bF_buf4), .Y(_abc_41234_new_n1818_));
AOI21X1 AOI21X1_98 ( .A(intcyc_bF_buf1), .B(_abc_41234_new_n1828_), .C(_abc_41234_new_n1631_), .Y(_abc_41234_new_n1829_));
AOI21X1 AOI21X1_99 ( .A(_abc_41234_new_n1833_), .B(_abc_41234_new_n1637_), .C(_abc_41234_new_n1840_), .Y(_abc_41234_new_n1841_));
AOI22X1 AOI22X1_1 ( .A(_abc_41234_new_n514_), .B(_abc_41234_new_n533_), .C(_abc_41234_new_n563_), .D(_abc_41234_new_n554_), .Y(_abc_41234_new_n564_));
AOI22X1 AOI22X1_10 ( .A(alu_res_2_), .B(_abc_41234_new_n613_), .C(rdatahold_2_), .D(_abc_41234_new_n650_), .Y(_abc_41234_new_n780_));
AOI22X1 AOI22X1_100 ( .A(regfil_4__5_), .B(_abc_41234_new_n2247_), .C(regfil_5__5_), .D(_abc_41234_new_n2248_), .Y(_abc_41234_new_n2323_));
AOI22X1 AOI22X1_101 ( .A(rdatahold_5_), .B(_abc_41234_new_n2263_), .C(alu_opra_5_), .D(_abc_41234_new_n2266_), .Y(_abc_41234_new_n2328_));
AOI22X1 AOI22X1_102 ( .A(regfil_0__6_), .B(_abc_41234_new_n2247_), .C(regfil_2__6_), .D(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2331_));
AOI22X1 AOI22X1_103 ( .A(regfil_4__6_), .B(_abc_41234_new_n2247_), .C(regfil_5__6_bF_buf1_), .D(_abc_41234_new_n2248_), .Y(_abc_41234_new_n2335_));
AOI22X1 AOI22X1_104 ( .A(rdatahold_6_), .B(_abc_41234_new_n2263_), .C(alu_opra_6_), .D(_abc_41234_new_n2266_), .Y(_abc_41234_new_n2340_));
AOI22X1 AOI22X1_105 ( .A(regfil_7__7_), .B(_abc_41234_new_n2201_), .C(_abc_41234_new_n2208_), .D(_abc_41234_new_n2349_), .Y(_abc_41234_new_n2350_));
AOI22X1 AOI22X1_106 ( .A(_abc_41234_new_n1006_), .B(_abc_41234_new_n2261_), .C(alu_opra_7_), .D(_abc_41234_new_n2266_), .Y(_abc_41234_new_n2351_));
AOI22X1 AOI22X1_107 ( .A(_abc_41234_new_n509_), .B(_abc_41234_new_n2367_), .C(alu_parity), .D(_abc_41234_new_n2362_), .Y(_abc_41234_new_n2368_));
AOI22X1 AOI22X1_108 ( .A(_abc_41234_new_n509_), .B(_abc_41234_new_n2373_), .C(alu_zout), .D(_abc_41234_new_n2362_), .Y(_abc_41234_new_n2374_));
AOI22X1 AOI22X1_109 ( .A(_abc_41234_new_n516__bF_buf5), .B(eienb), .C(_abc_41234_new_n2450_), .D(_abc_41234_new_n2452_), .Y(_abc_41234_new_n2453_));
AOI22X1 AOI22X1_11 ( .A(_abc_41234_new_n602_), .B(_abc_41234_new_n781_), .C(_abc_41234_new_n788_), .D(_abc_41234_new_n785_), .Y(_abc_41234_new_n789_));
AOI22X1 AOI22X1_110 ( .A(statesel_1_), .B(_abc_41234_new_n2530_), .C(_abc_41234_new_n660__bF_buf0), .D(_abc_41234_new_n2554_), .Y(_abc_41234_new_n2555_));
AOI22X1 AOI22X1_111 ( .A(statesel_1_), .B(_abc_41234_new_n2528_), .C(_abc_41234_new_n2560_), .D(_abc_41234_new_n2535_), .Y(_abc_41234_new_n2561_));
AOI22X1 AOI22X1_112 ( .A(statesel_2_), .B(_abc_41234_new_n2530_), .C(_abc_41234_new_n660__bF_buf7), .D(_abc_41234_new_n2575_), .Y(_abc_41234_new_n2576_));
AOI22X1 AOI22X1_113 ( .A(statesel_2_), .B(_abc_41234_new_n2528_), .C(_abc_41234_new_n2585_), .D(_abc_41234_new_n2584_), .Y(_abc_41234_new_n2586_));
AOI22X1 AOI22X1_114 ( .A(statesel_5_), .B(_abc_41234_new_n2636_), .C(_abc_41234_new_n660__bF_buf4), .D(_abc_41234_new_n2632_), .Y(_abc_41234_new_n2637_));
AOI22X1 AOI22X1_115 ( .A(statesel_5_), .B(_abc_41234_new_n2528_), .C(_abc_41234_new_n2641_), .D(_abc_41234_new_n2535_), .Y(_abc_41234_new_n2642_));
AOI22X1 AOI22X1_116 ( .A(_abc_41234_new_n1630_), .B(_abc_41234_new_n2684_), .C(_abc_41234_new_n2689_), .D(_abc_41234_new_n2687_), .Y(_abc_41234_new_n2690_));
AOI22X1 AOI22X1_117 ( .A(_abc_41234_new_n2695_), .B(alu_res_0_), .C(wdatahold2_0_), .D(_abc_41234_new_n2696__bF_buf4), .Y(_abc_41234_new_n2697_));
AOI22X1 AOI22X1_118 ( .A(_abc_41234_new_n1627_), .B(_abc_41234_new_n2706_), .C(_abc_41234_new_n1630_), .D(_abc_41234_new_n2708_), .Y(_abc_41234_new_n2709_));
AOI22X1 AOI22X1_119 ( .A(wdatahold2_1_), .B(_abc_41234_new_n2696__bF_buf3), .C(_abc_41234_new_n2725_), .D(_abc_41234_new_n2724_), .Y(_abc_41234_new_n2726_));
AOI22X1 AOI22X1_12 ( .A(regfil_7__1_), .B(_abc_41234_new_n559_), .C(_abc_41234_new_n752_), .D(_abc_41234_new_n797_), .Y(_abc_41234_new_n798_));
AOI22X1 AOI22X1_120 ( .A(_abc_41234_new_n2695_), .B(alu_res_1_), .C(rdatahold_1_), .D(_abc_41234_new_n2727_), .Y(_abc_41234_new_n2728_));
AOI22X1 AOI22X1_121 ( .A(_abc_41234_new_n536__bF_buf2), .B(_abc_41234_new_n2740_), .C(regfil_5__2_), .D(_abc_41234_new_n537__bF_buf1), .Y(_abc_41234_new_n2741_));
AOI22X1 AOI22X1_122 ( .A(_abc_41234_new_n581_), .B(_abc_41234_new_n2765_), .C(_abc_41234_new_n1627_), .D(_abc_41234_new_n2776_), .Y(_abc_41234_new_n2782_));
AOI22X1 AOI22X1_123 ( .A(_abc_41234_new_n2695_), .B(alu_res_3_), .C(wdatahold2_3_), .D(_abc_41234_new_n2696__bF_buf2), .Y(_abc_41234_new_n2788_));
AOI22X1 AOI22X1_124 ( .A(_abc_41234_new_n2695_), .B(alu_res_4_), .C(wdatahold2_4_), .D(_abc_41234_new_n2696__bF_buf1), .Y(_abc_41234_new_n2820_));
AOI22X1 AOI22X1_125 ( .A(_abc_41234_new_n2695_), .B(alu_res_5_), .C(wdatahold2_5_), .D(_abc_41234_new_n2696__bF_buf0), .Y(_abc_41234_new_n2847_));
AOI22X1 AOI22X1_126 ( .A(_abc_41234_new_n1630_), .B(_abc_41234_new_n2866_), .C(regfil_5__6_bF_buf3_), .D(_abc_41234_new_n1041_), .Y(_abc_41234_new_n2867_));
AOI22X1 AOI22X1_127 ( .A(_abc_41234_new_n2695_), .B(alu_res_6_), .C(wdatahold2_6_), .D(_abc_41234_new_n2696__bF_buf4), .Y(_abc_41234_new_n2877_));
AOI22X1 AOI22X1_128 ( .A(_abc_41234_new_n536__bF_buf3), .B(_abc_41234_new_n2890_), .C(regfil_5__7_), .D(_abc_41234_new_n537__bF_buf0), .Y(_abc_41234_new_n2891_));
AOI22X1 AOI22X1_129 ( .A(_abc_41234_new_n2727_), .B(rdatahold_7_), .C(wdatahold2_7_), .D(_abc_41234_new_n2696__bF_buf3), .Y(_abc_41234_new_n2906_));
AOI22X1 AOI22X1_13 ( .A(_abc_41234_new_n794_), .B(_abc_41234_new_n513_), .C(_abc_41234_new_n799_), .D(_abc_41234_new_n798_), .Y(_abc_41234_new_n800_));
AOI22X1 AOI22X1_130 ( .A(rdatahold2_1_), .B(_abc_41234_new_n2513_), .C(_abc_41234_new_n660__bF_buf4), .D(_abc_41234_new_n2984_), .Y(_abc_41234_new_n2985_));
AOI22X1 AOI22X1_131 ( .A(_abc_41234_new_n2988_), .B(_abc_41234_new_n2990_), .C(raddrhold_1_), .D(_abc_41234_new_n2913_), .Y(_abc_41234_new_n2991_));
AOI22X1 AOI22X1_132 ( .A(_abc_41234_new_n2996_), .B(_abc_41234_new_n2999_), .C(_abc_41234_new_n669__bF_buf0), .D(_abc_41234_new_n2997_), .Y(_abc_41234_new_n3000_));
AOI22X1 AOI22X1_133 ( .A(_abc_41234_new_n2990_), .B(_abc_41234_new_n3020_), .C(raddrhold_2_), .D(_abc_41234_new_n2913_), .Y(_abc_41234_new_n3021_));
AOI22X1 AOI22X1_134 ( .A(_abc_41234_new_n2996_), .B(_abc_41234_new_n3031_), .C(_abc_41234_new_n669__bF_buf3), .D(_abc_41234_new_n3029_), .Y(_abc_41234_new_n3032_));
AOI22X1 AOI22X1_135 ( .A(_abc_41234_new_n2996_), .B(_abc_41234_new_n3056_), .C(_abc_41234_new_n669__bF_buf2), .D(_abc_41234_new_n3054_), .Y(_abc_41234_new_n3057_));
AOI22X1 AOI22X1_136 ( .A(_abc_41234_new_n2996_), .B(_abc_41234_new_n3083_), .C(_abc_41234_new_n669__bF_buf1), .D(_abc_41234_new_n3081_), .Y(_abc_41234_new_n3084_));
AOI22X1 AOI22X1_137 ( .A(_abc_41234_new_n2996_), .B(_abc_41234_new_n3106_), .C(_abc_41234_new_n2854_), .D(_abc_41234_new_n2917_), .Y(_abc_41234_new_n3107_));
AOI22X1 AOI22X1_138 ( .A(_abc_41234_new_n1687_), .B(_abc_41234_new_n2996_), .C(_abc_41234_new_n2917_), .D(_abc_41234_new_n1680_), .Y(_abc_41234_new_n3182_));
AOI22X1 AOI22X1_139 ( .A(_abc_41234_new_n3208_), .B(_abc_41234_new_n2996_), .C(_abc_41234_new_n2917_), .D(_abc_41234_new_n1716_), .Y(_abc_41234_new_n3209_));
AOI22X1 AOI22X1_14 ( .A(_abc_41234_new_n707_), .B(alu_res_2_), .C(\data[2] ), .D(_abc_41234_new_n758_), .Y(_abc_41234_new_n801_));
AOI22X1 AOI22X1_140 ( .A(_abc_41234_new_n3228_), .B(_abc_41234_new_n2996_), .C(_abc_41234_new_n2917_), .D(_abc_41234_new_n1734_), .Y(_abc_41234_new_n3229_));
AOI22X1 AOI22X1_141 ( .A(_abc_41234_new_n3233_), .B(_abc_41234_new_n3234_), .C(_abc_41234_new_n3231_), .D(_abc_41234_new_n3230_), .Y(_abc_41234_new_n3235_));
AOI22X1 AOI22X1_142 ( .A(_abc_41234_new_n2996_), .B(_abc_41234_new_n3249_), .C(_abc_41234_new_n3250_), .D(_abc_41234_new_n3251_), .Y(_abc_41234_new_n3252_));
AOI22X1 AOI22X1_143 ( .A(_abc_41234_new_n3234_), .B(_abc_41234_new_n3259_), .C(raddrhold_12_), .D(_abc_41234_new_n3260_), .Y(_abc_41234_new_n3261_));
AOI22X1 AOI22X1_144 ( .A(raddrhold_14_), .B(_abc_41234_new_n2951__bF_buf2), .C(_abc_41234_new_n3306_), .D(_abc_41234_new_n3234_), .Y(_abc_41234_new_n3307_));
AOI22X1 AOI22X1_145 ( .A(raddrhold_15_), .B(_abc_41234_new_n2951__bF_buf1), .C(_abc_41234_new_n3329_), .D(_abc_41234_new_n3234_), .Y(_abc_41234_new_n3330_));
AOI22X1 AOI22X1_146 ( .A(rdatahold2_0_), .B(_abc_41234_new_n3353_), .C(_abc_41234_new_n3337_), .D(_abc_41234_new_n2696__bF_buf2), .Y(_abc_41234_new_n3354_));
AOI22X1 AOI22X1_147 ( .A(rdatahold2_1_), .B(_abc_41234_new_n3353_), .C(_abc_41234_new_n3376_), .D(_abc_41234_new_n2696__bF_buf1), .Y(_abc_41234_new_n3377_));
AOI22X1 AOI22X1_148 ( .A(rdatahold2_2_), .B(_abc_41234_new_n3353_), .C(_abc_41234_new_n3398_), .D(_abc_41234_new_n2696__bF_buf0), .Y(_abc_41234_new_n3399_));
AOI22X1 AOI22X1_149 ( .A(rdatahold2_3_), .B(_abc_41234_new_n3353_), .C(_abc_41234_new_n3416_), .D(_abc_41234_new_n3417_), .Y(_abc_41234_new_n3418_));
AOI22X1 AOI22X1_15 ( .A(alu_res_3_), .B(_abc_41234_new_n613_), .C(_abc_41234_new_n825_), .D(_abc_41234_new_n657_), .Y(_abc_41234_new_n826_));
AOI22X1 AOI22X1_150 ( .A(rdatahold2_4_), .B(_abc_41234_new_n3353_), .C(regfil_5__4_), .D(_abc_41234_new_n2695_), .Y(_abc_41234_new_n3438_));
AOI22X1 AOI22X1_151 ( .A(rdatahold2_5_), .B(_abc_41234_new_n3353_), .C(regfil_5__5_), .D(_abc_41234_new_n2695_), .Y(_abc_41234_new_n3460_));
AOI22X1 AOI22X1_152 ( .A(rdatahold2_6_), .B(_abc_41234_new_n3353_), .C(regfil_5__6_bF_buf0_), .D(_abc_41234_new_n2695_), .Y(_abc_41234_new_n3480_));
AOI22X1 AOI22X1_153 ( .A(rdatahold2_7_), .B(_abc_41234_new_n3353_), .C(regfil_5__7_), .D(_abc_41234_new_n2695_), .Y(_abc_41234_new_n3501_));
AOI22X1 AOI22X1_154 ( .A(rdatahold_0_), .B(_abc_41234_new_n3353_), .C(regfil_4__0_), .D(_abc_41234_new_n2695_), .Y(_abc_41234_new_n3519_));
AOI22X1 AOI22X1_155 ( .A(rdatahold_1_), .B(_abc_41234_new_n3353_), .C(regfil_4__1_bF_buf0_), .D(_abc_41234_new_n2695_), .Y(_abc_41234_new_n3541_));
AOI22X1 AOI22X1_156 ( .A(rdatahold_2_), .B(_abc_41234_new_n3353_), .C(regfil_4__2_bF_buf0_), .D(_abc_41234_new_n2695_), .Y(_abc_41234_new_n3562_));
AOI22X1 AOI22X1_157 ( .A(rdatahold_3_), .B(_abc_41234_new_n3353_), .C(regfil_4__3_), .D(_abc_41234_new_n2695_), .Y(_abc_41234_new_n3584_));
AOI22X1 AOI22X1_158 ( .A(waddrhold_12_), .B(_abc_41234_new_n3338_), .C(_abc_41234_new_n3611_), .D(_abc_41234_new_n3608_), .Y(_abc_41234_new_n3612_));
AOI22X1 AOI22X1_159 ( .A(waddrhold_14_), .B(_abc_41234_new_n3338_), .C(_abc_41234_new_n3609_), .D(_abc_41234_new_n3653_), .Y(_abc_41234_new_n3654_));
AOI22X1 AOI22X1_16 ( .A(_abc_41234_new_n707_), .B(alu_res_3_), .C(\data[3] ), .D(_abc_41234_new_n758_), .Y(_abc_41234_new_n843_));
AOI22X1 AOI22X1_160 ( .A(_abc_41234_new_n2458_), .B(_abc_41234_new_n2481_), .C(_abc_41234_new_n3657_), .D(_abc_41234_new_n3658_), .Y(_abc_41234_new_n3659_));
AOI22X1 AOI22X1_161 ( .A(wdatahold_0_), .B(_abc_41234_new_n3609_), .C(regfil_7__0_), .D(_abc_41234_new_n3677_), .Y(_abc_41234_new_n3678_));
AOI22X1 AOI22X1_162 ( .A(wdatahold_1_), .B(_abc_41234_new_n3609_), .C(regfil_7__1_), .D(_abc_41234_new_n3677_), .Y(_abc_41234_new_n3680_));
AOI22X1 AOI22X1_163 ( .A(wdatahold_2_), .B(_abc_41234_new_n3609_), .C(regfil_7__2_), .D(_abc_41234_new_n3677_), .Y(_abc_41234_new_n3682_));
AOI22X1 AOI22X1_164 ( .A(wdatahold_3_), .B(_abc_41234_new_n3609_), .C(regfil_7__3_), .D(_abc_41234_new_n3677_), .Y(_abc_41234_new_n3684_));
AOI22X1 AOI22X1_165 ( .A(wdatahold_4_), .B(_abc_41234_new_n3609_), .C(regfil_7__4_), .D(_abc_41234_new_n3677_), .Y(_abc_41234_new_n3686_));
AOI22X1 AOI22X1_166 ( .A(wdatahold_5_), .B(_abc_41234_new_n3609_), .C(regfil_7__5_), .D(_abc_41234_new_n3677_), .Y(_abc_41234_new_n3688_));
AOI22X1 AOI22X1_167 ( .A(wdatahold_6_), .B(_abc_41234_new_n3609_), .C(regfil_7__6_), .D(_abc_41234_new_n3677_), .Y(_abc_41234_new_n3690_));
AOI22X1 AOI22X1_168 ( .A(wdatahold_7_), .B(_abc_41234_new_n3609_), .C(regfil_7__7_), .D(_abc_41234_new_n3677_), .Y(_abc_41234_new_n3692_));
AOI22X1 AOI22X1_169 ( .A(_abc_41234_new_n555_), .B(_abc_41234_new_n3697_), .C(_abc_41234_new_n673_), .D(_abc_41234_new_n3698_), .Y(_abc_41234_new_n3699_));
AOI22X1 AOI22X1_17 ( .A(alu_res_4_), .B(_abc_41234_new_n613_), .C(rdatahold_4_), .D(_abc_41234_new_n650_), .Y(_abc_41234_new_n864_));
AOI22X1 AOI22X1_170 ( .A(_abc_41234_new_n515__bF_buf3), .B(_abc_41234_new_n3699_), .C(_abc_41234_new_n3695_), .D(_abc_41234_new_n3696_), .Y(_abc_41234_new_n3700_));
AOI22X1 AOI22X1_171 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n3697_), .C(_abc_41234_new_n654_), .D(_abc_41234_new_n3698_), .Y(_abc_41234_new_n3705_));
AOI22X1 AOI22X1_172 ( .A(_abc_41234_new_n515__bF_buf2), .B(_abc_41234_new_n3705_), .C(_abc_41234_new_n3704_), .D(_abc_41234_new_n3703_), .Y(_abc_41234_new_n3706_));
AOI22X1 AOI22X1_173 ( .A(_abc_41234_new_n536__bF_buf1), .B(_abc_41234_new_n3697_), .C(_abc_41234_new_n649_), .D(_abc_41234_new_n3698_), .Y(_abc_41234_new_n3711_));
AOI22X1 AOI22X1_174 ( .A(_abc_41234_new_n515__bF_buf1), .B(_abc_41234_new_n3711_), .C(_abc_41234_new_n3710_), .D(_abc_41234_new_n3709_), .Y(_abc_41234_new_n3712_));
AOI22X1 AOI22X1_175 ( .A(_abc_41234_new_n1200_), .B(_abc_41234_new_n3724_), .C(_abc_41234_new_n3721_), .D(_abc_41234_new_n1151_), .Y(_abc_41234_new_n3725_));
AOI22X1 AOI22X1_176 ( .A(rdatahold2_0_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n3718_), .D(_abc_41234_new_n3727_), .Y(_abc_41234_new_n3728_));
AOI22X1 AOI22X1_177 ( .A(rdatahold2_2_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n3758_), .D(_abc_41234_new_n3777_), .Y(_abc_41234_new_n3778_));
AOI22X1 AOI22X1_178 ( .A(_abc_41234_new_n1309_), .B(_abc_41234_new_n3792_), .C(_abc_41234_new_n3790_), .D(_abc_41234_new_n3789_), .Y(_abc_41234_new_n3793_));
AOI22X1 AOI22X1_179 ( .A(_abc_41234_new_n1206_), .B(_abc_41234_new_n3809_), .C(_abc_41234_new_n3822_), .D(_abc_41234_new_n3820_), .Y(_abc_41234_new_n3823_));
AOI22X1 AOI22X1_18 ( .A(_abc_41234_new_n602_), .B(_abc_41234_new_n865_), .C(_abc_41234_new_n874_), .D(_abc_41234_new_n877_), .Y(_abc_41234_new_n878_));
AOI22X1 AOI22X1_180 ( .A(_abc_41234_new_n1206_), .B(_abc_41234_new_n3877_), .C(_abc_41234_new_n3874_), .D(_abc_41234_new_n3870_), .Y(_abc_41234_new_n3878_));
AOI22X1 AOI22X1_181 ( .A(rdatahold2_7_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1055_), .D(_abc_41234_new_n3882_), .Y(_abc_41234_new_n3883_));
AOI22X1 AOI22X1_182 ( .A(_abc_41234_new_n3964_), .B(rdatahold2_2_), .C(_abc_41234_new_n3385_), .D(_abc_41234_new_n3963_), .Y(_abc_41234_new_n3965_));
AOI22X1 AOI22X1_183 ( .A(_abc_41234_new_n1106_), .B(regfil_5__3_bF_buf3_), .C(_abc_41234_new_n2462_), .D(_abc_41234_new_n3971_), .Y(_abc_41234_new_n3972_));
AOI22X1 AOI22X1_184 ( .A(_abc_41234_new_n2452_), .B(_abc_41234_new_n3977_), .C(_abc_41234_new_n3978_), .D(_abc_41234_new_n3980_), .Y(_abc_41234_new_n3981_));
AOI22X1 AOI22X1_185 ( .A(_abc_41234_new_n515__bF_buf3), .B(_abc_41234_new_n4044_), .C(sp_6_), .D(_abc_41234_new_n4012_), .Y(_abc_41234_new_n4045_));
AOI22X1 AOI22X1_186 ( .A(_abc_41234_new_n3469_), .B(_abc_41234_new_n3963_), .C(_abc_41234_new_n3960_), .D(_abc_41234_new_n4047_), .Y(_abc_41234_new_n4048_));
AOI22X1 AOI22X1_187 ( .A(rdatahold2_7_), .B(_abc_41234_new_n3964_), .C(_abc_41234_new_n3963_), .D(_abc_41234_new_n3490_), .Y(_abc_41234_new_n4075_));
AOI22X1 AOI22X1_188 ( .A(_abc_41234_new_n3508_), .B(_abc_41234_new_n3963_), .C(_abc_41234_new_n3960_), .D(_abc_41234_new_n4082_), .Y(_abc_41234_new_n4097_));
AOI22X1 AOI22X1_189 ( .A(regfil_4__1_bF_buf3_), .B(_abc_41234_new_n1106_), .C(_abc_41234_new_n2463_), .D(_abc_41234_new_n3530_), .Y(_abc_41234_new_n4111_));
AOI22X1 AOI22X1_19 ( .A(alu_res_4_), .B(_abc_41234_new_n707_), .C(regfil_7__4_), .D(_abc_41234_new_n703_), .Y(_abc_41234_new_n891_));
AOI22X1 AOI22X1_190 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n4114_), .C(sp_9_), .D(_abc_41234_new_n4112_), .Y(_abc_41234_new_n4115_));
AOI22X1 AOI22X1_191 ( .A(_abc_41234_new_n3530_), .B(_abc_41234_new_n3963_), .C(_abc_41234_new_n3960_), .D(_abc_41234_new_n4114_), .Y(_abc_41234_new_n4119_));
AOI22X1 AOI22X1_192 ( .A(sp_10_), .B(_abc_41234_new_n4012_), .C(_abc_41234_new_n1046__bF_buf2), .D(_abc_41234_new_n4137_), .Y(_abc_41234_new_n4138_));
AOI22X1 AOI22X1_193 ( .A(regfil_4__4_), .B(_abc_41234_new_n1106_), .C(_abc_41234_new_n2463_), .D(_abc_41234_new_n3595_), .Y(_abc_41234_new_n4181_));
AOI22X1 AOI22X1_194 ( .A(sp_12_), .B(_abc_41234_new_n4012_), .C(_abc_41234_new_n1046__bF_buf0), .D(_abc_41234_new_n4182_), .Y(_abc_41234_new_n4183_));
AOI22X1 AOI22X1_195 ( .A(rdatahold_4_), .B(_abc_41234_new_n3964_), .C(_abc_41234_new_n3963_), .D(_abc_41234_new_n3595_), .Y(_abc_41234_new_n4185_));
AOI22X1 AOI22X1_196 ( .A(_abc_41234_new_n3619_), .B(_abc_41234_new_n3963_), .C(_abc_41234_new_n3960_), .D(_abc_41234_new_n4198_), .Y(_abc_41234_new_n4206_));
AOI22X1 AOI22X1_197 ( .A(_abc_41234_new_n4299_), .B(_abc_41234_new_n515__bF_buf2), .C(_abc_41234_new_n1046__bF_buf7), .D(_abc_41234_new_n4315_), .Y(_abc_41234_new_n4316_));
AOI22X1 AOI22X1_198 ( .A(rdatahold2_0_), .B(_abc_41234_new_n4274__bF_buf2), .C(_abc_41234_new_n660__bF_buf1), .D(_abc_41234_new_n4317_), .Y(_abc_41234_new_n4318_));
AOI22X1 AOI22X1_199 ( .A(rdatahold2_1_), .B(_abc_41234_new_n4274__bF_buf1), .C(pc_1_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4336_));
AOI22X1 AOI22X1_2 ( .A(regfil_0__0_), .B(_abc_41234_new_n618_), .C(regfil_1__0_), .D(_abc_41234_new_n617_), .Y(_abc_41234_new_n619_));
AOI22X1 AOI22X1_20 ( .A(alu_res_5_), .B(_abc_41234_new_n613_), .C(rdatahold_5_), .D(_abc_41234_new_n650_), .Y(_abc_41234_new_n912_));
AOI22X1 AOI22X1_200 ( .A(rdatahold2_2_), .B(_abc_41234_new_n4274__bF_buf0), .C(pc_2_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4351_));
AOI22X1 AOI22X1_201 ( .A(_abc_41234_new_n2776_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n2773_), .D(_abc_41234_new_n4295_), .Y(_abc_41234_new_n4356_));
AOI22X1 AOI22X1_202 ( .A(rdatahold2_3_), .B(_abc_41234_new_n4274__bF_buf3), .C(pc_3_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4369_));
AOI22X1 AOI22X1_203 ( .A(_abc_41234_new_n2805_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n2801_), .D(_abc_41234_new_n4295_), .Y(_abc_41234_new_n4372_));
AOI22X1 AOI22X1_204 ( .A(rdatahold2_5_), .B(_abc_41234_new_n4274__bF_buf1), .C(pc_5_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4405_));
AOI22X1 AOI22X1_205 ( .A(_abc_41234_new_n2858_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n665__bF_buf2), .D(_abc_41234_new_n4410_), .Y(_abc_41234_new_n4411_));
AOI22X1 AOI22X1_206 ( .A(rdatahold2_6_), .B(_abc_41234_new_n4274__bF_buf0), .C(pc_6_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4424_));
AOI22X1 AOI22X1_207 ( .A(regfil_5__7_), .B(_abc_41234_new_n1303_), .C(_abc_41234_new_n4309_), .D(_abc_41234_new_n4430_), .Y(_abc_41234_new_n4431_));
AOI22X1 AOI22X1_208 ( .A(rdatahold2_7_), .B(_abc_41234_new_n4274__bF_buf3), .C(pc_7_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4443_));
AOI22X1 AOI22X1_209 ( .A(_abc_41234_new_n1624_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n4448_), .D(_abc_41234_new_n4295_), .Y(_abc_41234_new_n4449_));
AOI22X1 AOI22X1_21 ( .A(_abc_41234_new_n602_), .B(_abc_41234_new_n913_), .C(_abc_41234_new_n917_), .D(_abc_41234_new_n922_), .Y(_abc_41234_new_n923_));
AOI22X1 AOI22X1_210 ( .A(rdatahold_0_), .B(_abc_41234_new_n4274__bF_buf2), .C(pc_8_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4461_));
AOI22X1 AOI22X1_211 ( .A(_abc_41234_new_n1674_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n1680_), .D(_abc_41234_new_n4295_), .Y(_abc_41234_new_n4472_));
AOI22X1 AOI22X1_212 ( .A(rdatahold_1_), .B(_abc_41234_new_n4274__bF_buf1), .C(pc_9_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4478_));
AOI22X1 AOI22X1_213 ( .A(_abc_41234_new_n1716_), .B(_abc_41234_new_n4308_), .C(_abc_41234_new_n4301_), .D(_abc_41234_new_n4483_), .Y(_abc_41234_new_n4490_));
AOI22X1 AOI22X1_214 ( .A(rdatahold_2_), .B(_abc_41234_new_n4274__bF_buf0), .C(pc_10_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4497_));
AOI22X1 AOI22X1_215 ( .A(_abc_41234_new_n1728_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n1734_), .D(_abc_41234_new_n4295_), .Y(_abc_41234_new_n4503_));
AOI22X1 AOI22X1_216 ( .A(regfil_4__3_), .B(_abc_41234_new_n1303_), .C(pc_11_), .D(_abc_41234_new_n4312_), .Y(_abc_41234_new_n4510_));
AOI22X1 AOI22X1_217 ( .A(rdatahold_3_), .B(_abc_41234_new_n4274__bF_buf3), .C(pc_11_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4515_));
AOI22X1 AOI22X1_218 ( .A(_abc_41234_new_n1752_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n1756_), .D(_abc_41234_new_n4295_), .Y(_abc_41234_new_n4520_));
AOI22X1 AOI22X1_219 ( .A(rdatahold_4_), .B(_abc_41234_new_n4274__bF_buf2), .C(pc_12_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4535_));
AOI22X1 AOI22X1_22 ( .A(_abc_41234_new_n707_), .B(alu_res_5_), .C(\data[5] ), .D(_abc_41234_new_n758_), .Y(_abc_41234_new_n936_));
AOI22X1 AOI22X1_220 ( .A(_abc_41234_new_n1774_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n4295_), .D(_abc_41234_new_n1780_), .Y(_abc_41234_new_n4540_));
AOI22X1 AOI22X1_221 ( .A(regfil_4__5_), .B(_abc_41234_new_n1303_), .C(pc_13_), .D(_abc_41234_new_n4312_), .Y(_abc_41234_new_n4548_));
AOI22X1 AOI22X1_222 ( .A(rdatahold_5_), .B(_abc_41234_new_n4274__bF_buf1), .C(pc_13_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4553_));
AOI22X1 AOI22X1_223 ( .A(rdatahold_6_), .B(_abc_41234_new_n4274__bF_buf0), .C(pc_14_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4574_));
AOI22X1 AOI22X1_224 ( .A(regfil_4__7_), .B(_abc_41234_new_n1303_), .C(pc_15_), .D(_abc_41234_new_n4312_), .Y(_abc_41234_new_n4591_));
AOI22X1 AOI22X1_225 ( .A(rdatahold_7_), .B(_abc_41234_new_n4274__bF_buf3), .C(pc_15_), .D(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4597_));
AOI22X1 AOI22X1_226 ( .A(_abc_41234_new_n2358_), .B(pc_0_), .C(waddrhold_0_), .D(_abc_41234_new_n2696__bF_buf1), .Y(_abc_41234_new_n4616_));
AOI22X1 AOI22X1_227 ( .A(_abc_41234_new_n2358_), .B(pc_1_), .C(waddrhold_1_), .D(_abc_41234_new_n2696__bF_buf0), .Y(_abc_41234_new_n4621_));
AOI22X1 AOI22X1_228 ( .A(_abc_41234_new_n2358_), .B(pc_2_), .C(waddrhold_2_), .D(_abc_41234_new_n2696__bF_buf4), .Y(_abc_41234_new_n4626_));
AOI22X1 AOI22X1_229 ( .A(_abc_41234_new_n2358_), .B(pc_3_), .C(waddrhold_3_), .D(_abc_41234_new_n2696__bF_buf3), .Y(_abc_41234_new_n4631_));
AOI22X1 AOI22X1_23 ( .A(regfil_4__6_), .B(_abc_41234_new_n618_), .C(regfil_5__6_bF_buf3_), .D(_abc_41234_new_n617_), .Y(_abc_41234_new_n941_));
AOI22X1 AOI22X1_230 ( .A(_abc_41234_new_n2358_), .B(pc_4_), .C(waddrhold_4_), .D(_abc_41234_new_n2696__bF_buf2), .Y(_abc_41234_new_n4636_));
AOI22X1 AOI22X1_231 ( .A(_abc_41234_new_n2358_), .B(pc_5_), .C(waddrhold_5_), .D(_abc_41234_new_n2696__bF_buf1), .Y(_abc_41234_new_n4641_));
AOI22X1 AOI22X1_232 ( .A(_abc_41234_new_n2358_), .B(pc_6_), .C(waddrhold_6_), .D(_abc_41234_new_n2696__bF_buf0), .Y(_abc_41234_new_n4646_));
AOI22X1 AOI22X1_233 ( .A(_abc_41234_new_n2358_), .B(pc_7_), .C(waddrhold_7_), .D(_abc_41234_new_n2696__bF_buf4), .Y(_abc_41234_new_n4651_));
AOI22X1 AOI22X1_234 ( .A(_abc_41234_new_n660__bF_buf1), .B(_abc_41234_new_n4756_), .C(_abc_41234_new_n4735_), .D(_abc_41234_new_n2535_), .Y(_abc_41234_new_n4757_));
AOI22X1 AOI22X1_235 ( .A(_abc_41234_new_n4766_), .B(_abc_41234_new_n4729_), .C(_abc_41234_new_n4720_), .D(_abc_41234_new_n4768_), .Y(_abc_41234_new_n4769_));
AOI22X1 AOI22X1_236 ( .A(_abc_41234_new_n608_), .B(_abc_41234_new_n2427_), .C(_abc_41234_new_n4782_), .D(_abc_41234_new_n2634_), .Y(_abc_41234_new_n4783_));
AOI22X1 AOI22X1_237 ( .A(_abc_41234_new_n4793_), .B(_abc_41234_new_n4725_), .C(_abc_41234_new_n4720_), .D(_abc_41234_new_n4794_), .Y(_abc_41234_new_n4795_));
AOI22X1 AOI22X1_238 ( .A(_abc_41234_new_n2497_), .B(_abc_41234_new_n4736_), .C(_abc_41234_new_n664_), .D(_abc_41234_new_n2505_), .Y(_abc_41234_new_n4797_));
AOI22X1 AOI22X1_239 ( .A(_abc_41234_new_n4798_), .B(_abc_41234_new_n660__bF_buf0), .C(_abc_41234_new_n4796_), .D(_abc_41234_new_n2535_), .Y(_abc_41234_new_n4799_));
AOI22X1 AOI22X1_24 ( .A(regfil_7__6_), .B(_abc_41234_new_n545_), .C(regfil_6__6_), .D(_abc_41234_new_n621_), .Y(_abc_41234_new_n942_));
AOI22X1 AOI22X1_240 ( .A(_abc_41234_new_n4768_), .B(_abc_41234_new_n4803_), .C(_abc_41234_new_n4800_), .D(_abc_41234_new_n4760_), .Y(_abc_41234_new_n4804_));
AOI22X1 AOI22X1_241 ( .A(_abc_41234_new_n608_), .B(_abc_41234_new_n611_), .C(_abc_41234_new_n4782_), .D(_abc_41234_new_n682_), .Y(_abc_41234_new_n4807_));
AOI22X1 AOI22X1_242 ( .A(_abc_41234_new_n519_), .B(_abc_41234_new_n2518_), .C(_abc_41234_new_n4782_), .D(_abc_41234_new_n4600_), .Y(_abc_41234_new_n4813_));
AOI22X1 AOI22X1_243 ( .A(_abc_41234_new_n608_), .B(_abc_41234_new_n1033_), .C(_abc_41234_new_n4782_), .D(_abc_41234_new_n4831_), .Y(_abc_41234_new_n4832_));
AOI22X1 AOI22X1_244 ( .A(_abc_41234_new_n2429_), .B(_abc_41234_new_n4782_), .C(_abc_41234_new_n4780_), .D(_abc_41234_new_n4760_), .Y(_abc_41234_new_n4835_));
AOI22X1 AOI22X1_245 ( .A(_abc_41234_new_n507_), .B(_abc_41234_new_n2357_), .C(_abc_41234_new_n660__bF_buf7), .D(_abc_41234_new_n2951__bF_buf1), .Y(_abc_41234_new_n4841_));
AOI22X1 AOI22X1_246 ( .A(_abc_41234_new_n4860_), .B(_abc_41234_new_n4801_), .C(_abc_41234_new_n4715_), .D(_abc_41234_new_n4760_), .Y(_abc_41234_new_n4861_));
AOI22X1 AOI22X1_247 ( .A(alu__abc_40887_new_n38_), .B(alu__abc_40887_new_n40_), .C(alu__abc_40887_new_n141_), .D(alu__abc_40887_new_n135_), .Y(alu__abc_40887_new_n142_));
AOI22X1 AOI22X1_248 ( .A(alu_oprb_0_), .B(alu__abc_40887_new_n128_), .C(alu__abc_40887_new_n43_), .D(alu__abc_40887_new_n89_), .Y(alu__abc_40887_new_n149_));
AOI22X1 AOI22X1_249 ( .A(alu__abc_40887_new_n54_), .B(alu__abc_40887_new_n83_), .C(alu__abc_40887_new_n86_), .D(alu__abc_40887_new_n151_), .Y(alu__abc_40887_new_n152_));
AOI22X1 AOI22X1_25 ( .A(regfil_3__6_), .B(_abc_41234_new_n545_), .C(regfil_2__6_), .D(_abc_41234_new_n621_), .Y(_abc_41234_new_n946_));
AOI22X1 AOI22X1_250 ( .A(alu__abc_40887_new_n178_), .B(alu__abc_40887_new_n138_), .C(alu__abc_40887_new_n134_), .D(alu__abc_40887_new_n181_), .Y(alu__abc_40887_new_n182_));
AOI22X1 AOI22X1_251 ( .A(alu__abc_40887_new_n175_), .B(alu__abc_40887_new_n183_), .C(alu__abc_40887_new_n180_), .D(alu__abc_40887_new_n182_), .Y(alu__abc_40887_new_n184_));
AOI22X1 AOI22X1_252 ( .A(alu__abc_40887_new_n235_), .B(alu__abc_40887_new_n201_), .C(alu__abc_40887_new_n238_), .D(alu__abc_40887_new_n248_), .Y(alu__abc_40887_new_n249_));
AOI22X1 AOI22X1_253 ( .A(alu__abc_40887_new_n54_), .B(alu__abc_40887_new_n209_), .C(alu__abc_40887_new_n201_), .D(alu__abc_40887_new_n266_), .Y(alu__abc_40887_new_n267_));
AOI22X1 AOI22X1_26 ( .A(alu_res_6_), .B(_abc_41234_new_n613_), .C(rdatahold_6_), .D(_abc_41234_new_n650_), .Y(_abc_41234_new_n951_));
AOI22X1 AOI22X1_27 ( .A(_abc_41234_new_n602_), .B(_abc_41234_new_n952_), .C(_abc_41234_new_n957_), .D(_abc_41234_new_n961_), .Y(_abc_41234_new_n962_));
AOI22X1 AOI22X1_28 ( .A(_abc_41234_new_n707_), .B(alu_res_6_), .C(\data[6] ), .D(_abc_41234_new_n758_), .Y(_abc_41234_new_n979_));
AOI22X1 AOI22X1_29 ( .A(_abc_41234_new_n1004_), .B(_abc_41234_new_n1006_), .C(alu_res_7_), .D(_abc_41234_new_n613_), .Y(_abc_41234_new_n1007_));
AOI22X1 AOI22X1_3 ( .A(regfil_3__0_), .B(_abc_41234_new_n545_), .C(regfil_2__0_), .D(_abc_41234_new_n621_), .Y(_abc_41234_new_n622_));
AOI22X1 AOI22X1_30 ( .A(rdatahold_7_), .B(_abc_41234_new_n596_), .C(_abc_41234_new_n1008_), .D(_abc_41234_new_n602_), .Y(_abc_41234_new_n1009_));
AOI22X1 AOI22X1_31 ( .A(alu_res_7_), .B(_abc_41234_new_n707_), .C(rdatahold_7_), .D(_abc_41234_new_n513_), .Y(_abc_41234_new_n1017_));
AOI22X1 AOI22X1_32 ( .A(_abc_41234_new_n533_), .B(_abc_41234_new_n529_), .C(regfil_7__6_), .D(_abc_41234_new_n559_), .Y(_abc_41234_new_n1026_));
AOI22X1 AOI22X1_33 ( .A(rdatahold_0_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1055_), .D(_abc_41234_new_n1063_), .Y(_abc_41234_new_n1064_));
AOI22X1 AOI22X1_34 ( .A(_abc_41234_new_n1206_), .B(_abc_41234_new_n1232_), .C(_abc_41234_new_n1220_), .D(_abc_41234_new_n1216_), .Y(_abc_41234_new_n1233_));
AOI22X1 AOI22X1_35 ( .A(rdatahold_1_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1055_), .D(_abc_41234_new_n1237_), .Y(_abc_41234_new_n1238_));
AOI22X1 AOI22X1_36 ( .A(rdatahold_2_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1055_), .D(_abc_41234_new_n1288_), .Y(_abc_41234_new_n1289_));
AOI22X1 AOI22X1_37 ( .A(_abc_41234_new_n1108_), .B(_abc_41234_new_n1302_), .C(_abc_41234_new_n1338_), .D(_abc_41234_new_n1337_), .Y(_abc_41234_new_n1339_));
AOI22X1 AOI22X1_38 ( .A(_abc_41234_new_n1206_), .B(_abc_41234_new_n1295_), .C(_abc_41234_new_n1042_), .D(_abc_41234_new_n1339_), .Y(_abc_41234_new_n1340_));
AOI22X1 AOI22X1_39 ( .A(rdatahold_3_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1345_), .D(_abc_41234_new_n1343_), .Y(_abc_41234_new_n1346_));
AOI22X1 AOI22X1_4 ( .A(regfil_4__0_), .B(_abc_41234_new_n618_), .C(regfil_5__0_), .D(_abc_41234_new_n617_), .Y(_abc_41234_new_n624_));
AOI22X1 AOI22X1_40 ( .A(_abc_41234_new_n535_), .B(_abc_41234_new_n1369_), .C(_abc_41234_new_n1381_), .D(_abc_41234_new_n1373_), .Y(_abc_41234_new_n1382_));
AOI22X1 AOI22X1_41 ( .A(rdatahold_4_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1388_), .D(_abc_41234_new_n1387_), .Y(_abc_41234_new_n1389_));
AOI22X1 AOI22X1_42 ( .A(rdatahold_5_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1444_), .D(_abc_41234_new_n1445_), .Y(_abc_41234_new_n1446_));
AOI22X1 AOI22X1_43 ( .A(rdatahold_6_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1508_), .D(_abc_41234_new_n1510_), .Y(_abc_41234_new_n1511_));
AOI22X1 AOI22X1_44 ( .A(rdatahold_7_), .B(_abc_41234_new_n1037_), .C(_abc_41234_new_n1055_), .D(_abc_41234_new_n1560_), .Y(_abc_41234_new_n1561_));
AOI22X1 AOI22X1_45 ( .A(_abc_41234_new_n535_), .B(_abc_41234_new_n1039_), .C(_abc_41234_new_n1598_), .D(_abc_41234_new_n1600_), .Y(_abc_41234_new_n1601_));
AOI22X1 AOI22X1_46 ( .A(_abc_41234_new_n1039_), .B(_abc_41234_new_n1048_), .C(_abc_41234_new_n1565_), .D(_abc_41234_new_n1602_), .Y(_abc_41234_new_n1603_));
AOI22X1 AOI22X1_47 ( .A(_abc_41234_new_n1605_), .B(_abc_41234_new_n1644_), .C(_abc_41234_new_n1633_), .D(_abc_41234_new_n1662_), .Y(_abc_41234_new_n1663_));
AOI22X1 AOI22X1_48 ( .A(_abc_41234_new_n515__bF_buf2), .B(_abc_41234_new_n1612_), .C(_abc_41234_new_n1046__bF_buf5), .D(_abc_41234_new_n1663_), .Y(_abc_41234_new_n1664_));
AOI22X1 AOI22X1_49 ( .A(regfil_7__1_), .B(_abc_41234_new_n1684_), .C(_abc_41234_new_n536__bF_buf1), .D(_abc_41234_new_n1687_), .Y(_abc_41234_new_n1688_));
AOI22X1 AOI22X1_5 ( .A(regfil_7__0_), .B(_abc_41234_new_n545_), .C(regfil_6__0_), .D(_abc_41234_new_n621_), .Y(_abc_41234_new_n625_));
AOI22X1 AOI22X1_50 ( .A(_abc_41234_new_n1666_), .B(_abc_41234_new_n1644_), .C(_abc_41234_new_n1676_), .D(_abc_41234_new_n1693_), .Y(_abc_41234_new_n1694_));
AOI22X1 AOI22X1_51 ( .A(_abc_41234_new_n515__bF_buf1), .B(_abc_41234_new_n1668_), .C(_abc_41234_new_n1046__bF_buf4), .D(_abc_41234_new_n1694_), .Y(_abc_41234_new_n1695_));
AOI22X1 AOI22X1_52 ( .A(_abc_41234_new_n515__bF_buf0), .B(_abc_41234_new_n1699_), .C(_abc_41234_new_n1721_), .D(_abc_41234_new_n1720_), .Y(_abc_41234_new_n1722_));
AOI22X1 AOI22X1_53 ( .A(_abc_41234_new_n1639__bF_buf3), .B(_abc_41234_new_n1738_), .C(intcyc_bF_buf0), .D(_abc_41234_new_n1731_), .Y(_abc_41234_new_n1739_));
AOI22X1 AOI22X1_54 ( .A(_abc_41234_new_n515__bF_buf6), .B(_abc_41234_new_n1726_), .C(_abc_41234_new_n1742_), .D(_abc_41234_new_n1743_), .Y(_abc_41234_new_n1744_));
AOI22X1 AOI22X1_55 ( .A(_abc_41234_new_n1756_), .B(_abc_41234_new_n1637_), .C(_abc_41234_new_n1627_), .D(_abc_41234_new_n1752_), .Y(_abc_41234_new_n1757_));
AOI22X1 AOI22X1_56 ( .A(_abc_41234_new_n515__bF_buf5), .B(_abc_41234_new_n1748_), .C(_abc_41234_new_n1768_), .D(_abc_41234_new_n1767_), .Y(_abc_41234_new_n1769_));
AOI22X1 AOI22X1_57 ( .A(_abc_41234_new_n515__bF_buf4), .B(_abc_41234_new_n1773_), .C(_abc_41234_new_n1790_), .D(_abc_41234_new_n1789_), .Y(_abc_41234_new_n1791_));
AOI22X1 AOI22X1_58 ( .A(_abc_41234_new_n1800_), .B(_abc_41234_new_n1627_), .C(_abc_41234_new_n1637_), .D(_abc_41234_new_n1805_), .Y(_abc_41234_new_n1806_));
AOI22X1 AOI22X1_59 ( .A(_abc_41234_new_n515__bF_buf3), .B(_abc_41234_new_n1795_), .C(_abc_41234_new_n1818_), .D(_abc_41234_new_n1817_), .Y(_abc_41234_new_n1819_));
AOI22X1 AOI22X1_6 ( .A(_abc_41234_new_n631_), .B(_abc_41234_new_n644_), .C(rdatahold_0_), .D(_abc_41234_new_n633_), .Y(_abc_41234_new_n645_));
AOI22X1 AOI22X1_60 ( .A(_abc_41234_new_n515__bF_buf2), .B(_abc_41234_new_n1823_), .C(_abc_41234_new_n1843_), .D(_abc_41234_new_n1842_), .Y(_abc_41234_new_n1844_));
AOI22X1 AOI22X1_61 ( .A(rdatahold2_1_), .B(_abc_41234_new_n1855_), .C(_abc_41234_new_n1881_), .D(_abc_41234_new_n1877_), .Y(_abc_41234_new_n1882_));
AOI22X1 AOI22X1_62 ( .A(_abc_41234_new_n593_), .B(_abc_41234_new_n594_), .C(_abc_41234_new_n1977_), .D(_abc_41234_new_n600_), .Y(_abc_41234_new_n1978_));
AOI22X1 AOI22X1_63 ( .A(_abc_41234_new_n583_), .B(_abc_41234_new_n1987_), .C(_abc_41234_new_n631_), .D(_abc_41234_new_n1985_), .Y(_abc_41234_new_n1988_));
AOI22X1 AOI22X1_64 ( .A(_abc_41234_new_n583_), .B(_abc_41234_new_n1997_), .C(_abc_41234_new_n1994_), .D(_abc_41234_new_n631_), .Y(_abc_41234_new_n1998_));
AOI22X1 AOI22X1_65 ( .A(rdatahold_3_), .B(_abc_41234_new_n1855_), .C(_abc_41234_new_n2103_), .D(_abc_41234_new_n2102_), .Y(_abc_41234_new_n2104_));
AOI22X1 AOI22X1_66 ( .A(rdatahold_4_), .B(_abc_41234_new_n1855_), .C(_abc_41234_new_n2115_), .D(_abc_41234_new_n2114_), .Y(_abc_41234_new_n2116_));
AOI22X1 AOI22X1_67 ( .A(rdatahold_5_), .B(_abc_41234_new_n1855_), .C(_abc_41234_new_n2127_), .D(_abc_41234_new_n2126_), .Y(_abc_41234_new_n2128_));
AOI22X1 AOI22X1_68 ( .A(opcode_5_bF_buf0_), .B(_abc_41234_new_n2189__bF_buf4), .C(_abc_41234_new_n1046__bF_buf1), .D(_abc_41234_new_n2197_), .Y(_abc_41234_new_n2198_));
AOI22X1 AOI22X1_69 ( .A(_abc_41234_new_n516__bF_buf4), .B(_abc_41234_new_n2217_), .C(alu_oprb_0_), .D(_abc_41234_new_n2216_), .Y(_abc_41234_new_n2218_));
AOI22X1 AOI22X1_7 ( .A(alu_res_1_), .B(_abc_41234_new_n613_), .C(rdatahold_1_), .D(_abc_41234_new_n650_), .Y(_abc_41234_new_n736_));
AOI22X1 AOI22X1_70 ( .A(_abc_41234_new_n734_), .B(_abc_41234_new_n2224_), .C(rdatahold_1_), .D(_abc_41234_new_n2223_), .Y(_abc_41234_new_n2225_));
AOI22X1 AOI22X1_71 ( .A(_abc_41234_new_n778_), .B(_abc_41234_new_n2224_), .C(rdatahold_2_), .D(_abc_41234_new_n2223_), .Y(_abc_41234_new_n2228_));
AOI22X1 AOI22X1_72 ( .A(alu_oprb_3_), .B(_abc_41234_new_n2221_), .C(_abc_41234_new_n2189__bF_buf1), .D(_abc_41234_new_n825_), .Y(_abc_41234_new_n2230_));
AOI22X1 AOI22X1_73 ( .A(rdatahold_3_), .B(_abc_41234_new_n2223_), .C(alu_oprb_3_), .D(_abc_41234_new_n2216_), .Y(_abc_41234_new_n2231_));
AOI22X1 AOI22X1_74 ( .A(_abc_41234_new_n862_), .B(_abc_41234_new_n2224_), .C(rdatahold_4_), .D(_abc_41234_new_n2223_), .Y(_abc_41234_new_n2234_));
AOI22X1 AOI22X1_75 ( .A(_abc_41234_new_n910_), .B(_abc_41234_new_n2224_), .C(rdatahold_5_), .D(_abc_41234_new_n2223_), .Y(_abc_41234_new_n2237_));
AOI22X1 AOI22X1_76 ( .A(alu_oprb_6_), .B(_abc_41234_new_n2221_), .C(_abc_41234_new_n2189__bF_buf0), .D(_abc_41234_new_n949_), .Y(_abc_41234_new_n2239_));
AOI22X1 AOI22X1_77 ( .A(rdatahold_6_), .B(_abc_41234_new_n2223_), .C(alu_oprb_6_), .D(_abc_41234_new_n2216_), .Y(_abc_41234_new_n2240_));
AOI22X1 AOI22X1_78 ( .A(_abc_41234_new_n1002_), .B(_abc_41234_new_n2224_), .C(_abc_41234_new_n1006_), .D(_abc_41234_new_n2215_), .Y(_abc_41234_new_n2243_));
AOI22X1 AOI22X1_79 ( .A(regfil_4__0_), .B(_abc_41234_new_n2247_), .C(regfil_5__0_), .D(_abc_41234_new_n2248_), .Y(_abc_41234_new_n2249_));
AOI22X1 AOI22X1_8 ( .A(_abc_41234_new_n602_), .B(_abc_41234_new_n737_), .C(_abc_41234_new_n742_), .D(_abc_41234_new_n746_), .Y(_abc_41234_new_n747_));
AOI22X1 AOI22X1_80 ( .A(regfil_0__0_), .B(_abc_41234_new_n2247_), .C(regfil_2__0_), .D(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2256_));
AOI22X1 AOI22X1_81 ( .A(regfil_7__0_), .B(_abc_41234_new_n2201_), .C(_abc_41234_new_n2252_), .D(_abc_41234_new_n2259_), .Y(_abc_41234_new_n2260_));
AOI22X1 AOI22X1_82 ( .A(rdatahold_0_), .B(_abc_41234_new_n2263_), .C(alu_opra_0_), .D(_abc_41234_new_n2266_), .Y(_abc_41234_new_n2267_));
AOI22X1 AOI22X1_83 ( .A(regfil_4__1_bF_buf3_), .B(_abc_41234_new_n2247_), .C(regfil_5__1_), .D(_abc_41234_new_n2248_), .Y(_abc_41234_new_n2270_));
AOI22X1 AOI22X1_84 ( .A(regfil_0__1_), .B(_abc_41234_new_n2247_), .C(regfil_2__1_), .D(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2274_));
AOI22X1 AOI22X1_85 ( .A(regfil_7__1_), .B(_abc_41234_new_n2201_), .C(_abc_41234_new_n2272_), .D(_abc_41234_new_n2277_), .Y(_abc_41234_new_n2278_));
AOI22X1 AOI22X1_86 ( .A(rdatahold_1_), .B(_abc_41234_new_n2263_), .C(alu_opra_1_), .D(_abc_41234_new_n2266_), .Y(_abc_41234_new_n2279_));
AOI22X1 AOI22X1_87 ( .A(regfil_4__2_bF_buf3_), .B(_abc_41234_new_n2247_), .C(regfil_5__2_), .D(_abc_41234_new_n2248_), .Y(_abc_41234_new_n2282_));
AOI22X1 AOI22X1_88 ( .A(regfil_0__2_), .B(_abc_41234_new_n2247_), .C(regfil_2__2_), .D(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2286_));
AOI22X1 AOI22X1_89 ( .A(regfil_7__2_), .B(_abc_41234_new_n2201_), .C(_abc_41234_new_n2284_), .D(_abc_41234_new_n2289_), .Y(_abc_41234_new_n2290_));
AOI22X1 AOI22X1_9 ( .A(regfil_7__0_), .B(_abc_41234_new_n559_), .C(_abc_41234_new_n514_), .D(_abc_41234_new_n752_), .Y(_abc_41234_new_n753_));
AOI22X1 AOI22X1_90 ( .A(rdatahold_2_), .B(_abc_41234_new_n2263_), .C(alu_opra_2_), .D(_abc_41234_new_n2266_), .Y(_abc_41234_new_n2291_));
AOI22X1 AOI22X1_91 ( .A(regfil_4__3_), .B(_abc_41234_new_n2247_), .C(regfil_5__3_bF_buf1_), .D(_abc_41234_new_n2248_), .Y(_abc_41234_new_n2294_));
AOI22X1 AOI22X1_92 ( .A(regfil_0__3_), .B(_abc_41234_new_n2247_), .C(regfil_2__3_), .D(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2298_));
AOI22X1 AOI22X1_93 ( .A(regfil_7__3_), .B(_abc_41234_new_n2201_), .C(_abc_41234_new_n2296_), .D(_abc_41234_new_n2301_), .Y(_abc_41234_new_n2302_));
AOI22X1 AOI22X1_94 ( .A(rdatahold_3_), .B(_abc_41234_new_n2263_), .C(alu_opra_3_), .D(_abc_41234_new_n2266_), .Y(_abc_41234_new_n2303_));
AOI22X1 AOI22X1_95 ( .A(regfil_4__4_), .B(_abc_41234_new_n2247_), .C(regfil_5__4_), .D(_abc_41234_new_n2248_), .Y(_abc_41234_new_n2306_));
AOI22X1 AOI22X1_96 ( .A(regfil_0__4_), .B(_abc_41234_new_n2247_), .C(regfil_2__4_), .D(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2310_));
AOI22X1 AOI22X1_97 ( .A(regfil_7__4_), .B(_abc_41234_new_n2201_), .C(_abc_41234_new_n2308_), .D(_abc_41234_new_n2313_), .Y(_abc_41234_new_n2314_));
AOI22X1 AOI22X1_98 ( .A(rdatahold_4_), .B(_abc_41234_new_n2263_), .C(alu_opra_4_), .D(_abc_41234_new_n2266_), .Y(_abc_41234_new_n2315_));
AOI22X1 AOI22X1_99 ( .A(regfil_0__5_), .B(_abc_41234_new_n2247_), .C(regfil_2__5_), .D(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2318_));
BUFX2 BUFX2_1 ( .A(regfil_4__1_), .Y(regfil_4__1_bF_buf2_));
BUFX2 BUFX2_10 ( .A(_abc_41234_new_n525_), .Y(_abc_41234_new_n525__bF_buf2));
BUFX2 BUFX2_11 ( .A(_abc_41234_new_n525_), .Y(_abc_41234_new_n525__bF_buf1));
BUFX2 BUFX2_12 ( .A(_abc_41234_new_n525_), .Y(_abc_41234_new_n525__bF_buf0));
BUFX2 BUFX2_13 ( .A(sp_0_), .Y(sp_0_bF_buf0_));
BUFX2 BUFX2_14 ( .A(regfil_4__2_), .Y(regfil_4__2_bF_buf2_));
BUFX2 BUFX2_15 ( .A(regfil_4__2_), .Y(regfil_4__2_bF_buf1_));
BUFX2 BUFX2_16 ( .A(regfil_4__2_), .Y(regfil_4__2_bF_buf0_));
BUFX2 BUFX2_17 ( .A(_abc_41234_new_n2919_), .Y(_abc_41234_new_n2919__bF_buf2));
BUFX2 BUFX2_18 ( .A(_abc_41234_new_n2919_), .Y(_abc_41234_new_n2919__bF_buf1));
BUFX2 BUFX2_19 ( .A(_abc_41234_new_n2919_), .Y(_abc_41234_new_n2919__bF_buf0));
BUFX2 BUFX2_2 ( .A(regfil_4__1_), .Y(regfil_4__1_bF_buf1_));
BUFX2 BUFX2_20 ( .A(_abc_41234_new_n2190_), .Y(_abc_41234_new_n2190__bF_buf1));
BUFX2 BUFX2_21 ( .A(_abc_41234_new_n2190_), .Y(_abc_41234_new_n2190__bF_buf0));
BUFX2 BUFX2_22 ( .A(_abc_41234_new_n665_), .Y(_abc_41234_new_n665__bF_buf2));
BUFX2 BUFX2_23 ( .A(_abc_41234_new_n665_), .Y(_abc_41234_new_n665__bF_buf0));
BUFX2 BUFX2_24 ( .A(_abc_41234_new_n4274_), .Y(_abc_41234_new_n4274__bF_buf2));
BUFX2 BUFX2_25 ( .A(_auto_iopadmap_cc_368_execute_45628_0_), .Y(\addr[0] ));
BUFX2 BUFX2_26 ( .A(_auto_iopadmap_cc_368_execute_45628_1_), .Y(\addr[1] ));
BUFX2 BUFX2_27 ( .A(_auto_iopadmap_cc_368_execute_45628_2_), .Y(\addr[2] ));
BUFX2 BUFX2_28 ( .A(_auto_iopadmap_cc_368_execute_45628_3_), .Y(\addr[3] ));
BUFX2 BUFX2_29 ( .A(_auto_iopadmap_cc_368_execute_45628_4_), .Y(\addr[4] ));
BUFX2 BUFX2_3 ( .A(regfil_4__1_), .Y(regfil_4__1_bF_buf0_));
BUFX2 BUFX2_30 ( .A(_auto_iopadmap_cc_368_execute_45628_5_), .Y(\addr[5] ));
BUFX2 BUFX2_31 ( .A(_auto_iopadmap_cc_368_execute_45628_6_), .Y(\addr[6] ));
BUFX2 BUFX2_32 ( .A(_auto_iopadmap_cc_368_execute_45628_7_), .Y(\addr[7] ));
BUFX2 BUFX2_33 ( .A(_auto_iopadmap_cc_368_execute_45628_8_), .Y(\addr[8] ));
BUFX2 BUFX2_34 ( .A(_auto_iopadmap_cc_368_execute_45628_9_), .Y(\addr[9] ));
BUFX2 BUFX2_35 ( .A(_auto_iopadmap_cc_368_execute_45628_10_), .Y(\addr[10] ));
BUFX2 BUFX2_36 ( .A(_auto_iopadmap_cc_368_execute_45628_11_), .Y(\addr[11] ));
BUFX2 BUFX2_37 ( .A(_auto_iopadmap_cc_368_execute_45628_12_), .Y(\addr[12] ));
BUFX2 BUFX2_38 ( .A(_auto_iopadmap_cc_368_execute_45628_13_), .Y(\addr[13] ));
BUFX2 BUFX2_39 ( .A(_auto_iopadmap_cc_368_execute_45628_14_), .Y(\addr[14] ));
BUFX2 BUFX2_4 ( .A(regfil_5__6_), .Y(regfil_5__6_bF_buf0_));
BUFX2 BUFX2_40 ( .A(_auto_iopadmap_cc_368_execute_45628_15_), .Y(\addr[15] ));
BUFX2 BUFX2_41 ( .A(_auto_iopadmap_cc_368_execute_45645), .Y(inta));
BUFX2 BUFX2_42 ( .A(_auto_iopadmap_cc_368_execute_45647), .Y(readio));
BUFX2 BUFX2_43 ( .A(_auto_iopadmap_cc_368_execute_45649), .Y(readmem));
BUFX2 BUFX2_44 ( .A(_auto_iopadmap_cc_368_execute_45651), .Y(writeio));
BUFX2 BUFX2_45 ( .A(_auto_iopadmap_cc_368_execute_45653), .Y(writemem));
BUFX2 BUFX2_5 ( .A(regfil_5__3_), .Y(regfil_5__3_bF_buf1_));
BUFX2 BUFX2_6 ( .A(regfil_5__3_), .Y(regfil_5__3_bF_buf0_));
BUFX2 BUFX2_7 ( .A(_abc_41234_new_n1639_), .Y(_abc_41234_new_n1639__bF_buf1));
BUFX2 BUFX2_8 ( .A(opcode_3_), .Y(opcode_3_bF_buf2_));
BUFX2 BUFX2_9 ( .A(opcode_3_), .Y(opcode_3_bF_buf0_));
BUFX4 BUFX4_1 ( .A(clock_bF_buf13), .Y(clock_bF_buf13_bF_buf3));
BUFX4 BUFX4_10 ( .A(_abc_41234_new_n544_), .Y(_abc_41234_new_n544__bF_buf2));
BUFX4 BUFX4_100 ( .A(_abc_41234_new_n1066_), .Y(_abc_41234_new_n1066__bF_buf2));
BUFX4 BUFX4_101 ( .A(_abc_41234_new_n1066_), .Y(_abc_41234_new_n1066__bF_buf1));
BUFX4 BUFX4_102 ( .A(_abc_41234_new_n1066_), .Y(_abc_41234_new_n1066__bF_buf0));
BUFX4 BUFX4_103 ( .A(_abc_41234_new_n3914_), .Y(_abc_41234_new_n3914__bF_buf3));
BUFX4 BUFX4_104 ( .A(_abc_41234_new_n3914_), .Y(_abc_41234_new_n3914__bF_buf2));
BUFX4 BUFX4_105 ( .A(_abc_41234_new_n3914_), .Y(_abc_41234_new_n3914__bF_buf1));
BUFX4 BUFX4_106 ( .A(_abc_41234_new_n3914_), .Y(_abc_41234_new_n3914__bF_buf0));
BUFX4 BUFX4_107 ( .A(_abc_41234_new_n2415_), .Y(_abc_41234_new_n2415__bF_buf4));
BUFX4 BUFX4_108 ( .A(_abc_41234_new_n2415_), .Y(_abc_41234_new_n2415__bF_buf3));
BUFX4 BUFX4_109 ( .A(_abc_41234_new_n2415_), .Y(_abc_41234_new_n2415__bF_buf2));
BUFX4 BUFX4_11 ( .A(_abc_41234_new_n544_), .Y(_abc_41234_new_n544__bF_buf1));
BUFX4 BUFX4_110 ( .A(_abc_41234_new_n2415_), .Y(_abc_41234_new_n2415__bF_buf1));
BUFX4 BUFX4_111 ( .A(_abc_41234_new_n2415_), .Y(_abc_41234_new_n2415__bF_buf0));
BUFX4 BUFX4_112 ( .A(_abc_41234_new_n546_), .Y(_abc_41234_new_n546__bF_buf5));
BUFX4 BUFX4_113 ( .A(_abc_41234_new_n546_), .Y(_abc_41234_new_n546__bF_buf4));
BUFX4 BUFX4_114 ( .A(_abc_41234_new_n546_), .Y(_abc_41234_new_n546__bF_buf3));
BUFX4 BUFX4_115 ( .A(_abc_41234_new_n546_), .Y(_abc_41234_new_n546__bF_buf2));
BUFX4 BUFX4_116 ( .A(_abc_41234_new_n546_), .Y(_abc_41234_new_n546__bF_buf1));
BUFX4 BUFX4_117 ( .A(_abc_41234_new_n546_), .Y(_abc_41234_new_n546__bF_buf0));
BUFX4 BUFX4_118 ( .A(_abc_41234_new_n537_), .Y(_abc_41234_new_n537__bF_buf3));
BUFX4 BUFX4_119 ( .A(_abc_41234_new_n537_), .Y(_abc_41234_new_n537__bF_buf2));
BUFX4 BUFX4_12 ( .A(_abc_41234_new_n544_), .Y(_abc_41234_new_n544__bF_buf0));
BUFX4 BUFX4_120 ( .A(_abc_41234_new_n537_), .Y(_abc_41234_new_n537__bF_buf1));
BUFX4 BUFX4_121 ( .A(_abc_41234_new_n537_), .Y(_abc_41234_new_n537__bF_buf0));
BUFX4 BUFX4_122 ( .A(_abc_41234_new_n669_), .Y(_abc_41234_new_n669__bF_buf3));
BUFX4 BUFX4_123 ( .A(_abc_41234_new_n669_), .Y(_abc_41234_new_n669__bF_buf2));
BUFX4 BUFX4_124 ( .A(_abc_41234_new_n669_), .Y(_abc_41234_new_n669__bF_buf1));
BUFX4 BUFX4_125 ( .A(_abc_41234_new_n669_), .Y(_abc_41234_new_n669__bF_buf0));
BUFX4 BUFX4_126 ( .A(opcode_3_), .Y(opcode_3_bF_buf3_));
BUFX4 BUFX4_127 ( .A(opcode_3_), .Y(opcode_3_bF_buf1_));
BUFX4 BUFX4_128 ( .A(_abc_41234_new_n534_), .Y(_abc_41234_new_n534__bF_buf5));
BUFX4 BUFX4_129 ( .A(_abc_41234_new_n534_), .Y(_abc_41234_new_n534__bF_buf4));
BUFX4 BUFX4_13 ( .A(_abc_41234_new_n1049_), .Y(_abc_41234_new_n1049__bF_buf4));
BUFX4 BUFX4_130 ( .A(_abc_41234_new_n534_), .Y(_abc_41234_new_n534__bF_buf3));
BUFX4 BUFX4_131 ( .A(_abc_41234_new_n534_), .Y(_abc_41234_new_n534__bF_buf2));
BUFX4 BUFX4_132 ( .A(_abc_41234_new_n534_), .Y(_abc_41234_new_n534__bF_buf1));
BUFX4 BUFX4_133 ( .A(_abc_41234_new_n534_), .Y(_abc_41234_new_n534__bF_buf0));
BUFX4 BUFX4_134 ( .A(_abc_41234_new_n722_), .Y(_abc_41234_new_n722__bF_buf3));
BUFX4 BUFX4_135 ( .A(_abc_41234_new_n722_), .Y(_abc_41234_new_n722__bF_buf2));
BUFX4 BUFX4_136 ( .A(_abc_41234_new_n722_), .Y(_abc_41234_new_n722__bF_buf1));
BUFX4 BUFX4_137 ( .A(_abc_41234_new_n722_), .Y(_abc_41234_new_n722__bF_buf0));
BUFX4 BUFX4_138 ( .A(_abc_41234_new_n2185_), .Y(_abc_41234_new_n2185__bF_buf5));
BUFX4 BUFX4_139 ( .A(_abc_41234_new_n2185_), .Y(_abc_41234_new_n2185__bF_buf4));
BUFX4 BUFX4_14 ( .A(_abc_41234_new_n1049_), .Y(_abc_41234_new_n1049__bF_buf3));
BUFX4 BUFX4_140 ( .A(_abc_41234_new_n2185_), .Y(_abc_41234_new_n2185__bF_buf3));
BUFX4 BUFX4_141 ( .A(_abc_41234_new_n2185_), .Y(_abc_41234_new_n2185__bF_buf2));
BUFX4 BUFX4_142 ( .A(_abc_41234_new_n2185_), .Y(_abc_41234_new_n2185__bF_buf1));
BUFX4 BUFX4_143 ( .A(_abc_41234_new_n2185_), .Y(_abc_41234_new_n2185__bF_buf0));
BUFX4 BUFX4_144 ( .A(intcyc), .Y(intcyc_bF_buf3));
BUFX4 BUFX4_145 ( .A(intcyc), .Y(intcyc_bF_buf2));
BUFX4 BUFX4_146 ( .A(intcyc), .Y(intcyc_bF_buf1));
BUFX4 BUFX4_147 ( .A(intcyc), .Y(intcyc_bF_buf0));
BUFX4 BUFX4_148 ( .A(_abc_41234_new_n660_), .Y(_abc_41234_new_n660__bF_buf7));
BUFX4 BUFX4_149 ( .A(_abc_41234_new_n660_), .Y(_abc_41234_new_n660__bF_buf6));
BUFX4 BUFX4_15 ( .A(_abc_41234_new_n1049_), .Y(_abc_41234_new_n1049__bF_buf2));
BUFX4 BUFX4_150 ( .A(_abc_41234_new_n660_), .Y(_abc_41234_new_n660__bF_buf5));
BUFX4 BUFX4_151 ( .A(_abc_41234_new_n660_), .Y(_abc_41234_new_n660__bF_buf4));
BUFX4 BUFX4_152 ( .A(_abc_41234_new_n660_), .Y(_abc_41234_new_n660__bF_buf3));
BUFX4 BUFX4_153 ( .A(_abc_41234_new_n660_), .Y(_abc_41234_new_n660__bF_buf2));
BUFX4 BUFX4_154 ( .A(_abc_41234_new_n660_), .Y(_abc_41234_new_n660__bF_buf1));
BUFX4 BUFX4_155 ( .A(_abc_41234_new_n660_), .Y(_abc_41234_new_n660__bF_buf0));
BUFX4 BUFX4_156 ( .A(_abc_41234_new_n525_), .Y(_abc_41234_new_n525__bF_buf3));
BUFX4 BUFX4_157 ( .A(_abc_41234_new_n2696_), .Y(_abc_41234_new_n2696__bF_buf4));
BUFX4 BUFX4_158 ( .A(_abc_41234_new_n2696_), .Y(_abc_41234_new_n2696__bF_buf3));
BUFX4 BUFX4_159 ( .A(_abc_41234_new_n2696_), .Y(_abc_41234_new_n2696__bF_buf2));
BUFX4 BUFX4_16 ( .A(_abc_41234_new_n1049_), .Y(_abc_41234_new_n1049__bF_buf1));
BUFX4 BUFX4_160 ( .A(_abc_41234_new_n2696_), .Y(_abc_41234_new_n2696__bF_buf1));
BUFX4 BUFX4_161 ( .A(_abc_41234_new_n2696_), .Y(_abc_41234_new_n2696__bF_buf0));
BUFX4 BUFX4_162 ( .A(_abc_41234_new_n516_), .Y(_abc_41234_new_n516__bF_buf5));
BUFX4 BUFX4_163 ( .A(_abc_41234_new_n516_), .Y(_abc_41234_new_n516__bF_buf4));
BUFX4 BUFX4_164 ( .A(_abc_41234_new_n516_), .Y(_abc_41234_new_n516__bF_buf3));
BUFX4 BUFX4_165 ( .A(_abc_41234_new_n516_), .Y(_abc_41234_new_n516__bF_buf2));
BUFX4 BUFX4_166 ( .A(_abc_41234_new_n516_), .Y(_abc_41234_new_n516__bF_buf1));
BUFX4 BUFX4_167 ( .A(_abc_41234_new_n516_), .Y(_abc_41234_new_n516__bF_buf0));
BUFX4 BUFX4_168 ( .A(sp_0_), .Y(sp_0_bF_buf3_));
BUFX4 BUFX4_169 ( .A(sp_0_), .Y(sp_0_bF_buf2_));
BUFX4 BUFX4_17 ( .A(_abc_41234_new_n1049_), .Y(_abc_41234_new_n1049__bF_buf0));
BUFX4 BUFX4_170 ( .A(sp_0_), .Y(sp_0_bF_buf1_));
BUFX4 BUFX4_171 ( .A(_abc_41234_new_n1047_), .Y(_abc_41234_new_n1047__bF_buf4));
BUFX4 BUFX4_172 ( .A(_abc_41234_new_n1047_), .Y(_abc_41234_new_n1047__bF_buf3));
BUFX4 BUFX4_173 ( .A(_abc_41234_new_n1047_), .Y(_abc_41234_new_n1047__bF_buf2));
BUFX4 BUFX4_174 ( .A(_abc_41234_new_n1047_), .Y(_abc_41234_new_n1047__bF_buf1));
BUFX4 BUFX4_175 ( .A(_abc_41234_new_n1047_), .Y(_abc_41234_new_n1047__bF_buf0));
BUFX4 BUFX4_176 ( .A(regfil_4__2_), .Y(regfil_4__2_bF_buf3_));
BUFX4 BUFX4_177 ( .A(opcode_5_), .Y(opcode_5_bF_buf4_));
BUFX4 BUFX4_178 ( .A(opcode_5_), .Y(opcode_5_bF_buf3_));
BUFX4 BUFX4_179 ( .A(opcode_5_), .Y(opcode_5_bF_buf2_));
BUFX4 BUFX4_18 ( .A(clock), .Y(clock_bF_buf14));
BUFX4 BUFX4_180 ( .A(opcode_5_), .Y(opcode_5_bF_buf1_));
BUFX4 BUFX4_181 ( .A(opcode_5_), .Y(opcode_5_bF_buf0_));
BUFX4 BUFX4_182 ( .A(_abc_41234_new_n2919_), .Y(_abc_41234_new_n2919__bF_buf3));
BUFX4 BUFX4_183 ( .A(_abc_41234_new_n536_), .Y(_abc_41234_new_n536__bF_buf5));
BUFX4 BUFX4_184 ( .A(_abc_41234_new_n536_), .Y(_abc_41234_new_n536__bF_buf4));
BUFX4 BUFX4_185 ( .A(_abc_41234_new_n536_), .Y(_abc_41234_new_n536__bF_buf3));
BUFX4 BUFX4_186 ( .A(_abc_41234_new_n536_), .Y(_abc_41234_new_n536__bF_buf2));
BUFX4 BUFX4_187 ( .A(_abc_41234_new_n536_), .Y(_abc_41234_new_n536__bF_buf1));
BUFX4 BUFX4_188 ( .A(_abc_41234_new_n536_), .Y(_abc_41234_new_n536__bF_buf0));
BUFX4 BUFX4_189 ( .A(_abc_41234_new_n668_), .Y(_abc_41234_new_n668__bF_buf5));
BUFX4 BUFX4_19 ( .A(clock), .Y(clock_bF_buf13));
BUFX4 BUFX4_190 ( .A(_abc_41234_new_n668_), .Y(_abc_41234_new_n668__bF_buf4));
BUFX4 BUFX4_191 ( .A(_abc_41234_new_n668_), .Y(_abc_41234_new_n668__bF_buf3));
BUFX4 BUFX4_192 ( .A(_abc_41234_new_n668_), .Y(_abc_41234_new_n668__bF_buf2));
BUFX4 BUFX4_193 ( .A(_abc_41234_new_n668_), .Y(_abc_41234_new_n668__bF_buf1));
BUFX4 BUFX4_194 ( .A(_abc_41234_new_n668_), .Y(_abc_41234_new_n668__bF_buf0));
BUFX4 BUFX4_195 ( .A(_abc_41234_new_n2190_), .Y(_abc_41234_new_n2190__bF_buf3));
BUFX4 BUFX4_196 ( .A(_abc_41234_new_n2190_), .Y(_abc_41234_new_n2190__bF_buf2));
BUFX4 BUFX4_197 ( .A(_abc_41234_new_n665_), .Y(_abc_41234_new_n665__bF_buf3));
BUFX4 BUFX4_198 ( .A(_abc_41234_new_n665_), .Y(_abc_41234_new_n665__bF_buf1));
BUFX4 BUFX4_199 ( .A(_abc_41234_new_n2951_), .Y(_abc_41234_new_n2951__bF_buf3));
BUFX4 BUFX4_2 ( .A(clock_bF_buf13), .Y(clock_bF_buf13_bF_buf2));
BUFX4 BUFX4_20 ( .A(clock), .Y(clock_bF_buf12));
BUFX4 BUFX4_200 ( .A(_abc_41234_new_n2951_), .Y(_abc_41234_new_n2951__bF_buf2));
BUFX4 BUFX4_201 ( .A(_abc_41234_new_n2951_), .Y(_abc_41234_new_n2951__bF_buf1));
BUFX4 BUFX4_202 ( .A(_abc_41234_new_n2951_), .Y(_abc_41234_new_n2951__bF_buf0));
BUFX4 BUFX4_203 ( .A(_abc_41234_new_n4274_), .Y(_abc_41234_new_n4274__bF_buf3));
BUFX4 BUFX4_204 ( .A(_abc_41234_new_n4274_), .Y(_abc_41234_new_n4274__bF_buf1));
BUFX4 BUFX4_205 ( .A(_abc_41234_new_n4274_), .Y(_abc_41234_new_n4274__bF_buf0));
BUFX4 BUFX4_206 ( .A(_abc_41234_new_n1643_), .Y(_abc_41234_new_n1643__bF_buf5));
BUFX4 BUFX4_207 ( .A(_abc_41234_new_n1643_), .Y(_abc_41234_new_n1643__bF_buf4));
BUFX4 BUFX4_208 ( .A(_abc_41234_new_n1643_), .Y(_abc_41234_new_n1643__bF_buf3));
BUFX4 BUFX4_209 ( .A(_abc_41234_new_n1643_), .Y(_abc_41234_new_n1643__bF_buf2));
BUFX4 BUFX4_21 ( .A(clock), .Y(clock_bF_buf11));
BUFX4 BUFX4_210 ( .A(_abc_41234_new_n1643_), .Y(_abc_41234_new_n1643__bF_buf1));
BUFX4 BUFX4_211 ( .A(_abc_41234_new_n1643_), .Y(_abc_41234_new_n1643__bF_buf0));
BUFX4 BUFX4_212 ( .A(_abc_41234_new_n2942_), .Y(_abc_41234_new_n2942__bF_buf3));
BUFX4 BUFX4_213 ( .A(_abc_41234_new_n2942_), .Y(_abc_41234_new_n2942__bF_buf2));
BUFX4 BUFX4_214 ( .A(_abc_41234_new_n2942_), .Y(_abc_41234_new_n2942__bF_buf1));
BUFX4 BUFX4_215 ( .A(_abc_41234_new_n2942_), .Y(_abc_41234_new_n2942__bF_buf0));
BUFX4 BUFX4_216 ( .A(_abc_41234_new_n515_), .Y(_abc_41234_new_n515__bF_buf6));
BUFX4 BUFX4_217 ( .A(_abc_41234_new_n515_), .Y(_abc_41234_new_n515__bF_buf5));
BUFX4 BUFX4_218 ( .A(_abc_41234_new_n515_), .Y(_abc_41234_new_n515__bF_buf4));
BUFX4 BUFX4_219 ( .A(_abc_41234_new_n515_), .Y(_abc_41234_new_n515__bF_buf3));
BUFX4 BUFX4_22 ( .A(clock), .Y(clock_bF_buf10));
BUFX4 BUFX4_220 ( .A(_abc_41234_new_n515_), .Y(_abc_41234_new_n515__bF_buf2));
BUFX4 BUFX4_221 ( .A(_abc_41234_new_n515_), .Y(_abc_41234_new_n515__bF_buf1));
BUFX4 BUFX4_222 ( .A(_abc_41234_new_n515_), .Y(_abc_41234_new_n515__bF_buf0));
BUFX4 BUFX4_223 ( .A(_abc_41234_new_n4297_), .Y(_abc_41234_new_n4297__bF_buf3));
BUFX4 BUFX4_224 ( .A(_abc_41234_new_n4297_), .Y(_abc_41234_new_n4297__bF_buf2));
BUFX4 BUFX4_225 ( .A(_abc_41234_new_n4297_), .Y(_abc_41234_new_n4297__bF_buf1));
BUFX4 BUFX4_226 ( .A(_abc_41234_new_n4297_), .Y(_abc_41234_new_n4297__bF_buf0));
BUFX4 BUFX4_227 ( .A(reset), .Y(reset_bF_buf9));
BUFX4 BUFX4_228 ( .A(reset), .Y(reset_bF_buf8));
BUFX4 BUFX4_229 ( .A(reset), .Y(reset_bF_buf7));
BUFX4 BUFX4_23 ( .A(clock), .Y(clock_bF_buf9));
BUFX4 BUFX4_230 ( .A(reset), .Y(reset_bF_buf6));
BUFX4 BUFX4_231 ( .A(reset), .Y(reset_bF_buf5));
BUFX4 BUFX4_232 ( .A(reset), .Y(reset_bF_buf4));
BUFX4 BUFX4_233 ( .A(reset), .Y(reset_bF_buf3));
BUFX4 BUFX4_234 ( .A(reset), .Y(reset_bF_buf2));
BUFX4 BUFX4_235 ( .A(reset), .Y(reset_bF_buf1));
BUFX4 BUFX4_236 ( .A(reset), .Y(reset_bF_buf0));
BUFX4 BUFX4_24 ( .A(clock), .Y(clock_bF_buf8));
BUFX4 BUFX4_25 ( .A(clock), .Y(clock_bF_buf7));
BUFX4 BUFX4_26 ( .A(clock), .Y(clock_bF_buf6));
BUFX4 BUFX4_27 ( .A(clock), .Y(clock_bF_buf5));
BUFX4 BUFX4_28 ( .A(clock), .Y(clock_bF_buf4));
BUFX4 BUFX4_29 ( .A(clock), .Y(clock_bF_buf3));
BUFX4 BUFX4_3 ( .A(clock_bF_buf13), .Y(clock_bF_buf13_bF_buf1));
BUFX4 BUFX4_30 ( .A(clock), .Y(clock_bF_buf2));
BUFX4 BUFX4_31 ( .A(clock), .Y(clock_bF_buf1));
BUFX4 BUFX4_32 ( .A(clock), .Y(clock_bF_buf0));
BUFX4 BUFX4_33 ( .A(_abc_41234_new_n1105_), .Y(_abc_41234_new_n1105__bF_buf3));
BUFX4 BUFX4_34 ( .A(_abc_41234_new_n1105_), .Y(_abc_41234_new_n1105__bF_buf2));
BUFX4 BUFX4_35 ( .A(_abc_41234_new_n1105_), .Y(_abc_41234_new_n1105__bF_buf1));
BUFX4 BUFX4_36 ( .A(_abc_41234_new_n1105_), .Y(_abc_41234_new_n1105__bF_buf0));
BUFX4 BUFX4_37 ( .A(_abc_41234_new_n2959_), .Y(_abc_41234_new_n2959__bF_buf3));
BUFX4 BUFX4_38 ( .A(_abc_41234_new_n2959_), .Y(_abc_41234_new_n2959__bF_buf2));
BUFX4 BUFX4_39 ( .A(_abc_41234_new_n2959_), .Y(_abc_41234_new_n2959__bF_buf1));
BUFX4 BUFX4_4 ( .A(clock_bF_buf13), .Y(clock_bF_buf13_bF_buf0));
BUFX4 BUFX4_40 ( .A(_abc_41234_new_n2959_), .Y(_abc_41234_new_n2959__bF_buf0));
BUFX4 BUFX4_41 ( .A(_abc_41234_new_n1046_), .Y(_abc_41234_new_n1046__bF_buf7));
BUFX4 BUFX4_42 ( .A(_abc_41234_new_n1046_), .Y(_abc_41234_new_n1046__bF_buf6));
BUFX4 BUFX4_43 ( .A(_abc_41234_new_n1046_), .Y(_abc_41234_new_n1046__bF_buf5));
BUFX4 BUFX4_44 ( .A(_abc_41234_new_n1046_), .Y(_abc_41234_new_n1046__bF_buf4));
BUFX4 BUFX4_45 ( .A(_abc_41234_new_n1046_), .Y(_abc_41234_new_n1046__bF_buf3));
BUFX4 BUFX4_46 ( .A(_abc_41234_new_n1046_), .Y(_abc_41234_new_n1046__bF_buf2));
BUFX4 BUFX4_47 ( .A(_abc_41234_new_n1046_), .Y(_abc_41234_new_n1046__bF_buf1));
BUFX4 BUFX4_48 ( .A(_abc_41234_new_n1046_), .Y(_abc_41234_new_n1046__bF_buf0));
BUFX4 BUFX4_49 ( .A(regfil_4__1_), .Y(regfil_4__1_bF_buf3_));
BUFX4 BUFX4_5 ( .A(clock_bF_buf14), .Y(clock_bF_buf14_bF_buf3));
BUFX4 BUFX4_50 ( .A(opcode_4_), .Y(opcode_4_bF_buf6_));
BUFX4 BUFX4_51 ( .A(opcode_4_), .Y(opcode_4_bF_buf5_));
BUFX4 BUFX4_52 ( .A(opcode_4_), .Y(opcode_4_bF_buf4_));
BUFX4 BUFX4_53 ( .A(opcode_4_), .Y(opcode_4_bF_buf3_));
BUFX4 BUFX4_54 ( .A(opcode_4_), .Y(opcode_4_bF_buf2_));
BUFX4 BUFX4_55 ( .A(opcode_4_), .Y(opcode_4_bF_buf1_));
BUFX4 BUFX4_56 ( .A(opcode_4_), .Y(opcode_4_bF_buf0_));
BUFX4 BUFX4_57 ( .A(_abc_41234_new_n2189_), .Y(_abc_41234_new_n2189__bF_buf5));
BUFX4 BUFX4_58 ( .A(_abc_41234_new_n2189_), .Y(_abc_41234_new_n2189__bF_buf4));
BUFX4 BUFX4_59 ( .A(_abc_41234_new_n2189_), .Y(_abc_41234_new_n2189__bF_buf3));
BUFX4 BUFX4_6 ( .A(clock_bF_buf14), .Y(clock_bF_buf14_bF_buf2));
BUFX4 BUFX4_60 ( .A(_abc_41234_new_n2189_), .Y(_abc_41234_new_n2189__bF_buf2));
BUFX4 BUFX4_61 ( .A(_abc_41234_new_n2189_), .Y(_abc_41234_new_n2189__bF_buf1));
BUFX4 BUFX4_62 ( .A(_abc_41234_new_n2189_), .Y(_abc_41234_new_n2189__bF_buf0));
BUFX4 BUFX4_63 ( .A(_abc_41234_new_n2207_), .Y(_abc_41234_new_n2207__bF_buf3));
BUFX4 BUFX4_64 ( .A(_abc_41234_new_n2207_), .Y(_abc_41234_new_n2207__bF_buf2));
BUFX4 BUFX4_65 ( .A(_abc_41234_new_n2207_), .Y(_abc_41234_new_n2207__bF_buf1));
BUFX4 BUFX4_66 ( .A(_abc_41234_new_n2207_), .Y(_abc_41234_new_n2207__bF_buf0));
BUFX4 BUFX4_67 ( .A(_abc_41234_new_n1040_), .Y(_abc_41234_new_n1040__bF_buf4));
BUFX4 BUFX4_68 ( .A(_abc_41234_new_n1040_), .Y(_abc_41234_new_n1040__bF_buf3));
BUFX4 BUFX4_69 ( .A(_abc_41234_new_n1040_), .Y(_abc_41234_new_n1040__bF_buf2));
BUFX4 BUFX4_7 ( .A(clock_bF_buf14), .Y(clock_bF_buf14_bF_buf1));
BUFX4 BUFX4_70 ( .A(_abc_41234_new_n1040_), .Y(_abc_41234_new_n1040__bF_buf1));
BUFX4 BUFX4_71 ( .A(_abc_41234_new_n1040_), .Y(_abc_41234_new_n1040__bF_buf0));
BUFX4 BUFX4_72 ( .A(regfil_5__6_), .Y(regfil_5__6_bF_buf3_));
BUFX4 BUFX4_73 ( .A(regfil_5__6_), .Y(regfil_5__6_bF_buf2_));
BUFX4 BUFX4_74 ( .A(regfil_5__6_), .Y(regfil_5__6_bF_buf1_));
BUFX4 BUFX4_75 ( .A(_abc_41234_new_n2947_), .Y(_abc_41234_new_n2947__bF_buf3));
BUFX4 BUFX4_76 ( .A(_abc_41234_new_n2947_), .Y(_abc_41234_new_n2947__bF_buf2));
BUFX4 BUFX4_77 ( .A(_abc_41234_new_n2947_), .Y(_abc_41234_new_n2947__bF_buf1));
BUFX4 BUFX4_78 ( .A(_abc_41234_new_n2947_), .Y(_abc_41234_new_n2947__bF_buf0));
BUFX4 BUFX4_79 ( .A(_abc_41234_new_n526_), .Y(_abc_41234_new_n526__bF_buf3));
BUFX4 BUFX4_8 ( .A(clock_bF_buf14), .Y(clock_bF_buf14_bF_buf0));
BUFX4 BUFX4_80 ( .A(_abc_41234_new_n526_), .Y(_abc_41234_new_n526__bF_buf2));
BUFX4 BUFX4_81 ( .A(_abc_41234_new_n526_), .Y(_abc_41234_new_n526__bF_buf1));
BUFX4 BUFX4_82 ( .A(_abc_41234_new_n526_), .Y(_abc_41234_new_n526__bF_buf0));
BUFX4 BUFX4_83 ( .A(regfil_5__3_), .Y(regfil_5__3_bF_buf3_));
BUFX4 BUFX4_84 ( .A(regfil_5__3_), .Y(regfil_5__3_bF_buf2_));
BUFX4 BUFX4_85 ( .A(_abc_41234_new_n620_), .Y(_abc_41234_new_n620__bF_buf5));
BUFX4 BUFX4_86 ( .A(_abc_41234_new_n620_), .Y(_abc_41234_new_n620__bF_buf4));
BUFX4 BUFX4_87 ( .A(_abc_41234_new_n620_), .Y(_abc_41234_new_n620__bF_buf3));
BUFX4 BUFX4_88 ( .A(_abc_41234_new_n620_), .Y(_abc_41234_new_n620__bF_buf2));
BUFX4 BUFX4_89 ( .A(_abc_41234_new_n620_), .Y(_abc_41234_new_n620__bF_buf1));
BUFX4 BUFX4_9 ( .A(_abc_41234_new_n544_), .Y(_abc_41234_new_n544__bF_buf3));
BUFX4 BUFX4_90 ( .A(_abc_41234_new_n620_), .Y(_abc_41234_new_n620__bF_buf0));
BUFX4 BUFX4_91 ( .A(_abc_41234_new_n523_), .Y(_abc_41234_new_n523__bF_buf4));
BUFX4 BUFX4_92 ( .A(_abc_41234_new_n523_), .Y(_abc_41234_new_n523__bF_buf3));
BUFX4 BUFX4_93 ( .A(_abc_41234_new_n523_), .Y(_abc_41234_new_n523__bF_buf2));
BUFX4 BUFX4_94 ( .A(_abc_41234_new_n523_), .Y(_abc_41234_new_n523__bF_buf1));
BUFX4 BUFX4_95 ( .A(_abc_41234_new_n523_), .Y(_abc_41234_new_n523__bF_buf0));
BUFX4 BUFX4_96 ( .A(_abc_41234_new_n1639_), .Y(_abc_41234_new_n1639__bF_buf3));
BUFX4 BUFX4_97 ( .A(_abc_41234_new_n1639_), .Y(_abc_41234_new_n1639__bF_buf2));
BUFX4 BUFX4_98 ( .A(_abc_41234_new_n1639_), .Y(_abc_41234_new_n1639__bF_buf0));
BUFX4 BUFX4_99 ( .A(_abc_41234_new_n1066_), .Y(_abc_41234_new_n1066__bF_buf3));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock_bF_buf14_bF_buf3), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_0_), .Q(state_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock_bF_buf5), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_3_), .Q(regfil_4__3_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clock_bF_buf5), .D(_0sp_15_0__8_), .Q(sp_8_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clock_bF_buf4), .D(_0sp_15_0__9_), .Q(sp_9_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clock_bF_buf3), .D(_0sp_15_0__10_), .Q(sp_10_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clock_bF_buf2), .D(_0sp_15_0__11_), .Q(sp_11_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clock_bF_buf1), .D(_0sp_15_0__12_), .Q(sp_12_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clock_bF_buf0), .D(_0sp_15_0__13_), .Q(sp_13_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clock_bF_buf14_bF_buf0), .D(_0sp_15_0__14_), .Q(sp_14_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clock_bF_buf13_bF_buf0), .D(_0sp_15_0__15_), .Q(sp_15_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clock_bF_buf12), .D(_0regd_2_0__0_), .Q(regd_0_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clock_bF_buf11), .D(_0regd_2_0__1_), .Q(regd_1_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock_bF_buf4), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_4_), .Q(regfil_4__4_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clock_bF_buf10), .D(_0regd_2_0__2_), .Q(regd_2_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clock_bF_buf9), .D(_0datao_7_0__0_), .Q(\data[0] ));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clock_bF_buf8), .D(_0datao_7_0__1_), .Q(\data[1] ));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clock_bF_buf7), .D(_0datao_7_0__2_), .Q(\data[2] ));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clock_bF_buf6), .D(_0datao_7_0__3_), .Q(\data[3] ));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clock_bF_buf5), .D(_0datao_7_0__4_), .Q(\data[4] ));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clock_bF_buf4), .D(_0datao_7_0__5_), .Q(\data[5] ));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clock_bF_buf3), .D(_0datao_7_0__6_), .Q(\data[6] ));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clock_bF_buf2), .D(_0datao_7_0__7_), .Q(\data[7] ));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clock_bF_buf1), .D(_0waddrhold_15_0__0_), .Q(waddrhold_0_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock_bF_buf3), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_5_), .Q(regfil_4__5_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clock_bF_buf0), .D(_0waddrhold_15_0__1_), .Q(waddrhold_1_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clock_bF_buf14_bF_buf3), .D(_0waddrhold_15_0__2_), .Q(waddrhold_2_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clock_bF_buf13_bF_buf3), .D(_0waddrhold_15_0__3_), .Q(waddrhold_3_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clock_bF_buf12), .D(_0waddrhold_15_0__4_), .Q(waddrhold_4_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clock_bF_buf11), .D(_0waddrhold_15_0__5_), .Q(waddrhold_5_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clock_bF_buf10), .D(_0waddrhold_15_0__6_), .Q(waddrhold_6_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clock_bF_buf9), .D(_0waddrhold_15_0__7_), .Q(waddrhold_7_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clock_bF_buf8), .D(_0waddrhold_15_0__8_), .Q(waddrhold_8_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clock_bF_buf7), .D(_0waddrhold_15_0__9_), .Q(waddrhold_9_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clock_bF_buf6), .D(_0waddrhold_15_0__10_), .Q(waddrhold_10_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock_bF_buf2), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_6_), .Q(regfil_4__6_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clock_bF_buf5), .D(_0waddrhold_15_0__11_), .Q(waddrhold_11_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clock_bF_buf4), .D(_0waddrhold_15_0__12_), .Q(waddrhold_12_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clock_bF_buf3), .D(_0waddrhold_15_0__13_), .Q(waddrhold_13_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clock_bF_buf2), .D(_0waddrhold_15_0__14_), .Q(waddrhold_14_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clock_bF_buf1), .D(_0waddrhold_15_0__15_), .Q(waddrhold_15_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clock_bF_buf0), .D(_0raddrhold_15_0__0_), .Q(raddrhold_0_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clock_bF_buf14_bF_buf2), .D(_0raddrhold_15_0__1_), .Q(raddrhold_1_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clock_bF_buf13_bF_buf2), .D(_0raddrhold_15_0__2_), .Q(raddrhold_2_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clock_bF_buf12), .D(_0raddrhold_15_0__3_), .Q(raddrhold_3_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clock_bF_buf11), .D(_0raddrhold_15_0__4_), .Q(raddrhold_4_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock_bF_buf1), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_7_), .Q(regfil_4__7_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clock_bF_buf10), .D(_0raddrhold_15_0__5_), .Q(raddrhold_5_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clock_bF_buf9), .D(_0raddrhold_15_0__6_), .Q(raddrhold_6_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clock_bF_buf8), .D(_0raddrhold_15_0__7_), .Q(raddrhold_7_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clock_bF_buf7), .D(_0raddrhold_15_0__8_), .Q(raddrhold_8_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clock_bF_buf6), .D(_0raddrhold_15_0__9_), .Q(raddrhold_9_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clock_bF_buf5), .D(_0raddrhold_15_0__10_), .Q(raddrhold_10_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clock_bF_buf4), .D(_0raddrhold_15_0__11_), .Q(raddrhold_11_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clock_bF_buf3), .D(_0raddrhold_15_0__12_), .Q(raddrhold_12_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clock_bF_buf2), .D(_0raddrhold_15_0__13_), .Q(raddrhold_13_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clock_bF_buf1), .D(_0raddrhold_15_0__14_), .Q(raddrhold_14_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock_bF_buf0), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_0_), .Q(regfil_5__0_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clock_bF_buf0), .D(_0raddrhold_15_0__15_), .Q(raddrhold_15_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clock_bF_buf14_bF_buf1), .D(_0wdatahold_7_0__0_), .Q(wdatahold_0_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clock_bF_buf13_bF_buf1), .D(_0wdatahold_7_0__1_), .Q(wdatahold_1_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clock_bF_buf12), .D(_0wdatahold_7_0__2_), .Q(wdatahold_2_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clock_bF_buf11), .D(_0wdatahold_7_0__3_), .Q(wdatahold_3_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clock_bF_buf10), .D(_0wdatahold_7_0__4_), .Q(wdatahold_4_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clock_bF_buf9), .D(_0wdatahold_7_0__5_), .Q(wdatahold_5_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clock_bF_buf8), .D(_0wdatahold_7_0__6_), .Q(wdatahold_6_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clock_bF_buf7), .D(_0wdatahold_7_0__7_), .Q(wdatahold_7_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clock_bF_buf6), .D(_0wdatahold2_7_0__0_), .Q(wdatahold2_0_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock_bF_buf14_bF_buf2), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_1_), .Q(regfil_5__1_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clock_bF_buf5), .D(_0wdatahold2_7_0__1_), .Q(wdatahold2_1_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clock_bF_buf4), .D(_0wdatahold2_7_0__2_), .Q(wdatahold2_2_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clock_bF_buf3), .D(_0wdatahold2_7_0__3_), .Q(wdatahold2_3_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clock_bF_buf2), .D(_0wdatahold2_7_0__4_), .Q(wdatahold2_4_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clock_bF_buf1), .D(_0wdatahold2_7_0__5_), .Q(wdatahold2_5_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clock_bF_buf0), .D(_0wdatahold2_7_0__6_), .Q(wdatahold2_6_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clock_bF_buf14_bF_buf0), .D(_0wdatahold2_7_0__7_), .Q(wdatahold2_7_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clock_bF_buf13_bF_buf0), .D(_0rdatahold_7_0__0_), .Q(rdatahold_0_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clock_bF_buf12), .D(_0rdatahold_7_0__1_), .Q(rdatahold_1_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clock_bF_buf11), .D(_0rdatahold_7_0__2_), .Q(rdatahold_2_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock_bF_buf13_bF_buf2), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_2_), .Q(regfil_5__2_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clock_bF_buf10), .D(_0rdatahold_7_0__3_), .Q(rdatahold_3_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clock_bF_buf9), .D(_0rdatahold_7_0__4_), .Q(rdatahold_4_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clock_bF_buf8), .D(_0rdatahold_7_0__5_), .Q(rdatahold_5_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clock_bF_buf7), .D(_0rdatahold_7_0__6_), .Q(rdatahold_6_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clock_bF_buf6), .D(_0rdatahold_7_0__7_), .Q(rdatahold_7_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clock_bF_buf5), .D(_0rdatahold2_7_0__0_), .Q(rdatahold2_0_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clock_bF_buf4), .D(_0rdatahold2_7_0__1_), .Q(rdatahold2_1_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clock_bF_buf3), .D(_0rdatahold2_7_0__2_), .Q(rdatahold2_2_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clock_bF_buf2), .D(_0rdatahold2_7_0__3_), .Q(rdatahold2_3_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clock_bF_buf1), .D(_0rdatahold2_7_0__4_), .Q(rdatahold2_4_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock_bF_buf12), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_3_), .Q(regfil_5__3_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clock_bF_buf0), .D(_0rdatahold2_7_0__5_), .Q(rdatahold2_5_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clock_bF_buf14_bF_buf3), .D(_0rdatahold2_7_0__6_), .Q(rdatahold2_6_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clock_bF_buf13_bF_buf3), .D(_0rdatahold2_7_0__7_), .Q(rdatahold2_7_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clock_bF_buf12), .D(_0popdes_1_0__0_), .Q(popdes_0_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clock_bF_buf11), .D(_0popdes_1_0__1_), .Q(popdes_1_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clock_bF_buf10), .D(_0statesel_5_0__0_), .Q(statesel_0_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clock_bF_buf9), .D(_0statesel_5_0__1_), .Q(statesel_1_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clock_bF_buf8), .D(_0statesel_5_0__2_), .Q(statesel_2_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clock_bF_buf7), .D(_0statesel_5_0__3_), .Q(statesel_3_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clock_bF_buf6), .D(_0statesel_5_0__4_), .Q(statesel_4_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock_bF_buf11), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_4_), .Q(regfil_5__4_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clock_bF_buf5), .D(_0statesel_5_0__5_), .Q(statesel_5_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clock_bF_buf4), .D(_0eienb_0_0_), .Q(eienb));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clock_bF_buf3), .D(_0opcode_7_0__0_), .Q(opcode_0_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clock_bF_buf2), .D(_0opcode_7_0__1_), .Q(opcode_1_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clock_bF_buf1), .D(_0opcode_7_0__2_), .Q(opcode_2_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clock_bF_buf0), .D(_0opcode_7_0__3_), .Q(opcode_3_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clock_bF_buf14_bF_buf2), .D(_0opcode_7_0__4_), .Q(opcode_4_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clock_bF_buf13_bF_buf2), .D(_0opcode_7_0__5_), .Q(opcode_5_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clock_bF_buf12), .D(_0opcode_7_0__6_), .Q(opcode_6_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clock_bF_buf11), .D(_0opcode_7_0__7_), .Q(opcode_7_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock_bF_buf13_bF_buf3), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_1_), .Q(state_1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock_bF_buf10), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_5_), .Q(regfil_5__5_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clock_bF_buf10), .D(_0carry_0_0_), .Q(carry));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clock_bF_buf9), .D(_0auxcar_0_0_), .Q(auxcar));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clock_bF_buf8), .D(_0sign_0_0_), .Q(sign));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clock_bF_buf7), .D(_0zero_0_0_), .Q(zero));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clock_bF_buf6), .D(_0parity_0_0_), .Q(parity));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clock_bF_buf5), .D(_0ei_0_0_), .Q(ei));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clock_bF_buf4), .D(_0intcyc_0_0_), .Q(intcyc));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clock_bF_buf3), .D(_0aluopra_7_0__0_), .Q(alu_opra_0_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clock_bF_buf2), .D(_0aluopra_7_0__1_), .Q(alu_opra_1_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clock_bF_buf1), .D(_0aluopra_7_0__2_), .Q(alu_opra_2_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock_bF_buf9), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_6_), .Q(regfil_5__6_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clock_bF_buf0), .D(_0aluopra_7_0__3_), .Q(alu_opra_3_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clock_bF_buf14_bF_buf1), .D(_0aluopra_7_0__4_), .Q(alu_opra_4_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clock_bF_buf13_bF_buf1), .D(_0aluopra_7_0__5_), .Q(alu_opra_5_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clock_bF_buf12), .D(_0aluopra_7_0__6_), .Q(alu_opra_6_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clock_bF_buf11), .D(_0aluopra_7_0__7_), .Q(alu_opra_7_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clock_bF_buf10), .D(_0aluoprb_7_0__0_), .Q(alu_oprb_0_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clock_bF_buf9), .D(_0aluoprb_7_0__1_), .Q(alu_oprb_1_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clock_bF_buf8), .D(_0aluoprb_7_0__2_), .Q(alu_oprb_2_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clock_bF_buf7), .D(_0aluoprb_7_0__3_), .Q(alu_oprb_3_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clock_bF_buf6), .D(_0aluoprb_7_0__4_), .Q(alu_oprb_4_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock_bF_buf8), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_7_), .Q(regfil_5__7_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clock_bF_buf5), .D(_0aluoprb_7_0__5_), .Q(alu_oprb_5_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clock_bF_buf4), .D(_0aluoprb_7_0__6_), .Q(alu_oprb_6_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clock_bF_buf3), .D(_0aluoprb_7_0__7_), .Q(alu_oprb_7_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clock_bF_buf2), .D(_0alucin_0_0_), .Q(alu_cin));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clock_bF_buf1), .D(_0alusel_2_0__0_), .Q(alu_sel_0_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clock_bF_buf0), .D(_0alusel_2_0__1_), .Q(alu_sel_1_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clock_bF_buf14_bF_buf0), .D(_0alusel_2_0__2_), .Q(alu_sel_2_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clock_bF_buf13_bF_buf0), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_0_), .Q(regfil_7__0_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clock_bF_buf12), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_1_), .Q(regfil_7__1_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clock_bF_buf11), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_2_), .Q(regfil_7__2_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock_bF_buf7), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_0_), .Q(regfil_1__0_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clock_bF_buf10), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_3_), .Q(regfil_7__3_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clock_bF_buf9), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_4_), .Q(regfil_7__4_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clock_bF_buf8), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_5_), .Q(regfil_7__5_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clock_bF_buf7), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_6_), .Q(regfil_7__6_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clock_bF_buf6), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_7_), .Q(regfil_7__7_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clock_bF_buf5), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_0_), .Q(regfil_3__0_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clock_bF_buf4), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_1_), .Q(regfil_3__1_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clock_bF_buf3), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_2_), .Q(regfil_3__2_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clock_bF_buf2), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_3_), .Q(regfil_3__3_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clock_bF_buf1), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_4_), .Q(regfil_3__4_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock_bF_buf6), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_1_), .Q(regfil_1__1_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clock_bF_buf0), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_5_), .Q(regfil_3__5_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clock_bF_buf14_bF_buf3), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_6_), .Q(regfil_3__6_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clock_bF_buf13_bF_buf3), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_7_), .Q(regfil_3__7_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock_bF_buf5), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_2_), .Q(regfil_1__2_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock_bF_buf4), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_3_), .Q(regfil_1__3_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock_bF_buf3), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_4_), .Q(regfil_1__4_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock_bF_buf2), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_5_), .Q(regfil_1__5_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock_bF_buf1), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_6_), .Q(regfil_1__6_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock_bF_buf12), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_2_), .Q(state_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock_bF_buf0), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_7_), .Q(regfil_1__7_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock_bF_buf14_bF_buf1), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_0_), .Q(regfil_6__0_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock_bF_buf13_bF_buf1), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_1_), .Q(regfil_6__1_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock_bF_buf12), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_2_), .Q(regfil_6__2_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock_bF_buf11), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_3_), .Q(regfil_6__3_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock_bF_buf10), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_4_), .Q(regfil_6__4_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock_bF_buf9), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_5_), .Q(regfil_6__5_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock_bF_buf8), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_6_), .Q(regfil_6__6_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock_bF_buf7), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_7_), .Q(regfil_6__7_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock_bF_buf6), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_0_), .Q(regfil_2__0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock_bF_buf11), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_3_), .Q(state_3_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock_bF_buf5), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_1_), .Q(regfil_2__1_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock_bF_buf4), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_2_), .Q(regfil_2__2_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock_bF_buf3), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_3_), .Q(regfil_2__3_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock_bF_buf2), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_4_), .Q(regfil_2__4_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock_bF_buf1), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_5_), .Q(regfil_2__5_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock_bF_buf0), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_6_), .Q(regfil_2__6_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock_bF_buf14_bF_buf0), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_7_), .Q(regfil_2__7_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock_bF_buf13_bF_buf0), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_0_), .Q(regfil_0__0_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock_bF_buf12), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_1_), .Q(regfil_0__1_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock_bF_buf11), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_2_), .Q(regfil_0__2_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock_bF_buf10), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_4_), .Q(state_4_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock_bF_buf10), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_3_), .Q(regfil_0__3_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock_bF_buf9), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_4_), .Q(regfil_0__4_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock_bF_buf8), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_5_), .Q(regfil_0__5_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock_bF_buf7), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_6_), .Q(regfil_0__6_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock_bF_buf6), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_7_), .Q(regfil_0__7_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock_bF_buf5), .D(_0writeio_0_0_), .Q(_auto_iopadmap_cc_368_execute_45651));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock_bF_buf4), .D(_0inta_0_0_), .Q(_auto_iopadmap_cc_368_execute_45645));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock_bF_buf3), .D(_0readio_0_0_), .Q(_auto_iopadmap_cc_368_execute_45647));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock_bF_buf2), .D(_0addr_15_0__0_), .Q(_auto_iopadmap_cc_368_execute_45628_0_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock_bF_buf1), .D(_0addr_15_0__1_), .Q(_auto_iopadmap_cc_368_execute_45628_1_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock_bF_buf9), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_5_), .Q(state_5_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock_bF_buf0), .D(_0addr_15_0__2_), .Q(_auto_iopadmap_cc_368_execute_45628_2_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock_bF_buf14_bF_buf3), .D(_0addr_15_0__3_), .Q(_auto_iopadmap_cc_368_execute_45628_3_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock_bF_buf13_bF_buf3), .D(_0addr_15_0__4_), .Q(_auto_iopadmap_cc_368_execute_45628_4_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock_bF_buf12), .D(_0addr_15_0__5_), .Q(_auto_iopadmap_cc_368_execute_45628_5_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock_bF_buf11), .D(_0addr_15_0__6_), .Q(_auto_iopadmap_cc_368_execute_45628_6_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock_bF_buf10), .D(_0addr_15_0__7_), .Q(_auto_iopadmap_cc_368_execute_45628_7_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock_bF_buf9), .D(_0addr_15_0__8_), .Q(_auto_iopadmap_cc_368_execute_45628_8_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clock_bF_buf8), .D(_0addr_15_0__9_), .Q(_auto_iopadmap_cc_368_execute_45628_9_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clock_bF_buf7), .D(_0addr_15_0__10_), .Q(_auto_iopadmap_cc_368_execute_45628_10_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clock_bF_buf6), .D(_0addr_15_0__11_), .Q(_auto_iopadmap_cc_368_execute_45628_11_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock_bF_buf8), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_0_), .Q(regfil_4__0_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clock_bF_buf5), .D(_0addr_15_0__12_), .Q(_auto_iopadmap_cc_368_execute_45628_12_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clock_bF_buf4), .D(_0addr_15_0__13_), .Q(_auto_iopadmap_cc_368_execute_45628_13_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clock_bF_buf3), .D(_0addr_15_0__14_), .Q(_auto_iopadmap_cc_368_execute_45628_14_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clock_bF_buf2), .D(_0addr_15_0__15_), .Q(_auto_iopadmap_cc_368_execute_45628_15_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clock_bF_buf1), .D(_0readmem_0_0_), .Q(_auto_iopadmap_cc_368_execute_45649));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clock_bF_buf0), .D(_0writemem_0_0_), .Q(_auto_iopadmap_cc_368_execute_45653));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clock_bF_buf14_bF_buf2), .D(_0pc_15_0__0_), .Q(pc_0_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clock_bF_buf13_bF_buf2), .D(_0pc_15_0__1_), .Q(pc_1_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clock_bF_buf12), .D(_0pc_15_0__2_), .Q(pc_2_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clock_bF_buf11), .D(_0pc_15_0__3_), .Q(pc_3_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock_bF_buf7), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_1_), .Q(regfil_4__1_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clock_bF_buf10), .D(_0pc_15_0__4_), .Q(pc_4_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clock_bF_buf9), .D(_0pc_15_0__5_), .Q(pc_5_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clock_bF_buf8), .D(_0pc_15_0__6_), .Q(pc_6_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clock_bF_buf7), .D(_0pc_15_0__7_), .Q(pc_7_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clock_bF_buf6), .D(_0pc_15_0__8_), .Q(pc_8_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clock_bF_buf5), .D(_0pc_15_0__9_), .Q(pc_9_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clock_bF_buf4), .D(_0pc_15_0__10_), .Q(pc_10_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clock_bF_buf3), .D(_0pc_15_0__11_), .Q(pc_11_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clock_bF_buf2), .D(_0pc_15_0__12_), .Q(pc_12_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clock_bF_buf1), .D(_0pc_15_0__13_), .Q(pc_13_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock_bF_buf6), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_2_), .Q(regfil_4__2_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clock_bF_buf0), .D(_0pc_15_0__14_), .Q(pc_14_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clock_bF_buf14_bF_buf1), .D(_0pc_15_0__15_), .Q(pc_15_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clock_bF_buf13_bF_buf1), .D(_0sp_15_0__0_), .Q(sp_0_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clock_bF_buf12), .D(_0sp_15_0__1_), .Q(sp_1_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clock_bF_buf11), .D(_0sp_15_0__2_), .Q(sp_2_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clock_bF_buf10), .D(_0sp_15_0__3_), .Q(sp_3_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clock_bF_buf9), .D(_0sp_15_0__4_), .Q(sp_4_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clock_bF_buf8), .D(_0sp_15_0__5_), .Q(sp_5_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clock_bF_buf7), .D(_0sp_15_0__6_), .Q(sp_6_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clock_bF_buf6), .D(_0sp_15_0__7_), .Q(sp_7_));
INVX1 INVX1_1 ( .A(state_4_), .Y(_abc_41234_new_n501_));
INVX1 INVX1_10 ( .A(state_2_), .Y(_abc_41234_new_n589_));
INVX1 INVX1_100 ( .A(_abc_41234_new_n527_), .Y(_abc_41234_new_n1625_));
INVX1 INVX1_101 ( .A(_abc_41234_new_n1628_), .Y(_abc_41234_new_n1629_));
INVX1 INVX1_102 ( .A(wdatahold2_1_), .Y(_abc_41234_new_n1666_));
INVX1 INVX1_103 ( .A(_abc_41234_new_n1620_), .Y(_abc_41234_new_n1671_));
INVX1 INVX1_104 ( .A(_abc_41234_new_n1673_), .Y(_abc_41234_new_n1674_));
INVX1 INVX1_105 ( .A(_abc_41234_new_n1651_), .Y(_abc_41234_new_n1677_));
INVX1 INVX1_106 ( .A(_abc_41234_new_n581_), .Y(_abc_41234_new_n1682_));
INVX1 INVX1_107 ( .A(_abc_41234_new_n1686_), .Y(_abc_41234_new_n1687_));
INVX1 INVX1_108 ( .A(_abc_41234_new_n1692_), .Y(_abc_41234_new_n1693_));
INVX1 INVX1_109 ( .A(wdatahold2_2_), .Y(_abc_41234_new_n1697_));
INVX1 INVX1_11 ( .A(_abc_41234_new_n591_), .Y(_abc_41234_new_n592_));
INVX1 INVX1_110 ( .A(_abc_41234_new_n1706_), .Y(_abc_41234_new_n1707_));
INVX1 INVX1_111 ( .A(_abc_41234_new_n1709_), .Y(_abc_41234_new_n1710_));
INVX1 INVX1_112 ( .A(wdatahold2_3_), .Y(_abc_41234_new_n1724_));
INVX1 INVX1_113 ( .A(_abc_41234_new_n1730_), .Y(_abc_41234_new_n1731_));
INVX1 INVX1_114 ( .A(wdatahold2_4_), .Y(_abc_41234_new_n1746_));
INVX1 INVX1_115 ( .A(_abc_41234_new_n1755_), .Y(_abc_41234_new_n1756_));
INVX1 INVX1_116 ( .A(wdatahold2_5_), .Y(_abc_41234_new_n1771_));
INVX1 INVX1_117 ( .A(wdatahold2_6_), .Y(_abc_41234_new_n1793_));
INVX1 INVX1_118 ( .A(_abc_41234_new_n1804_), .Y(_abc_41234_new_n1805_));
INVX1 INVX1_119 ( .A(_abc_41234_new_n1809_), .Y(_abc_41234_new_n1810_));
INVX1 INVX1_12 ( .A(_abc_41234_new_n506_), .Y(_abc_41234_new_n603_));
INVX1 INVX1_120 ( .A(wdatahold2_7_), .Y(_abc_41234_new_n1821_));
INVX1 INVX1_121 ( .A(_abc_41234_new_n1853_), .Y(_abc_41234_new_n1854_));
INVX1 INVX1_122 ( .A(_abc_41234_new_n1857_), .Y(_abc_41234_new_n1864_));
INVX1 INVX1_123 ( .A(_abc_41234_new_n1902_), .Y(_abc_41234_new_n1903_));
INVX1 INVX1_124 ( .A(_abc_41234_new_n1912_), .Y(_abc_41234_new_n1913_));
INVX1 INVX1_125 ( .A(_abc_41234_new_n1925_), .Y(_abc_41234_new_n1926_));
INVX1 INVX1_126 ( .A(_abc_41234_new_n1929_), .Y(_abc_41234_new_n1930_));
INVX1 INVX1_127 ( .A(_abc_41234_new_n1943_), .Y(_abc_41234_new_n1944_));
INVX1 INVX1_128 ( .A(_abc_41234_new_n1957_), .Y(_abc_41234_new_n1958_));
INVX1 INVX1_129 ( .A(_abc_41234_new_n571_), .Y(_abc_41234_new_n1975_));
INVX1 INVX1_13 ( .A(_abc_41234_new_n604_), .Y(_abc_41234_new_n605_));
INVX1 INVX1_130 ( .A(_abc_41234_new_n636_), .Y(_abc_41234_new_n2002_));
INVX1 INVX1_131 ( .A(_abc_41234_new_n2019_), .Y(_abc_41234_new_n2021_));
INVX1 INVX1_132 ( .A(_abc_41234_new_n2027_), .Y(_abc_41234_new_n2028_));
INVX1 INVX1_133 ( .A(regfil_6__6_), .Y(_abc_41234_new_n2048_));
INVX1 INVX1_134 ( .A(_abc_41234_new_n2060_), .Y(_abc_41234_new_n2061_));
INVX1 INVX1_135 ( .A(_abc_41234_new_n2107_), .Y(_abc_41234_new_n2108_));
INVX1 INVX1_136 ( .A(_abc_41234_new_n2144_), .Y(_abc_41234_new_n2147_));
INVX1 INVX1_137 ( .A(_abc_41234_new_n2175_), .Y(_abc_41234_new_n2176_));
INVX1 INVX1_138 ( .A(alu_sel_1_), .Y(_abc_41234_new_n2184_));
INVX1 INVX1_139 ( .A(alu_sel_2_), .Y(_abc_41234_new_n2196_));
INVX1 INVX1_14 ( .A(_abc_41234_new_n613_), .Y(_abc_41234_new_n614_));
INVX1 INVX1_140 ( .A(_abc_41234_new_n627_), .Y(_abc_41234_new_n2205_));
INVX1 INVX1_141 ( .A(alu_oprb_0_), .Y(_abc_41234_new_n2206_));
INVX1 INVX1_142 ( .A(_abc_41234_new_n2208_), .Y(_abc_41234_new_n2209_));
INVX1 INVX1_143 ( .A(_abc_41234_new_n2212_), .Y(_abc_41234_new_n2213_));
INVX1 INVX1_144 ( .A(_abc_41234_new_n2214_), .Y(_abc_41234_new_n2215_));
INVX1 INVX1_145 ( .A(alu_oprb_1_), .Y(_abc_41234_new_n2220_));
INVX1 INVX1_146 ( .A(alu_oprb_2_), .Y(_abc_41234_new_n2227_));
INVX1 INVX1_147 ( .A(alu_oprb_4_), .Y(_abc_41234_new_n2233_));
INVX1 INVX1_148 ( .A(alu_oprb_5_), .Y(_abc_41234_new_n2236_));
INVX1 INVX1_149 ( .A(alu_oprb_7_), .Y(_abc_41234_new_n2242_));
INVX1 INVX1_15 ( .A(regfil_1__7_), .Y(_abc_41234_new_n637_));
INVX1 INVX1_150 ( .A(_abc_41234_new_n2258_), .Y(_abc_41234_new_n2259_));
INVX1 INVX1_151 ( .A(_abc_41234_new_n2261_), .Y(_abc_41234_new_n2262_));
INVX1 INVX1_152 ( .A(_abc_41234_new_n2276_), .Y(_abc_41234_new_n2277_));
INVX1 INVX1_153 ( .A(_abc_41234_new_n2288_), .Y(_abc_41234_new_n2289_));
INVX1 INVX1_154 ( .A(_abc_41234_new_n2300_), .Y(_abc_41234_new_n2301_));
INVX1 INVX1_155 ( .A(_abc_41234_new_n2312_), .Y(_abc_41234_new_n2313_));
INVX1 INVX1_156 ( .A(ei), .Y(_abc_41234_new_n2354_));
INVX1 INVX1_157 ( .A(intr), .Y(_abc_41234_new_n2355_));
INVX1 INVX1_158 ( .A(parity), .Y(_abc_41234_new_n2361_));
INVX1 INVX1_159 ( .A(_abc_41234_new_n2363_), .Y(_abc_41234_new_n2364_));
INVX1 INVX1_16 ( .A(regd_2_), .Y(_abc_41234_new_n649_));
INVX1 INVX1_160 ( .A(rdatahold2_2_), .Y(_abc_41234_new_n2365_));
INVX1 INVX1_161 ( .A(rdatahold2_7_), .Y(_abc_41234_new_n2377_));
INVX1 INVX1_162 ( .A(alu_sout), .Y(_abc_41234_new_n2379_));
INVX1 INVX1_163 ( .A(_abc_41234_new_n1546_), .Y(_abc_41234_new_n2396_));
INVX1 INVX1_164 ( .A(_abc_41234_new_n1323_), .Y(_abc_41234_new_n2398_));
INVX1 INVX1_165 ( .A(alu_cout), .Y(_abc_41234_new_n2418_));
INVX1 INVX1_166 ( .A(_abc_41234_new_n2428_), .Y(_abc_41234_new_n2429_));
INVX1 INVX1_167 ( .A(\data[1] ), .Y(_abc_41234_new_n2432_));
INVX1 INVX1_168 ( .A(\data[2] ), .Y(_abc_41234_new_n2435_));
INVX1 INVX1_169 ( .A(\data[3] ), .Y(_abc_41234_new_n2437_));
INVX1 INVX1_17 ( .A(regd_1_), .Y(_abc_41234_new_n654_));
INVX1 INVX1_170 ( .A(\data[5] ), .Y(_abc_41234_new_n2441_));
INVX1 INVX1_171 ( .A(\data[6] ), .Y(_abc_41234_new_n2443_));
INVX1 INVX1_172 ( .A(_abc_41234_new_n2449_), .Y(_abc_41234_new_n2450_));
INVX1 INVX1_173 ( .A(_abc_41234_new_n2460_), .Y(_abc_41234_new_n2461_));
INVX1 INVX1_174 ( .A(_abc_41234_new_n2474_), .Y(_abc_41234_new_n2475_));
INVX1 INVX1_175 ( .A(_abc_41234_new_n2476_), .Y(_abc_41234_new_n2477_));
INVX1 INVX1_176 ( .A(_abc_41234_new_n2486_), .Y(_abc_41234_new_n2487_));
INVX1 INVX1_177 ( .A(_abc_41234_new_n2502_), .Y(_abc_41234_new_n2503_));
INVX1 INVX1_178 ( .A(_abc_41234_new_n2528_), .Y(_abc_41234_new_n2529_));
INVX1 INVX1_179 ( .A(_abc_41234_new_n2530_), .Y(_abc_41234_new_n2531_));
INVX1 INVX1_18 ( .A(_abc_41234_new_n615_), .Y(_abc_41234_new_n657_));
INVX1 INVX1_180 ( .A(_abc_41234_new_n2543_), .Y(_abc_41234_new_n2544_));
INVX1 INVX1_181 ( .A(statesel_1_), .Y(_abc_41234_new_n2556_));
INVX1 INVX1_182 ( .A(_abc_41234_new_n2559_), .Y(_abc_41234_new_n2560_));
INVX1 INVX1_183 ( .A(_abc_41234_new_n2493_), .Y(_abc_41234_new_n2571_));
INVX1 INVX1_184 ( .A(_abc_41234_new_n2525_), .Y(_abc_41234_new_n2577_));
INVX1 INVX1_185 ( .A(_abc_41234_new_n2579_), .Y(_abc_41234_new_n2580_));
INVX1 INVX1_186 ( .A(_abc_41234_new_n2601_), .Y(_abc_41234_new_n2602_));
INVX1 INVX1_187 ( .A(_abc_41234_new_n2597_), .Y(_abc_41234_new_n2613_));
INVX1 INVX1_188 ( .A(_abc_41234_new_n2624_), .Y(_abc_41234_new_n2633_));
INVX1 INVX1_189 ( .A(_abc_41234_new_n2526_), .Y(_abc_41234_new_n2634_));
INVX1 INVX1_19 ( .A(_abc_41234_new_n521_), .Y(_abc_41234_new_n658_));
INVX1 INVX1_190 ( .A(_abc_41234_new_n2622_), .Y(_abc_41234_new_n2638_));
INVX1 INVX1_191 ( .A(_abc_41234_new_n2639_), .Y(_abc_41234_new_n2640_));
INVX1 INVX1_192 ( .A(rdatahold2_1_), .Y(_abc_41234_new_n2651_));
INVX1 INVX1_193 ( .A(rdatahold2_5_), .Y(_abc_41234_new_n2658_));
INVX1 INVX1_194 ( .A(wdatahold_0_), .Y(_abc_41234_new_n2670_));
INVX1 INVX1_195 ( .A(wdatahold_1_), .Y(_abc_41234_new_n2701_));
INVX1 INVX1_196 ( .A(_abc_41234_new_n2515_), .Y(_abc_41234_new_n2727_));
INVX1 INVX1_197 ( .A(wdatahold_2_), .Y(_abc_41234_new_n2731_));
INVX1 INVX1_198 ( .A(_abc_41234_new_n2737_), .Y(_abc_41234_new_n2738_));
INVX1 INVX1_199 ( .A(wdatahold_3_), .Y(_abc_41234_new_n2764_));
INVX1 INVX1_2 ( .A(state_3_), .Y(_abc_41234_new_n503_));
INVX1 INVX1_20 ( .A(_abc_41234_new_n666_), .Y(_abc_41234_new_n667_));
INVX1 INVX1_200 ( .A(_abc_41234_new_n2732_), .Y(_abc_41234_new_n2771_));
INVX1 INVX1_201 ( .A(wdatahold_4_), .Y(_abc_41234_new_n2792_));
INVX1 INVX1_202 ( .A(_abc_41234_new_n1616_), .Y(_abc_41234_new_n2803_));
INVX1 INVX1_203 ( .A(auxcar), .Y(_abc_41234_new_n2809_));
INVX1 INVX1_204 ( .A(wdatahold_5_), .Y(_abc_41234_new_n2824_));
INVX1 INVX1_205 ( .A(pc_5_), .Y(_abc_41234_new_n2831_));
INVX1 INVX1_206 ( .A(wdatahold_6_), .Y(_abc_41234_new_n2851_));
INVX1 INVX1_207 ( .A(_abc_41234_new_n2854_), .Y(_abc_41234_new_n2855_));
INVX1 INVX1_208 ( .A(_abc_41234_new_n1617_), .Y(_abc_41234_new_n2856_));
INVX1 INVX1_209 ( .A(wdatahold_7_), .Y(_abc_41234_new_n2881_));
INVX1 INVX1_21 ( .A(regd_0_), .Y(_abc_41234_new_n673_));
INVX1 INVX1_210 ( .A(_abc_41234_new_n2931_), .Y(_abc_41234_new_n2933_));
INVX1 INVX1_211 ( .A(_abc_41234_new_n2456_), .Y(_abc_41234_new_n2934_));
INVX1 INVX1_212 ( .A(_abc_41234_new_n2979_), .Y(_abc_41234_new_n2980_));
INVX1 INVX1_213 ( .A(_abc_41234_new_n2998_), .Y(_abc_41234_new_n2999_));
INVX1 INVX1_214 ( .A(_abc_41234_new_n3005_), .Y(_abc_41234_new_n3006_));
INVX1 INVX1_215 ( .A(_abc_41234_new_n3014_), .Y(_abc_41234_new_n3015_));
INVX1 INVX1_216 ( .A(_abc_41234_new_n3018_), .Y(_abc_41234_new_n3019_));
INVX1 INVX1_217 ( .A(_abc_41234_new_n3030_), .Y(_abc_41234_new_n3031_));
INVX1 INVX1_218 ( .A(_abc_41234_new_n3036_), .Y(_abc_41234_new_n3037_));
INVX1 INVX1_219 ( .A(_abc_41234_new_n3055_), .Y(_abc_41234_new_n3056_));
INVX1 INVX1_22 ( .A(waitr), .Y(_abc_41234_new_n681_));
INVX1 INVX1_220 ( .A(_abc_41234_new_n3061_), .Y(_abc_41234_new_n3062_));
INVX1 INVX1_221 ( .A(_abc_41234_new_n3082_), .Y(_abc_41234_new_n3083_));
INVX1 INVX1_222 ( .A(_abc_41234_new_n3088_), .Y(_abc_41234_new_n3089_));
INVX1 INVX1_223 ( .A(_abc_41234_new_n3105_), .Y(_abc_41234_new_n3106_));
INVX1 INVX1_224 ( .A(_abc_41234_new_n3114_), .Y(_abc_41234_new_n3115_));
INVX1 INVX1_225 ( .A(_abc_41234_new_n3186_), .Y(_abc_41234_new_n3187_));
INVX1 INVX1_226 ( .A(_abc_41234_new_n1701_), .Y(_abc_41234_new_n3208_));
INVX1 INVX1_227 ( .A(raddrhold_11_), .Y(_abc_41234_new_n3225_));
INVX1 INVX1_228 ( .A(_abc_41234_new_n1737_), .Y(_abc_41234_new_n3228_));
INVX1 INVX1_229 ( .A(raddrhold_12_), .Y(_abc_41234_new_n3248_));
INVX1 INVX1_23 ( .A(_abc_41234_new_n689_), .Y(_abc_41234_new_n690_));
INVX1 INVX1_230 ( .A(_abc_41234_new_n1761_), .Y(_abc_41234_new_n3249_));
INVX1 INVX1_231 ( .A(_abc_41234_new_n1780_), .Y(_abc_41234_new_n3273_));
INVX1 INVX1_232 ( .A(_abc_41234_new_n3234_), .Y(_abc_41234_new_n3283_));
INVX1 INVX1_233 ( .A(raddrhold_15_), .Y(_abc_41234_new_n3316_));
INVX1 INVX1_234 ( .A(_abc_41234_new_n3347_), .Y(_abc_41234_new_n3366_));
INVX1 INVX1_235 ( .A(_abc_41234_new_n3373_), .Y(_abc_41234_new_n3374_));
INVX1 INVX1_236 ( .A(_abc_41234_new_n3415_), .Y(_abc_41234_new_n3416_));
INVX1 INVX1_237 ( .A(waddrhold_4_), .Y(_abc_41234_new_n3422_));
INVX1 INVX1_238 ( .A(_abc_41234_new_n3439_), .Y(_abc_41234_new_n3440_));
INVX1 INVX1_239 ( .A(_abc_41234_new_n3447_), .Y(_abc_41234_new_n3448_));
INVX1 INVX1_24 ( .A(state_5_), .Y(_abc_41234_new_n691_));
INVX1 INVX1_240 ( .A(waddrhold_6_), .Y(_abc_41234_new_n3466_));
INVX1 INVX1_241 ( .A(_abc_41234_new_n3481_), .Y(_abc_41234_new_n3482_));
INVX1 INVX1_242 ( .A(_abc_41234_new_n3520_), .Y(_abc_41234_new_n3521_));
INVX1 INVX1_243 ( .A(_abc_41234_new_n3528_), .Y(_abc_41234_new_n3529_));
INVX1 INVX1_244 ( .A(waddrhold_10_), .Y(_abc_41234_new_n3547_));
INVX1 INVX1_245 ( .A(_abc_41234_new_n3489_), .Y(_abc_41234_new_n3548_));
INVX1 INVX1_246 ( .A(_abc_41234_new_n3563_), .Y(_abc_41234_new_n3564_));
INVX1 INVX1_247 ( .A(waddrhold_11_), .Y(_abc_41234_new_n3569_));
INVX1 INVX1_248 ( .A(_abc_41234_new_n3585_), .Y(_abc_41234_new_n3586_));
INVX1 INVX1_249 ( .A(waddrhold_14_), .Y(_abc_41234_new_n3644_));
INVX1 INVX1_25 ( .A(_abc_41234_new_n695_), .Y(_abc_41234_new_n696_));
INVX1 INVX1_250 ( .A(_abc_41234_new_n3714_), .Y(_abc_41234_new_n3716_));
INVX1 INVX1_251 ( .A(_abc_41234_new_n1158_), .Y(_abc_41234_new_n3722_));
INVX1 INVX1_252 ( .A(_abc_41234_new_n1074_), .Y(_abc_41234_new_n3734_));
INVX1 INVX1_253 ( .A(_abc_41234_new_n1157_), .Y(_abc_41234_new_n3738_));
INVX1 INVX1_254 ( .A(_abc_41234_new_n3739_), .Y(_abc_41234_new_n3740_));
INVX1 INVX1_255 ( .A(_abc_41234_new_n1120_), .Y(_abc_41234_new_n3744_));
INVX1 INVX1_256 ( .A(_abc_41234_new_n1225_), .Y(_abc_41234_new_n3795_));
INVX1 INVX1_257 ( .A(_abc_41234_new_n1133_), .Y(_abc_41234_new_n3811_));
INVX1 INVX1_258 ( .A(_abc_41234_new_n3813_), .Y(_abc_41234_new_n3814_));
INVX1 INVX1_259 ( .A(_abc_41234_new_n1138_), .Y(_abc_41234_new_n3857_));
INVX1 INVX1_26 ( .A(_abc_41234_new_n700_), .Y(_abc_41234_new_n701_));
INVX1 INVX1_260 ( .A(_abc_41234_new_n1176_), .Y(_abc_41234_new_n3864_));
INVX1 INVX1_261 ( .A(_abc_41234_new_n1079_), .Y(_abc_41234_new_n3871_));
INVX1 INVX1_262 ( .A(_abc_41234_new_n1230_), .Y(_abc_41234_new_n3875_));
INVX1 INVX1_263 ( .A(_abc_41234_new_n1083_), .Y(_abc_41234_new_n3901_));
INVX1 INVX1_264 ( .A(_abc_41234_new_n522_), .Y(_abc_41234_new_n3959_));
INVX1 INVX1_265 ( .A(_abc_41234_new_n3995_), .Y(_abc_41234_new_n3996_));
INVX1 INVX1_266 ( .A(_abc_41234_new_n4013_), .Y(_abc_41234_new_n4014_));
INVX1 INVX1_267 ( .A(_abc_41234_new_n4039_), .Y(_abc_41234_new_n4040_));
INVX1 INVX1_268 ( .A(_abc_41234_new_n4041_), .Y(_abc_41234_new_n4042_));
INVX1 INVX1_269 ( .A(_abc_41234_new_n4069_), .Y(_abc_41234_new_n4070_));
INVX1 INVX1_27 ( .A(_abc_41234_new_n710_), .Y(_abc_41234_new_n711_));
INVX1 INVX1_270 ( .A(_abc_41234_new_n4101_), .Y(_abc_41234_new_n4102_));
INVX1 INVX1_271 ( .A(_abc_41234_new_n4126_), .Y(_abc_41234_new_n4127_));
INVX1 INVX1_272 ( .A(_abc_41234_new_n4174_), .Y(_abc_41234_new_n4175_));
INVX1 INVX1_273 ( .A(_abc_41234_new_n3638_), .Y(_abc_41234_new_n4213_));
INVX1 INVX1_274 ( .A(_abc_41234_new_n4224_), .Y(_abc_41234_new_n4225_));
INVX1 INVX1_275 ( .A(_abc_41234_new_n2940_), .Y(_abc_41234_new_n4277_));
INVX1 INVX1_276 ( .A(_abc_41234_new_n4274__bF_buf2), .Y(_abc_41234_new_n4383_));
INVX1 INVX1_277 ( .A(_abc_41234_new_n2833_), .Y(_abc_41234_new_n4388_));
INVX1 INVX1_278 ( .A(_abc_41234_new_n2884_), .Y(_abc_41234_new_n4430_));
INVX1 INVX1_279 ( .A(_abc_41234_new_n2889_), .Y(_abc_41234_new_n4436_));
INVX1 INVX1_28 ( .A(opcode_1_), .Y(_abc_41234_new_n721_));
INVX1 INVX1_280 ( .A(_abc_41234_new_n1653_), .Y(_abc_41234_new_n4448_));
INVX1 INVX1_281 ( .A(_abc_41234_new_n4480_), .Y(_abc_41234_new_n4481_));
INVX1 INVX1_282 ( .A(_abc_41234_new_n4499_), .Y(_abc_41234_new_n4500_));
INVX1 INVX1_283 ( .A(_abc_41234_new_n1470_), .Y(_abc_41234_new_n4527_));
INVX1 INVX1_284 ( .A(_abc_41234_new_n4543_), .Y(_abc_41234_new_n4544_));
INVX1 INVX1_285 ( .A(_abc_41234_new_n4537_), .Y(_abc_41234_new_n4555_));
INVX1 INVX1_286 ( .A(_abc_41234_new_n4564_), .Y(_abc_41234_new_n4565_));
INVX1 INVX1_287 ( .A(_abc_41234_new_n4600_), .Y(_abc_41234_new_n4601_));
INVX1 INVX1_288 ( .A(_auto_iopadmap_cc_368_execute_45628_0_), .Y(_abc_41234_new_n4611_));
INVX1 INVX1_289 ( .A(_auto_iopadmap_cc_368_execute_45628_1_), .Y(_abc_41234_new_n4620_));
INVX1 INVX1_29 ( .A(regfil_6__1_), .Y(_abc_41234_new_n725_));
INVX1 INVX1_290 ( .A(_auto_iopadmap_cc_368_execute_45628_2_), .Y(_abc_41234_new_n4625_));
INVX1 INVX1_291 ( .A(_auto_iopadmap_cc_368_execute_45628_3_), .Y(_abc_41234_new_n4630_));
INVX1 INVX1_292 ( .A(_auto_iopadmap_cc_368_execute_45628_4_), .Y(_abc_41234_new_n4635_));
INVX1 INVX1_293 ( .A(_auto_iopadmap_cc_368_execute_45628_5_), .Y(_abc_41234_new_n4640_));
INVX1 INVX1_294 ( .A(_auto_iopadmap_cc_368_execute_45628_6_), .Y(_abc_41234_new_n4645_));
INVX1 INVX1_295 ( .A(_auto_iopadmap_cc_368_execute_45628_7_), .Y(_abc_41234_new_n4650_));
INVX1 INVX1_296 ( .A(_auto_iopadmap_cc_368_execute_45628_8_), .Y(_abc_41234_new_n4655_));
INVX1 INVX1_297 ( .A(_auto_iopadmap_cc_368_execute_45628_9_), .Y(_abc_41234_new_n4659_));
INVX1 INVX1_298 ( .A(_auto_iopadmap_cc_368_execute_45628_10_), .Y(_abc_41234_new_n4666_));
INVX1 INVX1_299 ( .A(_auto_iopadmap_cc_368_execute_45628_11_), .Y(_abc_41234_new_n4671_));
INVX1 INVX1_3 ( .A(state_1_), .Y(_abc_41234_new_n505_));
INVX1 INVX1_30 ( .A(_abc_41234_new_n734_), .Y(_abc_41234_new_n735_));
INVX1 INVX1_300 ( .A(_auto_iopadmap_cc_368_execute_45628_12_), .Y(_abc_41234_new_n4676_));
INVX1 INVX1_301 ( .A(_auto_iopadmap_cc_368_execute_45628_13_), .Y(_abc_41234_new_n4680_));
INVX1 INVX1_302 ( .A(_auto_iopadmap_cc_368_execute_45628_14_), .Y(_abc_41234_new_n4684_));
INVX1 INVX1_303 ( .A(_auto_iopadmap_cc_368_execute_45628_15_), .Y(_abc_41234_new_n4689_));
INVX1 INVX1_304 ( .A(_auto_iopadmap_cc_368_execute_45645), .Y(_abc_41234_new_n4698_));
INVX1 INVX1_305 ( .A(_abc_41234_new_n2356_), .Y(_abc_41234_new_n4699_));
INVX1 INVX1_306 ( .A(statesel_5_), .Y(_abc_41234_new_n4719_));
INVX1 INVX1_307 ( .A(_abc_41234_new_n4725_), .Y(_abc_41234_new_n4726_));
INVX1 INVX1_308 ( .A(_abc_41234_new_n4729_), .Y(_abc_41234_new_n4730_));
INVX1 INVX1_309 ( .A(_abc_41234_new_n4761_), .Y(_abc_41234_new_n4762_));
INVX1 INVX1_31 ( .A(regfil_0__1_), .Y(_abc_41234_new_n739_));
INVX1 INVX1_310 ( .A(_abc_41234_new_n4727_), .Y(_abc_41234_new_n4767_));
INVX1 INVX1_311 ( .A(_abc_41234_new_n4720_), .Y(_abc_41234_new_n4778_));
INVX1 INVX1_312 ( .A(_abc_41234_new_n4802_), .Y(_abc_41234_new_n4803_));
INVX1 INVX1_313 ( .A(_abc_41234_new_n4814_), .Y(_abc_41234_new_n4815_));
INVX1 INVX1_314 ( .A(_abc_41234_new_n4760_), .Y(_abc_41234_new_n4821_));
INVX1 INVX1_315 ( .A(_abc_41234_new_n4789_), .Y(_abc_41234_new_n4822_));
INVX1 INVX1_316 ( .A(_abc_41234_new_n4704_), .Y(_abc_41234_new_n4831_));
INVX1 INVX1_317 ( .A(_abc_41234_new_n4830_), .Y(_abc_41234_new_n4840_));
INVX1 INVX1_318 ( .A(_abc_41234_new_n4768_), .Y(_abc_41234_new_n4845_));
INVX1 INVX1_319 ( .A(_abc_41234_new_n4846_), .Y(_abc_41234_new_n4847_));
INVX1 INVX1_32 ( .A(_abc_41234_new_n586_), .Y(_abc_41234_new_n740_));
INVX1 INVX1_320 ( .A(_abc_41234_new_n4799_), .Y(_abc_41234_new_n4866_));
INVX1 INVX1_321 ( .A(_abc_41234_new_n4829_), .Y(_abc_41234_new_n4869_));
INVX1 INVX1_322 ( .A(_abc_41234_new_n3677_), .Y(_abc_41234_new_n4873_));
INVX1 INVX1_323 ( .A(alu__abc_40887_new_n34_), .Y(alu__abc_40887_new_n35_));
INVX1 INVX1_324 ( .A(alu__abc_40887_new_n39_), .Y(alu__abc_40887_new_n40_));
INVX1 INVX1_325 ( .A(alu__abc_40887_new_n41_), .Y(alu__abc_40887_new_n42_));
INVX1 INVX1_326 ( .A(alu__abc_40887_new_n60_), .Y(alu__abc_40887_new_n61_));
INVX1 INVX1_327 ( .A(alu__abc_40887_new_n68_), .Y(alu__abc_40887_new_n69_));
INVX1 INVX1_328 ( .A(alu__abc_40887_new_n65_), .Y(alu__abc_40887_new_n72_));
INVX1 INVX1_329 ( .A(alu__abc_40887_new_n56_), .Y(alu__abc_40887_new_n76_));
INVX1 INVX1_33 ( .A(_abc_41234_new_n743_), .Y(_abc_41234_new_n744_));
INVX1 INVX1_330 ( .A(alu_sel_1_), .Y(alu__abc_40887_new_n102_));
INVX1 INVX1_331 ( .A(alu_sel_2_), .Y(alu__abc_40887_new_n115_));
INVX1 INVX1_332 ( .A(alu_sel_0_), .Y(alu__abc_40887_new_n116_));
INVX1 INVX1_333 ( .A(alu_opra_3_), .Y(alu__abc_40887_new_n119_));
INVX1 INVX1_334 ( .A(alu__abc_40887_new_n120_), .Y(alu__abc_40887_new_n121_));
INVX1 INVX1_335 ( .A(alu_oprb_2_), .Y(alu__abc_40887_new_n122_));
INVX1 INVX1_336 ( .A(alu_opra_1_), .Y(alu__abc_40887_new_n125_));
INVX1 INVX1_337 ( .A(alu__abc_40887_new_n133_), .Y(alu__abc_40887_new_n134_));
INVX1 INVX1_338 ( .A(alu_opra_5_), .Y(alu__abc_40887_new_n136_));
INVX1 INVX1_339 ( .A(alu_opra_4_), .Y(alu__abc_40887_new_n137_));
INVX1 INVX1_34 ( .A(_abc_41234_new_n682_), .Y(_abc_41234_new_n755_));
INVX1 INVX1_340 ( .A(alu__abc_40887_new_n140_), .Y(alu__abc_40887_new_n141_));
INVX1 INVX1_341 ( .A(alu_opra_6_), .Y(alu__abc_40887_new_n143_));
INVX1 INVX1_342 ( .A(alu__abc_40887_new_n123_), .Y(alu__abc_40887_new_n146_));
INVX1 INVX1_343 ( .A(alu_opra_2_), .Y(alu__abc_40887_new_n150_));
INVX1 INVX1_344 ( .A(alu__abc_40887_new_n144_), .Y(alu__abc_40887_new_n156_));
INVX1 INVX1_345 ( .A(alu_cin), .Y(alu__abc_40887_new_n167_));
INVX1 INVX1_346 ( .A(alu__abc_40887_new_n168_), .Y(alu__abc_40887_new_n169_));
INVX1 INVX1_347 ( .A(alu__abc_40887_new_n62_), .Y(alu__abc_40887_new_n178_));
INVX1 INVX1_348 ( .A(alu__abc_40887_new_n199_), .Y(alu__abc_40887_new_n200_));
INVX1 INVX1_349 ( .A(alu__abc_40887_new_n202_), .Y(alu__abc_40887_new_n203_));
INVX1 INVX1_35 ( .A(regfil_6__2_), .Y(_abc_41234_new_n775_));
INVX1 INVX1_350 ( .A(alu__abc_40887_new_n33_), .Y(alu__abc_40887_new_n207_));
INVX1 INVX1_351 ( .A(alu__abc_40887_new_n74_), .Y(alu__abc_40887_new_n217_));
INVX1 INVX1_352 ( .A(alu__abc_40887_new_n230_), .Y(alu__abc_40887_new_n231_));
INVX1 INVX1_353 ( .A(alu__abc_40887_new_n45_), .Y(alu__abc_40887_new_n234_));
INVX1 INVX1_354 ( .A(alu__abc_40887_new_n205_), .Y(alu__abc_40887_new_n243_));
INVX1 INVX1_355 ( .A(alu__abc_40887_new_n118_), .Y(alu__abc_40887_new_n270_));
INVX1 INVX1_356 ( .A(alu__abc_40887_new_n276_), .Y(alu__abc_40887_new_n277_));
INVX1 INVX1_357 ( .A(alu__abc_40887_new_n201_), .Y(alu__abc_40887_new_n314_));
INVX1 INVX1_358 ( .A(alu__abc_40887_new_n195_), .Y(alu__abc_40887_new_n322_));
INVX1 INVX1_359 ( .A(alu__abc_40887_new_n331_), .Y(alu__abc_40887_new_n334_));
INVX1 INVX1_36 ( .A(_abc_41234_new_n741_), .Y(_abc_41234_new_n783_));
INVX1 INVX1_360 ( .A(alu__abc_40887_new_n249_), .Y(alu__abc_40887_new_n350_));
INVX1 INVX1_361 ( .A(alu_opra_7_), .Y(alu__abc_40887_new_n367_));
INVX1 INVX1_362 ( .A(alu__abc_40887_new_n186_), .Y(alu__abc_40887_new_n370_));
INVX1 INVX1_363 ( .A(alu__abc_40887_new_n105_), .Y(alu__abc_40887_new_n375_));
INVX1 INVX1_37 ( .A(regfil_0__3_), .Y(_abc_41234_new_n805_));
INVX1 INVX1_38 ( .A(_abc_41234_new_n806_), .Y(_abc_41234_new_n807_));
INVX1 INVX1_39 ( .A(regfil_6__3_), .Y(_abc_41234_new_n822_));
INVX1 INVX1_4 ( .A(_abc_41234_new_n518_), .Y(_abc_41234_new_n519_));
INVX1 INVX1_40 ( .A(regfil_6__4_), .Y(_abc_41234_new_n852_));
INVX1 INVX1_41 ( .A(_abc_41234_new_n862_), .Y(_abc_41234_new_n863_));
INVX1 INVX1_42 ( .A(_abc_41234_new_n870_), .Y(_abc_41234_new_n871_));
INVX1 INVX1_43 ( .A(regfil_1__5_), .Y(_abc_41234_new_n896_));
INVX1 INVX1_44 ( .A(regfil_6__5_), .Y(_abc_41234_new_n907_));
INVX1 INVX1_45 ( .A(_abc_41234_new_n910_), .Y(_abc_41234_new_n911_));
INVX1 INVX1_46 ( .A(regfil_0__5_), .Y(_abc_41234_new_n914_));
INVX1 INVX1_47 ( .A(_abc_41234_new_n882_), .Y(_abc_41234_new_n930_));
INVX1 INVX1_48 ( .A(_abc_41234_new_n946_), .Y(_abc_41234_new_n947_));
INVX1 INVX1_49 ( .A(_abc_41234_new_n949_), .Y(_abc_41234_new_n950_));
INVX1 INVX1_5 ( .A(state_0_), .Y(_abc_41234_new_n520_));
INVX1 INVX1_50 ( .A(_abc_41234_new_n931_), .Y(_abc_41234_new_n968_));
INVX1 INVX1_51 ( .A(regfil_6__7_), .Y(_abc_41234_new_n999_));
INVX1 INVX1_52 ( .A(_abc_41234_new_n598_), .Y(_abc_41234_new_n1038_));
INVX1 INVX1_53 ( .A(_abc_41234_new_n1040__bF_buf4), .Y(_abc_41234_new_n1041_));
INVX1 INVX1_54 ( .A(_abc_41234_new_n1052_), .Y(_abc_41234_new_n1053_));
INVX1 INVX1_55 ( .A(_abc_41234_new_n646_), .Y(_abc_41234_new_n1056_));
INVX1 INVX1_56 ( .A(_abc_41234_new_n1068_), .Y(_abc_41234_new_n1069_));
INVX1 INVX1_57 ( .A(_abc_41234_new_n1113_), .Y(_abc_41234_new_n1114_));
INVX1 INVX1_58 ( .A(_abc_41234_new_n1146_), .Y(_abc_41234_new_n1147_));
INVX1 INVX1_59 ( .A(_abc_41234_new_n1148_), .Y(_abc_41234_new_n1149_));
INVX1 INVX1_6 ( .A(_abc_41234_new_n540_), .Y(_abc_41234_new_n541_));
INVX1 INVX1_60 ( .A(_abc_41234_new_n530_), .Y(_abc_41234_new_n1150_));
INVX1 INVX1_61 ( .A(_abc_41234_new_n1155_), .Y(_abc_41234_new_n1156_));
INVX1 INVX1_62 ( .A(_abc_41234_new_n1162_), .Y(_abc_41234_new_n1168_));
INVX1 INVX1_63 ( .A(_abc_41234_new_n1192_), .Y(_abc_41234_new_n1193_));
INVX1 INVX1_64 ( .A(_abc_41234_new_n1197_), .Y(_abc_41234_new_n1198_));
INVX1 INVX1_65 ( .A(_abc_41234_new_n1210_), .Y(_abc_41234_new_n1211_));
INVX1 INVX1_66 ( .A(_abc_41234_new_n1214_), .Y(_abc_41234_new_n1215_));
INVX1 INVX1_67 ( .A(_abc_41234_new_n1195_), .Y(_abc_41234_new_n1274_));
INVX1 INVX1_68 ( .A(_abc_41234_new_n1299_), .Y(_abc_41234_new_n1300_));
INVX1 INVX1_69 ( .A(_abc_41234_new_n1051_), .Y(_abc_41234_new_n1305_));
INVX1 INVX1_7 ( .A(_abc_41234_new_n542_), .Y(_abc_41234_new_n543_));
INVX1 INVX1_70 ( .A(_abc_41234_new_n1306_), .Y(_abc_41234_new_n1307_));
INVX1 INVX1_71 ( .A(_abc_41234_new_n1316_), .Y(_abc_41234_new_n1317_));
INVX1 INVX1_72 ( .A(_abc_41234_new_n1272_), .Y(_abc_41234_new_n1326_));
INVX1 INVX1_73 ( .A(_abc_41234_new_n1327_), .Y(_abc_41234_new_n1328_));
INVX1 INVX1_74 ( .A(_abc_41234_new_n1331_), .Y(_abc_41234_new_n1332_));
INVX1 INVX1_75 ( .A(_abc_41234_new_n1349_), .Y(_abc_41234_new_n1350_));
INVX1 INVX1_76 ( .A(_abc_41234_new_n1376_), .Y(_abc_41234_new_n1377_));
INVX1 INVX1_77 ( .A(_abc_41234_new_n879_), .Y(_abc_41234_new_n1386_));
INVX1 INVX1_78 ( .A(_abc_41234_new_n1391_), .Y(_abc_41234_new_n1392_));
INVX1 INVX1_79 ( .A(_abc_41234_new_n1425_), .Y(_abc_41234_new_n1426_));
INVX1 INVX1_8 ( .A(_abc_41234_new_n552_), .Y(_abc_41234_new_n553_));
INVX1 INVX1_80 ( .A(_abc_41234_new_n1333_), .Y(_abc_41234_new_n1429_));
INVX1 INVX1_81 ( .A(_abc_41234_new_n1457_), .Y(_abc_41234_new_n1458_));
INVX1 INVX1_82 ( .A(_abc_41234_new_n1459_), .Y(_abc_41234_new_n1461_));
INVX1 INVX1_83 ( .A(_abc_41234_new_n1462_), .Y(_abc_41234_new_n1463_));
INVX1 INVX1_84 ( .A(_abc_41234_new_n1472_), .Y(_abc_41234_new_n1473_));
INVX1 INVX1_85 ( .A(_abc_41234_new_n1477_), .Y(_abc_41234_new_n1478_));
INVX1 INVX1_86 ( .A(_abc_41234_new_n1420_), .Y(_abc_41234_new_n1482_));
INVX1 INVX1_87 ( .A(_abc_41234_new_n1498_), .Y(_abc_41234_new_n1499_));
INVX1 INVX1_88 ( .A(_abc_41234_new_n1527_), .Y(_abc_41234_new_n1528_));
INVX1 INVX1_89 ( .A(_abc_41234_new_n1497_), .Y(_abc_41234_new_n1531_));
INVX1 INVX1_9 ( .A(_abc_41234_new_n577_), .Y(_abc_41234_new_n578_));
INVX1 INVX1_90 ( .A(_abc_41234_new_n1537_), .Y(_abc_41234_new_n1538_));
INVX1 INVX1_91 ( .A(_abc_41234_new_n1542_), .Y(_abc_41234_new_n1543_));
INVX1 INVX1_92 ( .A(_abc_41234_new_n1547_), .Y(_abc_41234_new_n1550_));
INVX1 INVX1_93 ( .A(_abc_41234_new_n1010_), .Y(_abc_41234_new_n1558_));
INVX1 INVX1_94 ( .A(_abc_41234_new_n1525_), .Y(_abc_41234_new_n1566_));
INVX1 INVX1_95 ( .A(_abc_41234_new_n1578_), .Y(_abc_41234_new_n1579_));
INVX1 INVX1_96 ( .A(_abc_41234_new_n1580_), .Y(_abc_41234_new_n1581_));
INVX1 INVX1_97 ( .A(_abc_41234_new_n1536_), .Y(_abc_41234_new_n1587_));
INVX1 INVX1_98 ( .A(_abc_41234_new_n1591_), .Y(_abc_41234_new_n1592_));
INVX1 INVX1_99 ( .A(wdatahold2_0_), .Y(_abc_41234_new_n1605_));
INVX2 INVX2_1 ( .A(regfil_7__1_), .Y(_abc_41234_new_n514_));
INVX2 INVX2_10 ( .A(_abc_41234_new_n583_), .Y(_abc_41234_new_n584_));
INVX2 INVX2_100 ( .A(_abc_41234_new_n2976_), .Y(_abc_41234_new_n2977_));
INVX2 INVX2_101 ( .A(_abc_41234_new_n2735_), .Y(_abc_41234_new_n2995_));
INVX2 INVX2_102 ( .A(raddrhold_2_), .Y(_abc_41234_new_n3003_));
INVX2 INVX2_103 ( .A(raddrhold_3_), .Y(_abc_41234_new_n3023_));
INVX2 INVX2_104 ( .A(raddrhold_4_), .Y(_abc_41234_new_n3049_));
INVX2 INVX2_105 ( .A(raddrhold_5_), .Y(_abc_41234_new_n3074_));
INVX2 INVX2_106 ( .A(raddrhold_8_), .Y(_abc_41234_new_n3151_));
INVX2 INVX2_107 ( .A(raddrhold_9_), .Y(_abc_41234_new_n3175_));
INVX2 INVX2_108 ( .A(raddrhold_10_), .Y(_abc_41234_new_n3200_));
INVX2 INVX2_109 ( .A(raddrhold_13_), .Y(_abc_41234_new_n3272_));
INVX2 INVX2_11 ( .A(regfil_0__0_), .Y(_abc_41234_new_n585_));
INVX2 INVX2_110 ( .A(sp_13_), .Y(_abc_41234_new_n3279_));
INVX2 INVX2_111 ( .A(raddrhold_14_), .Y(_abc_41234_new_n3294_));
INVX2 INVX2_112 ( .A(waddrhold_0_), .Y(_abc_41234_new_n3337_));
INVX2 INVX2_113 ( .A(waddrhold_1_), .Y(_abc_41234_new_n3358_));
INVX2 INVX2_114 ( .A(waddrhold_2_), .Y(_abc_41234_new_n3381_));
INVX2 INVX2_115 ( .A(_abc_41234_new_n3384_), .Y(_abc_41234_new_n3385_));
INVX2 INVX2_116 ( .A(waddrhold_3_), .Y(_abc_41234_new_n3403_));
INVX2 INVX2_117 ( .A(_abc_41234_new_n3424_), .Y(_abc_41234_new_n3425_));
INVX2 INVX2_118 ( .A(waddrhold_5_), .Y(_abc_41234_new_n3445_));
INVX2 INVX2_119 ( .A(waddrhold_7_), .Y(_abc_41234_new_n3487_));
INVX2 INVX2_12 ( .A(_abc_41234_new_n608_), .Y(_abc_41234_new_n609_));
INVX2 INVX2_120 ( .A(waddrhold_8_), .Y(_abc_41234_new_n3507_));
INVX2 INVX2_121 ( .A(waddrhold_9_), .Y(_abc_41234_new_n3526_));
INVX2 INVX2_122 ( .A(waddrhold_12_), .Y(_abc_41234_new_n3605_));
INVX2 INVX2_123 ( .A(_abc_41234_new_n3609_), .Y(_abc_41234_new_n3610_));
INVX2 INVX2_124 ( .A(waddrhold_13_), .Y(_abc_41234_new_n3624_));
INVX2 INVX2_125 ( .A(waddrhold_15_), .Y(_abc_41234_new_n3661_));
INVX2 INVX2_126 ( .A(_abc_41234_new_n2489_), .Y(_abc_41234_new_n3697_));
INVX2 INVX2_127 ( .A(_abc_41234_new_n1124_), .Y(_abc_41234_new_n3810_));
INVX2 INVX2_128 ( .A(_abc_41234_new_n3960_), .Y(_abc_41234_new_n3961_));
INVX2 INVX2_129 ( .A(_abc_41234_new_n3923_), .Y(_abc_41234_new_n3964_));
INVX2 INVX2_13 ( .A(_abc_41234_new_n611_), .Y(_abc_41234_new_n612_));
INVX2 INVX2_130 ( .A(_abc_41234_new_n4079_), .Y(_abc_41234_new_n4080_));
INVX2 INVX2_131 ( .A(_abc_41234_new_n4309_), .Y(_abc_41234_new_n4329_));
INVX2 INVX2_132 ( .A(_abc_41234_new_n4660_), .Y(_abc_41234_new_n4661_));
INVX2 INVX2_133 ( .A(_abc_41234_new_n2557_), .Y(_abc_41234_new_n4708_));
INVX2 INVX2_134 ( .A(_abc_41234_new_n4709_), .Y(_abc_41234_new_n4710_));
INVX2 INVX2_135 ( .A(_abc_41234_new_n2558_), .Y(_abc_41234_new_n4712_));
INVX2 INVX2_136 ( .A(_abc_41234_new_n4713_), .Y(_abc_41234_new_n4714_));
INVX2 INVX2_137 ( .A(_abc_41234_new_n4715_), .Y(_abc_41234_new_n4716_));
INVX2 INVX2_138 ( .A(alu__abc_40887_new_n36_), .Y(alu__abc_40887_new_n37_));
INVX2 INVX2_139 ( .A(alu_opra_0_), .Y(alu__abc_40887_new_n128_));
INVX2 INVX2_14 ( .A(opcode_0_), .Y(_abc_41234_new_n616_));
INVX2 INVX2_140 ( .A(alu__abc_40887_new_n208_), .Y(alu__abc_40887_new_n209_));
INVX2 INVX2_141 ( .A(alu__abc_40887_new_n210_), .Y(alu__abc_40887_new_n227_));
INVX2 INVX2_142 ( .A(alu__abc_40887_new_n104_), .Y(alu__abc_40887_new_n241_));
INVX2 INVX2_143 ( .A(alu__abc_40887_new_n166_), .Y(alu__abc_40887_new_n271_));
INVX2 INVX2_15 ( .A(_abc_41234_new_n620__bF_buf5), .Y(_abc_41234_new_n621_));
INVX2 INVX2_16 ( .A(_abc_41234_new_n596_), .Y(_abc_41234_new_n632_));
INVX2 INVX2_17 ( .A(regfil_1__2_), .Y(_abc_41234_new_n634_));
INVX2 INVX2_18 ( .A(regfil_1__6_), .Y(_abc_41234_new_n638_));
INVX2 INVX2_19 ( .A(opcode_6_), .Y(_abc_41234_new_n661_));
INVX2 INVX2_2 ( .A(_abc_41234_new_n523__bF_buf4), .Y(_abc_41234_new_n524_));
INVX2 INVX2_20 ( .A(regfil_7__0_), .Y(_abc_41234_new_n680_));
INVX2 INVX2_21 ( .A(_abc_41234_new_n533_), .Y(_abc_41234_new_n688_));
INVX2 INVX2_22 ( .A(_abc_41234_new_n692_), .Y(_abc_41234_new_n693_));
INVX2 INVX2_23 ( .A(_abc_41234_new_n697_), .Y(_abc_41234_new_n698_));
INVX2 INVX2_24 ( .A(_abc_41234_new_n702_), .Y(_abc_41234_new_n703_));
INVX2 INVX2_25 ( .A(\data[0] ), .Y(_abc_41234_new_n714_));
INVX2 INVX2_26 ( .A(rdatahold_1_), .Y(_abc_41234_new_n718_));
INVX2 INVX2_27 ( .A(regfil_3__1_), .Y(_abc_41234_new_n730_));
INVX2 INVX2_28 ( .A(regfil_0__2_), .Y(_abc_41234_new_n766_));
INVX2 INVX2_29 ( .A(_abc_41234_new_n790_), .Y(_abc_41234_new_n791_));
INVX2 INVX2_3 ( .A(_abc_41234_new_n538_), .Y(_abc_41234_new_n539_));
INVX2 INVX2_30 ( .A(rdatahold_2_), .Y(_abc_41234_new_n794_));
INVX2 INVX2_31 ( .A(regfil_5__3_bF_buf3_), .Y(_abc_41234_new_n818_));
INVX2 INVX2_32 ( .A(rdatahold_3_), .Y(_abc_41234_new_n832_));
INVX2 INVX2_33 ( .A(_abc_41234_new_n559_), .Y(_abc_41234_new_n839_));
INVX2 INVX2_34 ( .A(regfil_7__4_), .Y(_abc_41234_new_n851_));
INVX2 INVX2_35 ( .A(regfil_1__4_), .Y(_abc_41234_new_n855_));
INVX2 INVX2_36 ( .A(regfil_2__4_), .Y(_abc_41234_new_n859_));
INVX2 INVX2_37 ( .A(regfil_0__4_), .Y(_abc_41234_new_n866_));
INVX2 INVX2_38 ( .A(\data[4] ), .Y(_abc_41234_new_n890_));
INVX2 INVX2_39 ( .A(regfil_2__5_), .Y(_abc_41234_new_n900_));
INVX2 INVX2_4 ( .A(_abc_41234_new_n526__bF_buf2), .Y(_abc_41234_new_n545_));
INVX2 INVX2_40 ( .A(regfil_0__6_), .Y(_abc_41234_new_n944_));
INVX2 INVX2_41 ( .A(regfil_7__6_), .Y(_abc_41234_new_n967_));
INVX2 INVX2_42 ( .A(regfil_0__7_), .Y(_abc_41234_new_n983_));
INVX2 INVX2_43 ( .A(regfil_3__7_), .Y(_abc_41234_new_n992_));
INVX2 INVX2_44 ( .A(regfil_2__7_), .Y(_abc_41234_new_n993_));
INVX2 INVX2_45 ( .A(rdatahold_7_), .Y(_abc_41234_new_n1005_));
INVX2 INVX2_46 ( .A(carry), .Y(_abc_41234_new_n1013_));
INVX2 INVX2_47 ( .A(\data[7] ), .Y(_abc_41234_new_n1016_));
INVX2 INVX2_48 ( .A(_abc_41234_new_n1042_), .Y(_abc_41234_new_n1043_));
INVX2 INVX2_49 ( .A(_abc_41234_new_n1037_), .Y(_abc_41234_new_n1044_));
INVX2 INVX2_5 ( .A(regfil_7__7_), .Y(_abc_41234_new_n560_));
INVX2 INVX2_50 ( .A(opcode_7_), .Y(_abc_41234_new_n1045_));
INVX2 INVX2_51 ( .A(_abc_41234_new_n1108_), .Y(_abc_41234_new_n1109_));
INVX2 INVX2_52 ( .A(regfil_2__0_), .Y(_abc_41234_new_n1143_));
INVX2 INVX2_53 ( .A(_abc_41234_new_n1151_), .Y(_abc_41234_new_n1152_));
INVX2 INVX2_54 ( .A(_abc_41234_new_n1199_), .Y(_abc_41234_new_n1200_));
INVX2 INVX2_55 ( .A(_abc_41234_new_n1039_), .Y(_abc_41234_new_n1217_));
INVX2 INVX2_56 ( .A(_abc_41234_new_n1223_), .Y(_abc_41234_new_n1224_));
INVX2 INVX2_57 ( .A(_abc_41234_new_n1308_), .Y(_abc_41234_new_n1309_));
INVX2 INVX2_58 ( .A(_abc_41234_new_n1324_), .Y(_abc_41234_new_n1325_));
INVX2 INVX2_59 ( .A(_abc_41234_new_n1055_), .Y(_abc_41234_new_n1344_));
INVX2 INVX2_6 ( .A(rdatahold_0_), .Y(_abc_41234_new_n565_));
INVX2 INVX2_60 ( .A(sp_14_), .Y(_abc_41234_new_n1524_));
INVX2 INVX2_61 ( .A(regfil_2__6_), .Y(_abc_41234_new_n1535_));
INVX2 INVX2_62 ( .A(_abc_41234_new_n1303_), .Y(_abc_41234_new_n1575_));
INVX2 INVX2_63 ( .A(pc_3_), .Y(_abc_41234_new_n1613_));
INVX2 INVX2_64 ( .A(pc_2_), .Y(_abc_41234_new_n1614_));
INVX2 INVX2_65 ( .A(_abc_41234_new_n1639__bF_buf3), .Y(_abc_41234_new_n1640_));
INVX2 INVX2_66 ( .A(pc_0_), .Y(_abc_41234_new_n1647_));
INVX2 INVX2_67 ( .A(pc_12_), .Y(_abc_41234_new_n1750_));
INVX2 INVX2_68 ( .A(pc_15_), .Y(_abc_41234_new_n1828_));
INVX2 INVX2_69 ( .A(regfil_3__0_), .Y(_abc_41234_new_n1848_));
INVX2 INVX2_7 ( .A(regfil_1__3_), .Y(_abc_41234_new_n568_));
INVX2 INVX2_70 ( .A(_abc_41234_new_n1849_), .Y(_abc_41234_new_n1850_));
INVX2 INVX2_71 ( .A(popdes_1_), .Y(_abc_41234_new_n1851_));
INVX2 INVX2_72 ( .A(_abc_41234_new_n1873_), .Y(_abc_41234_new_n1874_));
INVX2 INVX2_73 ( .A(popdes_0_), .Y(_abc_41234_new_n1878_));
INVX2 INVX2_74 ( .A(_abc_41234_new_n1875_), .Y(_abc_41234_new_n1887_));
INVX2 INVX2_75 ( .A(regfil_3__6_), .Y(_abc_41234_new_n1936_));
INVX2 INVX2_76 ( .A(_abc_41234_new_n573_), .Y(_abc_41234_new_n1995_));
INVX2 INVX2_77 ( .A(_abc_41234_new_n2247_), .Y(_abc_41234_new_n2342_));
INVX2 INVX2_78 ( .A(_abc_41234_new_n517_), .Y(_abc_41234_new_n2353_));
INVX2 INVX2_79 ( .A(rdatahold2_6_), .Y(_abc_41234_new_n2371_));
INVX2 INVX2_8 ( .A(regfil_1__0_), .Y(_abc_41234_new_n569_));
INVX2 INVX2_80 ( .A(sign), .Y(_abc_41234_new_n2376_));
INVX2 INVX2_81 ( .A(rdatahold2_0_), .Y(_abc_41234_new_n2421_));
INVX2 INVX2_82 ( .A(statesel_0_), .Y(_abc_41234_new_n2455_));
INVX2 INVX2_83 ( .A(statesel_2_), .Y(_abc_41234_new_n2581_));
INVX2 INVX2_84 ( .A(_abc_41234_new_n2578_), .Y(_abc_41234_new_n2582_));
INVX2 INVX2_85 ( .A(statesel_3_), .Y(_abc_41234_new_n2588_));
INVX2 INVX2_86 ( .A(_abc_41234_new_n2603_), .Y(_abc_41234_new_n2604_));
INVX2 INVX2_87 ( .A(statesel_4_), .Y(_abc_41234_new_n2611_));
INVX2 INVX2_88 ( .A(_abc_41234_new_n2620_), .Y(_abc_41234_new_n2621_));
INVX2 INVX2_89 ( .A(rdatahold2_3_), .Y(_abc_41234_new_n2654_));
INVX2 INVX2_9 ( .A(_abc_41234_new_n579_), .Y(_abc_41234_new_n580_));
INVX2 INVX2_90 ( .A(rdatahold2_4_), .Y(_abc_41234_new_n2656_));
INVX2 INVX2_91 ( .A(_abc_41234_new_n2706_), .Y(_abc_41234_new_n2707_));
INVX2 INVX2_92 ( .A(_abc_41234_new_n2773_), .Y(_abc_41234_new_n2774_));
INVX2 INVX2_93 ( .A(_abc_41234_new_n2801_), .Y(_abc_41234_new_n2802_));
INVX2 INVX2_94 ( .A(_abc_41234_new_n2804_), .Y(_abc_41234_new_n2805_));
INVX2 INVX2_95 ( .A(pc_6_), .Y(_abc_41234_new_n2865_));
INVX2 INVX2_96 ( .A(pc_7_), .Y(_abc_41234_new_n2882_));
INVX2 INVX2_97 ( .A(raddrhold_0_), .Y(_abc_41234_new_n2910_));
INVX2 INVX2_98 ( .A(_abc_41234_new_n2915_), .Y(_abc_41234_new_n2916_));
INVX2 INVX2_99 ( .A(raddrhold_1_), .Y(_abc_41234_new_n2965_));
INVX4 INVX4_1 ( .A(_abc_41234_new_n508_), .Y(_abc_41234_new_n509_));
INVX4 INVX4_10 ( .A(regfil_2__1_), .Y(_abc_41234_new_n731_));
INVX4 INVX4_11 ( .A(regfil_7__2_), .Y(_abc_41234_new_n751_));
INVX4 INVX4_12 ( .A(_abc_41234_new_n756_), .Y(_abc_41234_new_n757_));
INVX4 INVX4_13 ( .A(regfil_3__2_), .Y(_abc_41234_new_n768_));
INVX4 INVX4_14 ( .A(regfil_2__2_), .Y(_abc_41234_new_n769_));
INVX4 INVX4_15 ( .A(regfil_5__2_), .Y(_abc_41234_new_n772_));
INVX4 INVX4_16 ( .A(regfil_4__2_bF_buf3_), .Y(_abc_41234_new_n773_));
INVX4 INVX4_17 ( .A(regfil_3__3_), .Y(_abc_41234_new_n814_));
INVX4 INVX4_18 ( .A(regfil_2__3_), .Y(_abc_41234_new_n815_));
INVX4 INVX4_19 ( .A(regfil_7__3_), .Y(_abc_41234_new_n821_));
INVX4 INVX4_2 ( .A(_abc_41234_new_n512_), .Y(_abc_41234_new_n513_));
INVX4 INVX4_20 ( .A(rdatahold_4_), .Y(_abc_41234_new_n847_));
INVX4 INVX4_21 ( .A(regfil_5__4_), .Y(_abc_41234_new_n848_));
INVX4 INVX4_22 ( .A(regfil_4__4_), .Y(_abc_41234_new_n849_));
INVX4 INVX4_23 ( .A(regfil_3__4_), .Y(_abc_41234_new_n858_));
INVX4 INVX4_24 ( .A(rdatahold_5_), .Y(_abc_41234_new_n895_));
INVX4 INVX4_25 ( .A(regfil_3__5_), .Y(_abc_41234_new_n899_));
INVX4 INVX4_26 ( .A(regfil_5__5_), .Y(_abc_41234_new_n903_));
INVX4 INVX4_27 ( .A(regfil_4__5_), .Y(_abc_41234_new_n904_));
INVX4 INVX4_28 ( .A(regfil_7__5_), .Y(_abc_41234_new_n906_));
INVX4 INVX4_29 ( .A(rdatahold_6_), .Y(_abc_41234_new_n940_));
INVX4 INVX4_3 ( .A(regfil_1__1_), .Y(_abc_41234_new_n570_));
INVX4 INVX4_30 ( .A(regfil_5__7_), .Y(_abc_41234_new_n996_));
INVX4 INVX4_31 ( .A(regfil_4__7_), .Y(_abc_41234_new_n997_));
INVX4 INVX4_32 ( .A(_abc_41234_new_n1035_), .Y(_abc_41234_new_n1036_));
INVX4 INVX4_33 ( .A(_abc_41234_new_n1060_), .Y(_abc_41234_new_n1061_));
INVX4 INVX4_34 ( .A(sp_3_), .Y(_abc_41234_new_n1067_));
INVX4 INVX4_35 ( .A(sp_2_), .Y(_abc_41234_new_n1071_));
INVX4 INVX4_36 ( .A(sp_7_), .Y(_abc_41234_new_n1080_));
INVX4 INVX4_37 ( .A(regfil_5__6_bF_buf2_), .Y(_abc_41234_new_n1084_));
INVX4 INVX4_38 ( .A(sp_6_), .Y(_abc_41234_new_n1085_));
INVX4 INVX4_39 ( .A(sp_4_), .Y(_abc_41234_new_n1090_));
INVX4 INVX4_4 ( .A(_abc_41234_new_n502_), .Y(_abc_41234_new_n607_));
INVX4 INVX4_40 ( .A(sp_5_), .Y(_abc_41234_new_n1094_));
INVX4 INVX4_41 ( .A(_abc_41234_new_n1106_), .Y(_abc_41234_new_n1107_));
INVX4 INVX4_42 ( .A(_abc_41234_new_n1218_), .Y(_abc_41234_new_n1219_));
INVX4 INVX4_43 ( .A(regfil_5__0_), .Y(_abc_41234_new_n1221_));
INVX4 INVX4_44 ( .A(sp_9_), .Y(_abc_41234_new_n1251_));
INVX4 INVX4_45 ( .A(sp_8_), .Y(_abc_41234_new_n1255_));
INVX4 INVX4_46 ( .A(_abc_41234_new_n1206_), .Y(_abc_41234_new_n1263_));
INVX4 INVX4_47 ( .A(_abc_41234_new_n531_), .Y(_abc_41234_new_n1322_));
INVX4 INVX4_48 ( .A(sp_10_), .Y(_abc_41234_new_n1358_));
INVX4 INVX4_49 ( .A(sp_11_), .Y(_abc_41234_new_n1362_));
INVX4 INVX4_5 ( .A(_abc_41234_new_n662_), .Y(_abc_41234_new_n663_));
INVX4 INVX4_50 ( .A(sp_12_), .Y(_abc_41234_new_n1408_));
INVX4 INVX4_51 ( .A(regfil_4__6_), .Y(_abc_41234_new_n1509_));
INVX4 INVX4_52 ( .A(sp_15_), .Y(_abc_41234_new_n1569_));
INVX4 INVX4_53 ( .A(pc_8_), .Y(_abc_41234_new_n1622_));
INVX4 INVX4_54 ( .A(_abc_41234_new_n1630_), .Y(_abc_41234_new_n1631_));
INVX4 INVX4_55 ( .A(pc_1_), .Y(_abc_41234_new_n1646_));
INVX4 INVX4_56 ( .A(pc_9_), .Y(_abc_41234_new_n1670_));
INVX4 INVX4_57 ( .A(_abc_41234_new_n1105__bF_buf1), .Y(_abc_41234_new_n1684_));
INVX4 INVX4_58 ( .A(pc_10_), .Y(_abc_41234_new_n1705_));
INVX4 INVX4_59 ( .A(pc_11_), .Y(_abc_41234_new_n1727_));
INVX4 INVX4_6 ( .A(_abc_41234_new_n678_), .Y(_abc_41234_new_n679_));
INVX4 INVX4_60 ( .A(intcyc_bF_buf1), .Y(_abc_41234_new_n1729_));
INVX4 INVX4_61 ( .A(pc_13_), .Y(_abc_41234_new_n1775_));
INVX4 INVX4_62 ( .A(pc_14_), .Y(_abc_41234_new_n1798_));
INVX4 INVX4_63 ( .A(_abc_41234_new_n2181_), .Y(_abc_41234_new_n2201_));
INVX4 INVX4_64 ( .A(_abc_41234_new_n2248_), .Y(_abc_41234_new_n2253_));
INVX4 INVX4_65 ( .A(_abc_41234_new_n2245_), .Y(_abc_41234_new_n2255_));
INVX4 INVX4_66 ( .A(_abc_41234_new_n2451_), .Y(_abc_41234_new_n2452_));
INVX4 INVX4_67 ( .A(_abc_41234_new_n2462_), .Y(_abc_41234_new_n2488_));
INVX4 INVX4_68 ( .A(_abc_41234_new_n2504_), .Y(_abc_41234_new_n2505_));
INVX4 INVX4_69 ( .A(_abc_41234_new_n2534_), .Y(_abc_41234_new_n2535_));
INVX4 INVX4_7 ( .A(regfil_5__1_), .Y(_abc_41234_new_n719_));
INVX4 INVX4_70 ( .A(pc_4_), .Y(_abc_41234_new_n2806_));
INVX4 INVX4_71 ( .A(_abc_41234_new_n2917_), .Y(_abc_41234_new_n2918_));
INVX4 INVX4_72 ( .A(_abc_41234_new_n2919__bF_buf3), .Y(_abc_41234_new_n2920_));
INVX4 INVX4_73 ( .A(_abc_41234_new_n2951__bF_buf2), .Y(_abc_41234_new_n2953_));
INVX4 INVX4_74 ( .A(sp_1_), .Y(_abc_41234_new_n2973_));
INVX4 INVX4_75 ( .A(_abc_41234_new_n2467_), .Y(_abc_41234_new_n2996_));
INVX4 INVX4_76 ( .A(raddrhold_6_), .Y(_abc_41234_new_n3101_));
INVX4 INVX4_77 ( .A(raddrhold_7_), .Y(_abc_41234_new_n3125_));
INVX4 INVX4_78 ( .A(_abc_41234_new_n3338_), .Y(_abc_41234_new_n3339_));
INVX4 INVX4_79 ( .A(_abc_41234_new_n2519_), .Y(_abc_41234_new_n3353_));
INVX4 INVX4_8 ( .A(regfil_4__1_bF_buf3_), .Y(_abc_41234_new_n720_));
INVX4 INVX4_80 ( .A(_abc_41234_new_n3916_), .Y(_abc_41234_new_n3917_));
INVX4 INVX4_81 ( .A(_abc_41234_new_n3935_), .Y(_abc_41234_new_n3936_));
INVX4 INVX4_82 ( .A(_abc_41234_new_n3962_), .Y(_abc_41234_new_n3963_));
INVX4 INVX4_83 ( .A(_abc_41234_new_n2564_), .Y(_abc_41234_new_n4301_));
INVX4 INVX4_84 ( .A(_abc_41234_new_n4297__bF_buf2), .Y(_abc_41234_new_n4322_));
INVX4 INVX4_85 ( .A(_abc_41234_new_n4312_), .Y(_abc_41234_new_n4326_));
INVX4 INVX4_86 ( .A(_abc_41234_new_n4308_), .Y(_abc_41234_new_n4328_));
INVX4 INVX4_87 ( .A(_abc_41234_new_n2358_), .Y(_abc_41234_new_n4605_));
INVX4 INVX4_9 ( .A(_abc_41234_new_n618_), .Y(_abc_41234_new_n723_));
INVX8 INVX8_1 ( .A(reset_bF_buf8), .Y(_abc_41234_new_n516_));
INVX8 INVX8_10 ( .A(_abc_41234_new_n1046__bF_buf7), .Y(_abc_41234_new_n1047_));
INVX8 INVX8_11 ( .A(_abc_41234_new_n1049__bF_buf2), .Y(_abc_41234_new_n1066_));
INVX8 INVX8_12 ( .A(regfil_4__0_), .Y(_abc_41234_new_n1144_));
INVX8 INVX8_13 ( .A(_abc_41234_new_n1608_), .Y(_abc_41234_new_n1610_));
INVX8 INVX8_14 ( .A(_abc_41234_new_n1626_), .Y(_abc_41234_new_n1627_));
INVX8 INVX8_15 ( .A(_abc_41234_new_n1643__bF_buf5), .Y(_abc_41234_new_n1644_));
INVX8 INVX8_16 ( .A(_abc_41234_new_n665__bF_buf1), .Y(_abc_41234_new_n2185_));
INVX8 INVX8_17 ( .A(_abc_41234_new_n2189__bF_buf5), .Y(_abc_41234_new_n2190_));
INVX8 INVX8_18 ( .A(_abc_41234_new_n2174_), .Y(_abc_41234_new_n2207_));
INVX8 INVX8_19 ( .A(_abc_41234_new_n660__bF_buf1), .Y(_abc_41234_new_n2415_));
INVX8 INVX8_2 ( .A(opcode_4_bF_buf6_), .Y(_abc_41234_new_n529_));
INVX8 INVX8_20 ( .A(_abc_41234_new_n2497_), .Y(_abc_41234_new_n2498_));
INVX8 INVX8_21 ( .A(_abc_41234_new_n2694_), .Y(_abc_41234_new_n2695_));
INVX8 INVX8_22 ( .A(_abc_41234_new_n2671_), .Y(_abc_41234_new_n2696_));
INVX8 INVX8_23 ( .A(_abc_41234_new_n2913_), .Y(_abc_41234_new_n2914_));
INVX8 INVX8_24 ( .A(sp_0_bF_buf2_), .Y(_abc_41234_new_n2947_));
INVX8 INVX8_25 ( .A(_abc_41234_new_n2513_), .Y(_abc_41234_new_n2958_));
INVX8 INVX8_26 ( .A(_abc_41234_new_n2911_), .Y(_abc_41234_new_n2959_));
INVX8 INVX8_27 ( .A(_abc_41234_new_n1606_), .Y(_abc_41234_new_n3914_));
INVX8 INVX8_3 ( .A(_abc_41234_new_n515__bF_buf5), .Y(_abc_41234_new_n534_));
INVX8 INVX8_4 ( .A(opcode_5_bF_buf2_), .Y(_abc_41234_new_n536_));
INVX8 INVX8_5 ( .A(_abc_41234_new_n537__bF_buf2), .Y(_abc_41234_new_n544_));
INVX8 INVX8_6 ( .A(opcode_2_), .Y(_abc_41234_new_n546_));
INVX8 INVX8_7 ( .A(opcode_3_bF_buf1_), .Y(_abc_41234_new_n555_));
INVX8 INVX8_8 ( .A(_abc_41234_new_n668__bF_buf5), .Y(_abc_41234_new_n669_));
INVX8 INVX8_9 ( .A(regfil_4__3_), .Y(_abc_41234_new_n819_));
MUX2X1 MUX2X1_1 ( .A(_abc_41234_new_n553_), .B(_abc_41234_new_n541_), .S(regfil_7__0_), .Y(_abc_41234_new_n554_));
MUX2X1 MUX2X1_10 ( .A(_abc_41234_new_n2376_), .B(_abc_41234_new_n2377_), .S(_abc_41234_new_n510_), .Y(_abc_41234_new_n2378_));
MUX2X1 MUX2X1_11 ( .A(auxcar), .B(rdatahold2_4_), .S(_abc_41234_new_n510_), .Y(_abc_41234_new_n2387_));
MUX2X1 MUX2X1_12 ( .A(_abc_41234_new_n616_), .B(_abc_41234_new_n714_), .S(_abc_41234_new_n2430_), .Y(_0opcode_7_0__0_));
MUX2X1 MUX2X1_13 ( .A(_abc_41234_new_n546__bF_buf0), .B(_abc_41234_new_n2435_), .S(_abc_41234_new_n2430_), .Y(_0opcode_7_0__2_));
MUX2X1 MUX2X1_14 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n890_), .S(_abc_41234_new_n2430_), .Y(_0opcode_7_0__4_));
MUX2X1 MUX2X1_15 ( .A(_abc_41234_new_n536__bF_buf5), .B(_abc_41234_new_n2441_), .S(_abc_41234_new_n2430_), .Y(_0opcode_7_0__5_));
MUX2X1 MUX2X1_16 ( .A(_abc_41234_new_n2532_), .B(_abc_41234_new_n2535_), .S(statesel_0_), .Y(_abc_41234_new_n2536_));
MUX2X1 MUX2X1_17 ( .A(_abc_41234_new_n2421_), .B(_abc_41234_new_n565_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold2_7_0__0_));
MUX2X1 MUX2X1_18 ( .A(_abc_41234_new_n2651_), .B(_abc_41234_new_n718_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold2_7_0__1_));
MUX2X1 MUX2X1_19 ( .A(_abc_41234_new_n2365_), .B(_abc_41234_new_n794_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold2_7_0__2_));
MUX2X1 MUX2X1_2 ( .A(_abc_41234_new_n654_), .B(_abc_41234_new_n529_), .S(_abc_41234_new_n615_), .Y(_abc_41234_new_n655_));
MUX2X1 MUX2X1_20 ( .A(_abc_41234_new_n2654_), .B(_abc_41234_new_n832_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold2_7_0__3_));
MUX2X1 MUX2X1_21 ( .A(_abc_41234_new_n2656_), .B(_abc_41234_new_n847_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold2_7_0__4_));
MUX2X1 MUX2X1_22 ( .A(_abc_41234_new_n2658_), .B(_abc_41234_new_n895_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold2_7_0__5_));
MUX2X1 MUX2X1_23 ( .A(_abc_41234_new_n2371_), .B(_abc_41234_new_n940_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold2_7_0__6_));
MUX2X1 MUX2X1_24 ( .A(_abc_41234_new_n2377_), .B(_abc_41234_new_n1005_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold2_7_0__7_));
MUX2X1 MUX2X1_25 ( .A(_abc_41234_new_n565_), .B(_abc_41234_new_n714_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold_7_0__0_));
MUX2X1 MUX2X1_26 ( .A(_abc_41234_new_n718_), .B(_abc_41234_new_n2432_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold_7_0__1_));
MUX2X1 MUX2X1_27 ( .A(_abc_41234_new_n794_), .B(_abc_41234_new_n2435_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold_7_0__2_));
MUX2X1 MUX2X1_28 ( .A(_abc_41234_new_n832_), .B(_abc_41234_new_n2437_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold_7_0__3_));
MUX2X1 MUX2X1_29 ( .A(_abc_41234_new_n847_), .B(_abc_41234_new_n890_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold_7_0__4_));
MUX2X1 MUX2X1_3 ( .A(regfil_1__4_), .B(_abc_41234_new_n879_), .S(_abc_41234_new_n1967_), .Y(_abc_41234_new_n2001_));
MUX2X1 MUX2X1_30 ( .A(_abc_41234_new_n895_), .B(_abc_41234_new_n2441_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold_7_0__5_));
MUX2X1 MUX2X1_31 ( .A(_abc_41234_new_n940_), .B(_abc_41234_new_n2443_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold_7_0__6_));
MUX2X1 MUX2X1_32 ( .A(_abc_41234_new_n1005_), .B(_abc_41234_new_n1016_), .S(_abc_41234_new_n2649_), .Y(_0rdatahold_7_0__7_));
MUX2X1 MUX2X1_33 ( .A(_abc_41234_new_n2707_), .B(_abc_41234_new_n1646_), .S(_abc_41234_new_n1729_), .Y(_abc_41234_new_n2708_));
MUX2X1 MUX2X1_34 ( .A(_abc_41234_new_n3466_), .B(_abc_41234_new_n1084_), .S(_abc_41234_new_n668__bF_buf3), .Y(_abc_41234_new_n3474_));
MUX2X1 MUX2X1_35 ( .A(alu__abc_40887_new_n333_), .B(alu__abc_40887_new_n136_), .S(alu__abc_40887_new_n204_), .Y(alu_res_5_));
MUX2X1 MUX2X1_4 ( .A(regfil_1__5_), .B(_abc_41234_new_n924_), .S(_abc_41234_new_n1967_), .Y(_abc_41234_new_n2008_));
MUX2X1 MUX2X1_5 ( .A(regfil_1__6_), .B(_abc_41234_new_n963_), .S(_abc_41234_new_n1967_), .Y(_abc_41234_new_n2017_));
MUX2X1 MUX2X1_6 ( .A(regfil_1__7_), .B(_abc_41234_new_n1010_), .S(_abc_41234_new_n1967_), .Y(_abc_41234_new_n2026_));
MUX2X1 MUX2X1_7 ( .A(regfil_2__4_), .B(_abc_41234_new_n879_), .S(_abc_41234_new_n2053_), .Y(_abc_41234_new_n2106_));
MUX2X1 MUX2X1_8 ( .A(regfil_2__5_), .B(_abc_41234_new_n924_), .S(_abc_41234_new_n2053_), .Y(_abc_41234_new_n2118_));
MUX2X1 MUX2X1_9 ( .A(_abc_41234_new_n2153_), .B(_abc_41234_new_n1509_), .S(_abc_41234_new_n2135_), .Y(_abc_41234_new_n2154_));
NAND2X1 NAND2X1_1 ( .A(state_2_), .B(_abc_41234_new_n503_), .Y(_abc_41234_new_n504_));
NAND2X1 NAND2X1_10 ( .A(opcode_1_), .B(opcode_0_), .Y(_abc_41234_new_n526_));
NAND2X1 NAND2X1_100 ( .A(_abc_41234_new_n1180_), .B(_abc_41234_new_n1183_), .Y(_abc_41234_new_n1184_));
NAND2X1 NAND2X1_101 ( .A(regfil_1__4_), .B(regfil_5__4_), .Y(_abc_41234_new_n1186_));
NAND2X1 NAND2X1_102 ( .A(regfil_1__5_), .B(regfil_5__5_), .Y(_abc_41234_new_n1187_));
NAND2X1 NAND2X1_103 ( .A(_abc_41234_new_n1189_), .B(_abc_41234_new_n1190_), .Y(_abc_41234_new_n1191_));
NAND2X1 NAND2X1_104 ( .A(_abc_41234_new_n1196_), .B(_abc_41234_new_n1193_), .Y(_abc_41234_new_n1197_));
NAND2X1 NAND2X1_105 ( .A(_abc_41234_new_n531_), .B(_abc_41234_new_n1052_), .Y(_abc_41234_new_n1199_));
NAND2X1 NAND2X1_106 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n1207_), .Y(_abc_41234_new_n1208_));
NAND2X1 NAND2X1_107 ( .A(_abc_41234_new_n848_), .B(_abc_41234_new_n1209_), .Y(_abc_41234_new_n1210_));
NAND2X1 NAND2X1_108 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n1211_), .Y(_abc_41234_new_n1212_));
NAND2X1 NAND2X1_109 ( .A(_abc_41234_new_n996_), .B(_abc_41234_new_n1213_), .Y(_abc_41234_new_n1214_));
NAND2X1 NAND2X1_11 ( .A(opcode_3_bF_buf3_), .B(opcode_2_), .Y(_abc_41234_new_n527_));
NAND2X1 NAND2X1_110 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1215_), .Y(_abc_41234_new_n1216_));
NAND2X1 NAND2X1_111 ( .A(regfil_5__2_), .B(_abc_41234_new_n1222_), .Y(_abc_41234_new_n1223_));
NAND2X1 NAND2X1_112 ( .A(regfil_5__3_bF_buf0_), .B(_abc_41234_new_n1224_), .Y(_abc_41234_new_n1225_));
NAND2X1 NAND2X1_113 ( .A(_abc_41234_new_n1228_), .B(_abc_41234_new_n1231_), .Y(_abc_41234_new_n1232_));
NAND2X1 NAND2X1_114 ( .A(_abc_41234_new_n748_), .B(_abc_41234_new_n1060_), .Y(_abc_41234_new_n1236_));
NAND2X1 NAND2X1_115 ( .A(_abc_41234_new_n1240_), .B(_abc_41234_new_n1215_), .Y(_abc_41234_new_n1241_));
NAND2X1 NAND2X1_116 ( .A(_abc_41234_new_n1256_), .B(_abc_41234_new_n1257_), .Y(_abc_41234_new_n1258_));
NAND2X1 NAND2X1_117 ( .A(_abc_41234_new_n1268_), .B(_abc_41234_new_n1151_), .Y(_abc_41234_new_n1269_));
NAND2X1 NAND2X1_118 ( .A(_abc_41234_new_n1196_), .B(_abc_41234_new_n1273_), .Y(_abc_41234_new_n1277_));
NAND2X1 NAND2X1_119 ( .A(_abc_41234_new_n1294_), .B(_abc_41234_new_n1293_), .Y(_abc_41234_new_n1295_));
NAND2X1 NAND2X1_12 ( .A(_abc_41234_new_n537__bF_buf3), .B(_abc_41234_new_n528_), .Y(_abc_41234_new_n538_));
NAND2X1 NAND2X1_120 ( .A(regfil_4__2_bF_buf1_), .B(sp_10_), .Y(_abc_41234_new_n1299_));
NAND2X1 NAND2X1_121 ( .A(_abc_41234_new_n1303_), .B(_abc_41234_new_n535_), .Y(_abc_41234_new_n1304_));
NAND2X1 NAND2X1_122 ( .A(_abc_41234_new_n530_), .B(_abc_41234_new_n1305_), .Y(_abc_41234_new_n1306_));
NAND2X1 NAND2X1_123 ( .A(_abc_41234_new_n535_), .B(_abc_41234_new_n1307_), .Y(_abc_41234_new_n1308_));
NAND2X1 NAND2X1_124 ( .A(_abc_41234_new_n1146_), .B(_abc_41234_new_n1266_), .Y(_abc_41234_new_n1310_));
NAND2X1 NAND2X1_125 ( .A(_abc_41234_new_n1323_), .B(_abc_41234_new_n535_), .Y(_abc_41234_new_n1324_));
NAND2X1 NAND2X1_126 ( .A(regfil_0__2_), .B(regfil_4__2_bF_buf2_), .Y(_abc_41234_new_n1331_));
NAND2X1 NAND2X1_127 ( .A(_abc_41234_new_n1333_), .B(_abc_41234_new_n1329_), .Y(_abc_41234_new_n1334_));
NAND2X1 NAND2X1_128 ( .A(_abc_41234_new_n1364_), .B(_abc_41234_new_n1360_), .Y(_abc_41234_new_n1365_));
NAND2X1 NAND2X1_129 ( .A(regfil_4__2_bF_buf0_), .B(_abc_41234_new_n537__bF_buf0), .Y(_abc_41234_new_n1368_));
NAND2X1 NAND2X1_13 ( .A(_abc_41234_new_n539_), .B(_abc_41234_new_n535_), .Y(_abc_41234_new_n540_));
NAND2X1 NAND2X1_130 ( .A(regfil_0__3_), .B(regfil_4__3_), .Y(_abc_41234_new_n1375_));
NAND2X1 NAND2X1_131 ( .A(_abc_41234_new_n1375_), .B(_abc_41234_new_n1377_), .Y(_abc_41234_new_n1378_));
NAND2X1 NAND2X1_132 ( .A(_abc_41234_new_n1060_), .B(_abc_41234_new_n1386_), .Y(_abc_41234_new_n1387_));
NAND2X1 NAND2X1_133 ( .A(_abc_41234_new_n849_), .B(_abc_41234_new_n1349_), .Y(_abc_41234_new_n1391_));
NAND2X1 NAND2X1_134 ( .A(_abc_41234_new_n1049__bF_buf1), .B(_abc_41234_new_n1394_), .Y(_abc_41234_new_n1395_));
NAND2X1 NAND2X1_135 ( .A(_abc_41234_new_n1301_), .B(_abc_41234_new_n1364_), .Y(_abc_41234_new_n1400_));
NAND2X1 NAND2X1_136 ( .A(regfil_0__4_), .B(regfil_4__4_), .Y(_abc_41234_new_n1425_));
NAND2X1 NAND2X1_137 ( .A(rdatahold_5_), .B(_abc_41234_new_n596_), .Y(_abc_41234_new_n1443_));
NAND2X1 NAND2X1_138 ( .A(_abc_41234_new_n1049__bF_buf4), .B(_abc_41234_new_n1450_), .Y(_abc_41234_new_n1451_));
NAND2X1 NAND2X1_139 ( .A(regfil_4__5_), .B(sp_13_), .Y(_abc_41234_new_n1457_));
NAND2X1 NAND2X1_14 ( .A(_abc_41234_new_n545_), .B(_abc_41234_new_n547_), .Y(_abc_41234_new_n548_));
NAND2X1 NAND2X1_140 ( .A(_abc_41234_new_n1410_), .B(_abc_41234_new_n1461_), .Y(_abc_41234_new_n1462_));
NAND2X1 NAND2X1_141 ( .A(_abc_41234_new_n1463_), .B(_abc_41234_new_n1406_), .Y(_abc_41234_new_n1464_));
NAND2X1 NAND2X1_142 ( .A(regfil_4__4_), .B(_abc_41234_new_n537__bF_buf3), .Y(_abc_41234_new_n1469_));
NAND2X1 NAND2X1_143 ( .A(regfil_0__5_), .B(regfil_4__5_), .Y(_abc_41234_new_n1472_));
NAND2X1 NAND2X1_144 ( .A(_abc_41234_new_n1427_), .B(_abc_41234_new_n1476_), .Y(_abc_41234_new_n1477_));
NAND2X1 NAND2X1_145 ( .A(_abc_41234_new_n1478_), .B(_abc_41234_new_n1433_), .Y(_abc_41234_new_n1479_));
NAND2X1 NAND2X1_146 ( .A(_abc_41234_new_n1479_), .B(_abc_41234_new_n1480_), .Y(_abc_41234_new_n1481_));
NAND2X1 NAND2X1_147 ( .A(regfil_5__7_), .B(_abc_41234_new_n992_), .Y(_abc_41234_new_n1487_));
NAND2X1 NAND2X1_148 ( .A(regfil_3__7_), .B(_abc_41234_new_n996_), .Y(_abc_41234_new_n1488_));
NAND2X1 NAND2X1_149 ( .A(_abc_41234_new_n1421_), .B(_abc_41234_new_n1496_), .Y(_abc_41234_new_n1497_));
NAND2X1 NAND2X1_15 ( .A(_abc_41234_new_n515__bF_buf4), .B(_abc_41234_new_n549_), .Y(_abc_41234_new_n550_));
NAND2X1 NAND2X1_150 ( .A(_abc_41234_new_n1420_), .B(_abc_41234_new_n1496_), .Y(_abc_41234_new_n1500_));
NAND2X1 NAND2X1_151 ( .A(rdatahold_6_), .B(_abc_41234_new_n596_), .Y(_abc_41234_new_n1507_));
NAND2X1 NAND2X1_152 ( .A(_abc_41234_new_n1509_), .B(_abc_41234_new_n1448_), .Y(_abc_41234_new_n1513_));
NAND2X1 NAND2X1_153 ( .A(_abc_41234_new_n1543_), .B(_abc_41234_new_n1479_), .Y(_abc_41234_new_n1544_));
NAND2X1 NAND2X1_154 ( .A(_abc_41234_new_n1571_), .B(_abc_41234_new_n1567_), .Y(_abc_41234_new_n1573_));
NAND2X1 NAND2X1_155 ( .A(regfil_0__7_), .B(regfil_4__7_), .Y(_abc_41234_new_n1578_));
NAND2X1 NAND2X1_156 ( .A(_abc_41234_new_n537__bF_buf2), .B(_abc_41234_new_n1608_), .Y(_abc_41234_new_n1609_));
NAND2X1 NAND2X1_157 ( .A(pc_5_), .B(pc_4_), .Y(_abc_41234_new_n1617_));
NAND2X1 NAND2X1_158 ( .A(pc_7_), .B(pc_6_), .Y(_abc_41234_new_n1618_));
NAND2X1 NAND2X1_159 ( .A(pc_8_), .B(_abc_41234_new_n1620_), .Y(_abc_41234_new_n1621_));
NAND2X1 NAND2X1_16 ( .A(opcode_2_), .B(_abc_41234_new_n555_), .Y(_abc_41234_new_n556_));
NAND2X1 NAND2X1_160 ( .A(_abc_41234_new_n1642_), .B(_abc_41234_new_n1638_), .Y(_abc_41234_new_n1643_));
NAND2X1 NAND2X1_161 ( .A(_abc_41234_new_n1615_), .B(_abc_41234_new_n1648_), .Y(_abc_41234_new_n1649_));
NAND2X1 NAND2X1_162 ( .A(pc_8_), .B(_abc_41234_new_n1651_), .Y(_abc_41234_new_n1652_));
NAND2X1 NAND2X1_163 ( .A(_abc_41234_new_n1650_), .B(_abc_41234_new_n1652_), .Y(_abc_41234_new_n1653_));
NAND2X1 NAND2X1_164 ( .A(opcode_4_bF_buf4_), .B(_abc_41234_new_n1143_), .Y(_abc_41234_new_n1655_));
NAND2X1 NAND2X1_165 ( .A(_abc_41234_new_n1669_), .B(_abc_41234_new_n1672_), .Y(_abc_41234_new_n1673_));
NAND2X1 NAND2X1_166 ( .A(opcode_4_bF_buf2_), .B(_abc_41234_new_n731_), .Y(_abc_41234_new_n1685_));
NAND2X1 NAND2X1_167 ( .A(intcyc_bF_buf0), .B(_abc_41234_new_n1675_), .Y(_abc_41234_new_n1689_));
NAND2X1 NAND2X1_168 ( .A(opcode_4_bF_buf0_), .B(_abc_41234_new_n769_), .Y(_abc_41234_new_n1700_));
NAND2X1 NAND2X1_169 ( .A(_abc_41234_new_n1708_), .B(_abc_41234_new_n1707_), .Y(_abc_41234_new_n1709_));
NAND2X1 NAND2X1_17 ( .A(_abc_41234_new_n536__bF_buf4), .B(_abc_41234_new_n557_), .Y(_abc_41234_new_n558_));
NAND2X1 NAND2X1_170 ( .A(opcode_4_bF_buf5_), .B(_abc_41234_new_n815_), .Y(_abc_41234_new_n1736_));
NAND2X1 NAND2X1_171 ( .A(_abc_41234_new_n1754_), .B(_abc_41234_new_n1753_), .Y(_abc_41234_new_n1755_));
NAND2X1 NAND2X1_172 ( .A(opcode_4_bF_buf3_), .B(_abc_41234_new_n859_), .Y(_abc_41234_new_n1760_));
NAND2X1 NAND2X1_173 ( .A(_abc_41234_new_n1775_), .B(_abc_41234_new_n1754_), .Y(_abc_41234_new_n1778_));
NAND2X1 NAND2X1_174 ( .A(intcyc_bF_buf0), .B(_abc_41234_new_n1776_), .Y(_abc_41234_new_n1781_));
NAND2X1 NAND2X1_175 ( .A(opcode_4_bF_buf1_), .B(_abc_41234_new_n900_), .Y(_abc_41234_new_n1782_));
NAND2X1 NAND2X1_176 ( .A(_abc_41234_new_n1639__bF_buf1), .B(_abc_41234_new_n1784_), .Y(_abc_41234_new_n1785_));
NAND2X1 NAND2X1_177 ( .A(pc_14_), .B(_abc_41234_new_n1796_), .Y(_abc_41234_new_n1797_));
NAND2X1 NAND2X1_178 ( .A(pc_14_), .B(_abc_41234_new_n1802_), .Y(_abc_41234_new_n1803_));
NAND2X1 NAND2X1_179 ( .A(_abc_41234_new_n1801_), .B(_abc_41234_new_n1803_), .Y(_abc_41234_new_n1804_));
NAND2X1 NAND2X1_18 ( .A(opcode_4_bF_buf3_), .B(carry), .Y(_abc_41234_new_n561_));
NAND2X1 NAND2X1_180 ( .A(regfil_7__6_), .B(_abc_41234_new_n1684_), .Y(_abc_41234_new_n1809_));
NAND2X1 NAND2X1_181 ( .A(opcode_4_bF_buf6_), .B(_abc_41234_new_n1535_), .Y(_abc_41234_new_n1811_));
NAND2X1 NAND2X1_182 ( .A(_abc_41234_new_n1825_), .B(_abc_41234_new_n1826_), .Y(_abc_41234_new_n1827_));
NAND2X1 NAND2X1_183 ( .A(_abc_41234_new_n1832_), .B(_abc_41234_new_n1831_), .Y(_abc_41234_new_n1833_));
NAND2X1 NAND2X1_184 ( .A(intcyc_bF_buf0), .B(_abc_41234_new_n1829_), .Y(_abc_41234_new_n1834_));
NAND2X1 NAND2X1_185 ( .A(opcode_4_bF_buf4_), .B(_abc_41234_new_n993_), .Y(_abc_41234_new_n1835_));
NAND2X1 NAND2X1_186 ( .A(_abc_41234_new_n1639__bF_buf3), .B(_abc_41234_new_n1837_), .Y(_abc_41234_new_n1838_));
NAND2X1 NAND2X1_187 ( .A(_abc_41234_new_n1049__bF_buf0), .B(_abc_41234_new_n1858_), .Y(_abc_41234_new_n1859_));
NAND2X1 NAND2X1_188 ( .A(_abc_41234_new_n1882_), .B(_abc_41234_new_n1869_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_1_));
NAND2X1 NAND2X1_189 ( .A(_abc_41234_new_n768_), .B(_abc_41234_new_n1871_), .Y(_abc_41234_new_n1888_));
NAND2X1 NAND2X1_19 ( .A(_abc_41234_new_n565_), .B(_abc_41234_new_n513_), .Y(_abc_41234_new_n566_));
NAND2X1 NAND2X1_190 ( .A(regfil_3__2_), .B(_abc_41234_new_n1870_), .Y(_abc_41234_new_n1892_));
NAND2X1 NAND2X1_191 ( .A(_abc_41234_new_n1891_), .B(_abc_41234_new_n1892_), .Y(_abc_41234_new_n1893_));
NAND2X1 NAND2X1_192 ( .A(_abc_41234_new_n814_), .B(_abc_41234_new_n1892_), .Y(_abc_41234_new_n1901_));
NAND2X1 NAND2X1_193 ( .A(_abc_41234_new_n1901_), .B(_abc_41234_new_n1903_), .Y(_abc_41234_new_n1904_));
NAND2X1 NAND2X1_194 ( .A(_abc_41234_new_n858_), .B(_abc_41234_new_n1911_), .Y(_abc_41234_new_n1912_));
NAND2X1 NAND2X1_195 ( .A(regfil_3__4_), .B(_abc_41234_new_n1902_), .Y(_abc_41234_new_n1917_));
NAND2X1 NAND2X1_196 ( .A(_abc_41234_new_n1916_), .B(_abc_41234_new_n1917_), .Y(_abc_41234_new_n1918_));
NAND2X1 NAND2X1_197 ( .A(_abc_41234_new_n899_), .B(_abc_41234_new_n1913_), .Y(_abc_41234_new_n1925_));
NAND2X1 NAND2X1_198 ( .A(_abc_41234_new_n1931_), .B(_abc_41234_new_n1930_), .Y(_abc_41234_new_n1932_));
NAND2X1 NAND2X1_199 ( .A(regfil_3__6_), .B(_abc_41234_new_n1929_), .Y(_abc_41234_new_n1943_));
NAND2X1 NAND2X1_2 ( .A(state_0_), .B(_abc_41234_new_n505_), .Y(_abc_41234_new_n506_));
NAND2X1 NAND2X1_20 ( .A(regfil_1__2_), .B(_abc_41234_new_n571_), .Y(_abc_41234_new_n572_));
NAND2X1 NAND2X1_200 ( .A(_abc_41234_new_n530_), .B(_abc_41234_new_n581_), .Y(_abc_41234_new_n1960_));
NAND2X1 NAND2X1_201 ( .A(rdatahold2_0_), .B(_abc_41234_new_n596_), .Y(_abc_41234_new_n1971_));
NAND2X1 NAND2X1_202 ( .A(_abc_41234_new_n569_), .B(_abc_41234_new_n570_), .Y(_abc_41234_new_n1976_));
NAND2X1 NAND2X1_203 ( .A(_abc_41234_new_n1976_), .B(_abc_41234_new_n1975_), .Y(_abc_41234_new_n1977_));
NAND2X1 NAND2X1_204 ( .A(rdatahold2_1_), .B(_abc_41234_new_n596_), .Y(_abc_41234_new_n1980_));
NAND2X1 NAND2X1_205 ( .A(_abc_41234_new_n1984_), .B(_abc_41234_new_n635_), .Y(_abc_41234_new_n1985_));
NAND2X1 NAND2X1_206 ( .A(rdatahold2_2_), .B(_abc_41234_new_n596_), .Y(_abc_41234_new_n1989_));
NAND2X1 NAND2X1_207 ( .A(_abc_41234_new_n1993_), .B(_abc_41234_new_n636_), .Y(_abc_41234_new_n1994_));
NAND2X1 NAND2X1_208 ( .A(rdatahold2_3_), .B(_abc_41234_new_n596_), .Y(_abc_41234_new_n1999_));
NAND2X1 NAND2X1_209 ( .A(_abc_41234_new_n639_), .B(_abc_41234_new_n2002_), .Y(_abc_41234_new_n2009_));
NAND2X1 NAND2X1_21 ( .A(regfil_1__5_), .B(regfil_1__4_), .Y(_abc_41234_new_n574_));
NAND2X1 NAND2X1_210 ( .A(_abc_41234_new_n577_), .B(_abc_41234_new_n583_), .Y(_abc_41234_new_n2031_));
NAND2X1 NAND2X1_211 ( .A(_abc_41234_new_n748_), .B(_abc_41234_new_n2035_), .Y(_abc_41234_new_n2038_));
NAND2X1 NAND2X1_212 ( .A(_abc_41234_new_n2035_), .B(_abc_41234_new_n791_), .Y(_abc_41234_new_n2040_));
NAND2X1 NAND2X1_213 ( .A(_abc_41234_new_n2035_), .B(_abc_41234_new_n829_), .Y(_abc_41234_new_n2042_));
NAND2X1 NAND2X1_214 ( .A(_abc_41234_new_n2035_), .B(_abc_41234_new_n879_), .Y(_abc_41234_new_n2044_));
NAND2X1 NAND2X1_215 ( .A(_abc_41234_new_n2035_), .B(_abc_41234_new_n924_), .Y(_abc_41234_new_n2046_));
NAND2X1 NAND2X1_216 ( .A(_abc_41234_new_n2035_), .B(_abc_41234_new_n963_), .Y(_abc_41234_new_n2049_));
NAND2X1 NAND2X1_217 ( .A(_abc_41234_new_n2035_), .B(_abc_41234_new_n1010_), .Y(_abc_41234_new_n2051_));
NAND2X1 NAND2X1_218 ( .A(_abc_41234_new_n992_), .B(_abc_41234_new_n1940_), .Y(_abc_41234_new_n2056_));
NAND2X1 NAND2X1_219 ( .A(regfil_2__0_), .B(_abc_41234_new_n1953_), .Y(_abc_41234_new_n2060_));
NAND2X1 NAND2X1_22 ( .A(regfil_1__7_), .B(regfil_1__6_), .Y(_abc_41234_new_n575_));
NAND2X1 NAND2X1_220 ( .A(_abc_41234_new_n2066_), .B(_abc_41234_new_n2055_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_0_));
NAND2X1 NAND2X1_221 ( .A(_abc_41234_new_n2071_), .B(_abc_41234_new_n1956_), .Y(_abc_41234_new_n2072_));
NAND2X1 NAND2X1_222 ( .A(_abc_41234_new_n2090_), .B(_abc_41234_new_n2081_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_2_));
NAND2X1 NAND2X1_223 ( .A(_abc_41234_new_n2093_), .B(_abc_41234_new_n2104_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_3_));
NAND2X1 NAND2X1_224 ( .A(_abc_41234_new_n859_), .B(_abc_41234_new_n2098_), .Y(_abc_41234_new_n2110_));
NAND2X1 NAND2X1_225 ( .A(_abc_41234_new_n2111_), .B(_abc_41234_new_n2110_), .Y(_abc_41234_new_n2112_));
NAND2X1 NAND2X1_226 ( .A(_abc_41234_new_n2121_), .B(_abc_41234_new_n2098_), .Y(_abc_41234_new_n2122_));
NAND2X1 NAND2X1_227 ( .A(regfil_2__5_), .B(_abc_41234_new_n2110_), .Y(_abc_41234_new_n2123_));
NAND2X1 NAND2X1_228 ( .A(_abc_41234_new_n2122_), .B(_abc_41234_new_n2123_), .Y(_abc_41234_new_n2124_));
NAND2X1 NAND2X1_229 ( .A(_abc_41234_new_n2142_), .B(_abc_41234_new_n1953_), .Y(_abc_41234_new_n2146_));
NAND2X1 NAND2X1_23 ( .A(_abc_41234_new_n576_), .B(_abc_41234_new_n573_), .Y(_abc_41234_new_n577_));
NAND2X1 NAND2X1_230 ( .A(_abc_41234_new_n940_), .B(_abc_41234_new_n2133_), .Y(_abc_41234_new_n2155_));
NAND2X1 NAND2X1_231 ( .A(rdatahold_6_), .B(_abc_41234_new_n1862_), .Y(_abc_41234_new_n2157_));
NAND2X1 NAND2X1_232 ( .A(_abc_41234_new_n2144_), .B(_abc_41234_new_n2143_), .Y(_abc_41234_new_n2166_));
NAND2X1 NAND2X1_233 ( .A(regfil_2__7_), .B(_abc_41234_new_n2167_), .Y(_abc_41234_new_n2168_));
NAND2X1 NAND2X1_234 ( .A(opcode_3_bF_buf3_), .B(_abc_41234_new_n524_), .Y(_abc_41234_new_n2182_));
NAND2X1 NAND2X1_235 ( .A(alu_sel_2_), .B(_abc_41234_new_n2177_), .Y(_abc_41234_new_n2195_));
NAND2X1 NAND2X1_236 ( .A(_abc_41234_new_n524_), .B(_abc_41234_new_n2201_), .Y(_abc_41234_new_n2202_));
NAND2X1 NAND2X1_237 ( .A(_abc_41234_new_n695_), .B(_abc_41234_new_n603_), .Y(_abc_41234_new_n2212_));
NAND2X1 NAND2X1_238 ( .A(regfil_6__0_), .B(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2251_));
NAND2X1 NAND2X1_239 ( .A(regfil_6__1_), .B(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2271_));
NAND2X1 NAND2X1_24 ( .A(_abc_41234_new_n531_), .B(_abc_41234_new_n581_), .Y(_abc_41234_new_n582_));
NAND2X1 NAND2X1_240 ( .A(regfil_6__2_), .B(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2283_));
NAND2X1 NAND2X1_241 ( .A(regfil_6__3_), .B(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2295_));
NAND2X1 NAND2X1_242 ( .A(regfil_6__4_), .B(_abc_41234_new_n2250_), .Y(_abc_41234_new_n2307_));
NAND2X1 NAND2X1_243 ( .A(opcode_4_bF_buf6_), .B(_abc_41234_new_n555_), .Y(_abc_41234_new_n2322_));
NAND2X1 NAND2X1_244 ( .A(_abc_41234_new_n2345_), .B(_abc_41234_new_n2348_), .Y(_abc_41234_new_n2349_));
NAND2X1 NAND2X1_245 ( .A(zero), .B(_abc_41234_new_n2363_), .Y(_abc_41234_new_n2370_));
NAND2X1 NAND2X1_246 ( .A(regfil_7__7_), .B(_abc_41234_new_n969_), .Y(_abc_41234_new_n2384_));
NAND2X1 NAND2X1_247 ( .A(auxcar), .B(_abc_41234_new_n550_), .Y(_abc_41234_new_n2385_));
NAND2X1 NAND2X1_248 ( .A(1'h0), .B(_abc_41234_new_n2362_), .Y(_abc_41234_new_n2388_));
NAND2X1 NAND2X1_249 ( .A(_abc_41234_new_n1537_), .B(_abc_41234_new_n1591_), .Y(_abc_41234_new_n2402_));
NAND2X1 NAND2X1_25 ( .A(state_3_), .B(_abc_41234_new_n589_), .Y(_abc_41234_new_n590_));
NAND2X1 NAND2X1_250 ( .A(_abc_41234_new_n1684_), .B(_abc_41234_new_n557_), .Y(_abc_41234_new_n2412_));
NAND2X1 NAND2X1_251 ( .A(_abc_41234_new_n690_), .B(_abc_41234_new_n699_), .Y(_abc_41234_new_n2419_));
NAND2X1 NAND2X1_252 ( .A(_abc_41234_new_n517_), .B(_abc_41234_new_n2427_), .Y(_abc_41234_new_n2428_));
NAND2X1 NAND2X1_253 ( .A(_abc_41234_new_n756_), .B(_abc_41234_new_n2429_), .Y(_abc_41234_new_n2430_));
NAND2X1 NAND2X1_254 ( .A(_abc_41234_new_n516__bF_buf0), .B(_abc_41234_new_n1046__bF_buf0), .Y(_abc_41234_new_n2449_));
NAND2X1 NAND2X1_255 ( .A(_abc_41234_new_n1684_), .B(_abc_41234_new_n598_), .Y(_abc_41234_new_n2451_));
NAND2X1 NAND2X1_256 ( .A(_abc_41234_new_n546__bF_buf5), .B(_abc_41234_new_n618_), .Y(_abc_41234_new_n2456_));
NAND2X1 NAND2X1_257 ( .A(_abc_41234_new_n1856_), .B(_abc_41234_new_n2458_), .Y(_abc_41234_new_n2459_));
NAND2X1 NAND2X1_258 ( .A(_abc_41234_new_n667_), .B(_abc_41234_new_n2469_), .Y(_abc_41234_new_n2470_));
NAND2X1 NAND2X1_259 ( .A(_abc_41234_new_n536__bF_buf4), .B(_abc_41234_new_n2469_), .Y(_abc_41234_new_n2471_));
NAND2X1 NAND2X1_26 ( .A(_abc_41234_new_n593_), .B(_abc_41234_new_n594_), .Y(_abc_41234_new_n595_));
NAND2X1 NAND2X1_260 ( .A(_abc_41234_new_n531_), .B(_abc_41234_new_n1608_), .Y(_abc_41234_new_n2474_));
NAND2X1 NAND2X1_261 ( .A(_abc_41234_new_n2464_), .B(_abc_41234_new_n2478_), .Y(_abc_41234_new_n2479_));
NAND2X1 NAND2X1_262 ( .A(_abc_41234_new_n2471_), .B(_abc_41234_new_n2491_), .Y(_abc_41234_new_n2492_));
NAND2X1 NAND2X1_263 ( .A(_abc_41234_new_n530_), .B(_abc_41234_new_n1608_), .Y(_abc_41234_new_n2496_));
NAND2X1 NAND2X1_264 ( .A(_abc_41234_new_n695_), .B(_abc_41234_new_n658_), .Y(_abc_41234_new_n2512_));
NAND2X1 NAND2X1_265 ( .A(_abc_41234_new_n502_), .B(_abc_41234_new_n2514_), .Y(_abc_41234_new_n2515_));
NAND2X1 NAND2X1_266 ( .A(_abc_41234_new_n502_), .B(_abc_41234_new_n2518_), .Y(_abc_41234_new_n2519_));
NAND2X1 NAND2X1_267 ( .A(_abc_41234_new_n692_), .B(_abc_41234_new_n705_), .Y(_abc_41234_new_n2521_));
NAND2X1 NAND2X1_268 ( .A(_abc_41234_new_n2511_), .B(_abc_41234_new_n2524_), .Y(_abc_41234_new_n2525_));
NAND2X1 NAND2X1_269 ( .A(_abc_41234_new_n502_), .B(_abc_41234_new_n522_), .Y(_abc_41234_new_n2526_));
NAND2X1 NAND2X1_27 ( .A(opcode_3_bF_buf3_), .B(_abc_41234_new_n546__bF_buf4), .Y(_abc_41234_new_n597_));
NAND2X1 NAND2X1_270 ( .A(_abc_41234_new_n2547_), .B(_abc_41234_new_n2542_), .Y(_abc_41234_new_n2548_));
NAND2X1 NAND2X1_271 ( .A(statesel_2_), .B(_abc_41234_new_n2578_), .Y(_abc_41234_new_n2579_));
NAND2X1 NAND2X1_272 ( .A(_abc_41234_new_n2613_), .B(_abc_41234_new_n2494_), .Y(_abc_41234_new_n2614_));
NAND2X1 NAND2X1_273 ( .A(_abc_41234_new_n515__bF_buf1), .B(_abc_41234_new_n2615_), .Y(_abc_41234_new_n2616_));
NAND2X1 NAND2X1_274 ( .A(statesel_4_), .B(_abc_41234_new_n2622_), .Y(_abc_41234_new_n2624_));
NAND2X1 NAND2X1_275 ( .A(_abc_41234_new_n2631_), .B(_abc_41234_new_n2629_), .Y(_abc_41234_new_n2632_));
NAND2X1 NAND2X1_276 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n1048_), .Y(_abc_41234_new_n2644_));
NAND2X1 NAND2X1_277 ( .A(popdes_0_), .B(_abc_41234_new_n2644_), .Y(_abc_41234_new_n2645_));
NAND2X1 NAND2X1_278 ( .A(popdes_1_), .B(_abc_41234_new_n2644_), .Y(_abc_41234_new_n2647_));
NAND2X1 NAND2X1_279 ( .A(_abc_41234_new_n756_), .B(_abc_41234_new_n2634_), .Y(_abc_41234_new_n2649_));
NAND2X1 NAND2X1_28 ( .A(_abc_41234_new_n531_), .B(_abc_41234_new_n598_), .Y(_abc_41234_new_n599_));
NAND2X1 NAND2X1_280 ( .A(_abc_41234_new_n517_), .B(_abc_41234_new_n2514_), .Y(_abc_41234_new_n2671_));
NAND2X1 NAND2X1_281 ( .A(opcode_4_bF_buf5_), .B(_abc_41234_new_n1848_), .Y(_abc_41234_new_n2685_));
NAND2X1 NAND2X1_282 ( .A(_abc_41234_new_n692_), .B(_abc_41234_new_n611_), .Y(_abc_41234_new_n2694_));
NAND2X1 NAND2X1_283 ( .A(_abc_41234_new_n662_), .B(_abc_41234_new_n2505_), .Y(_abc_41234_new_n2721_));
NAND2X1 NAND2X1_284 ( .A(pc_0_), .B(_abc_41234_new_n2732_), .Y(_abc_41234_new_n2733_));
NAND2X1 NAND2X1_285 ( .A(opcode_4_bF_buf2_), .B(_abc_41234_new_n768_), .Y(_abc_41234_new_n2740_));
NAND2X1 NAND2X1_286 ( .A(regfil_5__2_), .B(_abc_41234_new_n537__bF_buf0), .Y(_abc_41234_new_n2752_));
NAND2X1 NAND2X1_287 ( .A(wdatahold_2_), .B(_abc_41234_new_n2756_), .Y(_abc_41234_new_n2757_));
NAND2X1 NAND2X1_288 ( .A(_abc_41234_new_n1729_), .B(_abc_41234_new_n2776_), .Y(_abc_41234_new_n2777_));
NAND2X1 NAND2X1_289 ( .A(opcode_4_bF_buf1_), .B(_abc_41234_new_n814_), .Y(_abc_41234_new_n2779_));
NAND2X1 NAND2X1_29 ( .A(state_3_), .B(state_2_), .Y(_abc_41234_new_n604_));
NAND2X1 NAND2X1_290 ( .A(regfil_5__4_), .B(_abc_41234_new_n537__bF_buf1), .Y(_abc_41234_new_n2794_));
NAND2X1 NAND2X1_291 ( .A(opcode_4_bF_buf0_), .B(_abc_41234_new_n858_), .Y(_abc_41234_new_n2811_));
NAND2X1 NAND2X1_292 ( .A(opcode_4_bF_buf6_), .B(_abc_41234_new_n899_), .Y(_abc_41234_new_n2839_));
NAND2X1 NAND2X1_293 ( .A(_abc_41234_new_n2856_), .B(_abc_41234_new_n2803_), .Y(_abc_41234_new_n2857_));
NAND2X1 NAND2X1_294 ( .A(zero), .B(_abc_41234_new_n1684_), .Y(_abc_41234_new_n2860_));
NAND2X1 NAND2X1_295 ( .A(regfil_5__6_bF_buf0_), .B(_abc_41234_new_n537__bF_buf2), .Y(_abc_41234_new_n2861_));
NAND2X1 NAND2X1_296 ( .A(_abc_41234_new_n2875_), .B(_abc_41234_new_n2852_), .Y(_abc_41234_new_n2876_));
NAND2X1 NAND2X1_297 ( .A(opcode_4_bF_buf5_), .B(_abc_41234_new_n992_), .Y(_abc_41234_new_n2890_));
NAND2X1 NAND2X1_298 ( .A(_abc_41234_new_n2904_), .B(_abc_41234_new_n2897_), .Y(_abc_41234_new_n2905_));
NAND2X1 NAND2X1_299 ( .A(opcode_3_bF_buf2_), .B(_abc_41234_new_n1684_), .Y(_abc_41234_new_n2931_));
NAND2X1 NAND2X1_3 ( .A(_abc_41234_new_n502_), .B(_abc_41234_new_n507_), .Y(_abc_41234_new_n508_));
NAND2X1 NAND2X1_30 ( .A(_abc_41234_new_n605_), .B(_abc_41234_new_n603_), .Y(_abc_41234_new_n606_));
NAND2X1 NAND2X1_300 ( .A(_abc_41234_new_n2940_), .B(_abc_41234_new_n2938_), .Y(_abc_41234_new_n2941_));
NAND2X1 NAND2X1_301 ( .A(_abc_41234_new_n2942__bF_buf3), .B(_abc_41234_new_n2944_), .Y(_abc_41234_new_n2945_));
NAND2X1 NAND2X1_302 ( .A(_abc_41234_new_n662_), .B(_abc_41234_new_n665__bF_buf2), .Y(_abc_41234_new_n2950_));
NAND2X1 NAND2X1_303 ( .A(opcode_4_bF_buf3_), .B(_abc_41234_new_n730_), .Y(_abc_41234_new_n2963_));
NAND2X1 NAND2X1_304 ( .A(raddrhold_2_), .B(_abc_41234_new_n2987_), .Y(_abc_41234_new_n3018_));
NAND2X1 NAND2X1_305 ( .A(_abc_41234_new_n3075_), .B(_abc_41234_new_n3024_), .Y(_abc_41234_new_n3076_));
NAND2X1 NAND2X1_306 ( .A(raddrhold_4_), .B(_abc_41234_new_n3024_), .Y(_abc_41234_new_n3077_));
NAND2X1 NAND2X1_307 ( .A(opcode_4_bF_buf4_), .B(_abc_41234_new_n1936_), .Y(_abc_41234_new_n3104_));
NAND2X1 NAND2X1_308 ( .A(_abc_41234_new_n2189__bF_buf5), .B(_abc_41234_new_n3138_), .Y(_abc_41234_new_n3139_));
NAND2X1 NAND2X1_309 ( .A(_abc_41234_new_n2189__bF_buf4), .B(_abc_41234_new_n3163_), .Y(_abc_41234_new_n3164_));
NAND2X1 NAND2X1_31 ( .A(state_1_), .B(state_0_), .Y(_abc_41234_new_n610_));
NAND2X1 NAND2X1_310 ( .A(_abc_41234_new_n3204_), .B(_abc_41234_new_n3217_), .Y(_abc_41234_new_n3218_));
NAND2X1 NAND2X1_311 ( .A(raddrhold_10_), .B(_abc_41234_new_n3177_), .Y(_abc_41234_new_n3220_));
NAND2X1 NAND2X1_312 ( .A(_abc_41234_new_n2911_), .B(_abc_41234_new_n3220_), .Y(_abc_41234_new_n3221_));
NAND2X1 NAND2X1_313 ( .A(_abc_41234_new_n1046__bF_buf3), .B(_abc_41234_new_n3237_), .Y(_abc_41234_new_n3238_));
NAND2X1 NAND2X1_314 ( .A(_abc_41234_new_n849_), .B(_abc_41234_new_n669__bF_buf3), .Y(_abc_41234_new_n3250_));
NAND2X1 NAND2X1_315 ( .A(_abc_41234_new_n1046__bF_buf2), .B(_abc_41234_new_n3256_), .Y(_abc_41234_new_n3257_));
NAND2X1 NAND2X1_316 ( .A(_abc_41234_new_n1046__bF_buf1), .B(_abc_41234_new_n3280_), .Y(_abc_41234_new_n3281_));
NAND2X1 NAND2X1_317 ( .A(raddrhold_12_), .B(_abc_41234_new_n3267_), .Y(_abc_41234_new_n3289_));
NAND2X1 NAND2X1_318 ( .A(_abc_41234_new_n3300_), .B(_abc_41234_new_n3299_), .Y(_abc_41234_new_n3301_));
NAND2X1 NAND2X1_319 ( .A(_abc_41234_new_n2947__bF_buf2), .B(_abc_41234_new_n1643__bF_buf2), .Y(_abc_41234_new_n3340_));
NAND2X1 NAND2X1_32 ( .A(opcode_1_), .B(_abc_41234_new_n616_), .Y(_abc_41234_new_n620_));
NAND2X1 NAND2X1_320 ( .A(_abc_41234_new_n2458_), .B(_abc_41234_new_n2481_), .Y(_abc_41234_new_n3359_));
NAND2X1 NAND2X1_321 ( .A(_abc_41234_new_n2973_), .B(_abc_41234_new_n3359_), .Y(_abc_41234_new_n3360_));
NAND2X1 NAND2X1_322 ( .A(waddrhold_1_), .B(_abc_41234_new_n3343_), .Y(_abc_41234_new_n3364_));
NAND2X1 NAND2X1_323 ( .A(_abc_41234_new_n3337_), .B(_abc_41234_new_n3358_), .Y(_abc_41234_new_n3375_));
NAND2X1 NAND2X1_324 ( .A(_abc_41234_new_n515__bF_buf4), .B(_abc_41234_new_n2999_), .Y(_abc_41234_new_n3389_));
NAND2X1 NAND2X1_325 ( .A(waddrhold_2_), .B(_abc_41234_new_n3373_), .Y(_abc_41234_new_n3397_));
NAND2X1 NAND2X1_326 ( .A(_abc_41234_new_n515__bF_buf3), .B(_abc_41234_new_n3031_), .Y(_abc_41234_new_n3408_));
NAND2X1 NAND2X1_327 ( .A(_abc_41234_new_n1067_), .B(_abc_41234_new_n3382_), .Y(_abc_41234_new_n3423_));
NAND2X1 NAND2X1_328 ( .A(sp_4_), .B(_abc_41234_new_n3423_), .Y(_abc_41234_new_n3426_));
NAND2X1 NAND2X1_329 ( .A(_abc_41234_new_n3426_), .B(_abc_41234_new_n3425_), .Y(_abc_41234_new_n3427_));
NAND2X1 NAND2X1_33 ( .A(_abc_41234_new_n624_), .B(_abc_41234_new_n625_), .Y(_abc_41234_new_n626_));
NAND2X1 NAND2X1_330 ( .A(_abc_41234_new_n515__bF_buf2), .B(_abc_41234_new_n3056_), .Y(_abc_41234_new_n3431_));
NAND2X1 NAND2X1_331 ( .A(waddrhold_4_), .B(_abc_41234_new_n3415_), .Y(_abc_41234_new_n3439_));
NAND2X1 NAND2X1_332 ( .A(_abc_41234_new_n3446_), .B(_abc_41234_new_n3448_), .Y(_abc_41234_new_n3449_));
NAND2X1 NAND2X1_333 ( .A(_abc_41234_new_n515__bF_buf1), .B(_abc_41234_new_n3083_), .Y(_abc_41234_new_n3453_));
NAND2X1 NAND2X1_334 ( .A(_abc_41234_new_n1085_), .B(_abc_41234_new_n3447_), .Y(_abc_41234_new_n3467_));
NAND2X1 NAND2X1_335 ( .A(_abc_41234_new_n3468_), .B(_abc_41234_new_n3467_), .Y(_abc_41234_new_n3469_));
NAND2X1 NAND2X1_336 ( .A(_abc_41234_new_n515__bF_buf0), .B(_abc_41234_new_n3106_), .Y(_abc_41234_new_n3473_));
NAND2X1 NAND2X1_337 ( .A(waddrhold_6_), .B(_abc_41234_new_n3461_), .Y(_abc_41234_new_n3481_));
NAND2X1 NAND2X1_338 ( .A(_abc_41234_new_n3489_), .B(_abc_41234_new_n3488_), .Y(_abc_41234_new_n3490_));
NAND2X1 NAND2X1_339 ( .A(waddrhold_8_), .B(_abc_41234_new_n3502_), .Y(_abc_41234_new_n3520_));
NAND2X1 NAND2X1_34 ( .A(alu_res_0_), .B(_abc_41234_new_n613_), .Y(_abc_41234_new_n628_));
NAND2X1 NAND2X1_340 ( .A(_abc_41234_new_n515__bF_buf6), .B(_abc_41234_new_n1687_), .Y(_abc_41234_new_n3534_));
NAND2X1 NAND2X1_341 ( .A(_abc_41234_new_n3550_), .B(_abc_41234_new_n3549_), .Y(_abc_41234_new_n3551_));
NAND2X1 NAND2X1_342 ( .A(_abc_41234_new_n515__bF_buf5), .B(_abc_41234_new_n3208_), .Y(_abc_41234_new_n3555_));
NAND2X1 NAND2X1_343 ( .A(waddrhold_10_), .B(_abc_41234_new_n3542_), .Y(_abc_41234_new_n3563_));
NAND2X1 NAND2X1_344 ( .A(_abc_41234_new_n3528_), .B(_abc_41234_new_n3548_), .Y(_abc_41234_new_n3570_));
NAND2X1 NAND2X1_345 ( .A(_abc_41234_new_n515__bF_buf4), .B(_abc_41234_new_n3228_), .Y(_abc_41234_new_n3577_));
NAND2X1 NAND2X1_346 ( .A(_abc_41234_new_n1408_), .B(_abc_41234_new_n3592_), .Y(_abc_41234_new_n3593_));
NAND2X1 NAND2X1_347 ( .A(_abc_41234_new_n3594_), .B(_abc_41234_new_n3593_), .Y(_abc_41234_new_n3595_));
NAND2X1 NAND2X1_348 ( .A(waddrhold_12_), .B(_abc_41234_new_n3586_), .Y(_abc_41234_new_n3608_));
NAND2X1 NAND2X1_349 ( .A(_abc_41234_new_n3617_), .B(_abc_41234_new_n3592_), .Y(_abc_41234_new_n3618_));
NAND2X1 NAND2X1_35 ( .A(_abc_41234_new_n629_), .B(_abc_41234_new_n602_), .Y(_abc_41234_new_n630_));
NAND2X1 NAND2X1_350 ( .A(_abc_41234_new_n3618_), .B(_abc_41234_new_n3616_), .Y(_abc_41234_new_n3619_));
NAND2X1 NAND2X1_351 ( .A(_abc_41234_new_n1569_), .B(_abc_41234_new_n3638_), .Y(_abc_41234_new_n3658_));
NAND2X1 NAND2X1_352 ( .A(waddrhold_15_), .B(_abc_41234_new_n3338_), .Y(_abc_41234_new_n3674_));
NAND2X1 NAND2X1_353 ( .A(_abc_41234_new_n1221_), .B(_abc_41234_new_n2947__bF_buf1), .Y(_abc_41234_new_n3719_));
NAND2X1 NAND2X1_354 ( .A(_abc_41234_new_n1073_), .B(_abc_41234_new_n3734_), .Y(_abc_41234_new_n3735_));
NAND2X1 NAND2X1_355 ( .A(_abc_41234_new_n1118_), .B(_abc_41234_new_n3744_), .Y(_abc_41234_new_n3745_));
NAND2X1 NAND2X1_356 ( .A(_abc_41234_new_n768_), .B(_abc_41234_new_n1066__bF_buf1), .Y(_abc_41234_new_n3758_));
NAND2X1 NAND2X1_357 ( .A(_abc_41234_new_n1076_), .B(_abc_41234_new_n1077_), .Y(_abc_41234_new_n3763_));
NAND2X1 NAND2X1_358 ( .A(_abc_41234_new_n1166_), .B(_abc_41234_new_n1160_), .Y(_abc_41234_new_n3767_));
NAND2X1 NAND2X1_359 ( .A(_abc_41234_new_n3767_), .B(_abc_41234_new_n3766_), .Y(_abc_41234_new_n3768_));
NAND2X1 NAND2X1_36 ( .A(_abc_41234_new_n585_), .B(_abc_41234_new_n641_), .Y(_abc_41234_new_n642_));
NAND2X1 NAND2X1_360 ( .A(_abc_41234_new_n1121_), .B(_abc_41234_new_n1122_), .Y(_abc_41234_new_n3770_));
NAND2X1 NAND2X1_361 ( .A(_abc_41234_new_n3770_), .B(_abc_41234_new_n3771_), .Y(_abc_41234_new_n3772_));
NAND2X1 NAND2X1_362 ( .A(_abc_41234_new_n3765_), .B(_abc_41234_new_n3774_), .Y(_abc_41234_new_n3775_));
NAND2X1 NAND2X1_363 ( .A(_abc_41234_new_n3783_), .B(_abc_41234_new_n3798_), .Y(_abc_41234_new_n3799_));
NAND2X1 NAND2X1_364 ( .A(_abc_41234_new_n1049__bF_buf0), .B(_abc_41234_new_n3806_), .Y(_abc_41234_new_n3807_));
NAND2X1 NAND2X1_365 ( .A(_abc_41234_new_n3808_), .B(_abc_41234_new_n1229_), .Y(_abc_41234_new_n3809_));
NAND2X1 NAND2X1_366 ( .A(_abc_41234_new_n3811_), .B(_abc_41234_new_n3810_), .Y(_abc_41234_new_n3812_));
NAND2X1 NAND2X1_367 ( .A(_abc_41234_new_n1180_), .B(_abc_41234_new_n1170_), .Y(_abc_41234_new_n3816_));
NAND2X1 NAND2X1_368 ( .A(rdatahold2_5_), .B(_abc_41234_new_n1037_), .Y(_abc_41234_new_n3829_));
NAND2X1 NAND2X1_369 ( .A(_abc_41234_new_n1183_), .B(_abc_41234_new_n3837_), .Y(_abc_41234_new_n3839_));
NAND2X1 NAND2X1_37 ( .A(_abc_41234_new_n643_), .B(_abc_41234_new_n642_), .Y(_abc_41234_new_n644_));
NAND2X1 NAND2X1_370 ( .A(_abc_41234_new_n1325_), .B(_abc_41234_new_n3839_), .Y(_abc_41234_new_n3840_));
NAND2X1 NAND2X1_371 ( .A(rdatahold2_6_), .B(_abc_41234_new_n1037_), .Y(_abc_41234_new_n3854_));
NAND2X1 NAND2X1_372 ( .A(_abc_41234_new_n3859_), .B(_abc_41234_new_n3861_), .Y(_abc_41234_new_n3862_));
NAND2X1 NAND2X1_373 ( .A(_abc_41234_new_n3876_), .B(_abc_41234_new_n3875_), .Y(_abc_41234_new_n3877_));
NAND2X1 NAND2X1_374 ( .A(regfil_5__6_bF_buf2_), .B(_abc_41234_new_n1303_), .Y(_abc_41234_new_n3899_));
NAND2X1 NAND2X1_375 ( .A(_abc_41234_new_n1088_), .B(_abc_41234_new_n3872_), .Y(_abc_41234_new_n3902_));
NAND2X1 NAND2X1_376 ( .A(_abc_41234_new_n1684_), .B(_abc_41234_new_n2563_), .Y(_abc_41234_new_n3916_));
NAND2X1 NAND2X1_377 ( .A(_abc_41234_new_n517_), .B(_abc_41234_new_n3911_), .Y(_abc_41234_new_n3923_));
NAND2X1 NAND2X1_378 ( .A(_abc_41234_new_n1684_), .B(_abc_41234_new_n581_), .Y(_abc_41234_new_n3935_));
NAND2X1 NAND2X1_379 ( .A(sp_0_bF_buf3_), .B(_abc_41234_new_n3383_), .Y(_abc_41234_new_n3949_));
NAND2X1 NAND2X1_38 ( .A(_abc_41234_new_n632_), .B(_abc_41234_new_n647_), .Y(_abc_41234_new_n648_));
NAND2X1 NAND2X1_380 ( .A(_abc_41234_new_n3949_), .B(_abc_41234_new_n3936_), .Y(_abc_41234_new_n3950_));
NAND2X1 NAND2X1_381 ( .A(_abc_41234_new_n1071_), .B(_abc_41234_new_n3931_), .Y(_abc_41234_new_n3953_));
NAND2X1 NAND2X1_382 ( .A(_abc_41234_new_n3954_), .B(_abc_41234_new_n3953_), .Y(_abc_41234_new_n3955_));
NAND2X1 NAND2X1_383 ( .A(_abc_41234_new_n692_), .B(_abc_41234_new_n2427_), .Y(_abc_41234_new_n3962_));
NAND2X1 NAND2X1_384 ( .A(sp_3_), .B(_abc_41234_new_n3383_), .Y(_abc_41234_new_n3969_));
NAND2X1 NAND2X1_385 ( .A(_abc_41234_new_n1046__bF_buf7), .B(_abc_41234_new_n3972_), .Y(_abc_41234_new_n3973_));
NAND2X1 NAND2X1_386 ( .A(_abc_41234_new_n1067_), .B(_abc_41234_new_n3949_), .Y(_abc_41234_new_n3978_));
NAND2X1 NAND2X1_387 ( .A(_abc_41234_new_n3983_), .B(_abc_41234_new_n3975_), .Y(_abc_41234_new_n3984_));
NAND2X1 NAND2X1_388 ( .A(_abc_41234_new_n3404_), .B(_abc_41234_new_n3963_), .Y(_abc_41234_new_n3985_));
NAND2X1 NAND2X1_389 ( .A(sp_4_), .B(_abc_41234_new_n3979_), .Y(_abc_41234_new_n3995_));
NAND2X1 NAND2X1_39 ( .A(_abc_41234_new_n655_), .B(_abc_41234_new_n653_), .Y(_abc_41234_new_n656_));
NAND2X1 NAND2X1_390 ( .A(_abc_41234_new_n515__bF_buf5), .B(_abc_41234_new_n3916_), .Y(_abc_41234_new_n4009_));
NAND2X1 NAND2X1_391 ( .A(_abc_41234_new_n2947__bF_buf1), .B(_abc_41234_new_n3424_), .Y(_abc_41234_new_n4023_));
NAND2X1 NAND2X1_392 ( .A(_abc_41234_new_n515__bF_buf4), .B(_abc_41234_new_n4026_), .Y(_abc_41234_new_n4027_));
NAND2X1 NAND2X1_393 ( .A(_abc_41234_new_n4027_), .B(_abc_41234_new_n4020_), .Y(_abc_41234_new_n4028_));
NAND2X1 NAND2X1_394 ( .A(_abc_41234_new_n3963_), .B(_abc_41234_new_n3449_), .Y(_abc_41234_new_n4030_));
NAND2X1 NAND2X1_395 ( .A(_abc_41234_new_n3960_), .B(_abc_41234_new_n4016_), .Y(_abc_41234_new_n4032_));
NAND2X1 NAND2X1_396 ( .A(sp_6_), .B(_abc_41234_new_n4013_), .Y(_abc_41234_new_n4039_));
NAND2X1 NAND2X1_397 ( .A(sp_0_bF_buf2_), .B(_abc_41234_new_n4040_), .Y(_abc_41234_new_n4041_));
NAND2X1 NAND2X1_398 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n4047_), .Y(_abc_41234_new_n4051_));
NAND2X1 NAND2X1_399 ( .A(regfil_5__6_bF_buf1_), .B(_abc_41234_new_n1106_), .Y(_abc_41234_new_n4052_));
NAND2X1 NAND2X1_4 ( .A(popdes_0_), .B(popdes_1_), .Y(_abc_41234_new_n510_));
NAND2X1 NAND2X1_40 ( .A(_abc_41234_new_n517_), .B(_abc_41234_new_n658_), .Y(_abc_41234_new_n659_));
NAND2X1 NAND2X1_400 ( .A(_abc_41234_new_n516__bF_buf0), .B(_abc_41234_new_n4056_), .Y(_abc_41234_new_n4057_));
NAND2X1 NAND2X1_401 ( .A(_abc_41234_new_n4059_), .B(_abc_41234_new_n4060_), .Y(_abc_41234_new_n4061_));
NAND2X1 NAND2X1_402 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n4082_), .Y(_abc_41234_new_n4083_));
NAND2X1 NAND2X1_403 ( .A(_abc_41234_new_n1255_), .B(_abc_41234_new_n4069_), .Y(_abc_41234_new_n4092_));
NAND2X1 NAND2X1_404 ( .A(_abc_41234_new_n3936_), .B(_abc_41234_new_n4104_), .Y(_abc_41234_new_n4105_));
NAND2X1 NAND2X1_405 ( .A(_abc_41234_new_n515__bF_buf0), .B(_abc_41234_new_n4129_), .Y(_abc_41234_new_n4130_));
NAND2X1 NAND2X1_406 ( .A(sp_10_), .B(_abc_41234_new_n4101_), .Y(_abc_41234_new_n4131_));
NAND2X1 NAND2X1_407 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n4133_), .Y(_abc_41234_new_n4134_));
NAND2X1 NAND2X1_408 ( .A(regfil_4__2_bF_buf3_), .B(_abc_41234_new_n1106_), .Y(_abc_41234_new_n4135_));
NAND2X1 NAND2X1_409 ( .A(_abc_41234_new_n3960_), .B(_abc_41234_new_n4133_), .Y(_abc_41234_new_n4140_));
NAND2X1 NAND2X1_41 ( .A(_abc_41234_new_n676_), .B(_abc_41234_new_n672_), .Y(_abc_41234_new_n677_));
NAND2X1 NAND2X1_410 ( .A(rdatahold_2_), .B(_abc_41234_new_n3964_), .Y(_abc_41234_new_n4141_));
NAND2X1 NAND2X1_411 ( .A(_abc_41234_new_n3963_), .B(_abc_41234_new_n3551_), .Y(_abc_41234_new_n4142_));
NAND2X1 NAND2X1_412 ( .A(_abc_41234_new_n4146_), .B(_abc_41234_new_n4147_), .Y(_abc_41234_new_n4148_));
NAND2X1 NAND2X1_413 ( .A(_abc_41234_new_n3963_), .B(_abc_41234_new_n3573_), .Y(_abc_41234_new_n4164_));
NAND2X1 NAND2X1_414 ( .A(_abc_41234_new_n2947__bF_buf2), .B(_abc_41234_new_n3592_), .Y(_abc_41234_new_n4169_));
NAND2X1 NAND2X1_415 ( .A(_abc_41234_new_n515__bF_buf5), .B(_abc_41234_new_n4177_), .Y(_abc_41234_new_n4178_));
NAND2X1 NAND2X1_416 ( .A(_abc_41234_new_n4179_), .B(_abc_41234_new_n4175_), .Y(_abc_41234_new_n4180_));
NAND2X1 NAND2X1_417 ( .A(sp_13_), .B(_abc_41234_new_n4174_), .Y(_abc_41234_new_n4189_));
NAND2X1 NAND2X1_418 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n4219_), .Y(_abc_41234_new_n4220_));
NAND2X1 NAND2X1_419 ( .A(_abc_41234_new_n3960_), .B(_abc_41234_new_n4219_), .Y(_abc_41234_new_n4228_));
NAND2X1 NAND2X1_42 ( .A(_abc_41234_new_n549_), .B(_abc_41234_new_n535_), .Y(_abc_41234_new_n685_));
NAND2X1 NAND2X1_420 ( .A(rdatahold_6_), .B(_abc_41234_new_n3964_), .Y(_abc_41234_new_n4230_));
NAND2X1 NAND2X1_421 ( .A(sp_15_), .B(_abc_41234_new_n4211_), .Y(_abc_41234_new_n4234_));
NAND2X1 NAND2X1_422 ( .A(_abc_41234_new_n3657_), .B(_abc_41234_new_n3658_), .Y(_abc_41234_new_n4245_));
NAND2X1 NAND2X1_423 ( .A(_abc_41234_new_n3963_), .B(_abc_41234_new_n4245_), .Y(_abc_41234_new_n4252_));
NAND2X1 NAND2X1_424 ( .A(rdatahold_7_), .B(_abc_41234_new_n3964_), .Y(_abc_41234_new_n4253_));
NAND2X1 NAND2X1_425 ( .A(_abc_41234_new_n646_), .B(_abc_41234_new_n4257_), .Y(_abc_41234_new_n4258_));
NAND2X1 NAND2X1_426 ( .A(_abc_41234_new_n748_), .B(_abc_41234_new_n4257_), .Y(_abc_41234_new_n4260_));
NAND2X1 NAND2X1_427 ( .A(_abc_41234_new_n4257_), .B(_abc_41234_new_n791_), .Y(_abc_41234_new_n4262_));
NAND2X1 NAND2X1_428 ( .A(_abc_41234_new_n4257_), .B(_abc_41234_new_n829_), .Y(_abc_41234_new_n4264_));
NAND2X1 NAND2X1_429 ( .A(_abc_41234_new_n4257_), .B(_abc_41234_new_n879_), .Y(_abc_41234_new_n4266_));
NAND2X1 NAND2X1_43 ( .A(state_1_), .B(_abc_41234_new_n520_), .Y(_abc_41234_new_n694_));
NAND2X1 NAND2X1_430 ( .A(_abc_41234_new_n4257_), .B(_abc_41234_new_n924_), .Y(_abc_41234_new_n4268_));
NAND2X1 NAND2X1_431 ( .A(_abc_41234_new_n4257_), .B(_abc_41234_new_n963_), .Y(_abc_41234_new_n4270_));
NAND2X1 NAND2X1_432 ( .A(_abc_41234_new_n4257_), .B(_abc_41234_new_n1010_), .Y(_abc_41234_new_n4272_));
NAND2X1 NAND2X1_433 ( .A(pc_0_), .B(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4276_));
NAND2X1 NAND2X1_434 ( .A(_abc_41234_new_n1684_), .B(_abc_41234_new_n1628_), .Y(_abc_41234_new_n4288_));
NAND2X1 NAND2X1_435 ( .A(_abc_41234_new_n2458_), .B(_abc_41234_new_n4293_), .Y(_abc_41234_new_n4294_));
NAND2X1 NAND2X1_436 ( .A(_abc_41234_new_n4298_), .B(_abc_41234_new_n4296_), .Y(_abc_41234_new_n4299_));
NAND2X1 NAND2X1_437 ( .A(_abc_41234_new_n1305_), .B(_abc_41234_new_n2677_), .Y(_abc_41234_new_n4300_));
NAND2X1 NAND2X1_438 ( .A(pc_3_), .B(_abc_41234_new_n2732_), .Y(_abc_41234_new_n4353_));
NAND2X1 NAND2X1_439 ( .A(_abc_41234_new_n4354_), .B(_abc_41234_new_n4353_), .Y(_abc_41234_new_n4355_));
NAND2X1 NAND2X1_44 ( .A(_abc_41234_new_n516__bF_buf3), .B(_abc_41234_new_n699_), .Y(_abc_41234_new_n700_));
NAND2X1 NAND2X1_440 ( .A(_abc_41234_new_n1613_), .B(_abc_41234_new_n4297__bF_buf3), .Y(_abc_41234_new_n4358_));
NAND2X1 NAND2X1_441 ( .A(pc_4_), .B(_abc_41234_new_n4275_), .Y(_abc_41234_new_n4384_));
NAND2X1 NAND2X1_442 ( .A(pc_6_), .B(_abc_41234_new_n4407_), .Y(_abc_41234_new_n4408_));
NAND2X1 NAND2X1_443 ( .A(_abc_41234_new_n4301_), .B(_abc_41234_new_n4410_), .Y(_abc_41234_new_n4417_));
NAND2X1 NAND2X1_444 ( .A(_abc_41234_new_n1046__bF_buf2), .B(_abc_41234_new_n4420_), .Y(_abc_41234_new_n4421_));
NAND2X1 NAND2X1_445 ( .A(_abc_41234_new_n1046__bF_buf1), .B(_abc_41234_new_n4434_), .Y(_abc_41234_new_n4435_));
NAND2X1 NAND2X1_446 ( .A(pc_8_), .B(_abc_41234_new_n4427_), .Y(_abc_41234_new_n4446_));
NAND2X1 NAND2X1_447 ( .A(_abc_41234_new_n4446_), .B(_abc_41234_new_n4445_), .Y(_abc_41234_new_n4447_));
NAND2X1 NAND2X1_448 ( .A(_abc_41234_new_n1046__bF_buf0), .B(_abc_41234_new_n4457_), .Y(_abc_41234_new_n4458_));
NAND2X1 NAND2X1_449 ( .A(_abc_41234_new_n1670_), .B(_abc_41234_new_n4446_), .Y(_abc_41234_new_n4466_));
NAND2X1 NAND2X1_45 ( .A(_abc_41234_new_n517_), .B(_abc_41234_new_n705_), .Y(_abc_41234_new_n706_));
NAND2X1 NAND2X1_450 ( .A(_abc_41234_new_n4465_), .B(_abc_41234_new_n4466_), .Y(_abc_41234_new_n4467_));
NAND2X1 NAND2X1_451 ( .A(_abc_41234_new_n1670_), .B(_abc_41234_new_n4297__bF_buf3), .Y(_abc_41234_new_n4474_));
NAND2X1 NAND2X1_452 ( .A(_abc_41234_new_n665__bF_buf0), .B(_abc_41234_new_n4483_), .Y(_abc_41234_new_n4484_));
NAND2X1 NAND2X1_453 ( .A(_abc_41234_new_n1606_), .B(_abc_41234_new_n1716_), .Y(_abc_41234_new_n4494_));
NAND2X1 NAND2X1_454 ( .A(_abc_41234_new_n4494_), .B(_abc_41234_new_n4493_), .Y(_abc_41234_new_n4495_));
NAND2X1 NAND2X1_455 ( .A(_abc_41234_new_n4501_), .B(_abc_41234_new_n4500_), .Y(_abc_41234_new_n4502_));
NAND2X1 NAND2X1_456 ( .A(_abc_41234_new_n1734_), .B(_abc_41234_new_n4507_), .Y(_abc_41234_new_n4508_));
NAND2X1 NAND2X1_457 ( .A(_abc_41234_new_n660__bF_buf6), .B(_abc_41234_new_n4513_), .Y(_abc_41234_new_n4514_));
NAND2X1 NAND2X1_458 ( .A(pc_12_), .B(_abc_41234_new_n4499_), .Y(_abc_41234_new_n4518_));
NAND2X1 NAND2X1_459 ( .A(_abc_41234_new_n4518_), .B(_abc_41234_new_n4517_), .Y(_abc_41234_new_n4519_));
NAND2X1 NAND2X1_46 ( .A(opcode_0_), .B(_abc_41234_new_n721_), .Y(_abc_41234_new_n722_));
NAND2X1 NAND2X1_460 ( .A(_abc_41234_new_n4304_), .B(_abc_41234_new_n4307_), .Y(_abc_41234_new_n4528_));
NAND2X1 NAND2X1_461 ( .A(pc_12_), .B(_abc_41234_new_n4312_), .Y(_abc_41234_new_n4530_));
NAND2X1 NAND2X1_462 ( .A(_abc_41234_new_n4537_), .B(_abc_41234_new_n4538_), .Y(_abc_41234_new_n4539_));
NAND2X1 NAND2X1_463 ( .A(pc_14_), .B(_abc_41234_new_n4555_), .Y(_abc_41234_new_n4556_));
NAND2X1 NAND2X1_464 ( .A(_abc_41234_new_n4557_), .B(_abc_41234_new_n4556_), .Y(_abc_41234_new_n4558_));
NAND2X1 NAND2X1_465 ( .A(_abc_41234_new_n1606_), .B(_abc_41234_new_n1833_), .Y(_abc_41234_new_n4594_));
NAND2X1 NAND2X1_466 ( .A(_abc_41234_new_n660__bF_buf2), .B(_abc_41234_new_n4595_), .Y(_abc_41234_new_n4596_));
NAND2X1 NAND2X1_467 ( .A(_abc_41234_new_n2518_), .B(_abc_41234_new_n519_), .Y(_abc_41234_new_n4599_));
NAND2X1 NAND2X1_468 ( .A(_abc_41234_new_n502_), .B(_abc_41234_new_n705_), .Y(_abc_41234_new_n4612_));
NAND2X1 NAND2X1_469 ( .A(raddrhold_9_), .B(_abc_41234_new_n516__bF_buf1), .Y(_abc_41234_new_n4662_));
NAND2X1 NAND2X1_47 ( .A(regfil_0__1_), .B(_abc_41234_new_n618_), .Y(_abc_41234_new_n728_));
NAND2X1 NAND2X1_470 ( .A(raddrhold_10_), .B(_abc_41234_new_n516__bF_buf0), .Y(_abc_41234_new_n4667_));
NAND2X1 NAND2X1_471 ( .A(raddrhold_11_), .B(_abc_41234_new_n516__bF_buf5), .Y(_abc_41234_new_n4672_));
NAND2X1 NAND2X1_472 ( .A(raddrhold_14_), .B(_abc_41234_new_n2911_), .Y(_abc_41234_new_n4685_));
NAND2X1 NAND2X1_473 ( .A(_auto_iopadmap_cc_368_execute_45645), .B(_abc_41234_new_n4695_), .Y(_abc_41234_new_n4696_));
NAND2X1 NAND2X1_474 ( .A(_abc_41234_new_n1033_), .B(_abc_41234_new_n608_), .Y(_abc_41234_new_n4703_));
NAND2X1 NAND2X1_475 ( .A(_abc_41234_new_n502_), .B(_abc_41234_new_n3911_), .Y(_abc_41234_new_n4704_));
NAND2X1 NAND2X1_476 ( .A(_auto_iopadmap_cc_368_execute_45651), .B(_abc_41234_new_n516__bF_buf3), .Y(_abc_41234_new_n4706_));
NAND2X1 NAND2X1_477 ( .A(parity), .B(_abc_41234_new_n2248_), .Y(_abc_41234_new_n4751_));
NAND2X1 NAND2X1_478 ( .A(_abc_41234_new_n4763_), .B(_abc_41234_new_n4760_), .Y(_abc_41234_new_n4764_));
NAND2X1 NAND2X1_479 ( .A(_abc_41234_new_n4772_), .B(_abc_41234_new_n4771_), .Y(_abc_41234_new_n4773_));
NAND2X1 NAND2X1_48 ( .A(\data[1] ), .B(_abc_41234_new_n758_), .Y(_abc_41234_new_n759_));
NAND2X1 NAND2X1_480 ( .A(_abc_41234_new_n4757_), .B(_abc_41234_new_n4774_), .Y(_abc_41234_new_n4775_));
NAND2X1 NAND2X1_481 ( .A(_abc_41234_new_n4766_), .B(_abc_41234_new_n4760_), .Y(_abc_41234_new_n4776_));
NAND2X1 NAND2X1_482 ( .A(_abc_41234_new_n4780_), .B(_abc_41234_new_n4779_), .Y(_abc_41234_new_n4781_));
NAND2X1 NAND2X1_483 ( .A(_abc_41234_new_n535_), .B(_abc_41234_new_n4293_), .Y(_abc_41234_new_n4784_));
NAND2X1 NAND2X1_484 ( .A(_abc_41234_new_n4799_), .B(_abc_41234_new_n4804_), .Y(_abc_41234_new_n4805_));
NAND2X1 NAND2X1_485 ( .A(_abc_41234_new_n2557_), .B(_abc_41234_new_n2601_), .Y(_abc_41234_new_n4809_));
NAND2X1 NAND2X1_486 ( .A(_abc_41234_new_n4811_), .B(_abc_41234_new_n2535_), .Y(_abc_41234_new_n4812_));
NAND2X1 NAND2X1_487 ( .A(_abc_41234_new_n4817_), .B(_abc_41234_new_n4806_), .Y(_abc_41234_new_n4818_));
NAND2X1 NAND2X1_488 ( .A(_abc_41234_new_n2208_), .B(_abc_41234_new_n4823_), .Y(_abc_41234_new_n4824_));
NAND2X1 NAND2X1_489 ( .A(_abc_41234_new_n4832_), .B(_abc_41234_new_n4830_), .Y(_abc_41234_new_n4833_));
NAND2X1 NAND2X1_49 ( .A(rdatahold_2_), .B(_abc_41234_new_n596_), .Y(_abc_41234_new_n765_));
NAND2X1 NAND2X1_490 ( .A(_abc_41234_new_n4761_), .B(_abc_41234_new_n4803_), .Y(_abc_41234_new_n4834_));
NAND2X1 NAND2X1_491 ( .A(_abc_41234_new_n4846_), .B(_abc_41234_new_n4779_), .Y(_abc_41234_new_n4852_));
NAND2X1 NAND2X1_492 ( .A(_abc_41234_new_n4781_), .B(_abc_41234_new_n4771_), .Y(_abc_41234_new_n4858_));
NAND2X1 NAND2X1_493 ( .A(_abc_41234_new_n4849_), .B(_abc_41234_new_n2535_), .Y(_abc_41234_new_n4870_));
NAND2X1 NAND2X1_494 ( .A(_abc_41234_new_n4842_), .B(_abc_41234_new_n4875_), .Y(_abc_41234_new_n4876_));
NAND2X1 NAND2X1_495 ( .A(_abc_41234_new_n4789_), .B(_abc_41234_new_n4779_), .Y(_abc_41234_new_n4882_));
NAND2X1 NAND2X1_496 ( .A(_abc_41234_new_n3936_), .B(_abc_41234_new_n4054_), .Y(_abc_41234_new_n4890_));
NAND2X1 NAND2X1_497 ( .A(alu_oprb_7_), .B(alu_opra_7_), .Y(alu__abc_40887_new_n34_));
NAND2X1 NAND2X1_498 ( .A(alu_oprb_6_), .B(alu_opra_6_), .Y(alu__abc_40887_new_n38_));
NAND2X1 NAND2X1_499 ( .A(alu__abc_40887_new_n38_), .B(alu__abc_40887_new_n40_), .Y(alu__abc_40887_new_n41_));
NAND2X1 NAND2X1_5 ( .A(_abc_41234_new_n511_), .B(_abc_41234_new_n509_), .Y(_abc_41234_new_n512_));
NAND2X1 NAND2X1_50 ( .A(_abc_41234_new_n771_), .B(_abc_41234_new_n777_), .Y(_abc_41234_new_n778_));
NAND2X1 NAND2X1_500 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_40887_new_n43_));
NAND2X1 NAND2X1_501 ( .A(alu_oprb_0_), .B(alu_opra_0_), .Y(alu__abc_40887_new_n45_));
NAND2X1 NAND2X1_502 ( .A(alu_oprb_4_), .B(alu_opra_4_), .Y(alu__abc_40887_new_n56_));
NAND2X1 NAND2X1_503 ( .A(alu_oprb_5_), .B(alu_opra_5_), .Y(alu__abc_40887_new_n60_));
NAND2X1 NAND2X1_504 ( .A(alu__abc_40887_new_n58_), .B(alu__abc_40887_new_n62_), .Y(alu__abc_40887_new_n63_));
NAND2X1 NAND2X1_505 ( .A(alu__abc_40887_new_n55_), .B(alu__abc_40887_new_n53_), .Y(alu__abc_40887_new_n70_));
NAND2X1 NAND2X1_506 ( .A(alu__abc_40887_new_n66_), .B(alu__abc_40887_new_n73_), .Y(alu__abc_40887_new_n74_));
NAND2X1 NAND2X1_507 ( .A(alu__abc_40887_new_n58_), .B(alu__abc_40887_new_n70_), .Y(alu__abc_40887_new_n75_));
NAND2X1 NAND2X1_508 ( .A(alu__abc_40887_new_n76_), .B(alu__abc_40887_new_n62_), .Y(alu__abc_40887_new_n79_));
NAND2X1 NAND2X1_509 ( .A(alu_oprb_3_), .B(alu_opra_3_), .Y(alu__abc_40887_new_n83_));
NAND2X1 NAND2X1_51 ( .A(_abc_41234_new_n778_), .B(_abc_41234_new_n657_), .Y(_abc_41234_new_n779_));
NAND2X1 NAND2X1_510 ( .A(alu__abc_40887_new_n83_), .B(alu__abc_40887_new_n54_), .Y(alu__abc_40887_new_n84_));
NAND2X1 NAND2X1_511 ( .A(alu_oprb_2_), .B(alu_opra_2_), .Y(alu__abc_40887_new_n86_));
NAND2X1 NAND2X1_512 ( .A(alu__abc_40887_new_n49_), .B(alu__abc_40887_new_n46_), .Y(alu__abc_40887_new_n87_));
NAND2X1 NAND2X1_513 ( .A(alu__abc_40887_new_n43_), .B(alu__abc_40887_new_n89_), .Y(alu__abc_40887_new_n90_));
NAND2X1 NAND2X1_514 ( .A(alu__abc_40887_new_n56_), .B(alu__abc_40887_new_n57_), .Y(alu__abc_40887_new_n97_));
NAND2X1 NAND2X1_515 ( .A(alu__abc_40887_new_n97_), .B(alu__abc_40887_new_n78_), .Y(alu__abc_40887_new_n98_));
NAND2X1 NAND2X1_516 ( .A(alu_sel_0_), .B(alu__abc_40887_new_n102_), .Y(alu__abc_40887_new_n103_));
NAND2X1 NAND2X1_517 ( .A(alu__abc_40887_new_n38_), .B(alu__abc_40887_new_n66_), .Y(alu__abc_40887_new_n105_));
NAND2X1 NAND2X1_518 ( .A(alu__abc_40887_new_n107_), .B(alu__abc_40887_new_n106_), .Y(alu__abc_40887_new_n108_));
NAND2X1 NAND2X1_519 ( .A(alu__abc_40887_new_n108_), .B(alu__abc_40887_new_n112_), .Y(alu__abc_40887_new_n113_));
NAND2X1 NAND2X1_52 ( .A(_abc_41234_new_n780_), .B(_abc_41234_new_n779_), .Y(_abc_41234_new_n781_));
NAND2X1 NAND2X1_520 ( .A(alu_opra_2_), .B(alu__abc_40887_new_n122_), .Y(alu__abc_40887_new_n123_));
NAND2X1 NAND2X1_521 ( .A(alu_oprb_0_), .B(alu__abc_40887_new_n128_), .Y(alu__abc_40887_new_n129_));
NAND2X1 NAND2X1_522 ( .A(alu__abc_40887_new_n122_), .B(alu__abc_40887_new_n150_), .Y(alu__abc_40887_new_n151_));
NAND2X1 NAND2X1_523 ( .A(alu__abc_40887_new_n158_), .B(alu__abc_40887_new_n155_), .Y(alu__abc_40887_new_n159_));
NAND2X1 NAND2X1_524 ( .A(alu__abc_40887_new_n86_), .B(alu__abc_40887_new_n151_), .Y(alu__abc_40887_new_n162_));
NAND2X1 NAND2X1_525 ( .A(alu__abc_40887_new_n165_), .B(alu__abc_40887_new_n163_), .Y(alu__abc_40887_new_n166_));
NAND2X1 NAND2X1_526 ( .A(alu__abc_40887_new_n172_), .B(alu__abc_40887_new_n166_), .Y(alu__abc_40887_new_n173_));
NAND2X1 NAND2X1_527 ( .A(alu__abc_40887_new_n126_), .B(alu__abc_40887_new_n130_), .Y(alu__abc_40887_new_n176_));
NAND2X1 NAND2X1_528 ( .A(alu__abc_40887_new_n147_), .B(alu__abc_40887_new_n153_), .Y(alu__abc_40887_new_n181_));
NAND2X1 NAND2X1_529 ( .A(alu__abc_40887_new_n157_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n187_));
NAND2X1 NAND2X1_53 ( .A(_abc_41234_new_n766_), .B(_abc_41234_new_n743_), .Y(_abc_41234_new_n786_));
NAND2X1 NAND2X1_530 ( .A(alu__abc_40887_new_n183_), .B(alu__abc_40887_new_n175_), .Y(alu__abc_40887_new_n190_));
NAND2X1 NAND2X1_531 ( .A(alu__abc_40887_new_n164_), .B(alu__abc_40887_new_n161_), .Y(alu__abc_40887_new_n191_));
NAND2X1 NAND2X1_532 ( .A(alu_sel_2_), .B(alu__abc_40887_new_n117_), .Y(alu__abc_40887_new_n204_));
NAND2X1 NAND2X1_533 ( .A(alu_sel_2_), .B(alu__abc_40887_new_n202_), .Y(alu__abc_40887_new_n208_));
NAND2X1 NAND2X1_534 ( .A(alu_sel_2_), .B(alu__abc_40887_new_n199_), .Y(alu__abc_40887_new_n211_));
NAND2X1 NAND2X1_535 ( .A(alu__abc_40887_new_n213_), .B(alu__abc_40887_new_n206_), .Y(alu__abc_40887_new_n214_));
NAND2X1 NAND2X1_536 ( .A(alu__abc_40887_new_n217_), .B(alu__abc_40887_new_n218_), .Y(alu__abc_40887_new_n219_));
NAND2X1 NAND2X1_537 ( .A(alu__abc_40887_new_n130_), .B(alu__abc_40887_new_n171_), .Y(alu__abc_40887_new_n236_));
NAND2X1 NAND2X1_538 ( .A(alu__abc_40887_new_n45_), .B(alu__abc_40887_new_n91_), .Y(alu__abc_40887_new_n239_));
NAND2X1 NAND2X1_539 ( .A(alu__abc_40887_new_n88_), .B(alu__abc_40887_new_n85_), .Y(alu__abc_40887_new_n266_));
NAND2X1 NAND2X1_54 ( .A(regfil_7__1_), .B(_abc_41234_new_n795_), .Y(_abc_41234_new_n796_));
NAND2X1 NAND2X1_540 ( .A(alu__abc_40887_new_n193_), .B(alu__abc_40887_new_n271_), .Y(alu__abc_40887_new_n272_));
NAND2X1 NAND2X1_541 ( .A(alu__abc_40887_new_n205_), .B(alu__abc_40887_new_n271_), .Y(alu__abc_40887_new_n278_));
NAND2X1 NAND2X1_542 ( .A(alu__abc_40887_new_n201_), .B(alu__abc_40887_new_n279_), .Y(alu__abc_40887_new_n280_));
NAND2X1 NAND2X1_543 ( .A(alu__abc_40887_new_n194_), .B(alu__abc_40887_new_n191_), .Y(alu__abc_40887_new_n286_));
NAND2X1 NAND2X1_544 ( .A(alu__abc_40887_new_n282_), .B(alu__abc_40887_new_n280_), .Y(alu__abc_40887_new_n296_));
NAND2X1 NAND2X1_545 ( .A(alu__abc_40887_new_n300_), .B(alu__abc_40887_new_n304_), .Y(alu__abc_40887_new_n305_));
NAND2X1 NAND2X1_546 ( .A(alu__abc_40887_new_n75_), .B(alu__abc_40887_new_n98_), .Y(alu__abc_40887_new_n306_));
NAND2X1 NAND2X1_547 ( .A(alu__abc_40887_new_n139_), .B(alu__abc_40887_new_n180_), .Y(alu__abc_40887_new_n309_));
NAND2X1 NAND2X1_548 ( .A(alu__abc_40887_new_n201_), .B(alu__abc_40887_new_n110_), .Y(alu__abc_40887_new_n319_));
NAND2X1 NAND2X1_549 ( .A(alu__abc_40887_new_n334_), .B(alu__abc_40887_new_n333_), .Y(alu__abc_40887_new_n335_));
NAND2X1 NAND2X1_55 ( .A(regfil_0__3_), .B(_abc_41234_new_n618_), .Y(_abc_41234_new_n812_));
NAND2X1 NAND2X1_550 ( .A(alu__abc_40887_new_n337_), .B(alu__abc_40887_new_n338_), .Y(alu__abc_40887_new_n339_));
NAND2X1 NAND2X1_551 ( .A(alu__abc_40887_new_n331_), .B(alu__abc_40887_new_n333_), .Y(alu__abc_40887_new_n341_));
NAND2X1 NAND2X1_552 ( .A(alu__abc_40887_new_n348_), .B(alu__abc_40887_new_n343_), .Y(alu_parity));
NAND2X1 NAND2X1_553 ( .A(alu__abc_40887_new_n204_), .B(alu__abc_40887_new_n249_), .Y(alu__abc_40887_new_n356_));
NAND2X1 NAND2X1_554 ( .A(alu__abc_40887_new_n204_), .B(alu__abc_40887_new_n298_), .Y(alu__abc_40887_new_n358_));
NAND2X1 NAND2X1_555 ( .A(alu__abc_40887_new_n204_), .B(alu__abc_40887_new_n331_), .Y(alu__abc_40887_new_n362_));
NAND2X1 NAND2X1_556 ( .A(alu__abc_40887_new_n204_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n365_));
NAND2X1 NAND2X1_557 ( .A(alu__abc_40887_new_n204_), .B(alu_sout), .Y(alu__abc_40887_new_n368_));
NAND2X1 NAND2X1_56 ( .A(_abc_41234_new_n824_), .B(_abc_41234_new_n817_), .Y(_abc_41234_new_n825_));
NAND2X1 NAND2X1_57 ( .A(_abc_41234_new_n832_), .B(_abc_41234_new_n513_), .Y(_abc_41234_new_n833_));
NAND2X1 NAND2X1_58 ( .A(regfil_0__4_), .B(_abc_41234_new_n618_), .Y(_abc_41234_new_n856_));
NAND2X1 NAND2X1_59 ( .A(regfil_0__0_), .B(regfil_0__1_), .Y(_abc_41234_new_n867_));
NAND2X1 NAND2X1_6 ( .A(_abc_41234_new_n516__bF_buf5), .B(_abc_41234_new_n517_), .Y(_abc_41234_new_n518_));
NAND2X1 NAND2X1_60 ( .A(regfil_0__2_), .B(regfil_0__3_), .Y(_abc_41234_new_n868_));
NAND2X1 NAND2X1_61 ( .A(_abc_41234_new_n869_), .B(_abc_41234_new_n578_), .Y(_abc_41234_new_n870_));
NAND2X1 NAND2X1_62 ( .A(_abc_41234_new_n866_), .B(_abc_41234_new_n871_), .Y(_abc_41234_new_n872_));
NAND2X1 NAND2X1_63 ( .A(regfil_0__4_), .B(_abc_41234_new_n870_), .Y(_abc_41234_new_n873_));
NAND2X1 NAND2X1_64 ( .A(_abc_41234_new_n866_), .B(_abc_41234_new_n807_), .Y(_abc_41234_new_n875_));
NAND2X1 NAND2X1_65 ( .A(regfil_0__5_), .B(_abc_41234_new_n618_), .Y(_abc_41234_new_n897_));
NAND2X1 NAND2X1_66 ( .A(_abc_41234_new_n866_), .B(_abc_41234_new_n914_), .Y(_abc_41234_new_n918_));
NAND2X1 NAND2X1_67 ( .A(_abc_41234_new_n895_), .B(_abc_41234_new_n513_), .Y(_abc_41234_new_n927_));
NAND2X1 NAND2X1_68 ( .A(_abc_41234_new_n906_), .B(_abc_41234_new_n883_), .Y(_abc_41234_new_n933_));
NAND2X1 NAND2X1_69 ( .A(regfil_0__4_), .B(regfil_0__5_), .Y(_abc_41234_new_n953_));
NAND2X1 NAND2X1_7 ( .A(_abc_41234_new_n505_), .B(_abc_41234_new_n520_), .Y(_abc_41234_new_n521_));
NAND2X1 NAND2X1_70 ( .A(_abc_41234_new_n944_), .B(_abc_41234_new_n958_), .Y(_abc_41234_new_n959_));
NAND2X1 NAND2X1_71 ( .A(_abc_41234_new_n940_), .B(_abc_41234_new_n513_), .Y(_abc_41234_new_n966_));
NAND2X1 NAND2X1_72 ( .A(regfil_0__7_), .B(_abc_41234_new_n985_), .Y(_abc_41234_new_n986_));
NAND2X1 NAND2X1_73 ( .A(_abc_41234_new_n995_), .B(_abc_41234_new_n1001_), .Y(_abc_41234_new_n1002_));
NAND2X1 NAND2X1_74 ( .A(_abc_41234_new_n1002_), .B(_abc_41234_new_n657_), .Y(_abc_41234_new_n1003_));
NAND2X1 NAND2X1_75 ( .A(_abc_41234_new_n1007_), .B(_abc_41234_new_n1003_), .Y(_abc_41234_new_n1008_));
NAND2X1 NAND2X1_76 ( .A(_abc_41234_new_n560_), .B(_abc_41234_new_n976_), .Y(_abc_41234_new_n1014_));
NAND2X1 NAND2X1_77 ( .A(opcode_4_bF_buf0_), .B(_abc_41234_new_n533_), .Y(_abc_41234_new_n1020_));
NAND2X1 NAND2X1_78 ( .A(popdes_1_), .B(_abc_41234_new_n593_), .Y(_abc_41234_new_n1032_));
NAND2X1 NAND2X1_79 ( .A(_abc_41234_new_n519_), .B(_abc_41234_new_n1033_), .Y(_abc_41234_new_n1034_));
NAND2X1 NAND2X1_8 ( .A(_abc_41234_new_n519_), .B(_abc_41234_new_n522_), .Y(_abc_41234_new_n523_));
NAND2X1 NAND2X1_80 ( .A(_abc_41234_new_n537__bF_buf1), .B(_abc_41234_new_n581_), .Y(_abc_41234_new_n1040_));
NAND2X1 NAND2X1_81 ( .A(_abc_41234_new_n1039_), .B(_abc_41234_new_n1048_), .Y(_abc_41234_new_n1049_));
NAND2X1 NAND2X1_82 ( .A(_abc_41234_new_n1050_), .B(_abc_41234_new_n617_), .Y(_abc_41234_new_n1051_));
NAND2X1 NAND2X1_83 ( .A(_abc_41234_new_n655_), .B(_abc_41234_new_n602_), .Y(_abc_41234_new_n1057_));
NAND2X1 NAND2X1_84 ( .A(_abc_41234_new_n653_), .B(_abc_41234_new_n1057_), .Y(_abc_41234_new_n1058_));
NAND2X1 NAND2X1_85 ( .A(regfil_5__1_), .B(sp_1_), .Y(_abc_41234_new_n1073_));
NAND2X1 NAND2X1_86 ( .A(regfil_5__0_), .B(sp_0_bF_buf3_), .Y(_abc_41234_new_n1075_));
NAND2X1 NAND2X1_87 ( .A(_abc_41234_new_n1083_), .B(_abc_41234_new_n1088_), .Y(_abc_41234_new_n1089_));
NAND2X1 NAND2X1_88 ( .A(_abc_41234_new_n1093_), .B(_abc_41234_new_n1097_), .Y(_abc_41234_new_n1098_));
NAND2X1 NAND2X1_89 ( .A(opcode_4_bF_buf5_), .B(opcode_5_bF_buf4_), .Y(_abc_41234_new_n1105_));
NAND2X1 NAND2X1_9 ( .A(_abc_41234_new_n515__bF_buf6), .B(_abc_41234_new_n524_), .Y(_abc_41234_new_n525_));
NAND2X1 NAND2X1_90 ( .A(regfil_5__1_), .B(regfil_3__1_), .Y(_abc_41234_new_n1118_));
NAND2X1 NAND2X1_91 ( .A(regfil_3__0_), .B(regfil_5__0_), .Y(_abc_41234_new_n1119_));
NAND2X1 NAND2X1_92 ( .A(_abc_41234_new_n1116_), .B(_abc_41234_new_n1123_), .Y(_abc_41234_new_n1124_));
NAND2X1 NAND2X1_93 ( .A(_abc_41234_new_n1127_), .B(_abc_41234_new_n1130_), .Y(_abc_41234_new_n1131_));
NAND2X1 NAND2X1_94 ( .A(_abc_41234_new_n1132_), .B(_abc_41234_new_n1133_), .Y(_abc_41234_new_n1134_));
NAND2X1 NAND2X1_95 ( .A(regfil_5__4_), .B(regfil_3__4_), .Y(_abc_41234_new_n1136_));
NAND2X1 NAND2X1_96 ( .A(regfil_1__1_), .B(regfil_5__1_), .Y(_abc_41234_new_n1157_));
NAND2X1 NAND2X1_97 ( .A(regfil_1__0_), .B(regfil_5__0_), .Y(_abc_41234_new_n1158_));
NAND2X1 NAND2X1_98 ( .A(_abc_41234_new_n1169_), .B(_abc_41234_new_n1167_), .Y(_abc_41234_new_n1170_));
NAND2X1 NAND2X1_99 ( .A(_abc_41234_new_n1173_), .B(_abc_41234_new_n1176_), .Y(_abc_41234_new_n1177_));
NAND3X1 NAND3X1_1 ( .A(_abc_41234_new_n546__bF_buf3), .B(_abc_41234_new_n619_), .C(_abc_41234_new_n622_), .Y(_abc_41234_new_n623_));
NAND3X1 NAND3X1_10 ( .A(_abc_41234_new_n567_), .B(_abc_41234_new_n716_), .C(_abc_41234_new_n713_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_0_));
NAND3X1 NAND3X1_100 ( .A(auxcar), .B(_abc_41234_new_n523__bF_buf3), .C(_abc_41234_new_n2363_), .Y(_abc_41234_new_n2391_));
NAND3X1 NAND3X1_101 ( .A(carry), .B(_abc_41234_new_n700_), .C(_abc_41234_new_n2394_), .Y(_abc_41234_new_n2395_));
NAND3X1 NAND3X1_102 ( .A(_abc_41234_new_n1013_), .B(_abc_41234_new_n1684_), .C(_abc_41234_new_n528_), .Y(_abc_41234_new_n2404_));
NAND3X1 NAND3X1_103 ( .A(_abc_41234_new_n2400_), .B(_abc_41234_new_n2408_), .C(_abc_41234_new_n2410_), .Y(_abc_41234_new_n2411_));
NAND3X1 NAND3X1_104 ( .A(carry), .B(_abc_41234_new_n1051_), .C(_abc_41234_new_n1635_), .Y(_abc_41234_new_n2413_));
NAND3X1 NAND3X1_105 ( .A(_abc_41234_new_n515__bF_buf0), .B(_abc_41234_new_n2412_), .C(_abc_41234_new_n2413_), .Y(_abc_41234_new_n2414_));
NAND3X1 NAND3X1_106 ( .A(_abc_41234_new_n2467_), .B(_abc_41234_new_n582_), .C(_abc_41234_new_n1609_), .Y(_abc_41234_new_n2468_));
NAND3X1 NAND3X1_107 ( .A(_abc_41234_new_n2185__bF_buf2), .B(_abc_41234_new_n1040__bF_buf2), .C(_abc_41234_new_n1960_), .Y(_abc_41234_new_n2483_));
NAND3X1 NAND3X1_108 ( .A(_abc_41234_new_n2470_), .B(_abc_41234_new_n2499_), .C(_abc_41234_new_n2498_), .Y(_abc_41234_new_n2500_));
NAND3X1 NAND3X1_109 ( .A(_abc_41234_new_n2476_), .B(_abc_41234_new_n2564_), .C(_abc_41234_new_n2464_), .Y(_abc_41234_new_n2565_));
NAND3X1 NAND3X1_11 ( .A(_abc_41234_new_n766_), .B(_abc_41234_new_n805_), .C(_abc_41234_new_n743_), .Y(_abc_41234_new_n806_));
NAND3X1 NAND3X1_110 ( .A(_abc_41234_new_n2398_), .B(_abc_41234_new_n2456_), .C(_abc_41234_new_n2478_), .Y(_abc_41234_new_n2589_));
NAND3X1 NAND3X1_111 ( .A(_abc_41234_new_n1046__bF_buf4), .B(_abc_41234_new_n2717_), .C(_abc_41234_new_n1643__bF_buf4), .Y(_abc_41234_new_n2718_));
NAND3X1 NAND3X1_112 ( .A(_abc_41234_new_n2718_), .B(_abc_41234_new_n2723_), .C(_abc_41234_new_n2704_), .Y(_abc_41234_new_n2724_));
NAND3X1 NAND3X1_113 ( .A(_abc_41234_new_n662_), .B(_abc_41234_new_n778_), .C(_abc_41234_new_n2505_), .Y(_abc_41234_new_n2751_));
NAND3X1 NAND3X1_114 ( .A(_abc_41234_new_n2755_), .B(_abc_41234_new_n2757_), .C(_abc_41234_new_n2751_), .Y(_abc_41234_new_n2758_));
NAND3X1 NAND3X1_115 ( .A(_abc_41234_new_n2862_), .B(_abc_41234_new_n2860_), .C(_abc_41234_new_n2861_), .Y(_abc_41234_new_n2863_));
NAND3X1 NAND3X1_116 ( .A(_abc_41234_new_n2207__bF_buf0), .B(_abc_41234_new_n2467_), .C(_abc_41234_new_n2918_), .Y(_abc_41234_new_n2919_));
NAND3X1 NAND3X1_117 ( .A(_abc_41234_new_n2474_), .B(_abc_41234_new_n2564_), .C(_abc_41234_new_n2458_), .Y(_abc_41234_new_n2943_));
NAND3X1 NAND3X1_118 ( .A(_abc_41234_new_n516__bF_buf0), .B(_abc_41234_new_n691_), .C(_abc_41234_new_n697_), .Y(_abc_41234_new_n2989_));
NAND3X1 NAND3X1_119 ( .A(_abc_41234_new_n3103_), .B(_abc_41234_new_n3107_), .C(_abc_41234_new_n2919__bF_buf0), .Y(_abc_41234_new_n3108_));
NAND3X1 NAND3X1_12 ( .A(_abc_41234_new_n809_), .B(_abc_41234_new_n828_), .C(_abc_41234_new_n811_), .Y(_abc_41234_new_n829_));
NAND3X1 NAND3X1_120 ( .A(_abc_41234_new_n2911_), .B(_abc_41234_new_n3146_), .C(_abc_41234_new_n3145_), .Y(_abc_41234_new_n3147_));
NAND3X1 NAND3X1_121 ( .A(_abc_41234_new_n2911_), .B(_abc_41234_new_n3170_), .C(_abc_41234_new_n3169_), .Y(_abc_41234_new_n3171_));
NAND3X1 NAND3X1_122 ( .A(_abc_41234_new_n2919__bF_buf0), .B(_abc_41234_new_n3181_), .C(_abc_41234_new_n3182_), .Y(_abc_41234_new_n3183_));
NAND3X1 NAND3X1_123 ( .A(_abc_41234_new_n2919__bF_buf2), .B(_abc_41234_new_n3207_), .C(_abc_41234_new_n3209_), .Y(_abc_41234_new_n3210_));
NAND3X1 NAND3X1_124 ( .A(_abc_41234_new_n3238_), .B(_abc_41234_new_n3241_), .C(_abc_41234_new_n3235_), .Y(_abc_41234_new_n3242_));
NAND3X1 NAND3X1_125 ( .A(_abc_41234_new_n3257_), .B(_abc_41234_new_n3255_), .C(_abc_41234_new_n3261_), .Y(_abc_41234_new_n3262_));
NAND3X1 NAND3X1_126 ( .A(_abc_41234_new_n3075_), .B(_abc_41234_new_n3263_), .C(_abc_41234_new_n3024_), .Y(_abc_41234_new_n3264_));
NAND3X1 NAND3X1_127 ( .A(raddrhold_10_), .B(raddrhold_11_), .C(_abc_41234_new_n3265_), .Y(_abc_41234_new_n3266_));
NAND3X1 NAND3X1_128 ( .A(_abc_41234_new_n3281_), .B(_abc_41234_new_n3287_), .C(_abc_41234_new_n3278_), .Y(_abc_41234_new_n3288_));
NAND3X1 NAND3X1_129 ( .A(_abc_41234_new_n3307_), .B(_abc_41234_new_n3301_), .C(_abc_41234_new_n3304_), .Y(_abc_41234_new_n3308_));
NAND3X1 NAND3X1_13 ( .A(_abc_41234_new_n821_), .B(_abc_41234_new_n834_), .C(_abc_41234_new_n795_), .Y(_abc_41234_new_n837_));
NAND3X1 NAND3X1_130 ( .A(raddrhold_12_), .B(raddrhold_13_), .C(_abc_41234_new_n3267_), .Y(_abc_41234_new_n3309_));
NAND3X1 NAND3X1_131 ( .A(_abc_41234_new_n3330_), .B(_abc_41234_new_n3324_), .C(_abc_41234_new_n3327_), .Y(_abc_41234_new_n3331_));
NAND3X1 NAND3X1_132 ( .A(_abc_41234_new_n3364_), .B(_abc_41234_new_n3370_), .C(_abc_41234_new_n3363_), .Y(_abc_41234_new_n3371_));
NAND3X1 NAND3X1_133 ( .A(_abc_41234_new_n1080_), .B(_abc_41234_new_n1085_), .C(_abc_41234_new_n3447_), .Y(_abc_41234_new_n3489_));
NAND3X1 NAND3X1_134 ( .A(_abc_41234_new_n1358_), .B(_abc_41234_new_n3528_), .C(_abc_41234_new_n3548_), .Y(_abc_41234_new_n3549_));
NAND3X1 NAND3X1_135 ( .A(_abc_41234_new_n1358_), .B(_abc_41234_new_n1362_), .C(_abc_41234_new_n3528_), .Y(_abc_41234_new_n3572_));
NAND3X1 NAND3X1_136 ( .A(waddrhold_10_), .B(waddrhold_11_), .C(_abc_41234_new_n3542_), .Y(_abc_41234_new_n3585_));
NAND3X1 NAND3X1_137 ( .A(waddrhold_13_), .B(waddrhold_14_), .C(_abc_41234_new_n3632_), .Y(_abc_41234_new_n3653_));
NAND3X1 NAND3X1_138 ( .A(_abc_41234_new_n3671_), .B(_abc_41234_new_n3674_), .C(_abc_41234_new_n3673_), .Y(_0waddrhold_15_0__15_));
NAND3X1 NAND3X1_139 ( .A(_abc_41234_new_n1075_), .B(_abc_41234_new_n3719_), .C(_abc_41234_new_n1108_), .Y(_abc_41234_new_n3720_));
NAND3X1 NAND3X1_14 ( .A(_abc_41234_new_n600_), .B(_abc_41234_new_n873_), .C(_abc_41234_new_n872_), .Y(_abc_41234_new_n874_));
NAND3X1 NAND3X1_140 ( .A(_abc_41234_new_n3720_), .B(_abc_41234_new_n3726_), .C(_abc_41234_new_n3725_), .Y(_abc_41234_new_n3727_));
NAND3X1 NAND3X1_141 ( .A(_abc_41234_new_n3763_), .B(_abc_41234_new_n3764_), .C(_abc_41234_new_n1108_), .Y(_abc_41234_new_n3765_));
NAND3X1 NAND3X1_142 ( .A(_abc_41234_new_n1309_), .B(_abc_41234_new_n3812_), .C(_abc_41234_new_n3814_), .Y(_abc_41234_new_n3815_));
NAND3X1 NAND3X1_143 ( .A(_abc_41234_new_n3816_), .B(_abc_41234_new_n3817_), .C(_abc_41234_new_n1325_), .Y(_abc_41234_new_n3818_));
NAND3X1 NAND3X1_144 ( .A(_abc_41234_new_n1304_), .B(_abc_41234_new_n3818_), .C(_abc_41234_new_n3815_), .Y(_abc_41234_new_n3819_));
NAND3X1 NAND3X1_145 ( .A(_abc_41234_new_n3829_), .B(_abc_41234_new_n3828_), .C(_abc_41234_new_n3850_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_5_));
NAND3X1 NAND3X1_146 ( .A(_abc_41234_new_n3854_), .B(_abc_41234_new_n3879_), .C(_abc_41234_new_n3853_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_6_));
NAND3X1 NAND3X1_147 ( .A(_abc_41234_new_n1200_), .B(_abc_41234_new_n3894_), .C(_abc_41234_new_n3893_), .Y(_abc_41234_new_n3895_));
NAND3X1 NAND3X1_148 ( .A(_abc_41234_new_n1046__bF_buf6), .B(_abc_41234_new_n4010_), .C(_abc_41234_new_n2481_), .Y(_abc_41234_new_n4011_));
NAND3X1 NAND3X1_149 ( .A(_abc_41234_new_n3914__bF_buf2), .B(_abc_41234_new_n4009_), .C(_abc_41234_new_n4011_), .Y(_abc_41234_new_n4012_));
NAND3X1 NAND3X1_15 ( .A(regfil_0__4_), .B(_abc_41234_new_n914_), .C(_abc_41234_new_n871_), .Y(_abc_41234_new_n915_));
NAND3X1 NAND3X1_150 ( .A(_abc_41234_new_n4051_), .B(_abc_41234_new_n4052_), .C(_abc_41234_new_n4050_), .Y(_abc_41234_new_n4053_));
NAND3X1 NAND3X1_151 ( .A(sp_7_), .B(sp_6_), .C(_abc_41234_new_n4013_), .Y(_abc_41234_new_n4059_));
NAND3X1 NAND3X1_152 ( .A(sp_9_), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n4107_), .Y(_abc_41234_new_n4108_));
NAND3X1 NAND3X1_153 ( .A(_abc_41234_new_n1046__bF_buf3), .B(_abc_41234_new_n4111_), .C(_abc_41234_new_n4115_), .Y(_abc_41234_new_n4116_));
NAND3X1 NAND3X1_154 ( .A(sp_0_bF_buf3_), .B(sp_10_), .C(_abc_41234_new_n4101_), .Y(_abc_41234_new_n4126_));
NAND3X1 NAND3X1_155 ( .A(_abc_41234_new_n4135_), .B(_abc_41234_new_n4136_), .C(_abc_41234_new_n4134_), .Y(_abc_41234_new_n4137_));
NAND3X1 NAND3X1_156 ( .A(_abc_41234_new_n4141_), .B(_abc_41234_new_n4142_), .C(_abc_41234_new_n4140_), .Y(_abc_41234_new_n4143_));
NAND3X1 NAND3X1_157 ( .A(sp_10_), .B(sp_11_), .C(_abc_41234_new_n4101_), .Y(_abc_41234_new_n4146_));
NAND3X1 NAND3X1_158 ( .A(_abc_41234_new_n4149_), .B(_abc_41234_new_n4150_), .C(_abc_41234_new_n4152_), .Y(_abc_41234_new_n4153_));
NAND3X1 NAND3X1_159 ( .A(_abc_41234_new_n4160_), .B(_abc_41234_new_n4161_), .C(_abc_41234_new_n4153_), .Y(_abc_41234_new_n4162_));
NAND3X1 NAND3X1_16 ( .A(_abc_41234_new_n600_), .B(_abc_41234_new_n916_), .C(_abc_41234_new_n915_), .Y(_abc_41234_new_n917_));
NAND3X1 NAND3X1_160 ( .A(sp_13_), .B(_abc_41234_new_n4010_), .C(_abc_41234_new_n2481_), .Y(_abc_41234_new_n4200_));
NAND3X1 NAND3X1_161 ( .A(_abc_41234_new_n4200_), .B(_abc_41234_new_n4201_), .C(_abc_41234_new_n4199_), .Y(_abc_41234_new_n4202_));
NAND3X1 NAND3X1_162 ( .A(sp_13_), .B(sp_14_), .C(_abc_41234_new_n4174_), .Y(_abc_41234_new_n4210_));
NAND3X1 NAND3X1_163 ( .A(sp_14_), .B(_abc_41234_new_n4010_), .C(_abc_41234_new_n2481_), .Y(_abc_41234_new_n4222_));
NAND3X1 NAND3X1_164 ( .A(_abc_41234_new_n4222_), .B(_abc_41234_new_n4223_), .C(_abc_41234_new_n4221_), .Y(_abc_41234_new_n4224_));
NAND3X1 NAND3X1_165 ( .A(_abc_41234_new_n4229_), .B(_abc_41234_new_n4230_), .C(_abc_41234_new_n4228_), .Y(_abc_41234_new_n4231_));
NAND3X1 NAND3X1_166 ( .A(_abc_41234_new_n3936_), .B(_abc_41234_new_n4235_), .C(_abc_41234_new_n4234_), .Y(_abc_41234_new_n4236_));
NAND3X1 NAND3X1_167 ( .A(_abc_41234_new_n2947__bF_buf0), .B(sp_15_), .C(_abc_41234_new_n3638_), .Y(_abc_41234_new_n4238_));
NAND3X1 NAND3X1_168 ( .A(_abc_41234_new_n2452_), .B(_abc_41234_new_n4238_), .C(_abc_41234_new_n4237_), .Y(_abc_41234_new_n4239_));
NAND3X1 NAND3X1_169 ( .A(_abc_41234_new_n4239_), .B(_abc_41234_new_n4240_), .C(_abc_41234_new_n4236_), .Y(_abc_41234_new_n4241_));
NAND3X1 NAND3X1_17 ( .A(_abc_41234_new_n600_), .B(_abc_41234_new_n956_), .C(_abc_41234_new_n955_), .Y(_abc_41234_new_n957_));
NAND3X1 NAND3X1_170 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n4242_), .C(_abc_41234_new_n4243_), .Y(_abc_41234_new_n4244_));
NAND3X1 NAND3X1_171 ( .A(_abc_41234_new_n3960_), .B(_abc_41234_new_n4242_), .C(_abc_41234_new_n4243_), .Y(_abc_41234_new_n4251_));
NAND3X1 NAND3X1_172 ( .A(_abc_41234_new_n4252_), .B(_abc_41234_new_n4253_), .C(_abc_41234_new_n4251_), .Y(_abc_41234_new_n4254_));
NAND3X1 NAND3X1_173 ( .A(_abc_41234_new_n4290_), .B(_abc_41234_new_n4280_), .C(_abc_41234_new_n4285_), .Y(_abc_41234_new_n4291_));
NAND3X1 NAND3X1_174 ( .A(_abc_41234_new_n4288_), .B(_abc_41234_new_n3935_), .C(_abc_41234_new_n1306_), .Y(_abc_41234_new_n4305_));
NAND3X1 NAND3X1_175 ( .A(_abc_41234_new_n4302_), .B(_abc_41234_new_n4304_), .C(_abc_41234_new_n4307_), .Y(_abc_41234_new_n4308_));
NAND3X1 NAND3X1_176 ( .A(_abc_41234_new_n2564_), .B(_abc_41234_new_n4310_), .C(_abc_41234_new_n1645_), .Y(_abc_41234_new_n4311_));
NAND3X1 NAND3X1_177 ( .A(_abc_41234_new_n4300_), .B(_abc_41234_new_n4314_), .C(_abc_41234_new_n4313_), .Y(_abc_41234_new_n4315_));
NAND3X1 NAND3X1_178 ( .A(_abc_41234_new_n3899_), .B(_abc_41234_new_n4417_), .C(_abc_41234_new_n4416_), .Y(_abc_41234_new_n4418_));
NAND3X1 NAND3X1_179 ( .A(pc_8_), .B(pc_9_), .C(_abc_41234_new_n4427_), .Y(_abc_41234_new_n4465_));
NAND3X1 NAND3X1_18 ( .A(_abc_41234_new_n967_), .B(_abc_41234_new_n968_), .C(_abc_41234_new_n795_), .Y(_abc_41234_new_n971_));
NAND3X1 NAND3X1_180 ( .A(_abc_41234_new_n4508_), .B(_abc_41234_new_n4512_), .C(_abc_41234_new_n4506_), .Y(_abc_41234_new_n4513_));
NAND3X1 NAND3X1_181 ( .A(_abc_41234_new_n4527_), .B(_abc_41234_new_n4530_), .C(_abc_41234_new_n4529_), .Y(_abc_41234_new_n4531_));
NAND3X1 NAND3X1_182 ( .A(pc_12_), .B(pc_13_), .C(_abc_41234_new_n4499_), .Y(_abc_41234_new_n4537_));
NAND3X1 NAND3X1_183 ( .A(_abc_41234_new_n4301_), .B(_abc_41234_new_n4537_), .C(_abc_41234_new_n4538_), .Y(_abc_41234_new_n4546_));
NAND3X1 NAND3X1_184 ( .A(_abc_41234_new_n4546_), .B(_abc_41234_new_n4548_), .C(_abc_41234_new_n4547_), .Y(_abc_41234_new_n4549_));
NAND3X1 NAND3X1_185 ( .A(_abc_41234_new_n1799_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n1797_), .Y(_abc_41234_new_n4560_));
NAND3X1 NAND3X1_186 ( .A(_abc_41234_new_n1801_), .B(_abc_41234_new_n1803_), .C(_abc_41234_new_n4295_), .Y(_abc_41234_new_n4561_));
NAND3X1 NAND3X1_187 ( .A(_abc_41234_new_n4322_), .B(_abc_41234_new_n4560_), .C(_abc_41234_new_n4561_), .Y(_abc_41234_new_n4562_));
NAND3X1 NAND3X1_188 ( .A(_abc_41234_new_n1801_), .B(_abc_41234_new_n4308_), .C(_abc_41234_new_n1803_), .Y(_abc_41234_new_n4567_));
NAND3X1 NAND3X1_189 ( .A(_abc_41234_new_n4301_), .B(_abc_41234_new_n4557_), .C(_abc_41234_new_n4556_), .Y(_abc_41234_new_n4568_));
NAND3X1 NAND3X1_19 ( .A(_abc_41234_new_n839_), .B(_abc_41234_new_n971_), .C(_abc_41234_new_n970_), .Y(_abc_41234_new_n972_));
NAND3X1 NAND3X1_190 ( .A(_abc_41234_new_n4567_), .B(_abc_41234_new_n4568_), .C(_abc_41234_new_n4569_), .Y(_abc_41234_new_n4570_));
NAND3X1 NAND3X1_191 ( .A(pc_14_), .B(pc_15_), .C(_abc_41234_new_n1796_), .Y(_abc_41234_new_n4577_));
NAND3X1 NAND3X1_192 ( .A(_abc_41234_new_n4577_), .B(_abc_41234_new_n2915_), .C(_abc_41234_new_n4576_), .Y(_abc_41234_new_n4578_));
NAND3X1 NAND3X1_193 ( .A(pc_14_), .B(pc_15_), .C(_abc_41234_new_n4555_), .Y(_abc_41234_new_n4580_));
NAND3X1 NAND3X1_194 ( .A(_abc_41234_new_n665__bF_buf3), .B(_abc_41234_new_n4579_), .C(_abc_41234_new_n4580_), .Y(_abc_41234_new_n4581_));
NAND3X1 NAND3X1_195 ( .A(pc_14_), .B(pc_15_), .C(_abc_41234_new_n1802_), .Y(_abc_41234_new_n4583_));
NAND3X1 NAND3X1_196 ( .A(_abc_41234_new_n4583_), .B(_abc_41234_new_n4295_), .C(_abc_41234_new_n4582_), .Y(_abc_41234_new_n4584_));
NAND3X1 NAND3X1_197 ( .A(_abc_41234_new_n4581_), .B(_abc_41234_new_n4584_), .C(_abc_41234_new_n4578_), .Y(_abc_41234_new_n4585_));
NAND3X1 NAND3X1_198 ( .A(_abc_41234_new_n4301_), .B(_abc_41234_new_n4579_), .C(_abc_41234_new_n4580_), .Y(_abc_41234_new_n4589_));
NAND3X1 NAND3X1_199 ( .A(_abc_41234_new_n4583_), .B(_abc_41234_new_n4308_), .C(_abc_41234_new_n4582_), .Y(_abc_41234_new_n4590_));
NAND3X1 NAND3X1_2 ( .A(_abc_41234_new_n569_), .B(_abc_41234_new_n634_), .C(_abc_41234_new_n570_), .Y(_abc_41234_new_n635_));
NAND3X1 NAND3X1_20 ( .A(_abc_41234_new_n583_), .B(_abc_41234_new_n984_), .C(_abc_41234_new_n986_), .Y(_abc_41234_new_n987_));
NAND3X1 NAND3X1_200 ( .A(_abc_41234_new_n4591_), .B(_abc_41234_new_n4589_), .C(_abc_41234_new_n4590_), .Y(_abc_41234_new_n4592_));
NAND3X1 NAND3X1_201 ( .A(_abc_41234_new_n4594_), .B(_abc_41234_new_n4593_), .C(_abc_41234_new_n4587_), .Y(_abc_41234_new_n4595_));
NAND3X1 NAND3X1_202 ( .A(_abc_41234_new_n4724_), .B(_abc_41234_new_n4718_), .C(_abc_41234_new_n4734_), .Y(_abc_41234_new_n4735_));
NAND3X1 NAND3X1_203 ( .A(_abc_41234_new_n2564_), .B(_abc_41234_new_n2938_), .C(_abc_41234_new_n4738_), .Y(_abc_41234_new_n4739_));
NAND3X1 NAND3X1_204 ( .A(opcode_5_bF_buf3_), .B(_abc_41234_new_n2450_), .C(_abc_41234_new_n4752_), .Y(_abc_41234_new_n4753_));
NAND3X1 NAND3X1_205 ( .A(_abc_41234_new_n4737_), .B(_abc_41234_new_n4755_), .C(_abc_41234_new_n4749_), .Y(_abc_41234_new_n4756_));
NAND3X1 NAND3X1_206 ( .A(_abc_41234_new_n4285_), .B(_abc_41234_new_n2920_), .C(_abc_41234_new_n4786_), .Y(_abc_41234_new_n4787_));
NAND3X1 NAND3X1_207 ( .A(_abc_41234_new_n4783_), .B(_abc_41234_new_n4787_), .C(_abc_41234_new_n4781_), .Y(_abc_41234_new_n4788_));
NAND3X1 NAND3X1_208 ( .A(_abc_41234_new_n4713_), .B(_abc_41234_new_n4727_), .C(_abc_41234_new_n4720_), .Y(_abc_41234_new_n4810_));
NAND3X1 NAND3X1_209 ( .A(_abc_41234_new_n4813_), .B(_abc_41234_new_n4815_), .C(_abc_41234_new_n4812_), .Y(_abc_41234_new_n4816_));
NAND3X1 NAND3X1_21 ( .A(_abc_41234_new_n944_), .B(regfil_0__7_), .C(_abc_41234_new_n958_), .Y(_abc_41234_new_n988_));
NAND3X1 NAND3X1_210 ( .A(_abc_41234_new_n2989_), .B(_abc_41234_new_n4834_), .C(_abc_41234_new_n4835_), .Y(_abc_41234_new_n4836_));
NAND3X1 NAND3X1_211 ( .A(_abc_41234_new_n4826_), .B(_abc_41234_new_n4837_), .C(_abc_41234_new_n4838_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_1_));
NAND3X1 NAND3X1_212 ( .A(_abc_41234_new_n4806_), .B(_abc_41234_new_n4844_), .C(_abc_41234_new_n4856_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_2_));
NAND3X1 NAND3X1_213 ( .A(_abc_41234_new_n4859_), .B(_abc_41234_new_n4867_), .C(_abc_41234_new_n4865_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_3_));
NAND3X1 NAND3X1_214 ( .A(_abc_41234_new_n4783_), .B(_abc_41234_new_n4813_), .C(_abc_41234_new_n4807_), .Y(_abc_41234_new_n4871_));
NAND3X1 NAND3X1_215 ( .A(_abc_41234_new_n4870_), .B(_abc_41234_new_n4877_), .C(_abc_41234_new_n4869_), .Y(_abc_41234_new_n4878_));
NAND3X1 NAND3X1_216 ( .A(_abc_41234_new_n4757_), .B(_abc_41234_new_n4804_), .C(_abc_41234_new_n4880_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_4_));
NAND3X1 NAND3X1_217 ( .A(_abc_41234_new_n4882_), .B(_abc_41234_new_n4883_), .C(_abc_41234_new_n4887_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_5_));
NAND3X1 NAND3X1_218 ( .A(ei), .B(_abc_41234_new_n4605_), .C(_abc_41234_new_n4890_), .Y(_abc_41234_new_n4891_));
NAND3X1 NAND3X1_219 ( .A(alu__abc_40887_new_n49_), .B(alu__abc_40887_new_n46_), .C(alu__abc_40887_new_n52_), .Y(alu__abc_40887_new_n53_));
NAND3X1 NAND3X1_22 ( .A(_abc_41234_new_n631_), .B(_abc_41234_new_n988_), .C(_abc_41234_new_n989_), .Y(_abc_41234_new_n990_));
NAND3X1 NAND3X1_220 ( .A(alu__abc_40887_new_n37_), .B(alu__abc_40887_new_n38_), .C(alu__abc_40887_new_n66_), .Y(alu__abc_40887_new_n68_));
NAND3X1 NAND3X1_221 ( .A(alu__abc_40887_new_n58_), .B(alu__abc_40887_new_n62_), .C(alu__abc_40887_new_n70_), .Y(alu__abc_40887_new_n71_));
NAND3X1 NAND3X1_222 ( .A(alu__abc_40887_new_n41_), .B(alu__abc_40887_new_n72_), .C(alu__abc_40887_new_n71_), .Y(alu__abc_40887_new_n73_));
NAND3X1 NAND3X1_223 ( .A(alu__abc_40887_new_n86_), .B(alu__abc_40887_new_n52_), .C(alu__abc_40887_new_n87_), .Y(alu__abc_40887_new_n88_));
NAND3X1 NAND3X1_224 ( .A(alu_cin), .B(alu__abc_40887_new_n45_), .C(alu__abc_40887_new_n91_), .Y(alu__abc_40887_new_n92_));
NAND3X1 NAND3X1_225 ( .A(alu__abc_40887_new_n87_), .B(alu__abc_40887_new_n93_), .C(alu__abc_40887_new_n94_), .Y(alu__abc_40887_new_n95_));
NAND3X1 NAND3X1_226 ( .A(alu__abc_40887_new_n96_), .B(alu__abc_40887_new_n99_), .C(alu__abc_40887_new_n81_), .Y(alu__abc_40887_new_n100_));
NAND3X1 NAND3X1_227 ( .A(alu__abc_40887_new_n36_), .B(alu__abc_40887_new_n38_), .C(alu__abc_40887_new_n66_), .Y(alu__abc_40887_new_n107_));
NAND3X1 NAND3X1_228 ( .A(alu__abc_40887_new_n71_), .B(alu__abc_40887_new_n79_), .C(alu__abc_40887_new_n109_), .Y(alu__abc_40887_new_n110_));
NAND3X1 NAND3X1_229 ( .A(alu__abc_40887_new_n75_), .B(alu__abc_40887_new_n98_), .C(alu__abc_40887_new_n96_), .Y(alu__abc_40887_new_n111_));
NAND3X1 NAND3X1_23 ( .A(_abc_41234_new_n987_), .B(_abc_41234_new_n1009_), .C(_abc_41234_new_n990_), .Y(_abc_41234_new_n1010_));
NAND3X1 NAND3X1_230 ( .A(alu__abc_40887_new_n101_), .B(alu__abc_40887_new_n104_), .C(alu__abc_40887_new_n113_), .Y(alu__abc_40887_new_n114_));
NAND3X1 NAND3X1_231 ( .A(alu__abc_40887_new_n36_), .B(alu__abc_40887_new_n156_), .C(alu__abc_40887_new_n155_), .Y(alu__abc_40887_new_n157_));
NAND3X1 NAND3X1_232 ( .A(alu__abc_40887_new_n42_), .B(alu__abc_40887_new_n141_), .C(alu__abc_40887_new_n135_), .Y(alu__abc_40887_new_n158_));
NAND3X1 NAND3X1_233 ( .A(alu__abc_40887_new_n52_), .B(alu__abc_40887_new_n123_), .C(alu__abc_40887_new_n163_), .Y(alu__abc_40887_new_n164_));
NAND3X1 NAND3X1_234 ( .A(alu__abc_40887_new_n49_), .B(alu__abc_40887_new_n126_), .C(alu__abc_40887_new_n130_), .Y(alu__abc_40887_new_n165_));
NAND3X1 NAND3X1_235 ( .A(alu_oprb_0_), .B(alu__abc_40887_new_n128_), .C(alu__abc_40887_new_n170_), .Y(alu__abc_40887_new_n171_));
NAND3X1 NAND3X1_236 ( .A(alu__abc_40887_new_n58_), .B(alu__abc_40887_new_n147_), .C(alu__abc_40887_new_n153_), .Y(alu__abc_40887_new_n183_));
NAND3X1 NAND3X1_237 ( .A(alu__abc_40887_new_n174_), .B(alu__abc_40887_new_n184_), .C(alu__abc_40887_new_n159_), .Y(alu__abc_40887_new_n185_));
NAND3X1 NAND3X1_238 ( .A(alu__abc_40887_new_n194_), .B(alu__abc_40887_new_n190_), .C(alu__abc_40887_new_n191_), .Y(alu__abc_40887_new_n195_));
NAND3X1 NAND3X1_239 ( .A(alu__abc_40887_new_n205_), .B(alu__abc_40887_new_n157_), .C(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n206_));
NAND3X1 NAND3X1_24 ( .A(_abc_41234_new_n1049__bF_buf4), .B(_abc_41234_new_n1053_), .C(_abc_41234_new_n1044_), .Y(_abc_41234_new_n1054_));
NAND3X1 NAND3X1_240 ( .A(alu__abc_40887_new_n215_), .B(alu__abc_40887_new_n198_), .C(alu__abc_40887_new_n114_), .Y(alu_sout));
NAND3X1 NAND3X1_241 ( .A(alu__abc_40887_new_n104_), .B(alu__abc_40887_new_n220_), .C(alu__abc_40887_new_n219_), .Y(alu__abc_40887_new_n221_));
NAND3X1 NAND3X1_242 ( .A(alu__abc_40887_new_n155_), .B(alu__abc_40887_new_n158_), .C(alu__abc_40887_new_n196_), .Y(alu__abc_40887_new_n222_));
NAND3X1 NAND3X1_243 ( .A(alu__abc_40887_new_n118_), .B(alu__abc_40887_new_n223_), .C(alu__abc_40887_new_n222_), .Y(alu__abc_40887_new_n224_));
NAND3X1 NAND3X1_244 ( .A(alu__abc_40887_new_n66_), .B(alu__abc_40887_new_n201_), .C(alu__abc_40887_new_n73_), .Y(alu__abc_40887_new_n225_));
NAND3X1 NAND3X1_245 ( .A(alu__abc_40887_new_n158_), .B(alu__abc_40887_new_n205_), .C(alu__abc_40887_new_n155_), .Y(alu__abc_40887_new_n226_));
NAND3X1 NAND3X1_246 ( .A(alu__abc_40887_new_n229_), .B(alu__abc_40887_new_n226_), .C(alu__abc_40887_new_n225_), .Y(alu__abc_40887_new_n230_));
NAND3X1 NAND3X1_247 ( .A(alu__abc_40887_new_n231_), .B(alu__abc_40887_new_n221_), .C(alu__abc_40887_new_n224_), .Y(alu__abc_40887_new_n232_));
NAND3X1 NAND3X1_248 ( .A(alu__abc_40887_new_n88_), .B(alu__abc_40887_new_n85_), .C(alu__abc_40887_new_n95_), .Y(alu__abc_40887_new_n261_));
NAND3X1 NAND3X1_249 ( .A(alu__abc_40887_new_n205_), .B(alu__abc_40887_new_n164_), .C(alu__abc_40887_new_n161_), .Y(alu__abc_40887_new_n263_));
NAND3X1 NAND3X1_25 ( .A(_abc_41234_new_n1117_), .B(_abc_41234_new_n1121_), .C(_abc_41234_new_n1122_), .Y(_abc_41234_new_n1123_));
NAND3X1 NAND3X1_250 ( .A(alu__abc_40887_new_n263_), .B(alu__abc_40887_new_n265_), .C(alu__abc_40887_new_n267_), .Y(alu__abc_40887_new_n268_));
NAND3X1 NAND3X1_251 ( .A(alu__abc_40887_new_n104_), .B(alu__abc_40887_new_n275_), .C(alu__abc_40887_new_n95_), .Y(alu__abc_40887_new_n276_));
NAND3X1 NAND3X1_252 ( .A(alu__abc_40887_new_n280_), .B(alu__abc_40887_new_n282_), .C(alu__abc_40887_new_n278_), .Y(alu__abc_40887_new_n283_));
NAND3X1 NAND3X1_253 ( .A(alu__abc_40887_new_n260_), .B(alu__abc_40887_new_n269_), .C(alu__abc_40887_new_n284_), .Y(alu__abc_40887_new_n285_));
NAND3X1 NAND3X1_254 ( .A(alu__abc_40887_new_n93_), .B(alu__abc_40887_new_n279_), .C(alu__abc_40887_new_n266_), .Y(alu__abc_40887_new_n290_));
NAND3X1 NAND3X1_255 ( .A(alu__abc_40887_new_n104_), .B(alu__abc_40887_new_n261_), .C(alu__abc_40887_new_n290_), .Y(alu__abc_40887_new_n291_));
NAND3X1 NAND3X1_256 ( .A(alu__abc_40887_new_n292_), .B(alu__abc_40887_new_n267_), .C(alu__abc_40887_new_n291_), .Y(alu__abc_40887_new_n293_));
NAND3X1 NAND3X1_257 ( .A(alu__abc_40887_new_n295_), .B(alu__abc_40887_new_n276_), .C(alu__abc_40887_new_n297_), .Y(alu__abc_40887_new_n298_));
NAND3X1 NAND3X1_258 ( .A(alu__abc_40887_new_n299_), .B(alu__abc_40887_new_n285_), .C(alu__abc_40887_new_n258_), .Y(alu__abc_40887_new_n300_));
NAND3X1 NAND3X1_259 ( .A(alu__abc_40887_new_n104_), .B(alu__abc_40887_new_n307_), .C(alu__abc_40887_new_n100_), .Y(alu__abc_40887_new_n308_));
NAND3X1 NAND3X1_26 ( .A(_abc_41234_new_n1163_), .B(_abc_41234_new_n1160_), .C(_abc_41234_new_n1166_), .Y(_abc_41234_new_n1167_));
NAND3X1 NAND3X1_260 ( .A(alu__abc_40887_new_n190_), .B(alu__abc_40887_new_n174_), .C(alu__abc_40887_new_n189_), .Y(alu__abc_40887_new_n311_));
NAND3X1 NAND3X1_261 ( .A(alu__abc_40887_new_n118_), .B(alu__abc_40887_new_n310_), .C(alu__abc_40887_new_n311_), .Y(alu__abc_40887_new_n312_));
NAND3X1 NAND3X1_262 ( .A(alu__abc_40887_new_n317_), .B(alu__abc_40887_new_n312_), .C(alu__abc_40887_new_n308_), .Y(alu__abc_40887_new_n318_));
NAND3X1 NAND3X1_263 ( .A(alu__abc_40887_new_n330_), .B(alu__abc_40887_new_n321_), .C(alu__abc_40887_new_n324_), .Y(alu__abc_40887_new_n331_));
NAND3X1 NAND3X1_264 ( .A(alu__abc_40887_new_n319_), .B(alu__abc_40887_new_n331_), .C(alu__abc_40887_new_n318_), .Y(alu__abc_40887_new_n332_));
NAND3X1 NAND3X1_265 ( .A(alu__abc_40887_new_n332_), .B(alu__abc_40887_new_n335_), .C(alu__abc_40887_new_n305_), .Y(alu__abc_40887_new_n336_));
NAND3X1 NAND3X1_266 ( .A(alu__abc_40887_new_n299_), .B(alu__abc_40887_new_n285_), .C(alu__abc_40887_new_n301_), .Y(alu__abc_40887_new_n337_));
NAND3X1 NAND3X1_267 ( .A(alu__abc_40887_new_n318_), .B(alu__abc_40887_new_n319_), .C(alu__abc_40887_new_n334_), .Y(alu__abc_40887_new_n340_));
NAND3X1 NAND3X1_268 ( .A(alu__abc_40887_new_n340_), .B(alu__abc_40887_new_n341_), .C(alu__abc_40887_new_n339_), .Y(alu__abc_40887_new_n342_));
NAND3X1 NAND3X1_269 ( .A(alu__abc_40887_new_n336_), .B(alu__abc_40887_new_n342_), .C(alu__abc_40887_new_n233_), .Y(alu__abc_40887_new_n343_));
NAND3X1 NAND3X1_27 ( .A(_abc_41234_new_n1188_), .B(_abc_41234_new_n1173_), .C(_abc_41234_new_n1176_), .Y(_abc_41234_new_n1189_));
NAND3X1 NAND3X1_270 ( .A(alu__abc_40887_new_n350_), .B(alu__abc_40887_new_n257_), .C(alu__abc_40887_new_n302_), .Y(alu__abc_40887_new_n351_));
NAND3X1 NAND3X1_271 ( .A(alu__abc_40887_new_n374_), .B(alu__abc_40887_new_n377_), .C(alu__abc_40887_new_n373_), .Y(alu_cout));
NAND3X1 NAND3X1_28 ( .A(_abc_41234_new_n1042_), .B(_abc_41234_new_n1111_), .C(_abc_41234_new_n1204_), .Y(_abc_41234_new_n1205_));
NAND3X1 NAND3X1_29 ( .A(regfil_5__5_), .B(regfil_5__4_), .C(_abc_41234_new_n1226_), .Y(_abc_41234_new_n1227_));
NAND3X1 NAND3X1_3 ( .A(_abc_41234_new_n637_), .B(_abc_41234_new_n638_), .C(_abc_41234_new_n639_), .Y(_abc_41234_new_n640_));
NAND3X1 NAND3X1_30 ( .A(regfil_5__4_), .B(regfil_5__3_bF_buf3_), .C(_abc_41234_new_n1224_), .Y(_abc_41234_new_n1229_));
NAND3X1 NAND3X1_31 ( .A(regfil_4__0_), .B(regfil_5__7_), .C(_abc_41234_new_n1230_), .Y(_abc_41234_new_n1231_));
NAND3X1 NAND3X1_32 ( .A(regfil_4__1_bF_buf0_), .B(regfil_4__2_bF_buf3_), .C(_abc_41234_new_n1246_), .Y(_abc_41234_new_n1294_));
NAND3X1 NAND3X1_33 ( .A(_abc_41234_new_n1309_), .B(_abc_41234_new_n1318_), .C(_abc_41234_new_n1320_), .Y(_abc_41234_new_n1321_));
NAND3X1 NAND3X1_34 ( .A(_abc_41234_new_n1325_), .B(_abc_41234_new_n1334_), .C(_abc_41234_new_n1335_), .Y(_abc_41234_new_n1336_));
NAND3X1 NAND3X1_35 ( .A(_abc_41234_new_n1304_), .B(_abc_41234_new_n1336_), .C(_abc_41234_new_n1321_), .Y(_abc_41234_new_n1337_));
NAND3X1 NAND3X1_36 ( .A(_abc_41234_new_n773_), .B(_abc_41234_new_n819_), .C(_abc_41234_new_n1240_), .Y(_abc_41234_new_n1348_));
NAND3X1 NAND3X1_37 ( .A(_abc_41234_new_n1218_), .B(_abc_41234_new_n1350_), .C(_abc_41234_new_n1351_), .Y(_abc_41234_new_n1352_));
NAND3X1 NAND3X1_38 ( .A(_abc_41234_new_n1108_), .B(_abc_41234_new_n1365_), .C(_abc_41234_new_n1366_), .Y(_abc_41234_new_n1367_));
NAND3X1 NAND3X1_39 ( .A(_abc_41234_new_n1357_), .B(_abc_41234_new_n1382_), .C(_abc_41234_new_n1367_), .Y(_abc_41234_new_n1383_));
NAND3X1 NAND3X1_4 ( .A(_abc_41234_new_n588_), .B(_abc_41234_new_n645_), .C(_abc_41234_new_n630_), .Y(_abc_41234_new_n646_));
NAND3X1 NAND3X1_40 ( .A(regfil_4__3_), .B(regfil_4__4_), .C(_abc_41234_new_n1353_), .Y(_abc_41234_new_n1397_));
NAND3X1 NAND3X1_41 ( .A(_abc_41234_new_n1146_), .B(_abc_41234_new_n1266_), .C(_abc_41234_new_n1413_), .Y(_abc_41234_new_n1414_));
NAND3X1 NAND3X1_42 ( .A(_abc_41234_new_n1196_), .B(_abc_41234_new_n1273_), .C(_abc_41234_new_n1430_), .Y(_abc_41234_new_n1432_));
NAND3X1 NAND3X1_43 ( .A(_abc_41234_new_n1443_), .B(_abc_41234_new_n1060_), .C(_abc_41234_new_n923_), .Y(_abc_41234_new_n1444_));
NAND3X1 NAND3X1_44 ( .A(_abc_41234_new_n1132_), .B(_abc_41234_new_n1133_), .C(_abc_41234_new_n1490_), .Y(_abc_41234_new_n1491_));
NAND3X1 NAND3X1_45 ( .A(_abc_41234_new_n1151_), .B(_abc_41234_new_n1500_), .C(_abc_41234_new_n1499_), .Y(_abc_41234_new_n1501_));
NAND3X1 NAND3X1_46 ( .A(_abc_41234_new_n1263_), .B(_abc_41234_new_n1468_), .C(_abc_41234_new_n1503_), .Y(_abc_41234_new_n1504_));
NAND3X1 NAND3X1_47 ( .A(_abc_41234_new_n1507_), .B(_abc_41234_new_n1060_), .C(_abc_41234_new_n962_), .Y(_abc_41234_new_n1508_));
NAND3X1 NAND3X1_48 ( .A(_abc_41234_new_n1108_), .B(_abc_41234_new_n1526_), .C(_abc_41234_new_n1529_), .Y(_abc_41234_new_n1530_));
NAND3X1 NAND3X1_49 ( .A(_abc_41234_new_n1263_), .B(_abc_41234_new_n1530_), .C(_abc_41234_new_n1554_), .Y(_abc_41234_new_n1555_));
NAND3X1 NAND3X1_5 ( .A(_abc_41234_new_n660__bF_buf7), .B(_abc_41234_new_n664_), .C(_abc_41234_new_n670_), .Y(_abc_41234_new_n671_));
NAND3X1 NAND3X1_50 ( .A(_abc_41234_new_n1108_), .B(_abc_41234_new_n1573_), .C(_abc_41234_new_n1572_), .Y(_abc_41234_new_n1574_));
NAND3X1 NAND3X1_51 ( .A(_abc_41234_new_n1547_), .B(_abc_41234_new_n1581_), .C(_abc_41234_new_n1544_), .Y(_abc_41234_new_n1584_));
NAND3X1 NAND3X1_52 ( .A(_abc_41234_new_n1583_), .B(_abc_41234_new_n1585_), .C(_abc_41234_new_n1584_), .Y(_abc_41234_new_n1586_));
NAND3X1 NAND3X1_53 ( .A(regfil_4__6_), .B(regfil_4__7_), .C(_abc_41234_new_n1517_), .Y(_abc_41234_new_n1598_));
NAND3X1 NAND3X1_54 ( .A(regfil_4__5_), .B(regfil_4__6_), .C(_abc_41234_new_n1452_), .Y(_abc_41234_new_n1599_));
NAND3X1 NAND3X1_55 ( .A(_abc_41234_new_n1574_), .B(_abc_41234_new_n1601_), .C(_abc_41234_new_n1597_), .Y(_abc_41234_new_n1602_));
NAND3X1 NAND3X1_56 ( .A(pc_8_), .B(pc_9_), .C(_abc_41234_new_n1620_), .Y(_abc_41234_new_n1669_));
NAND3X1 NAND3X1_57 ( .A(pc_8_), .B(pc_9_), .C(_abc_41234_new_n1651_), .Y(_abc_41234_new_n1679_));
NAND3X1 NAND3X1_58 ( .A(_abc_41234_new_n1681_), .B(_abc_41234_new_n1691_), .C(_abc_41234_new_n1643__bF_buf4), .Y(_abc_41234_new_n1692_));
NAND3X1 NAND3X1_59 ( .A(_abc_41234_new_n1643__bF_buf3), .B(_abc_41234_new_n1704_), .C(_abc_41234_new_n1719_), .Y(_abc_41234_new_n1720_));
NAND3X1 NAND3X1_6 ( .A(_abc_41234_new_n657_), .B(_abc_41234_new_n671_), .C(_abc_41234_new_n602_), .Y(_abc_41234_new_n672_));
NAND3X1 NAND3X1_60 ( .A(_abc_41234_new_n1732_), .B(_abc_41234_new_n1643__bF_buf2), .C(_abc_41234_new_n1741_), .Y(_abc_41234_new_n1742_));
NAND3X1 NAND3X1_61 ( .A(pc_11_), .B(pc_12_), .C(_abc_41234_new_n1706_), .Y(_abc_41234_new_n1749_));
NAND3X1 NAND3X1_62 ( .A(pc_11_), .B(pc_12_), .C(_abc_41234_new_n1733_), .Y(_abc_41234_new_n1754_));
NAND3X1 NAND3X1_63 ( .A(_abc_41234_new_n1757_), .B(_abc_41234_new_n1759_), .C(_abc_41234_new_n1766_), .Y(_abc_41234_new_n1767_));
NAND3X1 NAND3X1_64 ( .A(_abc_41234_new_n1643__bF_buf1), .B(_abc_41234_new_n1777_), .C(_abc_41234_new_n1788_), .Y(_abc_41234_new_n1789_));
NAND3X1 NAND3X1_65 ( .A(_abc_41234_new_n1816_), .B(_abc_41234_new_n1808_), .C(_abc_41234_new_n1806_), .Y(_abc_41234_new_n1817_));
NAND3X1 NAND3X1_66 ( .A(pc_14_), .B(_abc_41234_new_n1828_), .C(_abc_41234_new_n1802_), .Y(_abc_41234_new_n1832_));
NAND3X1 NAND3X1_67 ( .A(_abc_41234_new_n1643__bF_buf0), .B(_abc_41234_new_n1841_), .C(_abc_41234_new_n1830_), .Y(_abc_41234_new_n1842_));
NAND3X1 NAND3X1_68 ( .A(popdes_0_), .B(_abc_41234_new_n516__bF_buf2), .C(_abc_41234_new_n1851_), .Y(_abc_41234_new_n1852_));
NAND3X1 NAND3X1_69 ( .A(_abc_41234_new_n1863_), .B(_abc_41234_new_n1866_), .C(_abc_41234_new_n1861_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_0_));
NAND3X1 NAND3X1_7 ( .A(_abc_41234_new_n516__bF_buf4), .B(_abc_41234_new_n681_), .C(_abc_41234_new_n682_), .Y(_abc_41234_new_n683_));
NAND3X1 NAND3X1_70 ( .A(_abc_41234_new_n1886_), .B(_abc_41234_new_n1895_), .C(_abc_41234_new_n1885_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_2_));
NAND3X1 NAND3X1_71 ( .A(_abc_41234_new_n1899_), .B(_abc_41234_new_n1906_), .C(_abc_41234_new_n1898_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_3_));
NAND3X1 NAND3X1_72 ( .A(_abc_41234_new_n1910_), .B(_abc_41234_new_n1920_), .C(_abc_41234_new_n1909_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_4_));
NAND3X1 NAND3X1_73 ( .A(_abc_41234_new_n1924_), .B(_abc_41234_new_n1934_), .C(_abc_41234_new_n1923_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_5_));
NAND3X1 NAND3X1_74 ( .A(_abc_41234_new_n1939_), .B(_abc_41234_new_n1947_), .C(_abc_41234_new_n1938_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_6_));
NAND3X1 NAND3X1_75 ( .A(_abc_41234_new_n1951_), .B(_abc_41234_new_n1964_), .C(_abc_41234_new_n1950_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_7_));
NAND3X1 NAND3X1_76 ( .A(_abc_41234_new_n569_), .B(_abc_41234_new_n595_), .C(_abc_41234_new_n601_), .Y(_abc_41234_new_n1970_));
NAND3X1 NAND3X1_77 ( .A(_abc_41234_new_n1970_), .B(_abc_41234_new_n1971_), .C(_abc_41234_new_n1969_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_0_));
NAND3X1 NAND3X1_78 ( .A(_abc_41234_new_n1979_), .B(_abc_41234_new_n1980_), .C(_abc_41234_new_n1974_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_1_));
NAND3X1 NAND3X1_79 ( .A(_abc_41234_new_n1988_), .B(_abc_41234_new_n1989_), .C(_abc_41234_new_n1983_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_2_));
NAND3X1 NAND3X1_8 ( .A(_abc_41234_new_n540_), .B(_abc_41234_new_n683_), .C(_abc_41234_new_n686_), .Y(_abc_41234_new_n687_));
NAND3X1 NAND3X1_80 ( .A(_abc_41234_new_n1998_), .B(_abc_41234_new_n1999_), .C(_abc_41234_new_n1992_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_3_));
NAND3X1 NAND3X1_81 ( .A(_abc_41234_new_n2070_), .B(_abc_41234_new_n2078_), .C(_abc_41234_new_n2069_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_1_));
NAND3X1 NAND3X1_82 ( .A(regfil_2__1_), .B(regfil_2__2_), .C(_abc_41234_new_n2061_), .Y(_abc_41234_new_n2086_));
NAND3X1 NAND3X1_83 ( .A(_abc_41234_new_n1875_), .B(_abc_41234_new_n2085_), .C(_abc_41234_new_n2086_), .Y(_abc_41234_new_n2087_));
NAND3X1 NAND3X1_84 ( .A(_abc_41234_new_n769_), .B(_abc_41234_new_n815_), .C(_abc_41234_new_n2071_), .Y(_abc_41234_new_n2097_));
NAND3X1 NAND3X1_85 ( .A(regfil_2__3_), .B(regfil_2__4_), .C(_abc_41234_new_n2095_), .Y(_abc_41234_new_n2107_));
NAND3X1 NAND3X1_86 ( .A(popdes_0_), .B(_abc_41234_new_n1851_), .C(_abc_41234_new_n509_), .Y(_abc_41234_new_n2132_));
NAND3X1 NAND3X1_87 ( .A(_abc_41234_new_n516__bF_buf1), .B(_abc_41234_new_n660__bF_buf6), .C(_abc_41234_new_n2134_), .Y(_abc_41234_new_n2135_));
NAND3X1 NAND3X1_88 ( .A(_abc_41234_new_n515__bF_buf1), .B(_abc_41234_new_n660__bF_buf5), .C(_abc_41234_new_n1954_), .Y(_abc_41234_new_n2136_));
NAND3X1 NAND3X1_89 ( .A(_abc_41234_new_n516__bF_buf0), .B(_abc_41234_new_n660__bF_buf4), .C(_abc_41234_new_n2138_), .Y(_abc_41234_new_n2139_));
NAND3X1 NAND3X1_9 ( .A(_abc_41234_new_n688_), .B(_abc_41234_new_n708_), .C(_abc_41234_new_n704_), .Y(_abc_41234_new_n709_));
NAND3X1 NAND3X1_90 ( .A(_abc_41234_new_n1535_), .B(_abc_41234_new_n2144_), .C(_abc_41234_new_n2143_), .Y(_abc_41234_new_n2145_));
NAND3X1 NAND3X1_91 ( .A(_abc_41234_new_n2131_), .B(_abc_41234_new_n2157_), .C(_abc_41234_new_n2156_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_6_));
NAND3X1 NAND3X1_92 ( .A(_abc_41234_new_n1961_), .B(_abc_41234_new_n2169_), .C(_abc_41234_new_n2168_), .Y(_abc_41234_new_n2170_));
NAND3X1 NAND3X1_93 ( .A(_abc_41234_new_n2160_), .B(_abc_41234_new_n2161_), .C(_abc_41234_new_n2172_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_7_));
NAND3X1 NAND3X1_94 ( .A(_abc_41234_new_n2249_), .B(_abc_41234_new_n2251_), .C(_abc_41234_new_n2246_), .Y(_abc_41234_new_n2252_));
NAND3X1 NAND3X1_95 ( .A(_abc_41234_new_n2270_), .B(_abc_41234_new_n2271_), .C(_abc_41234_new_n2269_), .Y(_abc_41234_new_n2272_));
NAND3X1 NAND3X1_96 ( .A(_abc_41234_new_n2282_), .B(_abc_41234_new_n2283_), .C(_abc_41234_new_n2281_), .Y(_abc_41234_new_n2284_));
NAND3X1 NAND3X1_97 ( .A(_abc_41234_new_n2294_), .B(_abc_41234_new_n2295_), .C(_abc_41234_new_n2293_), .Y(_abc_41234_new_n2296_));
NAND3X1 NAND3X1_98 ( .A(_abc_41234_new_n2306_), .B(_abc_41234_new_n2307_), .C(_abc_41234_new_n2305_), .Y(_abc_41234_new_n2308_));
NAND3X1 NAND3X1_99 ( .A(_abc_41234_new_n501_), .B(alu_res_7_), .C(_abc_41234_new_n611_), .Y(_abc_41234_new_n2380_));
NOR2X1 NOR2X1_1 ( .A(state_5_), .B(_abc_41234_new_n501_), .Y(_abc_41234_new_n502_));
NOR2X1 NOR2X1_10 ( .A(_abc_41234_new_n532_), .B(_abc_41234_new_n525__bF_buf3), .Y(_abc_41234_new_n533_));
NOR2X1 NOR2X1_100 ( .A(_abc_41234_new_n1051_), .B(_abc_41234_new_n525__bF_buf0), .Y(_abc_41234_new_n1052_));
NOR2X1 NOR2X1_101 ( .A(_abc_41234_new_n1043_), .B(_abc_41234_new_n1054_), .Y(_abc_41234_new_n1055_));
NOR2X1 NOR2X1_102 ( .A(_abc_41234_new_n1058_), .B(_abc_41234_new_n1059_), .Y(_abc_41234_new_n1060_));
NOR2X1 NOR2X1_103 ( .A(_abc_41234_new_n818_), .B(_abc_41234_new_n1067_), .Y(_abc_41234_new_n1068_));
NOR2X1 NOR2X1_104 ( .A(regfil_5__3_bF_buf2_), .B(sp_3_), .Y(_abc_41234_new_n1070_));
NOR2X1 NOR2X1_105 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n1071_), .Y(_abc_41234_new_n1072_));
NOR2X1 NOR2X1_106 ( .A(regfil_5__1_), .B(sp_1_), .Y(_abc_41234_new_n1074_));
NOR2X1 NOR2X1_107 ( .A(_abc_41234_new_n996_), .B(_abc_41234_new_n1080_), .Y(_abc_41234_new_n1081_));
NOR2X1 NOR2X1_108 ( .A(regfil_5__7_), .B(sp_7_), .Y(_abc_41234_new_n1082_));
NOR2X1 NOR2X1_109 ( .A(_abc_41234_new_n1082_), .B(_abc_41234_new_n1081_), .Y(_abc_41234_new_n1083_));
NOR2X1 NOR2X1_11 ( .A(_abc_41234_new_n534__bF_buf5), .B(_abc_41234_new_n523__bF_buf3), .Y(_abc_41234_new_n535_));
NOR2X1 NOR2X1_110 ( .A(_abc_41234_new_n1084_), .B(_abc_41234_new_n1085_), .Y(_abc_41234_new_n1086_));
NOR2X1 NOR2X1_111 ( .A(regfil_5__6_bF_buf1_), .B(sp_6_), .Y(_abc_41234_new_n1087_));
NOR2X1 NOR2X1_112 ( .A(_abc_41234_new_n1087_), .B(_abc_41234_new_n1086_), .Y(_abc_41234_new_n1088_));
NOR2X1 NOR2X1_113 ( .A(_abc_41234_new_n848_), .B(_abc_41234_new_n1090_), .Y(_abc_41234_new_n1091_));
NOR2X1 NOR2X1_114 ( .A(regfil_5__4_), .B(sp_4_), .Y(_abc_41234_new_n1092_));
NOR2X1 NOR2X1_115 ( .A(_abc_41234_new_n1092_), .B(_abc_41234_new_n1091_), .Y(_abc_41234_new_n1093_));
NOR2X1 NOR2X1_116 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n1094_), .Y(_abc_41234_new_n1095_));
NOR2X1 NOR2X1_117 ( .A(regfil_5__5_), .B(sp_5_), .Y(_abc_41234_new_n1096_));
NOR2X1 NOR2X1_118 ( .A(_abc_41234_new_n1096_), .B(_abc_41234_new_n1095_), .Y(_abc_41234_new_n1097_));
NOR2X1 NOR2X1_119 ( .A(_abc_41234_new_n1089_), .B(_abc_41234_new_n1098_), .Y(_abc_41234_new_n1099_));
NOR2X1 NOR2X1_12 ( .A(opcode_4_bF_buf4_), .B(_abc_41234_new_n536__bF_buf5), .Y(_abc_41234_new_n537_));
NOR2X1 NOR2X1_120 ( .A(_abc_41234_new_n1105__bF_buf3), .B(_abc_41234_new_n1051_), .Y(_abc_41234_new_n1106_));
NOR2X1 NOR2X1_121 ( .A(_abc_41234_new_n1107_), .B(_abc_41234_new_n525__bF_buf3), .Y(_abc_41234_new_n1108_));
NOR2X1 NOR2X1_122 ( .A(regfil_5__3_bF_buf0_), .B(regfil_3__3_), .Y(_abc_41234_new_n1113_));
NOR2X1 NOR2X1_123 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n768_), .Y(_abc_41234_new_n1115_));
NOR2X1 NOR2X1_124 ( .A(_abc_41234_new_n1113_), .B(_abc_41234_new_n1112_), .Y(_abc_41234_new_n1117_));
NOR2X1 NOR2X1_125 ( .A(regfil_5__1_), .B(regfil_3__1_), .Y(_abc_41234_new_n1120_));
NOR2X1 NOR2X1_126 ( .A(regfil_5__7_), .B(regfil_3__7_), .Y(_abc_41234_new_n1126_));
NOR2X1 NOR2X1_127 ( .A(_abc_41234_new_n1126_), .B(_abc_41234_new_n1125_), .Y(_abc_41234_new_n1127_));
NOR2X1 NOR2X1_128 ( .A(regfil_5__6_bF_buf3_), .B(regfil_3__6_), .Y(_abc_41234_new_n1129_));
NOR2X1 NOR2X1_129 ( .A(_abc_41234_new_n1129_), .B(_abc_41234_new_n1128_), .Y(_abc_41234_new_n1130_));
NOR2X1 NOR2X1_13 ( .A(opcode_3_bF_buf2_), .B(_abc_41234_new_n546__bF_buf5), .Y(_abc_41234_new_n547_));
NOR2X1 NOR2X1_130 ( .A(_abc_41234_new_n1131_), .B(_abc_41234_new_n1134_), .Y(_abc_41234_new_n1135_));
NOR2X1 NOR2X1_131 ( .A(regfil_2__0_), .B(regfil_4__0_), .Y(_abc_41234_new_n1142_));
NOR2X1 NOR2X1_132 ( .A(_abc_41234_new_n1143_), .B(_abc_41234_new_n1144_), .Y(_abc_41234_new_n1145_));
NOR2X1 NOR2X1_133 ( .A(_abc_41234_new_n1142_), .B(_abc_41234_new_n1145_), .Y(_abc_41234_new_n1146_));
NOR2X1 NOR2X1_134 ( .A(_abc_41234_new_n1147_), .B(_abc_41234_new_n1141_), .Y(_abc_41234_new_n1148_));
NOR2X1 NOR2X1_135 ( .A(_abc_41234_new_n1150_), .B(_abc_41234_new_n1053_), .Y(_abc_41234_new_n1151_));
NOR2X1 NOR2X1_136 ( .A(_abc_41234_new_n544__bF_buf1), .B(_abc_41234_new_n1053_), .Y(_abc_41234_new_n1155_));
NOR2X1 NOR2X1_137 ( .A(regfil_1__1_), .B(regfil_5__1_), .Y(_abc_41234_new_n1159_));
NOR2X1 NOR2X1_138 ( .A(regfil_1__3_), .B(regfil_5__3_bF_buf2_), .Y(_abc_41234_new_n1162_));
NOR2X1 NOR2X1_139 ( .A(_abc_41234_new_n1162_), .B(_abc_41234_new_n1161_), .Y(_abc_41234_new_n1163_));
NOR2X1 NOR2X1_14 ( .A(_abc_41234_new_n544__bF_buf3), .B(_abc_41234_new_n548_), .Y(_abc_41234_new_n549_));
NOR2X1 NOR2X1_140 ( .A(regfil_1__2_), .B(regfil_5__2_), .Y(_abc_41234_new_n1165_));
NOR2X1 NOR2X1_141 ( .A(_abc_41234_new_n1165_), .B(_abc_41234_new_n1164_), .Y(_abc_41234_new_n1166_));
NOR2X1 NOR2X1_142 ( .A(regfil_1__7_), .B(regfil_5__7_), .Y(_abc_41234_new_n1172_));
NOR2X1 NOR2X1_143 ( .A(_abc_41234_new_n1172_), .B(_abc_41234_new_n1171_), .Y(_abc_41234_new_n1173_));
NOR2X1 NOR2X1_144 ( .A(regfil_1__6_), .B(regfil_5__6_bF_buf1_), .Y(_abc_41234_new_n1175_));
NOR2X1 NOR2X1_145 ( .A(_abc_41234_new_n1175_), .B(_abc_41234_new_n1174_), .Y(_abc_41234_new_n1176_));
NOR2X1 NOR2X1_146 ( .A(regfil_1__4_), .B(regfil_5__4_), .Y(_abc_41234_new_n1179_));
NOR2X1 NOR2X1_147 ( .A(_abc_41234_new_n1179_), .B(_abc_41234_new_n1178_), .Y(_abc_41234_new_n1180_));
NOR2X1 NOR2X1_148 ( .A(regfil_1__5_), .B(regfil_5__5_), .Y(_abc_41234_new_n1182_));
NOR2X1 NOR2X1_149 ( .A(_abc_41234_new_n1182_), .B(_abc_41234_new_n1181_), .Y(_abc_41234_new_n1183_));
NOR2X1 NOR2X1_15 ( .A(_abc_41234_new_n523__bF_buf2), .B(_abc_41234_new_n550_), .Y(_abc_41234_new_n551_));
NOR2X1 NOR2X1_150 ( .A(_abc_41234_new_n1177_), .B(_abc_41234_new_n1184_), .Y(_abc_41234_new_n1185_));
NOR2X1 NOR2X1_151 ( .A(regfil_0__0_), .B(regfil_4__0_), .Y(_abc_41234_new_n1194_));
NOR2X1 NOR2X1_152 ( .A(_abc_41234_new_n585_), .B(_abc_41234_new_n1144_), .Y(_abc_41234_new_n1195_));
NOR2X1 NOR2X1_153 ( .A(_abc_41234_new_n1194_), .B(_abc_41234_new_n1195_), .Y(_abc_41234_new_n1196_));
NOR2X1 NOR2X1_154 ( .A(_abc_41234_new_n1040__bF_buf3), .B(_abc_41234_new_n525__bF_buf2), .Y(_abc_41234_new_n1206_));
NOR2X1 NOR2X1_155 ( .A(regfil_5__0_), .B(regfil_5__1_), .Y(_abc_41234_new_n1207_));
NOR2X1 NOR2X1_156 ( .A(regfil_5__3_bF_buf1_), .B(_abc_41234_new_n1208_), .Y(_abc_41234_new_n1209_));
NOR2X1 NOR2X1_157 ( .A(regfil_5__6_bF_buf0_), .B(_abc_41234_new_n1212_), .Y(_abc_41234_new_n1213_));
NOR2X1 NOR2X1_158 ( .A(_abc_41234_new_n1217_), .B(_abc_41234_new_n525__bF_buf1), .Y(_abc_41234_new_n1218_));
NOR2X1 NOR2X1_159 ( .A(_abc_41234_new_n1221_), .B(_abc_41234_new_n719_), .Y(_abc_41234_new_n1222_));
NOR2X1 NOR2X1_16 ( .A(_abc_41234_new_n526__bF_buf1), .B(_abc_41234_new_n556_), .Y(_abc_41234_new_n557_));
NOR2X1 NOR2X1_160 ( .A(_abc_41234_new_n996_), .B(_abc_41234_new_n1084_), .Y(_abc_41234_new_n1226_));
NOR2X1 NOR2X1_161 ( .A(regfil_4__0_), .B(regfil_4__1_bF_buf2_), .Y(_abc_41234_new_n1240_));
NOR2X1 NOR2X1_162 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1245_), .Y(_abc_41234_new_n1246_));
NOR2X1 NOR2X1_163 ( .A(regfil_4__1_bF_buf0_), .B(_abc_41234_new_n1246_), .Y(_abc_41234_new_n1247_));
NOR2X1 NOR2X1_164 ( .A(regfil_4__1_bF_buf3_), .B(sp_9_), .Y(_abc_41234_new_n1250_));
NOR2X1 NOR2X1_165 ( .A(_abc_41234_new_n720_), .B(_abc_41234_new_n1251_), .Y(_abc_41234_new_n1252_));
NOR2X1 NOR2X1_166 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1255_), .Y(_abc_41234_new_n1256_));
NOR2X1 NOR2X1_167 ( .A(_abc_41234_new_n1250_), .B(_abc_41234_new_n1252_), .Y(_abc_41234_new_n1257_));
NOR2X1 NOR2X1_168 ( .A(_abc_41234_new_n1104_), .B(_abc_41234_new_n1103_), .Y(_abc_41234_new_n1260_));
NOR2X1 NOR2X1_169 ( .A(_abc_41234_new_n731_), .B(_abc_41234_new_n720_), .Y(_abc_41234_new_n1264_));
NOR2X1 NOR2X1_17 ( .A(_abc_41234_new_n558_), .B(_abc_41234_new_n525__bF_buf2), .Y(_abc_41234_new_n559_));
NOR2X1 NOR2X1_170 ( .A(regfil_2__1_), .B(regfil_4__1_bF_buf2_), .Y(_abc_41234_new_n1265_));
NOR2X1 NOR2X1_171 ( .A(_abc_41234_new_n1265_), .B(_abc_41234_new_n1264_), .Y(_abc_41234_new_n1266_));
NOR2X1 NOR2X1_172 ( .A(_abc_41234_new_n1145_), .B(_abc_41234_new_n1266_), .Y(_abc_41234_new_n1267_));
NOR2X1 NOR2X1_173 ( .A(regfil_0__1_), .B(regfil_4__1_bF_buf1_), .Y(_abc_41234_new_n1271_));
NOR2X1 NOR2X1_174 ( .A(_abc_41234_new_n739_), .B(_abc_41234_new_n720_), .Y(_abc_41234_new_n1272_));
NOR2X1 NOR2X1_175 ( .A(_abc_41234_new_n1271_), .B(_abc_41234_new_n1272_), .Y(_abc_41234_new_n1273_));
NOR2X1 NOR2X1_176 ( .A(_abc_41234_new_n1273_), .B(_abc_41234_new_n1275_), .Y(_abc_41234_new_n1276_));
NOR2X1 NOR2X1_177 ( .A(regfil_4__2_bF_buf2_), .B(sp_10_), .Y(_abc_41234_new_n1298_));
NOR2X1 NOR2X1_178 ( .A(_abc_41234_new_n1298_), .B(_abc_41234_new_n1300_), .Y(_abc_41234_new_n1301_));
NOR2X1 NOR2X1_179 ( .A(_abc_41234_new_n544__bF_buf0), .B(_abc_41234_new_n1051_), .Y(_abc_41234_new_n1303_));
NOR2X1 NOR2X1_18 ( .A(_abc_41234_new_n569_), .B(_abc_41234_new_n570_), .Y(_abc_41234_new_n571_));
NOR2X1 NOR2X1_180 ( .A(_abc_41234_new_n1310_), .B(_abc_41234_new_n1141_), .Y(_abc_41234_new_n1311_));
NOR2X1 NOR2X1_181 ( .A(regfil_2__2_), .B(regfil_4__2_bF_buf0_), .Y(_abc_41234_new_n1314_));
NOR2X1 NOR2X1_182 ( .A(_abc_41234_new_n769_), .B(_abc_41234_new_n773_), .Y(_abc_41234_new_n1315_));
NOR2X1 NOR2X1_183 ( .A(_abc_41234_new_n1313_), .B(_abc_41234_new_n1311_), .Y(_abc_41234_new_n1319_));
NOR2X1 NOR2X1_184 ( .A(_abc_41234_new_n1322_), .B(_abc_41234_new_n1051_), .Y(_abc_41234_new_n1323_));
NOR2X1 NOR2X1_185 ( .A(regfil_0__2_), .B(regfil_4__2_bF_buf3_), .Y(_abc_41234_new_n1330_));
NOR2X1 NOR2X1_186 ( .A(_abc_41234_new_n1330_), .B(_abc_41234_new_n1332_), .Y(_abc_41234_new_n1333_));
NOR2X1 NOR2X1_187 ( .A(_abc_41234_new_n1348_), .B(_abc_41234_new_n1214_), .Y(_abc_41234_new_n1349_));
NOR2X1 NOR2X1_188 ( .A(regfil_4__3_), .B(_abc_41234_new_n1353_), .Y(_abc_41234_new_n1354_));
NOR2X1 NOR2X1_189 ( .A(_abc_41234_new_n819_), .B(_abc_41234_new_n1294_), .Y(_abc_41234_new_n1355_));
NOR2X1 NOR2X1_19 ( .A(_abc_41234_new_n568_), .B(_abc_41234_new_n572_), .Y(_abc_41234_new_n573_));
NOR2X1 NOR2X1_190 ( .A(regfil_4__3_), .B(sp_11_), .Y(_abc_41234_new_n1361_));
NOR2X1 NOR2X1_191 ( .A(_abc_41234_new_n819_), .B(_abc_41234_new_n1362_), .Y(_abc_41234_new_n1363_));
NOR2X1 NOR2X1_192 ( .A(_abc_41234_new_n1361_), .B(_abc_41234_new_n1363_), .Y(_abc_41234_new_n1364_));
NOR2X1 NOR2X1_193 ( .A(_abc_41234_new_n1368_), .B(_abc_41234_new_n1051_), .Y(_abc_41234_new_n1369_));
NOR2X1 NOR2X1_194 ( .A(regfil_0__3_), .B(regfil_4__3_), .Y(_abc_41234_new_n1376_));
NOR2X1 NOR2X1_195 ( .A(_abc_41234_new_n849_), .B(_abc_41234_new_n1349_), .Y(_abc_41234_new_n1393_));
NOR2X1 NOR2X1_196 ( .A(regfil_4__4_), .B(_abc_41234_new_n1355_), .Y(_abc_41234_new_n1396_));
NOR2X1 NOR2X1_197 ( .A(_abc_41234_new_n1400_), .B(_abc_41234_new_n1296_), .Y(_abc_41234_new_n1402_));
NOR2X1 NOR2X1_198 ( .A(_abc_41234_new_n1404_), .B(_abc_41234_new_n1402_), .Y(_abc_41234_new_n1405_));
NOR2X1 NOR2X1_199 ( .A(regfil_4__4_), .B(sp_12_), .Y(_abc_41234_new_n1407_));
NOR2X1 NOR2X1_2 ( .A(_abc_41234_new_n504_), .B(_abc_41234_new_n506_), .Y(_abc_41234_new_n507_));
NOR2X1 NOR2X1_20 ( .A(_abc_41234_new_n574_), .B(_abc_41234_new_n575_), .Y(_abc_41234_new_n576_));
NOR2X1 NOR2X1_200 ( .A(_abc_41234_new_n849_), .B(_abc_41234_new_n1408_), .Y(_abc_41234_new_n1409_));
NOR2X1 NOR2X1_201 ( .A(_abc_41234_new_n1407_), .B(_abc_41234_new_n1409_), .Y(_abc_41234_new_n1410_));
NOR2X1 NOR2X1_202 ( .A(_abc_41234_new_n1371_), .B(_abc_41234_new_n1316_), .Y(_abc_41234_new_n1413_));
NOR2X1 NOR2X1_203 ( .A(regfil_2__4_), .B(regfil_4__4_), .Y(_abc_41234_new_n1419_));
NOR2X1 NOR2X1_204 ( .A(_abc_41234_new_n859_), .B(_abc_41234_new_n849_), .Y(_abc_41234_new_n1420_));
NOR2X1 NOR2X1_205 ( .A(_abc_41234_new_n1419_), .B(_abc_41234_new_n1420_), .Y(_abc_41234_new_n1421_));
NOR2X1 NOR2X1_206 ( .A(regfil_0__4_), .B(regfil_4__4_), .Y(_abc_41234_new_n1424_));
NOR2X1 NOR2X1_207 ( .A(_abc_41234_new_n1424_), .B(_abc_41234_new_n1426_), .Y(_abc_41234_new_n1427_));
NOR2X1 NOR2X1_208 ( .A(_abc_41234_new_n1378_), .B(_abc_41234_new_n1429_), .Y(_abc_41234_new_n1430_));
NOR2X1 NOR2X1_209 ( .A(regfil_4__5_), .B(_abc_41234_new_n1391_), .Y(_abc_41234_new_n1448_));
NOR2X1 NOR2X1_21 ( .A(opcode_3_bF_buf0_), .B(opcode_2_), .Y(_abc_41234_new_n579_));
NOR2X1 NOR2X1_210 ( .A(_abc_41234_new_n904_), .B(_abc_41234_new_n1392_), .Y(_abc_41234_new_n1449_));
NOR2X1 NOR2X1_211 ( .A(regfil_4__5_), .B(_abc_41234_new_n1452_), .Y(_abc_41234_new_n1453_));
NOR2X1 NOR2X1_212 ( .A(regfil_4__5_), .B(sp_13_), .Y(_abc_41234_new_n1456_));
NOR2X1 NOR2X1_213 ( .A(_abc_41234_new_n1465_), .B(_abc_41234_new_n1109_), .Y(_abc_41234_new_n1466_));
NOR2X1 NOR2X1_214 ( .A(_abc_41234_new_n1469_), .B(_abc_41234_new_n1051_), .Y(_abc_41234_new_n1470_));
NOR2X1 NOR2X1_215 ( .A(regfil_0__5_), .B(regfil_4__5_), .Y(_abc_41234_new_n1471_));
NOR2X1 NOR2X1_216 ( .A(_abc_41234_new_n1474_), .B(_abc_41234_new_n1434_), .Y(_abc_41234_new_n1475_));
NOR2X1 NOR2X1_217 ( .A(_abc_41234_new_n1471_), .B(_abc_41234_new_n1473_), .Y(_abc_41234_new_n1476_));
NOR2X1 NOR2X1_218 ( .A(regfil_2__5_), .B(regfil_4__5_), .Y(_abc_41234_new_n1483_));
NOR2X1 NOR2X1_219 ( .A(_abc_41234_new_n900_), .B(_abc_41234_new_n904_), .Y(_abc_41234_new_n1484_));
NOR2X1 NOR2X1_22 ( .A(_abc_41234_new_n526__bF_buf0), .B(_abc_41234_new_n580_), .Y(_abc_41234_new_n581_));
NOR2X1 NOR2X1_220 ( .A(_abc_41234_new_n1310_), .B(_abc_41234_new_n1493_), .Y(_abc_41234_new_n1494_));
NOR2X1 NOR2X1_221 ( .A(_abc_41234_new_n1483_), .B(_abc_41234_new_n1484_), .Y(_abc_41234_new_n1496_));
NOR2X1 NOR2X1_222 ( .A(_abc_41234_new_n904_), .B(_abc_41234_new_n1397_), .Y(_abc_41234_new_n1517_));
NOR2X1 NOR2X1_223 ( .A(regfil_4__6_), .B(sp_14_), .Y(_abc_41234_new_n1523_));
NOR2X1 NOR2X1_224 ( .A(_abc_41234_new_n1509_), .B(_abc_41234_new_n1524_), .Y(_abc_41234_new_n1525_));
NOR2X1 NOR2X1_225 ( .A(_abc_41234_new_n1523_), .B(_abc_41234_new_n1525_), .Y(_abc_41234_new_n1527_));
NOR2X1 NOR2X1_226 ( .A(regfil_2__6_), .B(regfil_4__6_), .Y(_abc_41234_new_n1534_));
NOR2X1 NOR2X1_227 ( .A(_abc_41234_new_n1535_), .B(_abc_41234_new_n1509_), .Y(_abc_41234_new_n1536_));
NOR2X1 NOR2X1_228 ( .A(_abc_41234_new_n1534_), .B(_abc_41234_new_n1536_), .Y(_abc_41234_new_n1537_));
NOR2X1 NOR2X1_229 ( .A(_abc_41234_new_n1538_), .B(_abc_41234_new_n1533_), .Y(_abc_41234_new_n1539_));
NOR2X1 NOR2X1_23 ( .A(_abc_41234_new_n582_), .B(_abc_41234_new_n525__bF_buf1), .Y(_abc_41234_new_n583_));
NOR2X1 NOR2X1_230 ( .A(regfil_0__6_), .B(regfil_4__6_), .Y(_abc_41234_new_n1545_));
NOR2X1 NOR2X1_231 ( .A(_abc_41234_new_n944_), .B(_abc_41234_new_n1509_), .Y(_abc_41234_new_n1546_));
NOR2X1 NOR2X1_232 ( .A(_abc_41234_new_n1545_), .B(_abc_41234_new_n1546_), .Y(_abc_41234_new_n1547_));
NOR2X1 NOR2X1_233 ( .A(_abc_41234_new_n1547_), .B(_abc_41234_new_n1544_), .Y(_abc_41234_new_n1548_));
NOR2X1 NOR2X1_234 ( .A(_abc_41234_new_n997_), .B(_abc_41234_new_n1513_), .Y(_abc_41234_new_n1564_));
NOR2X1 NOR2X1_235 ( .A(regfil_4__7_), .B(sp_15_), .Y(_abc_41234_new_n1568_));
NOR2X1 NOR2X1_236 ( .A(_abc_41234_new_n997_), .B(_abc_41234_new_n1569_), .Y(_abc_41234_new_n1570_));
NOR2X1 NOR2X1_237 ( .A(_abc_41234_new_n1568_), .B(_abc_41234_new_n1570_), .Y(_abc_41234_new_n1571_));
NOR2X1 NOR2X1_238 ( .A(_abc_41234_new_n1509_), .B(_abc_41234_new_n1575_), .Y(_abc_41234_new_n1576_));
NOR2X1 NOR2X1_239 ( .A(regfil_0__7_), .B(regfil_4__7_), .Y(_abc_41234_new_n1577_));
NOR2X1 NOR2X1_24 ( .A(_abc_41234_new_n585_), .B(_abc_41234_new_n577_), .Y(_abc_41234_new_n586_));
NOR2X1 NOR2X1_240 ( .A(_abc_41234_new_n1546_), .B(_abc_41234_new_n1581_), .Y(_abc_41234_new_n1582_));
NOR2X1 NOR2X1_241 ( .A(regfil_2__7_), .B(regfil_4__7_), .Y(_abc_41234_new_n1589_));
NOR2X1 NOR2X1_242 ( .A(_abc_41234_new_n993_), .B(_abc_41234_new_n997_), .Y(_abc_41234_new_n1590_));
NOR2X1 NOR2X1_243 ( .A(_abc_41234_new_n1589_), .B(_abc_41234_new_n1590_), .Y(_abc_41234_new_n1591_));
NOR2X1 NOR2X1_244 ( .A(_abc_41234_new_n515__bF_buf3), .B(_abc_41234_new_n1046__bF_buf6), .Y(_abc_41234_new_n1606_));
NOR2X1 NOR2X1_245 ( .A(_abc_41234_new_n1606_), .B(_abc_41234_new_n523__bF_buf0), .Y(_abc_41234_new_n1607_));
NOR2X1 NOR2X1_246 ( .A(_abc_41234_new_n620__bF_buf3), .B(_abc_41234_new_n580_), .Y(_abc_41234_new_n1608_));
NOR2X1 NOR2X1_247 ( .A(_abc_41234_new_n1613_), .B(_abc_41234_new_n1614_), .Y(_abc_41234_new_n1615_));
NOR2X1 NOR2X1_248 ( .A(_abc_41234_new_n1619_), .B(_abc_41234_new_n1616_), .Y(_abc_41234_new_n1620_));
NOR2X1 NOR2X1_249 ( .A(_abc_41234_new_n527_), .B(_abc_41234_new_n722__bF_buf2), .Y(_abc_41234_new_n1628_));
NOR2X1 NOR2X1_25 ( .A(_abc_41234_new_n586_), .B(_abc_41234_new_n584_), .Y(_abc_41234_new_n587_));
NOR2X1 NOR2X1_250 ( .A(_abc_41234_new_n1322_), .B(_abc_41234_new_n1629_), .Y(_abc_41234_new_n1630_));
NOR2X1 NOR2X1_251 ( .A(opcode_5_bF_buf3_), .B(_abc_41234_new_n548_), .Y(_abc_41234_new_n1634_));
NOR2X1 NOR2X1_252 ( .A(_abc_41234_new_n1627_), .B(_abc_41234_new_n1637_), .Y(_abc_41234_new_n1638_));
NOR2X1 NOR2X1_253 ( .A(_abc_41234_new_n556_), .B(_abc_41234_new_n722__bF_buf1), .Y(_abc_41234_new_n1639_));
NOR2X1 NOR2X1_254 ( .A(_abc_41234_new_n1041_), .B(_abc_41234_new_n1641_), .Y(_abc_41234_new_n1642_));
NOR2X1 NOR2X1_255 ( .A(_abc_41234_new_n539_), .B(_abc_41234_new_n1636_), .Y(_abc_41234_new_n1645_));
NOR2X1 NOR2X1_256 ( .A(_abc_41234_new_n1646_), .B(_abc_41234_new_n1647_), .Y(_abc_41234_new_n1648_));
NOR2X1 NOR2X1_257 ( .A(_abc_41234_new_n1619_), .B(_abc_41234_new_n1649_), .Y(_abc_41234_new_n1651_));
NOR2X1 NOR2X1_258 ( .A(opcode_5_bF_buf2_), .B(_abc_41234_new_n1656_), .Y(_abc_41234_new_n1657_));
NOR2X1 NOR2X1_259 ( .A(_abc_41234_new_n1661_), .B(_abc_41234_new_n1644_), .Y(_abc_41234_new_n1662_));
NOR2X1 NOR2X1_26 ( .A(_abc_41234_new_n590_), .B(_abc_41234_new_n521_), .Y(_abc_41234_new_n591_));
NOR2X1 NOR2X1_260 ( .A(opcode_5_bF_buf1_), .B(_abc_41234_new_n1701_), .Y(_abc_41234_new_n1702_));
NOR2X1 NOR2X1_261 ( .A(_abc_41234_new_n1705_), .B(_abc_41234_new_n1669_), .Y(_abc_41234_new_n1706_));
NOR2X1 NOR2X1_262 ( .A(_abc_41234_new_n1718_), .B(_abc_41234_new_n1713_), .Y(_abc_41234_new_n1719_));
NOR2X1 NOR2X1_263 ( .A(_abc_41234_new_n1705_), .B(_abc_41234_new_n1679_), .Y(_abc_41234_new_n1733_));
NOR2X1 NOR2X1_264 ( .A(opcode_5_bF_buf4_), .B(_abc_41234_new_n1761_), .Y(_abc_41234_new_n1762_));
NOR2X1 NOR2X1_265 ( .A(_abc_41234_new_n1765_), .B(_abc_41234_new_n1644_), .Y(_abc_41234_new_n1766_));
NOR2X1 NOR2X1_266 ( .A(_abc_41234_new_n1775_), .B(_abc_41234_new_n1749_), .Y(_abc_41234_new_n1796_));
NOR2X1 NOR2X1_267 ( .A(_abc_41234_new_n1775_), .B(_abc_41234_new_n1754_), .Y(_abc_41234_new_n1802_));
NOR2X1 NOR2X1_268 ( .A(_abc_41234_new_n1815_), .B(_abc_41234_new_n1644_), .Y(_abc_41234_new_n1816_));
NOR2X1 NOR2X1_269 ( .A(_abc_41234_new_n506_), .B(_abc_41234_new_n590_), .Y(_abc_41234_new_n1849_));
NOR2X1 NOR2X1_27 ( .A(reset_bF_buf7), .B(popdes_0_), .Y(_abc_41234_new_n593_));
NOR2X1 NOR2X1_270 ( .A(_abc_41234_new_n1852_), .B(_abc_41234_new_n508_), .Y(_abc_41234_new_n1853_));
NOR2X1 NOR2X1_271 ( .A(_abc_41234_new_n1856_), .B(_abc_41234_new_n525__bF_buf3), .Y(_abc_41234_new_n1857_));
NOR2X1 NOR2X1_272 ( .A(_abc_41234_new_n1857_), .B(_abc_41234_new_n1855_), .Y(_abc_41234_new_n1858_));
NOR2X1 NOR2X1_273 ( .A(_abc_41234_new_n518_), .B(_abc_41234_new_n1850_), .Y(_abc_41234_new_n1862_));
NOR2X1 NOR2X1_274 ( .A(_abc_41234_new_n1848_), .B(_abc_41234_new_n730_), .Y(_abc_41234_new_n1870_));
NOR2X1 NOR2X1_275 ( .A(regfil_3__0_), .B(regfil_3__1_), .Y(_abc_41234_new_n1871_));
NOR2X1 NOR2X1_276 ( .A(_abc_41234_new_n1871_), .B(_abc_41234_new_n1870_), .Y(_abc_41234_new_n1872_));
NOR2X1 NOR2X1_277 ( .A(_abc_41234_new_n555_), .B(_abc_41234_new_n1864_), .Y(_abc_41234_new_n1873_));
NOR2X1 NOR2X1_278 ( .A(opcode_3_bF_buf0_), .B(_abc_41234_new_n1864_), .Y(_abc_41234_new_n1875_));
NOR2X1 NOR2X1_279 ( .A(reset_bF_buf0), .B(_abc_41234_new_n1878_), .Y(_abc_41234_new_n1879_));
NOR2X1 NOR2X1_28 ( .A(popdes_1_), .B(_abc_41234_new_n508_), .Y(_abc_41234_new_n594_));
NOR2X1 NOR2X1_280 ( .A(_abc_41234_new_n814_), .B(_abc_41234_new_n1892_), .Y(_abc_41234_new_n1902_));
NOR2X1 NOR2X1_281 ( .A(regfil_3__3_), .B(_abc_41234_new_n1888_), .Y(_abc_41234_new_n1911_));
NOR2X1 NOR2X1_282 ( .A(_abc_41234_new_n858_), .B(_abc_41234_new_n1911_), .Y(_abc_41234_new_n1914_));
NOR2X1 NOR2X1_283 ( .A(_abc_41234_new_n899_), .B(_abc_41234_new_n1913_), .Y(_abc_41234_new_n1927_));
NOR2X1 NOR2X1_284 ( .A(_abc_41234_new_n899_), .B(_abc_41234_new_n1917_), .Y(_abc_41234_new_n1929_));
NOR2X1 NOR2X1_285 ( .A(regfil_3__6_), .B(_abc_41234_new_n1925_), .Y(_abc_41234_new_n1940_));
NOR2X1 NOR2X1_286 ( .A(_abc_41234_new_n1936_), .B(_abc_41234_new_n1926_), .Y(_abc_41234_new_n1941_));
NOR2X1 NOR2X1_287 ( .A(_abc_41234_new_n992_), .B(_abc_41234_new_n1943_), .Y(_abc_41234_new_n1953_));
NOR2X1 NOR2X1_288 ( .A(_abc_41234_new_n1150_), .B(_abc_41234_new_n1038_), .Y(_abc_41234_new_n1954_));
NOR2X1 NOR2X1_289 ( .A(_abc_41234_new_n1960_), .B(_abc_41234_new_n525__bF_buf2), .Y(_abc_41234_new_n1961_));
NOR2X1 NOR2X1_29 ( .A(_abc_41234_new_n526__bF_buf3), .B(_abc_41234_new_n597_), .Y(_abc_41234_new_n598_));
NOR2X1 NOR2X1_290 ( .A(_abc_41234_new_n574_), .B(_abc_41234_new_n1995_), .Y(_abc_41234_new_n2019_));
NOR2X1 NOR2X1_291 ( .A(regfil_1__6_), .B(_abc_41234_new_n2019_), .Y(_abc_41234_new_n2020_));
NOR2X1 NOR2X1_292 ( .A(_abc_41234_new_n656_), .B(_abc_41234_new_n1059_), .Y(_abc_41234_new_n2035_));
NOR2X1 NOR2X1_293 ( .A(regfil_6__0_), .B(_abc_41234_new_n2035_), .Y(_abc_41234_new_n2036_));
NOR2X1 NOR2X1_294 ( .A(regfil_2__0_), .B(_abc_41234_new_n2056_), .Y(_abc_41234_new_n2057_));
NOR2X1 NOR2X1_295 ( .A(_abc_41234_new_n1143_), .B(_abc_41234_new_n1956_), .Y(_abc_41234_new_n2058_));
NOR2X1 NOR2X1_296 ( .A(_abc_41234_new_n1887_), .B(_abc_41234_new_n2061_), .Y(_abc_41234_new_n2062_));
NOR2X1 NOR2X1_297 ( .A(regfil_2__0_), .B(regfil_2__1_), .Y(_abc_41234_new_n2071_));
NOR2X1 NOR2X1_298 ( .A(regfil_2__1_), .B(_abc_41234_new_n2061_), .Y(_abc_41234_new_n2075_));
NOR2X1 NOR2X1_299 ( .A(regfil_2__2_), .B(_abc_41234_new_n2072_), .Y(_abc_41234_new_n2082_));
NOR2X1 NOR2X1_3 ( .A(reset_bF_buf9), .B(_abc_41234_new_n510_), .Y(_abc_41234_new_n511_));
NOR2X1 NOR2X1_30 ( .A(_abc_41234_new_n596_), .B(_abc_41234_new_n601_), .Y(_abc_41234_new_n602_));
NOR2X1 NOR2X1_300 ( .A(_abc_41234_new_n815_), .B(_abc_41234_new_n2086_), .Y(_abc_41234_new_n2094_));
NOR2X1 NOR2X1_301 ( .A(_abc_41234_new_n2097_), .B(_abc_41234_new_n2056_), .Y(_abc_41234_new_n2098_));
NOR2X1 NOR2X1_302 ( .A(_abc_41234_new_n815_), .B(_abc_41234_new_n2082_), .Y(_abc_41234_new_n2099_));
NOR2X1 NOR2X1_303 ( .A(_abc_41234_new_n900_), .B(_abc_41234_new_n2107_), .Y(_abc_41234_new_n2119_));
NOR2X1 NOR2X1_304 ( .A(regfil_2__4_), .B(regfil_2__5_), .Y(_abc_41234_new_n2121_));
NOR2X1 NOR2X1_305 ( .A(reset_bF_buf9), .B(_abc_41234_new_n2132_), .Y(_abc_41234_new_n2133_));
NOR2X1 NOR2X1_306 ( .A(_abc_41234_new_n1047__bF_buf2), .B(_abc_41234_new_n1217_), .Y(_abc_41234_new_n2134_));
NOR2X1 NOR2X1_307 ( .A(reset_bF_buf8), .B(_abc_41234_new_n2136_), .Y(_abc_41234_new_n2137_));
NOR2X1 NOR2X1_308 ( .A(_abc_41234_new_n534__bF_buf4), .B(_abc_41234_new_n1960_), .Y(_abc_41234_new_n2138_));
NOR2X1 NOR2X1_309 ( .A(_abc_41234_new_n1143_), .B(_abc_41234_new_n731_), .Y(_abc_41234_new_n2140_));
NOR2X1 NOR2X1_31 ( .A(reset_bF_buf6), .B(_abc_41234_new_n607_), .Y(_abc_41234_new_n608_));
NOR2X1 NOR2X1_310 ( .A(_abc_41234_new_n769_), .B(_abc_41234_new_n815_), .Y(_abc_41234_new_n2141_));
NOR2X1 NOR2X1_311 ( .A(_abc_41234_new_n859_), .B(_abc_41234_new_n900_), .Y(_abc_41234_new_n2144_));
NOR2X1 NOR2X1_312 ( .A(_abc_41234_new_n1535_), .B(_abc_41234_new_n2122_), .Y(_abc_41234_new_n2150_));
NOR2X1 NOR2X1_313 ( .A(regfil_2__6_), .B(_abc_41234_new_n2122_), .Y(_abc_41234_new_n2163_));
NOR2X1 NOR2X1_314 ( .A(_abc_41234_new_n1535_), .B(_abc_41234_new_n2166_), .Y(_abc_41234_new_n2167_));
NOR2X1 NOR2X1_315 ( .A(opcode_1_), .B(_abc_41234_new_n546__bF_buf3), .Y(_abc_41234_new_n2174_));
NOR2X1 NOR2X1_316 ( .A(_abc_41234_new_n2178_), .B(_abc_41234_new_n523__bF_buf1), .Y(_abc_41234_new_n2179_));
NOR2X1 NOR2X1_317 ( .A(opcode_4_bF_buf2_), .B(_abc_41234_new_n2185__bF_buf5), .Y(_abc_41234_new_n2186_));
NOR2X1 NOR2X1_318 ( .A(_abc_41234_new_n2187_), .B(_abc_41234_new_n2186_), .Y(_abc_41234_new_n2188_));
NOR2X1 NOR2X1_319 ( .A(opcode_6_), .B(_abc_41234_new_n1045_), .Y(_abc_41234_new_n2189_));
NOR2X1 NOR2X1_32 ( .A(_abc_41234_new_n610_), .B(_abc_41234_new_n504_), .Y(_abc_41234_new_n611_));
NOR2X1 NOR2X1_320 ( .A(_abc_41234_new_n534__bF_buf1), .B(_abc_41234_new_n2207__bF_buf3), .Y(_abc_41234_new_n2208_));
NOR2X1 NOR2X1_321 ( .A(_abc_41234_new_n565_), .B(_abc_41234_new_n2214_), .Y(_abc_41234_new_n2217_));
NOR2X1 NOR2X1_322 ( .A(reset_bF_buf7), .B(_abc_41234_new_n2214_), .Y(_abc_41234_new_n2223_));
NOR2X1 NOR2X1_323 ( .A(_abc_41234_new_n2190__bF_buf2), .B(_abc_41234_new_n523__bF_buf3), .Y(_abc_41234_new_n2224_));
NOR2X1 NOR2X1_324 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n555_), .Y(_abc_41234_new_n2245_));
NOR2X1 NOR2X1_325 ( .A(opcode_4_bF_buf1_), .B(opcode_3_bF_buf2_), .Y(_abc_41234_new_n2247_));
NOR2X1 NOR2X1_326 ( .A(opcode_4_bF_buf0_), .B(_abc_41234_new_n555_), .Y(_abc_41234_new_n2248_));
NOR2X1 NOR2X1_327 ( .A(opcode_3_bF_buf1_), .B(_abc_41234_new_n529_), .Y(_abc_41234_new_n2250_));
NOR2X1 NOR2X1_328 ( .A(reset_bF_buf6), .B(_abc_41234_new_n2262_), .Y(_abc_41234_new_n2263_));
NOR2X1 NOR2X1_329 ( .A(_abc_41234_new_n2317_), .B(_abc_41234_new_n2319_), .Y(_abc_41234_new_n2320_));
NOR2X1 NOR2X1_33 ( .A(_abc_41234_new_n518_), .B(_abc_41234_new_n612_), .Y(_abc_41234_new_n613_));
NOR2X1 NOR2X1_330 ( .A(_abc_41234_new_n2320_), .B(_abc_41234_new_n2325_), .Y(_abc_41234_new_n2326_));
NOR2X1 NOR2X1_331 ( .A(_abc_41234_new_n2330_), .B(_abc_41234_new_n2332_), .Y(_abc_41234_new_n2333_));
NOR2X1 NOR2X1_332 ( .A(_abc_41234_new_n2333_), .B(_abc_41234_new_n2337_), .Y(_abc_41234_new_n2338_));
NOR2X1 NOR2X1_333 ( .A(_abc_41234_new_n2354_), .B(_abc_41234_new_n2355_), .Y(_abc_41234_new_n2356_));
NOR2X1 NOR2X1_334 ( .A(_abc_41234_new_n2353_), .B(_abc_41234_new_n2356_), .Y(_abc_41234_new_n2357_));
NOR2X1 NOR2X1_335 ( .A(_abc_41234_new_n2353_), .B(_abc_41234_new_n2212_), .Y(_abc_41234_new_n2358_));
NOR2X1 NOR2X1_336 ( .A(_abc_41234_new_n1577_), .B(_abc_41234_new_n2398_), .Y(_abc_41234_new_n2399_));
NOR2X1 NOR2X1_337 ( .A(_abc_41234_new_n1568_), .B(_abc_41234_new_n1107_), .Y(_abc_41234_new_n2409_));
NOR2X1 NOR2X1_338 ( .A(_abc_41234_new_n610_), .B(_abc_41234_new_n696_), .Y(_abc_41234_new_n2427_));
NOR2X1 NOR2X1_339 ( .A(_abc_41234_new_n1627_), .B(_abc_41234_new_n1630_), .Y(_abc_41234_new_n2458_));
NOR2X1 NOR2X1_34 ( .A(opcode_1_), .B(_abc_41234_new_n616_), .Y(_abc_41234_new_n617_));
NOR2X1 NOR2X1_340 ( .A(_abc_41234_new_n2457_), .B(_abc_41234_new_n2459_), .Y(_abc_41234_new_n2460_));
NOR2X1 NOR2X1_341 ( .A(_abc_41234_new_n722__bF_buf0), .B(_abc_41234_new_n580_), .Y(_abc_41234_new_n2462_));
NOR2X1 NOR2X1_342 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n2463_), .Y(_abc_41234_new_n2464_));
NOR2X1 NOR2X1_343 ( .A(_abc_41234_new_n597_), .B(_abc_41234_new_n620__bF_buf5), .Y(_abc_41234_new_n2466_));
NOR2X1 NOR2X1_344 ( .A(opcode_2_), .B(_abc_41234_new_n620__bF_buf4), .Y(_abc_41234_new_n2469_));
NOR2X1 NOR2X1_345 ( .A(_abc_41234_new_n2475_), .B(_abc_41234_new_n2473_), .Y(_abc_41234_new_n2476_));
NOR2X1 NOR2X1_346 ( .A(_abc_41234_new_n2465_), .B(_abc_41234_new_n2477_), .Y(_abc_41234_new_n2478_));
NOR2X1 NOR2X1_347 ( .A(_abc_41234_new_n1639__bF_buf2), .B(_abc_41234_new_n1637_), .Y(_abc_41234_new_n2481_));
NOR2X1 NOR2X1_348 ( .A(_abc_41234_new_n2483_), .B(_abc_41234_new_n2482_), .Y(_abc_41234_new_n2484_));
NOR2X1 NOR2X1_349 ( .A(_abc_41234_new_n2487_), .B(_abc_41234_new_n2492_), .Y(_abc_41234_new_n2493_));
NOR2X1 NOR2X1_35 ( .A(opcode_1_), .B(opcode_0_), .Y(_abc_41234_new_n618_));
NOR2X1 NOR2X1_350 ( .A(_abc_41234_new_n2261_), .B(_abc_41234_new_n1004_), .Y(_abc_41234_new_n2511_));
NOR2X1 NOR2X1_351 ( .A(_abc_41234_new_n693_), .B(_abc_41234_new_n2512_), .Y(_abc_41234_new_n2513_));
NOR2X1 NOR2X1_352 ( .A(_abc_41234_new_n604_), .B(_abc_41234_new_n694_), .Y(_abc_41234_new_n2514_));
NOR2X1 NOR2X1_353 ( .A(_abc_41234_new_n2513_), .B(_abc_41234_new_n2516_), .Y(_abc_41234_new_n2517_));
NOR2X1 NOR2X1_354 ( .A(_abc_41234_new_n604_), .B(_abc_41234_new_n610_), .Y(_abc_41234_new_n2518_));
NOR2X1 NOR2X1_355 ( .A(_abc_41234_new_n2522_), .B(_abc_41234_new_n2520_), .Y(_abc_41234_new_n2523_));
NOR2X1 NOR2X1_356 ( .A(_abc_41234_new_n681_), .B(_abc_41234_new_n2526_), .Y(_abc_41234_new_n2530_));
NOR2X1 NOR2X1_357 ( .A(waitr), .B(_abc_41234_new_n2526_), .Y(_abc_41234_new_n2533_));
NOR2X1 NOR2X1_358 ( .A(_abc_41234_new_n2461_), .B(_abc_41234_new_n2479_), .Y(_abc_41234_new_n2538_));
NOR2X1 NOR2X1_359 ( .A(_abc_41234_new_n2207__bF_buf2), .B(_abc_41234_new_n669__bF_buf0), .Y(_abc_41234_new_n2541_));
NOR2X1 NOR2X1_36 ( .A(_abc_41234_new_n599_), .B(_abc_41234_new_n525__bF_buf2), .Y(_abc_41234_new_n631_));
NOR2X1 NOR2X1_360 ( .A(_abc_41234_new_n2545_), .B(_abc_41234_new_n2544_), .Y(_abc_41234_new_n2546_));
NOR2X1 NOR2X1_361 ( .A(statesel_0_), .B(_abc_41234_new_n2556_), .Y(_abc_41234_new_n2557_));
NOR2X1 NOR2X1_362 ( .A(statesel_1_), .B(_abc_41234_new_n2455_), .Y(_abc_41234_new_n2558_));
NOR2X1 NOR2X1_363 ( .A(_abc_41234_new_n2557_), .B(_abc_41234_new_n2558_), .Y(_abc_41234_new_n2559_));
NOR2X1 NOR2X1_364 ( .A(opcode_2_), .B(_abc_41234_new_n526__bF_buf2), .Y(_abc_41234_new_n2563_));
NOR2X1 NOR2X1_365 ( .A(_abc_41234_new_n2455_), .B(_abc_41234_new_n2556_), .Y(_abc_41234_new_n2578_));
NOR2X1 NOR2X1_366 ( .A(_abc_41234_new_n2591_), .B(_abc_41234_new_n2544_), .Y(_abc_41234_new_n2592_));
NOR2X1 NOR2X1_367 ( .A(_abc_41234_new_n2533_), .B(_abc_41234_new_n2525_), .Y(_abc_41234_new_n2600_));
NOR2X1 NOR2X1_368 ( .A(statesel_3_), .B(_abc_41234_new_n2581_), .Y(_abc_41234_new_n2601_));
NOR2X1 NOR2X1_369 ( .A(_abc_41234_new_n2602_), .B(_abc_41234_new_n2582_), .Y(_abc_41234_new_n2603_));
NOR2X1 NOR2X1_37 ( .A(regfil_1__5_), .B(regfil_1__4_), .Y(_abc_41234_new_n639_));
NOR2X1 NOR2X1_370 ( .A(_abc_41234_new_n2580_), .B(_abc_41234_new_n2577_), .Y(_abc_41234_new_n2605_));
NOR2X1 NOR2X1_371 ( .A(_abc_41234_new_n2581_), .B(_abc_41234_new_n2588_), .Y(_abc_41234_new_n2620_));
NOR2X1 NOR2X1_372 ( .A(_abc_41234_new_n2582_), .B(_abc_41234_new_n2621_), .Y(_abc_41234_new_n2622_));
NOR2X1 NOR2X1_373 ( .A(statesel_4_), .B(_abc_41234_new_n2622_), .Y(_abc_41234_new_n2623_));
NOR2X1 NOR2X1_374 ( .A(statesel_5_), .B(_abc_41234_new_n2611_), .Y(_abc_41234_new_n2639_));
NOR2X1 NOR2X1_375 ( .A(_abc_41234_new_n2640_), .B(_abc_41234_new_n2638_), .Y(_abc_41234_new_n2641_));
NOR2X1 NOR2X1_376 ( .A(_abc_41234_new_n2672_), .B(_abc_41234_new_n2673_), .Y(_abc_41234_new_n2674_));
NOR2X1 NOR2X1_377 ( .A(reset_bF_buf2), .B(_abc_41234_new_n2674_), .Y(_abc_41234_new_n2675_));
NOR2X1 NOR2X1_378 ( .A(_abc_41234_new_n1221_), .B(_abc_41234_new_n544__bF_buf3), .Y(_abc_41234_new_n2677_));
NOR2X1 NOR2X1_379 ( .A(_abc_41234_new_n2504_), .B(_abc_41234_new_n2205_), .Y(_abc_41234_new_n2681_));
NOR2X1 NOR2X1_38 ( .A(_abc_41234_new_n640_), .B(_abc_41234_new_n636_), .Y(_abc_41234_new_n641_));
NOR2X1 NOR2X1_380 ( .A(_abc_41234_new_n1047__bF_buf2), .B(_abc_41234_new_n1643__bF_buf5), .Y(_abc_41234_new_n2702_));
NOR2X1 NOR2X1_381 ( .A(pc_1_), .B(pc_0_), .Y(_abc_41234_new_n2705_));
NOR2X1 NOR2X1_382 ( .A(opcode_4_bF_buf4_), .B(_abc_41234_new_n1682_), .Y(_abc_41234_new_n2710_));
NOR2X1 NOR2X1_383 ( .A(_abc_41234_new_n570_), .B(_abc_41234_new_n1322_), .Y(_abc_41234_new_n2711_));
NOR2X1 NOR2X1_384 ( .A(_abc_41234_new_n1614_), .B(_abc_41234_new_n1646_), .Y(_abc_41234_new_n2732_));
NOR2X1 NOR2X1_385 ( .A(pc_2_), .B(pc_1_), .Y(_abc_41234_new_n2737_));
NOR2X1 NOR2X1_386 ( .A(_abc_41234_new_n818_), .B(_abc_41234_new_n544__bF_buf2), .Y(_abc_41234_new_n2765_));
NOR2X1 NOR2X1_387 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n544__bF_buf1), .Y(_abc_41234_new_n2825_));
NOR2X1 NOR2X1_388 ( .A(_abc_41234_new_n2865_), .B(_abc_41234_new_n1729_), .Y(_abc_41234_new_n2866_));
NOR2X1 NOR2X1_389 ( .A(_abc_41234_new_n2887_), .B(_abc_41234_new_n2894_), .Y(_abc_41234_new_n2895_));
NOR2X1 NOR2X1_39 ( .A(_abc_41234_new_n583_), .B(_abc_41234_new_n631_), .Y(_abc_41234_new_n647_));
NOR2X1 NOR2X1_390 ( .A(_abc_41234_new_n2881_), .B(_abc_41234_new_n1608_), .Y(_abc_41234_new_n2899_));
NOR2X1 NOR2X1_391 ( .A(_abc_41234_new_n2504_), .B(_abc_41234_new_n1002_), .Y(_abc_41234_new_n2901_));
NOR2X1 NOR2X1_392 ( .A(_abc_41234_new_n607_), .B(_abc_41234_new_n698_), .Y(_abc_41234_new_n2911_));
NOR2X1 NOR2X1_393 ( .A(regfil_5__0_), .B(_abc_41234_new_n668__bF_buf5), .Y(_abc_41234_new_n2922_));
NOR2X1 NOR2X1_394 ( .A(_abc_41234_new_n2207__bF_buf3), .B(_abc_41234_new_n2922_), .Y(_abc_41234_new_n2923_));
NOR2X1 NOR2X1_395 ( .A(_abc_41234_new_n2925_), .B(_abc_41234_new_n2920_), .Y(_abc_41234_new_n2926_));
NOR2X1 NOR2X1_396 ( .A(_abc_41234_new_n2933_), .B(_abc_41234_new_n2935_), .Y(_abc_41234_new_n2936_));
NOR2X1 NOR2X1_397 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n1323_), .Y(_abc_41234_new_n2938_));
NOR2X1 NOR2X1_398 ( .A(opcode_5_bF_buf2_), .B(_abc_41234_new_n2456_), .Y(_abc_41234_new_n2939_));
NOR2X1 NOR2X1_399 ( .A(_abc_41234_new_n2941_), .B(_abc_41234_new_n2937_), .Y(_abc_41234_new_n2942_));
NOR2X1 NOR2X1_4 ( .A(opcode_6_), .B(opcode_7_), .Y(_abc_41234_new_n515_));
NOR2X1 NOR2X1_40 ( .A(_abc_41234_new_n606_), .B(_abc_41234_new_n609_), .Y(_abc_41234_new_n650_));
NOR2X1 NOR2X1_400 ( .A(_abc_41234_new_n2473_), .B(_abc_41234_new_n2943_), .Y(_abc_41234_new_n2944_));
NOR2X1 NOR2X1_401 ( .A(_abc_41234_new_n2910_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n2946_));
NOR2X1 NOR2X1_402 ( .A(_abc_41234_new_n668__bF_buf4), .B(_abc_41234_new_n2950_), .Y(_abc_41234_new_n2951_));
NOR2X1 NOR2X1_403 ( .A(_abc_41234_new_n2951__bF_buf3), .B(_abc_41234_new_n2930_), .Y(_abc_41234_new_n2952_));
NOR2X1 NOR2X1_404 ( .A(_abc_41234_new_n2968_), .B(_abc_41234_new_n2920_), .Y(_abc_41234_new_n2969_));
NOR2X1 NOR2X1_405 ( .A(_abc_41234_new_n2965_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n2972_));
NOR2X1 NOR2X1_406 ( .A(raddrhold_0_), .B(raddrhold_1_), .Y(_abc_41234_new_n2986_));
NOR2X1 NOR2X1_407 ( .A(_abc_41234_new_n2910_), .B(_abc_41234_new_n2965_), .Y(_abc_41234_new_n2987_));
NOR2X1 NOR2X1_408 ( .A(_abc_41234_new_n2986_), .B(_abc_41234_new_n2987_), .Y(_abc_41234_new_n2988_));
NOR2X1 NOR2X1_409 ( .A(_abc_41234_new_n501_), .B(_abc_41234_new_n2989_), .Y(_abc_41234_new_n2990_));
NOR2X1 NOR2X1_41 ( .A(_abc_41234_new_n652_), .B(_abc_41234_new_n648_), .Y(_abc_41234_new_n653_));
NOR2X1 NOR2X1_410 ( .A(regfil_5__2_), .B(_abc_41234_new_n668__bF_buf0), .Y(_abc_41234_new_n2993_));
NOR2X1 NOR2X1_411 ( .A(_abc_41234_new_n2207__bF_buf0), .B(_abc_41234_new_n2993_), .Y(_abc_41234_new_n2997_));
NOR2X1 NOR2X1_412 ( .A(_abc_41234_new_n3003_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3010_));
NOR2X1 NOR2X1_413 ( .A(raddrhold_2_), .B(_abc_41234_new_n2987_), .Y(_abc_41234_new_n3017_));
NOR2X1 NOR2X1_414 ( .A(_abc_41234_new_n3017_), .B(_abc_41234_new_n3019_), .Y(_abc_41234_new_n3020_));
NOR2X1 NOR2X1_415 ( .A(_abc_41234_new_n3023_), .B(_abc_41234_new_n3018_), .Y(_abc_41234_new_n3024_));
NOR2X1 NOR2X1_416 ( .A(_abc_41234_new_n3024_), .B(_abc_41234_new_n3025_), .Y(_abc_41234_new_n3026_));
NOR2X1 NOR2X1_417 ( .A(regfil_5__3_bF_buf0_), .B(_abc_41234_new_n668__bF_buf5), .Y(_abc_41234_new_n3027_));
NOR2X1 NOR2X1_418 ( .A(_abc_41234_new_n2207__bF_buf2), .B(_abc_41234_new_n3027_), .Y(_abc_41234_new_n3029_));
NOR2X1 NOR2X1_419 ( .A(_abc_41234_new_n3023_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3041_));
NOR2X1 NOR2X1_42 ( .A(_abc_41234_new_n504_), .B(_abc_41234_new_n659_), .Y(_abc_41234_new_n660_));
NOR2X1 NOR2X1_420 ( .A(regfil_5__4_), .B(_abc_41234_new_n668__bF_buf4), .Y(_abc_41234_new_n3052_));
NOR2X1 NOR2X1_421 ( .A(_abc_41234_new_n2207__bF_buf0), .B(_abc_41234_new_n3052_), .Y(_abc_41234_new_n3054_));
NOR2X1 NOR2X1_422 ( .A(_abc_41234_new_n3049_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3066_));
NOR2X1 NOR2X1_423 ( .A(_abc_41234_new_n3049_), .B(_abc_41234_new_n3074_), .Y(_abc_41234_new_n3075_));
NOR2X1 NOR2X1_424 ( .A(regfil_5__5_), .B(_abc_41234_new_n668__bF_buf3), .Y(_abc_41234_new_n3079_));
NOR2X1 NOR2X1_425 ( .A(_abc_41234_new_n2207__bF_buf2), .B(_abc_41234_new_n3079_), .Y(_abc_41234_new_n3081_));
NOR2X1 NOR2X1_426 ( .A(_abc_41234_new_n3074_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3093_));
NOR2X1 NOR2X1_427 ( .A(_abc_41234_new_n3101_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3110_));
NOR2X1 NOR2X1_428 ( .A(regfil_5__7_), .B(_abc_41234_new_n668__bF_buf0), .Y(_abc_41234_new_n3127_));
NOR2X1 NOR2X1_429 ( .A(_abc_41234_new_n2207__bF_buf0), .B(_abc_41234_new_n3127_), .Y(_abc_41234_new_n3128_));
NOR2X1 NOR2X1_43 ( .A(opcode_7_), .B(_abc_41234_new_n661_), .Y(_abc_41234_new_n662_));
NOR2X1 NOR2X1_430 ( .A(_abc_41234_new_n3130_), .B(_abc_41234_new_n2920_), .Y(_abc_41234_new_n3131_));
NOR2X1 NOR2X1_431 ( .A(_abc_41234_new_n3125_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3134_));
NOR2X1 NOR2X1_432 ( .A(regfil_4__0_), .B(_abc_41234_new_n668__bF_buf5), .Y(_abc_41234_new_n3152_));
NOR2X1 NOR2X1_433 ( .A(_abc_41234_new_n2207__bF_buf3), .B(_abc_41234_new_n3152_), .Y(_abc_41234_new_n3153_));
NOR2X1 NOR2X1_434 ( .A(_abc_41234_new_n3155_), .B(_abc_41234_new_n2920_), .Y(_abc_41234_new_n3156_));
NOR2X1 NOR2X1_435 ( .A(_abc_41234_new_n3151_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3159_));
NOR2X1 NOR2X1_436 ( .A(_abc_41234_new_n3175_), .B(_abc_41234_new_n3169_), .Y(_abc_41234_new_n3177_));
NOR2X1 NOR2X1_437 ( .A(_abc_41234_new_n2959__bF_buf0), .B(_abc_41234_new_n3177_), .Y(_abc_41234_new_n3178_));
NOR2X1 NOR2X1_438 ( .A(regfil_4__1_bF_buf2_), .B(_abc_41234_new_n668__bF_buf4), .Y(_abc_41234_new_n3179_));
NOR2X1 NOR2X1_439 ( .A(_abc_41234_new_n2207__bF_buf2), .B(_abc_41234_new_n3179_), .Y(_abc_41234_new_n3180_));
NOR2X1 NOR2X1_44 ( .A(reset_bF_buf5), .B(_abc_41234_new_n663_), .Y(_abc_41234_new_n664_));
NOR2X1 NOR2X1_440 ( .A(_abc_41234_new_n3175_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3191_));
NOR2X1 NOR2X1_441 ( .A(_abc_41234_new_n3200_), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3201_));
NOR2X1 NOR2X1_442 ( .A(regfil_4__2_bF_buf2_), .B(_abc_41234_new_n668__bF_buf3), .Y(_abc_41234_new_n3205_));
NOR2X1 NOR2X1_443 ( .A(_abc_41234_new_n2207__bF_buf1), .B(_abc_41234_new_n3205_), .Y(_abc_41234_new_n3206_));
NOR2X1 NOR2X1_444 ( .A(_abc_41234_new_n2190__bF_buf1), .B(_abc_41234_new_n3213_), .Y(_abc_41234_new_n3214_));
NOR2X1 NOR2X1_445 ( .A(raddrhold_10_), .B(_abc_41234_new_n3177_), .Y(_abc_41234_new_n3219_));
NOR2X1 NOR2X1_446 ( .A(regfil_4__3_), .B(_abc_41234_new_n668__bF_buf2), .Y(_abc_41234_new_n3226_));
NOR2X1 NOR2X1_447 ( .A(_abc_41234_new_n534__bF_buf0), .B(_abc_41234_new_n2920_), .Y(_abc_41234_new_n3231_));
NOR2X1 NOR2X1_448 ( .A(_abc_41234_new_n1047__bF_buf0), .B(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3239_));
NOR2X1 NOR2X1_449 ( .A(_abc_41234_new_n3248_), .B(_abc_41234_new_n2919__bF_buf0), .Y(_abc_41234_new_n3254_));
NOR2X1 NOR2X1_45 ( .A(_abc_41234_new_n546__bF_buf1), .B(_abc_41234_new_n620__bF_buf4), .Y(_abc_41234_new_n665_));
NOR2X1 NOR2X1_450 ( .A(_abc_41234_new_n3101_), .B(_abc_41234_new_n3125_), .Y(_abc_41234_new_n3263_));
NOR2X1 NOR2X1_451 ( .A(_abc_41234_new_n3151_), .B(_abc_41234_new_n3175_), .Y(_abc_41234_new_n3265_));
NOR2X1 NOR2X1_452 ( .A(_abc_41234_new_n3266_), .B(_abc_41234_new_n3264_), .Y(_abc_41234_new_n3267_));
NOR2X1 NOR2X1_453 ( .A(_abc_41234_new_n2918_), .B(_abc_41234_new_n3273_), .Y(_abc_41234_new_n3274_));
NOR2X1 NOR2X1_454 ( .A(regfil_4__5_), .B(_abc_41234_new_n668__bF_buf0), .Y(_abc_41234_new_n3275_));
NOR2X1 NOR2X1_455 ( .A(regfil_4__6_), .B(_abc_41234_new_n668__bF_buf5), .Y(_abc_41234_new_n3295_));
NOR2X1 NOR2X1_456 ( .A(_abc_41234_new_n3297_), .B(_abc_41234_new_n2920_), .Y(_abc_41234_new_n3298_));
NOR2X1 NOR2X1_457 ( .A(_abc_41234_new_n2944_), .B(_abc_41234_new_n1804_), .Y(_abc_41234_new_n3302_));
NOR2X1 NOR2X1_458 ( .A(raddrhold_14_), .B(_abc_41234_new_n3309_), .Y(_abc_41234_new_n3310_));
NOR2X1 NOR2X1_459 ( .A(regfil_4__7_), .B(_abc_41234_new_n668__bF_buf4), .Y(_abc_41234_new_n3318_));
NOR2X1 NOR2X1_46 ( .A(_abc_41234_new_n665__bF_buf3), .B(_abc_41234_new_n669__bF_buf3), .Y(_abc_41234_new_n670_));
NOR2X1 NOR2X1_460 ( .A(_abc_41234_new_n2207__bF_buf3), .B(_abc_41234_new_n3318_), .Y(_abc_41234_new_n3319_));
NOR2X1 NOR2X1_461 ( .A(_abc_41234_new_n3294_), .B(_abc_41234_new_n3309_), .Y(_abc_41234_new_n3332_));
NOR2X1 NOR2X1_462 ( .A(_abc_41234_new_n3358_), .B(_abc_41234_new_n1643__bF_buf0), .Y(_abc_41234_new_n3362_));
NOR2X1 NOR2X1_463 ( .A(_abc_41234_new_n534__bF_buf5), .B(_abc_41234_new_n2964_), .Y(_abc_41234_new_n3365_));
NOR2X1 NOR2X1_464 ( .A(_abc_41234_new_n3337_), .B(_abc_41234_new_n3358_), .Y(_abc_41234_new_n3373_));
NOR2X1 NOR2X1_465 ( .A(sp_2_), .B(sp_1_), .Y(_abc_41234_new_n3382_));
NOR2X1 NOR2X1_466 ( .A(_abc_41234_new_n1071_), .B(_abc_41234_new_n2973_), .Y(_abc_41234_new_n3383_));
NOR2X1 NOR2X1_467 ( .A(_abc_41234_new_n3382_), .B(_abc_41234_new_n3383_), .Y(_abc_41234_new_n3384_));
NOR2X1 NOR2X1_468 ( .A(_abc_41234_new_n3403_), .B(_abc_41234_new_n3397_), .Y(_abc_41234_new_n3415_));
NOR2X1 NOR2X1_469 ( .A(sp_4_), .B(_abc_41234_new_n3423_), .Y(_abc_41234_new_n3424_));
NOR2X1 NOR2X1_47 ( .A(_abc_41234_new_n675_), .B(_abc_41234_new_n648_), .Y(_abc_41234_new_n676_));
NOR2X1 NOR2X1_470 ( .A(sp_5_), .B(_abc_41234_new_n3425_), .Y(_abc_41234_new_n3447_));
NOR2X1 NOR2X1_471 ( .A(_abc_41234_new_n3445_), .B(_abc_41234_new_n3439_), .Y(_abc_41234_new_n3461_));
NOR2X1 NOR2X1_472 ( .A(_abc_41234_new_n3487_), .B(_abc_41234_new_n3481_), .Y(_abc_41234_new_n3502_));
NOR2X1 NOR2X1_473 ( .A(sp_8_), .B(sp_9_), .Y(_abc_41234_new_n3528_));
NOR2X1 NOR2X1_474 ( .A(_abc_41234_new_n3526_), .B(_abc_41234_new_n3520_), .Y(_abc_41234_new_n3542_));
NOR2X1 NOR2X1_475 ( .A(_abc_41234_new_n3572_), .B(_abc_41234_new_n3489_), .Y(_abc_41234_new_n3592_));
NOR2X1 NOR2X1_476 ( .A(_abc_41234_new_n534__bF_buf2), .B(_abc_41234_new_n1761_), .Y(_abc_41234_new_n3600_));
NOR2X1 NOR2X1_477 ( .A(reset_bF_buf8), .B(_abc_41234_new_n2671_), .Y(_abc_41234_new_n3609_));
NOR2X1 NOR2X1_478 ( .A(sp_12_), .B(sp_13_), .Y(_abc_41234_new_n3617_));
NOR2X1 NOR2X1_479 ( .A(_abc_41234_new_n3605_), .B(_abc_41234_new_n3585_), .Y(_abc_41234_new_n3632_));
NOR2X1 NOR2X1_48 ( .A(_abc_41234_new_n656_), .B(_abc_41234_new_n677_), .Y(_abc_41234_new_n678_));
NOR2X1 NOR2X1_480 ( .A(sp_14_), .B(_abc_41234_new_n3618_), .Y(_abc_41234_new_n3638_));
NOR2X1 NOR2X1_481 ( .A(waddrhold_14_), .B(_abc_41234_new_n3633_), .Y(_abc_41234_new_n3652_));
NOR2X1 NOR2X1_482 ( .A(_abc_41234_new_n1850_), .B(_abc_41234_new_n609_), .Y(_abc_41234_new_n3677_));
NOR2X1 NOR2X1_483 ( .A(_abc_41234_new_n663_), .B(_abc_41234_new_n2186_), .Y(_abc_41234_new_n3704_));
NOR2X1 NOR2X1_484 ( .A(_abc_41234_new_n646_), .B(_abc_41234_new_n3714_), .Y(_abc_41234_new_n3715_));
NOR2X1 NOR2X1_485 ( .A(regfil_1__0_), .B(regfil_5__0_), .Y(_abc_41234_new_n3723_));
NOR2X1 NOR2X1_486 ( .A(_abc_41234_new_n3723_), .B(_abc_41234_new_n3722_), .Y(_abc_41234_new_n3724_));
NOR2X1 NOR2X1_487 ( .A(_abc_41234_new_n1207_), .B(_abc_41234_new_n1222_), .Y(_abc_41234_new_n3732_));
NOR2X1 NOR2X1_488 ( .A(_abc_41234_new_n1159_), .B(_abc_41234_new_n3738_), .Y(_abc_41234_new_n3739_));
NOR2X1 NOR2X1_489 ( .A(_abc_41234_new_n3742_), .B(_abc_41234_new_n3741_), .Y(_abc_41234_new_n3743_));
NOR2X1 NOR2X1_49 ( .A(_abc_41234_new_n607_), .B(_abc_41234_new_n592_), .Y(_abc_41234_new_n682_));
NOR2X1 NOR2X1_490 ( .A(_abc_41234_new_n3746_), .B(_abc_41234_new_n1308_), .Y(_abc_41234_new_n3747_));
NOR2X1 NOR2X1_491 ( .A(_abc_41234_new_n3747_), .B(_abc_41234_new_n3743_), .Y(_abc_41234_new_n3748_));
NOR2X1 NOR2X1_492 ( .A(_abc_41234_new_n3737_), .B(_abc_41234_new_n3749_), .Y(_abc_41234_new_n3750_));
NOR2X1 NOR2X1_493 ( .A(_abc_41234_new_n3751_), .B(_abc_41234_new_n3750_), .Y(_abc_41234_new_n3752_));
NOR2X1 NOR2X1_494 ( .A(regfil_5__2_), .B(_abc_41234_new_n3716_), .Y(_abc_41234_new_n3756_));
NOR2X1 NOR2X1_495 ( .A(regfil_5__2_), .B(_abc_41234_new_n1222_), .Y(_abc_41234_new_n3761_));
NOR2X1 NOR2X1_496 ( .A(_abc_41234_new_n3768_), .B(_abc_41234_new_n1324_), .Y(_abc_41234_new_n3769_));
NOR2X1 NOR2X1_497 ( .A(_abc_41234_new_n1070_), .B(_abc_41234_new_n1068_), .Y(_abc_41234_new_n3784_));
NOR2X1 NOR2X1_498 ( .A(regfil_5__3_bF_buf1_), .B(_abc_41234_new_n1224_), .Y(_abc_41234_new_n3796_));
NOR2X1 NOR2X1_499 ( .A(_abc_41234_new_n848_), .B(_abc_41234_new_n1209_), .Y(_abc_41234_new_n3805_));
NOR2X1 NOR2X1_5 ( .A(state_5_), .B(state_4_), .Y(_abc_41234_new_n517_));
NOR2X1 NOR2X1_50 ( .A(auxcar), .B(_abc_41234_new_n543_), .Y(_abc_41234_new_n684_));
NOR2X1 NOR2X1_500 ( .A(_abc_41234_new_n3811_), .B(_abc_41234_new_n3810_), .Y(_abc_41234_new_n3813_));
NOR2X1 NOR2X1_501 ( .A(_abc_41234_new_n1183_), .B(_abc_41234_new_n3837_), .Y(_abc_41234_new_n3838_));
NOR2X1 NOR2X1_502 ( .A(_abc_41234_new_n3834_), .B(_abc_41234_new_n3843_), .Y(_abc_41234_new_n3844_));
NOR2X1 NOR2X1_503 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n1229_), .Y(_abc_41234_new_n3845_));
NOR2X1 NOR2X1_504 ( .A(_abc_41234_new_n3848_), .B(_abc_41234_new_n3844_), .Y(_abc_41234_new_n3849_));
NOR2X1 NOR2X1_505 ( .A(_abc_41234_new_n1134_), .B(_abc_41234_new_n3810_), .Y(_abc_41234_new_n3858_));
NOR2X1 NOR2X1_506 ( .A(_abc_41234_new_n3857_), .B(_abc_41234_new_n3858_), .Y(_abc_41234_new_n3860_));
NOR2X1 NOR2X1_507 ( .A(_abc_41234_new_n1308_), .B(_abc_41234_new_n3862_), .Y(_abc_41234_new_n3863_));
NOR2X1 NOR2X1_508 ( .A(_abc_41234_new_n1188_), .B(_abc_41234_new_n3865_), .Y(_abc_41234_new_n3866_));
NOR2X1 NOR2X1_509 ( .A(regfil_5__7_), .B(_abc_41234_new_n1230_), .Y(_abc_41234_new_n3888_));
NOR2X1 NOR2X1_51 ( .A(state_4_), .B(_abc_41234_new_n691_), .Y(_abc_41234_new_n692_));
NOR2X1 NOR2X1_510 ( .A(_abc_41234_new_n3864_), .B(_abc_41234_new_n3866_), .Y(_abc_41234_new_n3891_));
NOR2X1 NOR2X1_511 ( .A(_abc_41234_new_n1174_), .B(_abc_41234_new_n3891_), .Y(_abc_41234_new_n3892_));
NOR2X1 NOR2X1_512 ( .A(_abc_41234_new_n610_), .B(_abc_41234_new_n590_), .Y(_abc_41234_new_n3911_));
NOR2X1 NOR2X1_513 ( .A(_abc_41234_new_n3915_), .B(_abc_41234_new_n3919_), .Y(_abc_41234_new_n3920_));
NOR2X1 NOR2X1_514 ( .A(sp_1_), .B(sp_0_bF_buf0_), .Y(_abc_41234_new_n3931_));
NOR2X1 NOR2X1_515 ( .A(_abc_41234_new_n2973_), .B(_abc_41234_new_n2947__bF_buf3), .Y(_abc_41234_new_n3932_));
NOR2X1 NOR2X1_516 ( .A(_abc_41234_new_n3931_), .B(_abc_41234_new_n3932_), .Y(_abc_41234_new_n3934_));
NOR2X1 NOR2X1_517 ( .A(_abc_41234_new_n693_), .B(_abc_41234_new_n3959_), .Y(_abc_41234_new_n3960_));
NOR2X1 NOR2X1_518 ( .A(_abc_41234_new_n2947__bF_buf2), .B(_abc_41234_new_n3969_), .Y(_abc_41234_new_n3979_));
NOR2X1 NOR2X1_519 ( .A(_abc_41234_new_n3935_), .B(_abc_41234_new_n3979_), .Y(_abc_41234_new_n3980_));
NOR2X1 NOR2X1_52 ( .A(state_3_), .B(state_2_), .Y(_abc_41234_new_n695_));
NOR2X1 NOR2X1_520 ( .A(_abc_41234_new_n3990_), .B(_abc_41234_new_n3961_), .Y(_abc_41234_new_n4004_));
NOR2X1 NOR2X1_521 ( .A(_abc_41234_new_n2462_), .B(_abc_41234_new_n1106_), .Y(_abc_41234_new_n4010_));
NOR2X1 NOR2X1_522 ( .A(_abc_41234_new_n1094_), .B(_abc_41234_new_n3995_), .Y(_abc_41234_new_n4021_));
NOR2X1 NOR2X1_523 ( .A(sp_0_bF_buf3_), .B(_abc_41234_new_n3467_), .Y(_abc_41234_new_n4036_));
NOR2X1 NOR2X1_524 ( .A(sp_6_), .B(_abc_41234_new_n4013_), .Y(_abc_41234_new_n4046_));
NOR2X1 NOR2X1_525 ( .A(_abc_41234_new_n4046_), .B(_abc_41234_new_n4040_), .Y(_abc_41234_new_n4047_));
NOR2X1 NOR2X1_526 ( .A(_abc_41234_new_n1047__bF_buf2), .B(_abc_41234_new_n2415__bF_buf3), .Y(_abc_41234_new_n4054_));
NOR2X1 NOR2X1_527 ( .A(sp_0_bF_buf1_), .B(_abc_41234_new_n3489_), .Y(_abc_41234_new_n4069_));
NOR2X1 NOR2X1_528 ( .A(_abc_41234_new_n1255_), .B(_abc_41234_new_n4059_), .Y(_abc_41234_new_n4079_));
NOR2X1 NOR2X1_529 ( .A(_abc_41234_new_n2947__bF_buf0), .B(_abc_41234_new_n4102_), .Y(_abc_41234_new_n4103_));
NOR2X1 NOR2X1_53 ( .A(_abc_41234_new_n694_), .B(_abc_41234_new_n696_), .Y(_abc_41234_new_n697_));
NOR2X1 NOR2X1_530 ( .A(_abc_41234_new_n1106_), .B(_abc_41234_new_n2482_), .Y(_abc_41234_new_n4112_));
NOR2X1 NOR2X1_531 ( .A(sp_0_bF_buf0_), .B(_abc_41234_new_n3549_), .Y(_abc_41234_new_n4123_));
NOR2X1 NOR2X1_532 ( .A(_abc_41234_new_n1362_), .B(_abc_41234_new_n4126_), .Y(_abc_41234_new_n4159_));
NOR2X1 NOR2X1_533 ( .A(_abc_41234_new_n3961_), .B(_abc_41234_new_n4148_), .Y(_abc_41234_new_n4163_));
NOR2X1 NOR2X1_534 ( .A(_abc_41234_new_n4163_), .B(_abc_41234_new_n4165_), .Y(_abc_41234_new_n4166_));
NOR2X1 NOR2X1_535 ( .A(sp_12_), .B(_abc_41234_new_n4169_), .Y(_abc_41234_new_n4170_));
NOR2X1 NOR2X1_536 ( .A(_abc_41234_new_n1408_), .B(_abc_41234_new_n4146_), .Y(_abc_41234_new_n4174_));
NOR2X1 NOR2X1_537 ( .A(_abc_41234_new_n2947__bF_buf0), .B(_abc_41234_new_n4175_), .Y(_abc_41234_new_n4176_));
NOR2X1 NOR2X1_538 ( .A(_abc_41234_new_n2947__bF_buf3), .B(_abc_41234_new_n4189_), .Y(_abc_41234_new_n4190_));
NOR2X1 NOR2X1_539 ( .A(_abc_41234_new_n4204_), .B(_abc_41234_new_n4203_), .Y(_abc_41234_new_n4205_));
NOR2X1 NOR2X1_54 ( .A(_abc_41234_new_n693_), .B(_abc_41234_new_n698_), .Y(_abc_41234_new_n699_));
NOR2X1 NOR2X1_540 ( .A(_abc_41234_new_n2947__bF_buf2), .B(_abc_41234_new_n4210_), .Y(_abc_41234_new_n4211_));
NOR2X1 NOR2X1_541 ( .A(_abc_41234_new_n1966_), .B(_abc_41234_new_n1059_), .Y(_abc_41234_new_n4257_));
NOR2X1 NOR2X1_542 ( .A(_abc_41234_new_n660__bF_buf2), .B(_abc_41234_new_n4274__bF_buf3), .Y(_abc_41234_new_n4275_));
NOR2X1 NOR2X1_543 ( .A(_abc_41234_new_n4284_), .B(_abc_41234_new_n4282_), .Y(_abc_41234_new_n4285_));
NOR2X1 NOR2X1_544 ( .A(_abc_41234_new_n549_), .B(_abc_41234_new_n4292_), .Y(_abc_41234_new_n4293_));
NOR2X1 NOR2X1_545 ( .A(_abc_41234_new_n2456_), .B(_abc_41234_new_n2931_), .Y(_abc_41234_new_n4297_));
NOR2X1 NOR2X1_546 ( .A(_abc_41234_new_n2936_), .B(_abc_41234_new_n2932_), .Y(_abc_41234_new_n4302_));
NOR2X1 NOR2X1_547 ( .A(_abc_41234_new_n4277_), .B(_abc_41234_new_n4303_), .Y(_abc_41234_new_n4304_));
NOR2X1 NOR2X1_548 ( .A(_abc_41234_new_n4305_), .B(_abc_41234_new_n4306_), .Y(_abc_41234_new_n4307_));
NOR2X1 NOR2X1_549 ( .A(_abc_41234_new_n1303_), .B(_abc_41234_new_n4309_), .Y(_abc_41234_new_n4310_));
NOR2X1 NOR2X1_55 ( .A(_abc_41234_new_n559_), .B(_abc_41234_new_n703_), .Y(_abc_41234_new_n704_));
NOR2X1 NOR2X1_550 ( .A(_abc_41234_new_n4308_), .B(_abc_41234_new_n4311_), .Y(_abc_41234_new_n4312_));
NOR2X1 NOR2X1_551 ( .A(_abc_41234_new_n1646_), .B(_abc_41234_new_n4326_), .Y(_abc_41234_new_n4327_));
NOR2X1 NOR2X1_552 ( .A(_abc_41234_new_n2737_), .B(_abc_41234_new_n2732_), .Y(_abc_41234_new_n4338_));
NOR2X1 NOR2X1_553 ( .A(_abc_41234_new_n4342_), .B(_abc_41234_new_n4341_), .Y(_abc_41234_new_n4343_));
NOR2X1 NOR2X1_554 ( .A(_abc_41234_new_n1614_), .B(_abc_41234_new_n4326_), .Y(_abc_41234_new_n4344_));
NOR2X1 NOR2X1_555 ( .A(_abc_41234_new_n534__bF_buf5), .B(_abc_41234_new_n4359_), .Y(_abc_41234_new_n4360_));
NOR2X1 NOR2X1_556 ( .A(_abc_41234_new_n2774_), .B(_abc_41234_new_n4328_), .Y(_abc_41234_new_n4361_));
NOR2X1 NOR2X1_557 ( .A(_abc_41234_new_n3914__bF_buf0), .B(_abc_41234_new_n2802_), .Y(_abc_41234_new_n4376_));
NOR2X1 NOR2X1_558 ( .A(_abc_41234_new_n4297__bF_buf3), .B(_abc_41234_new_n4392_), .Y(_abc_41234_new_n4393_));
NOR2X1 NOR2X1_559 ( .A(_abc_41234_new_n2831_), .B(_abc_41234_new_n4326_), .Y(_abc_41234_new_n4396_));
NOR2X1 NOR2X1_56 ( .A(_abc_41234_new_n504_), .B(_abc_41234_new_n694_), .Y(_abc_41234_new_n705_));
NOR2X1 NOR2X1_560 ( .A(_abc_41234_new_n2564_), .B(_abc_41234_new_n4391_), .Y(_abc_41234_new_n4397_));
NOR2X1 NOR2X1_561 ( .A(_abc_41234_new_n1617_), .B(_abc_41234_new_n4353_), .Y(_abc_41234_new_n4407_));
NOR2X1 NOR2X1_562 ( .A(_abc_41234_new_n4414_), .B(_abc_41234_new_n4413_), .Y(_abc_41234_new_n4415_));
NOR2X1 NOR2X1_563 ( .A(_abc_41234_new_n3914__bF_buf1), .B(_abc_41234_new_n2889_), .Y(_abc_41234_new_n4426_));
NOR2X1 NOR2X1_564 ( .A(_abc_41234_new_n4427_), .B(_abc_41234_new_n4428_), .Y(_abc_41234_new_n4429_));
NOR2X1 NOR2X1_565 ( .A(_abc_41234_new_n4454_), .B(_abc_41234_new_n4455_), .Y(_abc_41234_new_n4456_));
NOR2X1 NOR2X1_566 ( .A(_abc_41234_new_n4329_), .B(_abc_41234_new_n1673_), .Y(_abc_41234_new_n4464_));
NOR2X1 NOR2X1_567 ( .A(_abc_41234_new_n1705_), .B(_abc_41234_new_n4465_), .Y(_abc_41234_new_n4480_));
NOR2X1 NOR2X1_568 ( .A(_abc_41234_new_n1705_), .B(_abc_41234_new_n4326_), .Y(_abc_41234_new_n4489_));
NOR2X1 NOR2X1_569 ( .A(_abc_41234_new_n1727_), .B(_abc_41234_new_n4322_), .Y(_abc_41234_new_n4505_));
NOR2X1 NOR2X1_57 ( .A(reset_bF_buf4), .B(_abc_41234_new_n706_), .Y(_abc_41234_new_n707_));
NOR2X1 NOR2X1_570 ( .A(_abc_41234_new_n4297__bF_buf1), .B(_abc_41234_new_n4521_), .Y(_abc_41234_new_n4522_));
NOR2X1 NOR2X1_571 ( .A(_abc_41234_new_n4523_), .B(_abc_41234_new_n4522_), .Y(_abc_41234_new_n4524_));
NOR2X1 NOR2X1_572 ( .A(_abc_41234_new_n2564_), .B(_abc_41234_new_n4519_), .Y(_abc_41234_new_n4526_));
NOR2X1 NOR2X1_573 ( .A(_abc_41234_new_n2185__bF_buf1), .B(_abc_41234_new_n4558_), .Y(_abc_41234_new_n4559_));
NOR2X1 NOR2X1_574 ( .A(_abc_41234_new_n1828_), .B(_abc_41234_new_n4322_), .Y(_abc_41234_new_n4586_));
NOR2X1 NOR2X1_575 ( .A(_abc_41234_new_n607_), .B(_abc_41234_new_n2512_), .Y(_abc_41234_new_n4600_));
NOR2X1 NOR2X1_576 ( .A(_abc_41234_new_n518_), .B(_abc_41234_new_n2212_), .Y(_abc_41234_new_n4660_));
NOR2X1 NOR2X1_577 ( .A(_abc_41234_new_n4604_), .B(_abc_41234_new_n4606_), .Y(_abc_41234_new_n4695_));
NOR2X1 NOR2X1_578 ( .A(_abc_41234_new_n1729_), .B(_abc_41234_new_n2959__bF_buf0), .Y(_abc_41234_new_n4697_));
NOR2X1 NOR2X1_579 ( .A(waitr), .B(_abc_41234_new_n4704_), .Y(_abc_41234_new_n4705_));
NOR2X1 NOR2X1_58 ( .A(_abc_41234_new_n707_), .B(_abc_41234_new_n513_), .Y(_abc_41234_new_n708_));
NOR2X1 NOR2X1_580 ( .A(statesel_2_), .B(_abc_41234_new_n2588_), .Y(_abc_41234_new_n4709_));
NOR2X1 NOR2X1_581 ( .A(statesel_2_), .B(statesel_3_), .Y(_abc_41234_new_n4713_));
NOR2X1 NOR2X1_582 ( .A(_abc_41234_new_n4712_), .B(_abc_41234_new_n2602_), .Y(_abc_41234_new_n4715_));
NOR2X1 NOR2X1_583 ( .A(statesel_4_), .B(_abc_41234_new_n4719_), .Y(_abc_41234_new_n4720_));
NOR2X1 NOR2X1_584 ( .A(_abc_41234_new_n2601_), .B(_abc_41234_new_n4721_), .Y(_abc_41234_new_n4722_));
NOR2X1 NOR2X1_585 ( .A(_abc_41234_new_n2611_), .B(_abc_41234_new_n4719_), .Y(_abc_41234_new_n4725_));
NOR2X1 NOR2X1_586 ( .A(statesel_0_), .B(statesel_1_), .Y(_abc_41234_new_n4727_));
NOR2X1 NOR2X1_587 ( .A(statesel_4_), .B(statesel_5_), .Y(_abc_41234_new_n4729_));
NOR2X1 NOR2X1_588 ( .A(statesel_0_), .B(_abc_41234_new_n4730_), .Y(_abc_41234_new_n4731_));
NOR2X1 NOR2X1_589 ( .A(_abc_41234_new_n4733_), .B(_abc_41234_new_n2641_), .Y(_abc_41234_new_n4734_));
NOR2X1 NOR2X1_59 ( .A(_abc_41234_new_n687_), .B(_abc_41234_new_n709_), .Y(_abc_41234_new_n710_));
NOR2X1 NOR2X1_590 ( .A(reset_bF_buf9), .B(_abc_41234_new_n534__bF_buf1), .Y(_abc_41234_new_n4736_));
NOR2X1 NOR2X1_591 ( .A(_abc_41234_new_n1630_), .B(_abc_41234_new_n2710_), .Y(_abc_41234_new_n4738_));
NOR2X1 NOR2X1_592 ( .A(opcode_5_bF_buf0_), .B(carry), .Y(_abc_41234_new_n4741_));
NOR2X1 NOR2X1_593 ( .A(_abc_41234_new_n2501_), .B(_abc_41234_new_n2415__bF_buf2), .Y(_abc_41234_new_n4758_));
NOR2X1 NOR2X1_594 ( .A(_abc_41234_new_n4726_), .B(_abc_41234_new_n2534_), .Y(_abc_41234_new_n4760_));
NOR2X1 NOR2X1_595 ( .A(_abc_41234_new_n4710_), .B(_abc_41234_new_n2582_), .Y(_abc_41234_new_n4761_));
NOR2X1 NOR2X1_596 ( .A(_abc_41234_new_n4712_), .B(_abc_41234_new_n4710_), .Y(_abc_41234_new_n4766_));
NOR2X1 NOR2X1_597 ( .A(_abc_41234_new_n4767_), .B(_abc_41234_new_n2621_), .Y(_abc_41234_new_n4768_));
NOR2X1 NOR2X1_598 ( .A(_abc_41234_new_n4769_), .B(_abc_41234_new_n2534_), .Y(_abc_41234_new_n4770_));
NOR2X1 NOR2X1_599 ( .A(_abc_41234_new_n3677_), .B(_abc_41234_new_n4770_), .Y(_abc_41234_new_n4771_));
NOR2X1 NOR2X1_6 ( .A(_abc_41234_new_n504_), .B(_abc_41234_new_n521_), .Y(_abc_41234_new_n522_));
NOR2X1 NOR2X1_60 ( .A(_abc_41234_new_n726_), .B(_abc_41234_new_n724_), .Y(_abc_41234_new_n727_));
NOR2X1 NOR2X1_600 ( .A(_abc_41234_new_n4660_), .B(_abc_41234_new_n551_), .Y(_abc_41234_new_n4772_));
NOR2X1 NOR2X1_601 ( .A(_abc_41234_new_n4765_), .B(_abc_41234_new_n4773_), .Y(_abc_41234_new_n4774_));
NOR2X1 NOR2X1_602 ( .A(_abc_41234_new_n4778_), .B(_abc_41234_new_n2534_), .Y(_abc_41234_new_n4779_));
NOR2X1 NOR2X1_603 ( .A(_abc_41234_new_n4714_), .B(_abc_41234_new_n2582_), .Y(_abc_41234_new_n4780_));
NOR2X1 NOR2X1_604 ( .A(reset_bF_buf7), .B(_abc_41234_new_n681_), .Y(_abc_41234_new_n4782_));
NOR2X1 NOR2X1_605 ( .A(_abc_41234_new_n4784_), .B(_abc_41234_new_n4785_), .Y(_abc_41234_new_n4786_));
NOR2X1 NOR2X1_606 ( .A(_abc_41234_new_n4712_), .B(_abc_41234_new_n2621_), .Y(_abc_41234_new_n4789_));
NOR2X1 NOR2X1_607 ( .A(statesel_4_), .B(_abc_41234_new_n4789_), .Y(_abc_41234_new_n4790_));
NOR2X1 NOR2X1_608 ( .A(statesel_1_), .B(_abc_41234_new_n2621_), .Y(_abc_41234_new_n4791_));
NOR2X1 NOR2X1_609 ( .A(_abc_41234_new_n4767_), .B(_abc_41234_new_n2602_), .Y(_abc_41234_new_n4800_));
NOR2X1 NOR2X1_61 ( .A(regfil_0__1_), .B(_abc_41234_new_n586_), .Y(_abc_41234_new_n738_));
NOR2X1 NOR2X1_610 ( .A(reset_bF_buf6), .B(_abc_41234_new_n4730_), .Y(_abc_41234_new_n4801_));
NOR2X1 NOR2X1_611 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n4704_), .Y(_abc_41234_new_n4814_));
NOR2X1 NOR2X1_612 ( .A(_abc_41234_new_n4808_), .B(_abc_41234_new_n4816_), .Y(_abc_41234_new_n4817_));
NOR2X1 NOR2X1_613 ( .A(_abc_41234_new_n4775_), .B(_abc_41234_new_n4818_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_0_));
NOR2X1 NOR2X1_614 ( .A(reset_bF_buf5), .B(_abc_41234_new_n4612_), .Y(_abc_41234_new_n4820_));
NOR2X1 NOR2X1_615 ( .A(_abc_41234_new_n4750_), .B(_abc_41234_new_n2415__bF_buf1), .Y(_abc_41234_new_n4823_));
NOR2X1 NOR2X1_616 ( .A(_abc_41234_new_n4820_), .B(_abc_41234_new_n4825_), .Y(_abc_41234_new_n4826_));
NOR2X1 NOR2X1_617 ( .A(_abc_41234_new_n4714_), .B(_abc_41234_new_n4708_), .Y(_abc_41234_new_n4827_));
NOR2X1 NOR2X1_618 ( .A(_abc_41234_new_n4828_), .B(_abc_41234_new_n2534_), .Y(_abc_41234_new_n4829_));
NOR2X1 NOR2X1_619 ( .A(_abc_41234_new_n3609_), .B(_abc_41234_new_n4829_), .Y(_abc_41234_new_n4830_));
NOR2X1 NOR2X1_62 ( .A(_abc_41234_new_n739_), .B(_abc_41234_new_n740_), .Y(_abc_41234_new_n741_));
NOR2X1 NOR2X1_620 ( .A(_abc_41234_new_n4833_), .B(_abc_41234_new_n4836_), .Y(_abc_41234_new_n4837_));
NOR2X1 NOR2X1_621 ( .A(_abc_41234_new_n4805_), .B(_abc_41234_new_n4775_), .Y(_abc_41234_new_n4838_));
NOR2X1 NOR2X1_622 ( .A(_abc_41234_new_n4814_), .B(_abc_41234_new_n4820_), .Y(_abc_41234_new_n4842_));
NOR2X1 NOR2X1_623 ( .A(_abc_41234_new_n4843_), .B(_abc_41234_new_n4840_), .Y(_abc_41234_new_n4844_));
NOR2X1 NOR2X1_624 ( .A(_abc_41234_new_n4767_), .B(_abc_41234_new_n4710_), .Y(_abc_41234_new_n4846_));
NOR2X1 NOR2X1_625 ( .A(_abc_41234_new_n4854_), .B(_abc_41234_new_n4855_), .Y(_abc_41234_new_n4856_));
NOR2X1 NOR2X1_626 ( .A(_abc_41234_new_n4808_), .B(_abc_41234_new_n4858_), .Y(_abc_41234_new_n4859_));
NOR2X1 NOR2X1_627 ( .A(_abc_41234_new_n2604_), .B(_abc_41234_new_n2600_), .Y(_abc_41234_new_n4860_));
NOR2X1 NOR2X1_628 ( .A(_abc_41234_new_n4862_), .B(_abc_41234_new_n4863_), .Y(_abc_41234_new_n4864_));
NOR2X1 NOR2X1_629 ( .A(_abc_41234_new_n4866_), .B(_abc_41234_new_n4833_), .Y(_abc_41234_new_n4867_));
NOR2X1 NOR2X1_63 ( .A(regfil_0__1_), .B(_abc_41234_new_n642_), .Y(_abc_41234_new_n743_));
NOR2X1 NOR2X1_630 ( .A(_abc_41234_new_n4872_), .B(_abc_41234_new_n4874_), .Y(_abc_41234_new_n4875_));
NOR2X1 NOR2X1_631 ( .A(_abc_41234_new_n4871_), .B(_abc_41234_new_n4876_), .Y(_abc_41234_new_n4877_));
NOR2X1 NOR2X1_632 ( .A(_abc_41234_new_n4878_), .B(_abc_41234_new_n4879_), .Y(_abc_41234_new_n4880_));
NOR2X1 NOR2X1_633 ( .A(alu_oprb_7_), .B(alu_opra_7_), .Y(alu__abc_40887_new_n33_));
NOR2X1 NOR2X1_634 ( .A(alu__abc_40887_new_n33_), .B(alu__abc_40887_new_n35_), .Y(alu__abc_40887_new_n36_));
NOR2X1 NOR2X1_635 ( .A(alu_oprb_6_), .B(alu_opra_6_), .Y(alu__abc_40887_new_n39_));
NOR2X1 NOR2X1_636 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_40887_new_n44_));
NOR2X1 NOR2X1_637 ( .A(alu_oprb_2_), .B(alu_opra_2_), .Y(alu__abc_40887_new_n48_));
NOR2X1 NOR2X1_638 ( .A(alu__abc_40887_new_n48_), .B(alu__abc_40887_new_n47_), .Y(alu__abc_40887_new_n49_));
NOR2X1 NOR2X1_639 ( .A(alu_oprb_3_), .B(alu_opra_3_), .Y(alu__abc_40887_new_n51_));
NOR2X1 NOR2X1_64 ( .A(_abc_41234_new_n748_), .B(_abc_41234_new_n679_), .Y(_abc_41234_new_n749_));
NOR2X1 NOR2X1_640 ( .A(alu__abc_40887_new_n51_), .B(alu__abc_40887_new_n50_), .Y(alu__abc_40887_new_n52_));
NOR2X1 NOR2X1_641 ( .A(alu_oprb_5_), .B(alu_opra_5_), .Y(alu__abc_40887_new_n59_));
NOR2X1 NOR2X1_642 ( .A(alu__abc_40887_new_n59_), .B(alu__abc_40887_new_n61_), .Y(alu__abc_40887_new_n62_));
NOR2X1 NOR2X1_643 ( .A(alu__abc_40887_new_n76_), .B(alu__abc_40887_new_n62_), .Y(alu__abc_40887_new_n77_));
NOR2X1 NOR2X1_644 ( .A(alu__abc_40887_new_n90_), .B(alu__abc_40887_new_n92_), .Y(alu__abc_40887_new_n93_));
NOR2X1 NOR2X1_645 ( .A(alu_sel_2_), .B(alu__abc_40887_new_n103_), .Y(alu__abc_40887_new_n104_));
NOR2X1 NOR2X1_646 ( .A(alu__abc_40887_new_n102_), .B(alu__abc_40887_new_n116_), .Y(alu__abc_40887_new_n117_));
NOR2X1 NOR2X1_647 ( .A(alu_oprb_3_), .B(alu__abc_40887_new_n119_), .Y(alu__abc_40887_new_n120_));
NOR2X1 NOR2X1_648 ( .A(alu_oprb_4_), .B(alu__abc_40887_new_n137_), .Y(alu__abc_40887_new_n138_));
NOR2X1 NOR2X1_649 ( .A(alu_oprb_6_), .B(alu__abc_40887_new_n143_), .Y(alu__abc_40887_new_n144_));
NOR2X1 NOR2X1_65 ( .A(reset_bF_buf3), .B(waitr), .Y(_abc_41234_new_n756_));
NOR2X1 NOR2X1_650 ( .A(alu_oprb_1_), .B(alu__abc_40887_new_n125_), .Y(alu__abc_40887_new_n148_));
NOR2X1 NOR2X1_651 ( .A(alu__abc_40887_new_n44_), .B(alu__abc_40887_new_n127_), .Y(alu__abc_40887_new_n170_));
NOR2X1 NOR2X1_652 ( .A(alu__abc_40887_new_n138_), .B(alu__abc_40887_new_n178_), .Y(alu__abc_40887_new_n179_));
NOR2X1 NOR2X1_653 ( .A(alu__abc_40887_new_n129_), .B(alu__abc_40887_new_n90_), .Y(alu__abc_40887_new_n192_));
NOR2X1 NOR2X1_654 ( .A(alu__abc_40887_new_n189_), .B(alu__abc_40887_new_n195_), .Y(alu__abc_40887_new_n196_));
NOR2X1 NOR2X1_655 ( .A(alu_sel_1_), .B(alu_sel_0_), .Y(alu__abc_40887_new_n199_));
NOR2X1 NOR2X1_656 ( .A(alu_sel_2_), .B(alu__abc_40887_new_n200_), .Y(alu__abc_40887_new_n201_));
NOR2X1 NOR2X1_657 ( .A(alu_sel_0_), .B(alu__abc_40887_new_n102_), .Y(alu__abc_40887_new_n202_));
NOR2X1 NOR2X1_658 ( .A(alu__abc_40887_new_n110_), .B(alu__abc_40887_new_n111_), .Y(alu__abc_40887_new_n218_));
NOR2X1 NOR2X1_659 ( .A(alu__abc_40887_new_n168_), .B(alu__abc_40887_new_n236_), .Y(alu__abc_40887_new_n237_));
NOR2X1 NOR2X1_66 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n755_), .Y(_abc_41234_new_n758_));
NOR2X1 NOR2X1_660 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n93_), .Y(alu__abc_40887_new_n242_));
NOR2X1 NOR2X1_661 ( .A(alu__abc_40887_new_n201_), .B(alu__abc_40887_new_n227_), .Y(alu__abc_40887_new_n250_));
NOR2X1 NOR2X1_662 ( .A(alu__abc_40887_new_n251_), .B(alu__abc_40887_new_n256_), .Y(alu__abc_40887_new_n257_));
NOR2X1 NOR2X1_663 ( .A(alu__abc_40887_new_n194_), .B(alu__abc_40887_new_n191_), .Y(alu__abc_40887_new_n259_));
NOR2X1 NOR2X1_664 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n96_), .Y(alu__abc_40887_new_n262_));
NOR2X1 NOR2X1_665 ( .A(alu__abc_40887_new_n83_), .B(alu__abc_40887_new_n211_), .Y(alu__abc_40887_new_n264_));
NOR2X1 NOR2X1_666 ( .A(alu__abc_40887_new_n49_), .B(alu__abc_40887_new_n46_), .Y(alu__abc_40887_new_n274_));
NOR2X1 NOR2X1_667 ( .A(alu__abc_40887_new_n274_), .B(alu__abc_40887_new_n82_), .Y(alu__abc_40887_new_n279_));
NOR2X1 NOR2X1_668 ( .A(alu__abc_40887_new_n172_), .B(alu__abc_40887_new_n166_), .Y(alu__abc_40887_new_n294_));
NOR2X1 NOR2X1_669 ( .A(alu__abc_40887_new_n190_), .B(alu__abc_40887_new_n174_), .Y(alu__abc_40887_new_n323_));
NOR2X1 NOR2X1_67 ( .A(_abc_41234_new_n754_), .B(_abc_41234_new_n762_), .Y(_abc_41234_new_n763_));
NOR2X1 NOR2X1_670 ( .A(alu__abc_40887_new_n56_), .B(alu__abc_40887_new_n211_), .Y(alu__abc_40887_new_n327_));
NOR2X1 NOR2X1_671 ( .A(alu__abc_40887_new_n327_), .B(alu__abc_40887_new_n326_), .Y(alu__abc_40887_new_n328_));
NOR2X1 NOR2X1_672 ( .A(alu__abc_40887_new_n232_), .B(alu_sout), .Y(alu__abc_40887_new_n344_));
NOR2X1 NOR2X1_673 ( .A(alu__abc_40887_new_n351_), .B(alu__abc_40887_new_n335_), .Y(alu__abc_40887_new_n352_));
NOR2X1 NOR2X1_68 ( .A(regfil_0__2_), .B(_abc_41234_new_n741_), .Y(_abc_41234_new_n782_));
NOR2X1 NOR2X1_69 ( .A(_abc_41234_new_n766_), .B(_abc_41234_new_n783_), .Y(_abc_41234_new_n784_));
NOR2X1 NOR2X1_7 ( .A(_abc_41234_new_n526__bF_buf3), .B(_abc_41234_new_n527_), .Y(_abc_41234_new_n528_));
NOR2X1 NOR2X1_70 ( .A(_abc_41234_new_n679_), .B(_abc_41234_new_n791_), .Y(_abc_41234_new_n792_));
NOR2X1 NOR2X1_71 ( .A(_abc_41234_new_n684_), .B(_abc_41234_new_n685_), .Y(_abc_41234_new_n795_));
NOR2X1 NOR2X1_72 ( .A(_abc_41234_new_n802_), .B(_abc_41234_new_n800_), .Y(_abc_41234_new_n803_));
NOR2X1 NOR2X1_73 ( .A(_abc_41234_new_n826_), .B(_abc_41234_new_n648_), .Y(_abc_41234_new_n827_));
NOR2X1 NOR2X1_74 ( .A(_abc_41234_new_n679_), .B(_abc_41234_new_n829_), .Y(_abc_41234_new_n830_));
NOR2X1 NOR2X1_75 ( .A(regfil_7__2_), .B(regfil_7__1_), .Y(_abc_41234_new_n834_));
NOR2X1 NOR2X1_76 ( .A(_abc_41234_new_n853_), .B(_abc_41234_new_n850_), .Y(_abc_41234_new_n854_));
NOR2X1 NOR2X1_77 ( .A(_abc_41234_new_n867_), .B(_abc_41234_new_n868_), .Y(_abc_41234_new_n869_));
NOR2X1 NOR2X1_78 ( .A(_abc_41234_new_n879_), .B(_abc_41234_new_n679_), .Y(_abc_41234_new_n880_));
NOR2X1 NOR2X1_79 ( .A(_abc_41234_new_n851_), .B(_abc_41234_new_n542_), .Y(_abc_41234_new_n882_));
NOR2X1 NOR2X1_8 ( .A(opcode_5_bF_buf4_), .B(_abc_41234_new_n529_), .Y(_abc_41234_new_n530_));
NOR2X1 NOR2X1_80 ( .A(_abc_41234_new_n882_), .B(_abc_41234_new_n686_), .Y(_abc_41234_new_n883_));
NOR2X1 NOR2X1_81 ( .A(_abc_41234_new_n892_), .B(_abc_41234_new_n889_), .Y(_abc_41234_new_n893_));
NOR2X1 NOR2X1_82 ( .A(_abc_41234_new_n901_), .B(_abc_41234_new_n898_), .Y(_abc_41234_new_n902_));
NOR2X1 NOR2X1_83 ( .A(_abc_41234_new_n679_), .B(_abc_41234_new_n924_), .Y(_abc_41234_new_n925_));
NOR2X1 NOR2X1_84 ( .A(_abc_41234_new_n906_), .B(_abc_41234_new_n930_), .Y(_abc_41234_new_n931_));
NOR2X1 NOR2X1_85 ( .A(_abc_41234_new_n918_), .B(_abc_41234_new_n806_), .Y(_abc_41234_new_n958_));
NOR2X1 NOR2X1_86 ( .A(_abc_41234_new_n679_), .B(_abc_41234_new_n963_), .Y(_abc_41234_new_n964_));
NOR2X1 NOR2X1_87 ( .A(_abc_41234_new_n967_), .B(_abc_41234_new_n968_), .Y(_abc_41234_new_n969_));
NOR2X1 NOR2X1_88 ( .A(regfil_7__6_), .B(regfil_7__5_), .Y(_abc_41234_new_n976_));
NOR2X1 NOR2X1_89 ( .A(_abc_41234_new_n967_), .B(_abc_41234_new_n906_), .Y(_abc_41234_new_n977_));
NOR2X1 NOR2X1_9 ( .A(opcode_4_bF_buf5_), .B(opcode_5_bF_buf3_), .Y(_abc_41234_new_n531_));
NOR2X1 NOR2X1_90 ( .A(_abc_41234_new_n944_), .B(_abc_41234_new_n954_), .Y(_abc_41234_new_n985_));
NOR2X1 NOR2X1_91 ( .A(_abc_41234_new_n607_), .B(_abc_41234_new_n606_), .Y(_abc_41234_new_n1004_));
NOR2X1 NOR2X1_92 ( .A(reset_bF_buf2), .B(_abc_41234_new_n1005_), .Y(_abc_41234_new_n1006_));
NOR2X1 NOR2X1_93 ( .A(_abc_41234_new_n1010_), .B(_abc_41234_new_n679_), .Y(_abc_41234_new_n1011_));
NOR2X1 NOR2X1_94 ( .A(regfil_7__7_), .B(_abc_41234_new_n1022_), .Y(_abc_41234_new_n1023_));
NOR2X1 NOR2X1_95 ( .A(_abc_41234_new_n590_), .B(_abc_41234_new_n694_), .Y(_abc_41234_new_n1033_));
NOR2X1 NOR2X1_96 ( .A(_abc_41234_new_n544__bF_buf2), .B(_abc_41234_new_n1038_), .Y(_abc_41234_new_n1039_));
NOR2X1 NOR2X1_97 ( .A(_abc_41234_new_n661_), .B(_abc_41234_new_n1045_), .Y(_abc_41234_new_n1046_));
NOR2X1 NOR2X1_98 ( .A(_abc_41234_new_n1047__bF_buf4), .B(_abc_41234_new_n523__bF_buf1), .Y(_abc_41234_new_n1048_));
NOR2X1 NOR2X1_99 ( .A(opcode_2_), .B(_abc_41234_new_n555_), .Y(_abc_41234_new_n1050_));
NOR3X1 NOR3X1_1 ( .A(_abc_41234_new_n1084_), .B(_abc_41234_new_n903_), .C(_abc_41234_new_n1229_), .Y(_abc_41234_new_n1230_));
NOR3X1 NOR3X1_10 ( .A(_abc_41234_new_n1705_), .B(_abc_41234_new_n1727_), .C(_abc_41234_new_n4465_), .Y(_abc_41234_new_n4499_));
NOR3X1 NOR3X1_11 ( .A(_abc_41234_new_n4525_), .B(_abc_41234_new_n4526_), .C(_abc_41234_new_n4531_), .Y(_abc_41234_new_n4532_));
NOR3X1 NOR3X1_12 ( .A(_abc_41234_new_n4777_), .B(_abc_41234_new_n4788_), .C(_abc_41234_new_n4805_), .Y(_abc_41234_new_n4806_));
NOR3X1 NOR3X1_13 ( .A(alu__abc_40887_new_n110_), .B(alu__abc_40887_new_n111_), .C(alu__abc_40887_new_n74_), .Y(alu__abc_40887_new_n112_));
NOR3X1 NOR3X1_14 ( .A(alu__abc_40887_new_n277_), .B(alu__abc_40887_new_n283_), .C(alu__abc_40887_new_n273_), .Y(alu__abc_40887_new_n284_));
NOR3X1 NOR3X1_15 ( .A(alu__abc_40887_new_n289_), .B(alu__abc_40887_new_n298_), .C(alu__abc_40887_new_n293_), .Y(alu__abc_40887_new_n302_));
NOR3X1 NOR3X1_2 ( .A(_abc_41234_new_n720_), .B(_abc_41234_new_n773_), .C(_abc_41234_new_n1231_), .Y(_abc_41234_new_n1353_));
NOR3X1 NOR3X1_3 ( .A(_abc_41234_new_n819_), .B(_abc_41234_new_n849_), .C(_abc_41234_new_n1294_), .Y(_abc_41234_new_n1452_));
NOR3X1 NOR3X1_4 ( .A(_abc_41234_new_n1152_), .B(_abc_41234_new_n1539_), .C(_abc_41234_new_n1540_), .Y(_abc_41234_new_n1541_));
NOR3X1 NOR3X1_5 ( .A(_abc_41234_new_n731_), .B(_abc_41234_new_n769_), .C(_abc_41234_new_n2060_), .Y(_abc_41234_new_n2095_));
NOR3X1 NOR3X1_6 ( .A(_abc_41234_new_n1094_), .B(_abc_41234_new_n1090_), .C(_abc_41234_new_n3969_), .Y(_abc_41234_new_n4013_));
NOR3X1 NOR3X1_7 ( .A(_abc_41234_new_n1255_), .B(_abc_41234_new_n1251_), .C(_abc_41234_new_n4059_), .Y(_abc_41234_new_n4101_));
NOR3X1 NOR3X1_8 ( .A(_abc_41234_new_n4279_), .B(_abc_41234_new_n4278_), .C(_abc_41234_new_n4277_), .Y(_abc_41234_new_n4280_));
NOR3X1 NOR3X1_9 ( .A(_abc_41234_new_n1617_), .B(_abc_41234_new_n1618_), .C(_abc_41234_new_n4353_), .Y(_abc_41234_new_n4427_));
OAI21X1 OAI21X1_1 ( .A(_abc_41234_new_n531_), .B(_abc_41234_new_n530_), .C(_abc_41234_new_n528_), .Y(_abc_41234_new_n532_));
OAI21X1 OAI21X1_10 ( .A(_abc_41234_new_n546__bF_buf2), .B(_abc_41234_new_n626_), .C(_abc_41234_new_n623_), .Y(_abc_41234_new_n627_));
OAI21X1 OAI21X1_100 ( .A(_abc_41234_new_n1039_), .B(_abc_41234_new_n1041_), .C(_abc_41234_new_n535_), .Y(_abc_41234_new_n1042_));
OAI21X1 OAI21X1_1000 ( .A(_abc_41234_new_n2488_), .B(_abc_41234_new_n3385_), .C(_abc_41234_new_n1046__bF_buf0), .Y(_abc_41234_new_n3945_));
OAI21X1 OAI21X1_1001 ( .A(_abc_41234_new_n1071_), .B(_abc_41234_new_n3927_), .C(_abc_41234_new_n3947_), .Y(_abc_41234_new_n3948_));
OAI21X1 OAI21X1_1002 ( .A(_abc_41234_new_n1071_), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n3950_), .Y(_abc_41234_new_n3951_));
OAI21X1 OAI21X1_1003 ( .A(sp_2_), .B(_abc_41234_new_n3932_), .C(_abc_41234_new_n3951_), .Y(_abc_41234_new_n3952_));
OAI21X1 OAI21X1_1004 ( .A(sp_1_), .B(sp_0_bF_buf2_), .C(sp_2_), .Y(_abc_41234_new_n3954_));
OAI21X1 OAI21X1_1005 ( .A(sp_2_), .B(_abc_41234_new_n3914__bF_buf1), .C(_abc_41234_new_n660__bF_buf2), .Y(_abc_41234_new_n3957_));
OAI21X1 OAI21X1_1006 ( .A(_abc_41234_new_n3385_), .B(_abc_41234_new_n3961_), .C(_abc_41234_new_n3965_), .Y(_abc_41234_new_n3966_));
OAI21X1 OAI21X1_1007 ( .A(_abc_41234_new_n1071_), .B(_abc_41234_new_n2973_), .C(_abc_41234_new_n1067_), .Y(_abc_41234_new_n3970_));
OAI21X1 OAI21X1_1008 ( .A(_abc_41234_new_n1067_), .B(_abc_41234_new_n3927_), .C(_abc_41234_new_n3974_), .Y(_abc_41234_new_n3975_));
OAI21X1 OAI21X1_1009 ( .A(sp_3_), .B(_abc_41234_new_n3914__bF_buf0), .C(_abc_41234_new_n660__bF_buf1), .Y(_abc_41234_new_n3982_));
OAI21X1 OAI21X1_101 ( .A(_abc_41234_new_n675_), .B(_abc_41234_new_n648_), .C(_abc_41234_new_n672_), .Y(_abc_41234_new_n1059_));
OAI21X1 OAI21X1_1010 ( .A(_abc_41234_new_n2654_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n3985_), .Y(_abc_41234_new_n3986_));
OAI21X1 OAI21X1_1011 ( .A(_abc_41234_new_n1090_), .B(_abc_41234_new_n3927_), .C(_abc_41234_new_n3993_), .Y(_abc_41234_new_n3994_));
OAI21X1 OAI21X1_1012 ( .A(sp_4_), .B(_abc_41234_new_n3979_), .C(_abc_41234_new_n3997_), .Y(_abc_41234_new_n3998_));
OAI21X1 OAI21X1_1013 ( .A(sp_0_bF_buf1_), .B(_abc_41234_new_n3423_), .C(sp_4_), .Y(_abc_41234_new_n3999_));
OAI21X1 OAI21X1_1014 ( .A(sp_0_bF_buf0_), .B(_abc_41234_new_n3425_), .C(_abc_41234_new_n3999_), .Y(_abc_41234_new_n4000_));
OAI21X1 OAI21X1_1015 ( .A(sp_4_), .B(_abc_41234_new_n3914__bF_buf3), .C(_abc_41234_new_n660__bF_buf0), .Y(_abc_41234_new_n4002_));
OAI21X1 OAI21X1_1016 ( .A(_abc_41234_new_n2656_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n4005_), .Y(_abc_41234_new_n4006_));
OAI21X1 OAI21X1_1017 ( .A(_abc_41234_new_n1090_), .B(_abc_41234_new_n3969_), .C(_abc_41234_new_n1094_), .Y(_abc_41234_new_n4015_));
OAI21X1 OAI21X1_1018 ( .A(_abc_41234_new_n1639__bF_buf2), .B(_abc_41234_new_n1637_), .C(_abc_41234_new_n3449_), .Y(_abc_41234_new_n4018_));
OAI21X1 OAI21X1_1019 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n1107_), .C(_abc_41234_new_n4018_), .Y(_abc_41234_new_n4019_));
OAI21X1 OAI21X1_102 ( .A(_abc_41234_new_n1058_), .B(_abc_41234_new_n1059_), .C(regfil_4__0_), .Y(_abc_41234_new_n1062_));
OAI21X1 OAI21X1_1020 ( .A(_abc_41234_new_n4017_), .B(_abc_41234_new_n4019_), .C(_abc_41234_new_n1046__bF_buf5), .Y(_abc_41234_new_n4020_));
OAI21X1 OAI21X1_1021 ( .A(sp_5_), .B(_abc_41234_new_n3996_), .C(_abc_41234_new_n3936_), .Y(_abc_41234_new_n4022_));
OAI21X1 OAI21X1_1022 ( .A(_abc_41234_new_n1094_), .B(_abc_41234_new_n4023_), .C(_abc_41234_new_n4024_), .Y(_abc_41234_new_n4025_));
OAI21X1 OAI21X1_1023 ( .A(_abc_41234_new_n4021_), .B(_abc_41234_new_n4022_), .C(_abc_41234_new_n4025_), .Y(_abc_41234_new_n4026_));
OAI21X1 OAI21X1_1024 ( .A(_abc_41234_new_n2415__bF_buf4), .B(_abc_41234_new_n4029_), .C(_abc_41234_new_n4030_), .Y(_abc_41234_new_n4031_));
OAI21X1 OAI21X1_1025 ( .A(_abc_41234_new_n2658_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n4032_), .Y(_abc_41234_new_n4033_));
OAI21X1 OAI21X1_1026 ( .A(_abc_41234_new_n4033_), .B(_abc_41234_new_n4031_), .C(_abc_41234_new_n516__bF_buf1), .Y(_abc_41234_new_n4034_));
OAI21X1 OAI21X1_1027 ( .A(_abc_41234_new_n1094_), .B(_abc_41234_new_n3913_), .C(_abc_41234_new_n4034_), .Y(_0sp_15_0__5_));
OAI21X1 OAI21X1_1028 ( .A(_abc_41234_new_n4037_), .B(_abc_41234_new_n4036_), .C(_abc_41234_new_n2452_), .Y(_abc_41234_new_n4038_));
OAI21X1 OAI21X1_1029 ( .A(sp_6_), .B(_abc_41234_new_n4021_), .C(_abc_41234_new_n3936_), .Y(_abc_41234_new_n4043_));
OAI21X1 OAI21X1_103 ( .A(_abc_41234_new_n1056_), .B(_abc_41234_new_n1061_), .C(_abc_41234_new_n1062_), .Y(_abc_41234_new_n1063_));
OAI21X1 OAI21X1_1030 ( .A(_abc_41234_new_n4043_), .B(_abc_41234_new_n4042_), .C(_abc_41234_new_n4038_), .Y(_abc_41234_new_n4044_));
OAI21X1 OAI21X1_1031 ( .A(_abc_41234_new_n2371_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n4048_), .Y(_abc_41234_new_n4049_));
OAI21X1 OAI21X1_1032 ( .A(_abc_41234_new_n1639__bF_buf1), .B(_abc_41234_new_n1637_), .C(_abc_41234_new_n3469_), .Y(_abc_41234_new_n4050_));
OAI21X1 OAI21X1_1033 ( .A(_abc_41234_new_n2415__bF_buf2), .B(_abc_41234_new_n4045_), .C(_abc_41234_new_n4055_), .Y(_abc_41234_new_n4056_));
OAI21X1 OAI21X1_1034 ( .A(_abc_41234_new_n1085_), .B(_abc_41234_new_n3913_), .C(_abc_41234_new_n4057_), .Y(_0sp_15_0__6_));
OAI21X1 OAI21X1_1035 ( .A(_abc_41234_new_n1085_), .B(_abc_41234_new_n4014_), .C(_abc_41234_new_n1080_), .Y(_abc_41234_new_n4060_));
OAI21X1 OAI21X1_1036 ( .A(_abc_41234_new_n2488_), .B(_abc_41234_new_n4061_), .C(_abc_41234_new_n4062_), .Y(_abc_41234_new_n4063_));
OAI21X1 OAI21X1_1037 ( .A(_abc_41234_new_n1080_), .B(_abc_41234_new_n3927_), .C(_abc_41234_new_n4064_), .Y(_abc_41234_new_n4065_));
OAI21X1 OAI21X1_1038 ( .A(_abc_41234_new_n2947__bF_buf3), .B(_abc_41234_new_n4059_), .C(_abc_41234_new_n4066_), .Y(_abc_41234_new_n4067_));
OAI21X1 OAI21X1_1039 ( .A(_abc_41234_new_n555_), .B(_abc_41234_new_n4036_), .C(_abc_41234_new_n3917_), .Y(_abc_41234_new_n4068_));
OAI21X1 OAI21X1_104 ( .A(regfil_2__0_), .B(_abc_41234_new_n1049__bF_buf3), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1065_));
OAI21X1 OAI21X1_1040 ( .A(_abc_41234_new_n2451_), .B(_abc_41234_new_n4070_), .C(_abc_41234_new_n515__bF_buf2), .Y(_abc_41234_new_n4071_));
OAI21X1 OAI21X1_1041 ( .A(sp_7_), .B(_abc_41234_new_n3914__bF_buf1), .C(_abc_41234_new_n660__bF_buf7), .Y(_abc_41234_new_n4073_));
OAI21X1 OAI21X1_1042 ( .A(_abc_41234_new_n3961_), .B(_abc_41234_new_n4061_), .C(_abc_41234_new_n4075_), .Y(_abc_41234_new_n4076_));
OAI21X1 OAI21X1_1043 ( .A(_abc_41234_new_n1080_), .B(_abc_41234_new_n4039_), .C(_abc_41234_new_n1255_), .Y(_abc_41234_new_n4081_));
OAI21X1 OAI21X1_1044 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1107_), .C(_abc_41234_new_n1046__bF_buf4), .Y(_abc_41234_new_n4084_));
OAI21X1 OAI21X1_1045 ( .A(_abc_41234_new_n1255_), .B(_abc_41234_new_n3927_), .C(_abc_41234_new_n4086_), .Y(_abc_41234_new_n4087_));
OAI21X1 OAI21X1_1046 ( .A(_abc_41234_new_n2947__bF_buf2), .B(_abc_41234_new_n4059_), .C(_abc_41234_new_n1255_), .Y(_abc_41234_new_n4088_));
OAI21X1 OAI21X1_1047 ( .A(_abc_41234_new_n2947__bF_buf1), .B(_abc_41234_new_n4080_), .C(_abc_41234_new_n4089_), .Y(_abc_41234_new_n4090_));
OAI21X1 OAI21X1_1048 ( .A(_abc_41234_new_n555_), .B(_abc_41234_new_n4069_), .C(_abc_41234_new_n3917_), .Y(_abc_41234_new_n4091_));
OAI21X1 OAI21X1_1049 ( .A(_abc_41234_new_n2451_), .B(_abc_41234_new_n4092_), .C(_abc_41234_new_n515__bF_buf1), .Y(_abc_41234_new_n4093_));
OAI21X1 OAI21X1_105 ( .A(_abc_41234_new_n1075_), .B(_abc_41234_new_n1074_), .C(_abc_41234_new_n1073_), .Y(_abc_41234_new_n1076_));
OAI21X1 OAI21X1_1050 ( .A(sp_8_), .B(_abc_41234_new_n3914__bF_buf0), .C(_abc_41234_new_n660__bF_buf6), .Y(_abc_41234_new_n4095_));
OAI21X1 OAI21X1_1051 ( .A(_abc_41234_new_n565_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n4097_), .Y(_abc_41234_new_n4098_));
OAI21X1 OAI21X1_1052 ( .A(_abc_41234_new_n2947__bF_buf3), .B(_abc_41234_new_n4080_), .C(_abc_41234_new_n1251_), .Y(_abc_41234_new_n4104_));
OAI21X1 OAI21X1_1053 ( .A(_abc_41234_new_n2451_), .B(_abc_41234_new_n4092_), .C(_abc_41234_new_n1251_), .Y(_abc_41234_new_n4106_));
OAI21X1 OAI21X1_1054 ( .A(sp_8_), .B(_abc_41234_new_n4070_), .C(_abc_41234_new_n2452_), .Y(_abc_41234_new_n4107_));
OAI21X1 OAI21X1_1055 ( .A(_abc_41234_new_n4103_), .B(_abc_41234_new_n4105_), .C(_abc_41234_new_n4109_), .Y(_abc_41234_new_n4110_));
OAI21X1 OAI21X1_1056 ( .A(_abc_41234_new_n1255_), .B(_abc_41234_new_n4059_), .C(_abc_41234_new_n1251_), .Y(_abc_41234_new_n4113_));
OAI21X1 OAI21X1_1057 ( .A(_abc_41234_new_n718_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n4119_), .Y(_abc_41234_new_n4120_));
OAI21X1 OAI21X1_1058 ( .A(_abc_41234_new_n4124_), .B(_abc_41234_new_n4123_), .C(_abc_41234_new_n2452_), .Y(_abc_41234_new_n4125_));
OAI21X1 OAI21X1_1059 ( .A(sp_10_), .B(_abc_41234_new_n4103_), .C(_abc_41234_new_n3936_), .Y(_abc_41234_new_n4128_));
OAI21X1 OAI21X1_106 ( .A(_abc_41234_new_n1070_), .B(_abc_41234_new_n1078_), .C(_abc_41234_new_n1069_), .Y(_abc_41234_new_n1079_));
OAI21X1 OAI21X1_1060 ( .A(_abc_41234_new_n4127_), .B(_abc_41234_new_n4128_), .C(_abc_41234_new_n4125_), .Y(_abc_41234_new_n4129_));
OAI21X1 OAI21X1_1061 ( .A(_abc_41234_new_n1251_), .B(_abc_41234_new_n4080_), .C(_abc_41234_new_n1358_), .Y(_abc_41234_new_n4132_));
OAI21X1 OAI21X1_1062 ( .A(_abc_41234_new_n1637_), .B(_abc_41234_new_n1639__bF_buf0), .C(_abc_41234_new_n3551_), .Y(_abc_41234_new_n4136_));
OAI21X1 OAI21X1_1063 ( .A(_abc_41234_new_n4143_), .B(_abc_41234_new_n4139_), .C(_abc_41234_new_n516__bF_buf5), .Y(_abc_41234_new_n4144_));
OAI21X1 OAI21X1_1064 ( .A(_abc_41234_new_n1358_), .B(_abc_41234_new_n3913_), .C(_abc_41234_new_n4144_), .Y(_0sp_15_0__10_));
OAI21X1 OAI21X1_1065 ( .A(_abc_41234_new_n1358_), .B(_abc_41234_new_n4102_), .C(_abc_41234_new_n1362_), .Y(_abc_41234_new_n4147_));
OAI21X1 OAI21X1_1066 ( .A(_abc_41234_new_n1637_), .B(_abc_41234_new_n1639__bF_buf3), .C(_abc_41234_new_n3573_), .Y(_abc_41234_new_n4150_));
OAI21X1 OAI21X1_1067 ( .A(_abc_41234_new_n819_), .B(_abc_41234_new_n1107_), .C(_abc_41234_new_n1046__bF_buf1), .Y(_abc_41234_new_n4151_));
OAI21X1 OAI21X1_1068 ( .A(sp_0_bF_buf2_), .B(_abc_41234_new_n3549_), .C(sp_11_), .Y(_abc_41234_new_n4154_));
OAI21X1 OAI21X1_1069 ( .A(sp_0_bF_buf1_), .B(_abc_41234_new_n3615_), .C(_abc_41234_new_n4154_), .Y(_abc_41234_new_n4155_));
OAI21X1 OAI21X1_107 ( .A(_abc_41234_new_n1089_), .B(_abc_41234_new_n1101_), .C(_abc_41234_new_n1100_), .Y(_abc_41234_new_n1102_));
OAI21X1 OAI21X1_1070 ( .A(_abc_41234_new_n1362_), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n515__bF_buf6), .Y(_abc_41234_new_n4156_));
OAI21X1 OAI21X1_1071 ( .A(sp_11_), .B(_abc_41234_new_n4127_), .C(_abc_41234_new_n3936_), .Y(_abc_41234_new_n4158_));
OAI21X1 OAI21X1_1072 ( .A(_abc_41234_new_n4158_), .B(_abc_41234_new_n4159_), .C(_abc_41234_new_n4157_), .Y(_abc_41234_new_n4160_));
OAI21X1 OAI21X1_1073 ( .A(_abc_41234_new_n832_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n4164_), .Y(_abc_41234_new_n4165_));
OAI21X1 OAI21X1_1074 ( .A(_abc_41234_new_n4171_), .B(_abc_41234_new_n4170_), .C(_abc_41234_new_n2452_), .Y(_abc_41234_new_n4172_));
OAI21X1 OAI21X1_1075 ( .A(sp_12_), .B(_abc_41234_new_n4159_), .C(_abc_41234_new_n3936_), .Y(_abc_41234_new_n4173_));
OAI21X1 OAI21X1_1076 ( .A(_abc_41234_new_n4173_), .B(_abc_41234_new_n4176_), .C(_abc_41234_new_n4172_), .Y(_abc_41234_new_n4177_));
OAI21X1 OAI21X1_1077 ( .A(_abc_41234_new_n1362_), .B(_abc_41234_new_n4131_), .C(_abc_41234_new_n1408_), .Y(_abc_41234_new_n4179_));
OAI21X1 OAI21X1_1078 ( .A(_abc_41234_new_n2488_), .B(_abc_41234_new_n4180_), .C(_abc_41234_new_n4181_), .Y(_abc_41234_new_n4182_));
OAI21X1 OAI21X1_1079 ( .A(_abc_41234_new_n3961_), .B(_abc_41234_new_n4180_), .C(_abc_41234_new_n4185_), .Y(_abc_41234_new_n4186_));
OAI21X1 OAI21X1_108 ( .A(_abc_41234_new_n1103_), .B(_abc_41234_new_n1104_), .C(_abc_41234_new_n1110_), .Y(_abc_41234_new_n1111_));
OAI21X1 OAI21X1_1080 ( .A(_abc_41234_new_n4186_), .B(_abc_41234_new_n4184_), .C(_abc_41234_new_n516__bF_buf4), .Y(_abc_41234_new_n4187_));
OAI21X1 OAI21X1_1081 ( .A(_abc_41234_new_n1408_), .B(_abc_41234_new_n3913_), .C(_abc_41234_new_n4187_), .Y(_0sp_15_0__12_));
OAI21X1 OAI21X1_1082 ( .A(sp_13_), .B(_abc_41234_new_n4176_), .C(_abc_41234_new_n3936_), .Y(_abc_41234_new_n4191_));
OAI21X1 OAI21X1_1083 ( .A(sp_12_), .B(_abc_41234_new_n4169_), .C(sp_13_), .Y(_abc_41234_new_n4192_));
OAI21X1 OAI21X1_1084 ( .A(sp_0_bF_buf0_), .B(_abc_41234_new_n3618_), .C(_abc_41234_new_n4192_), .Y(_abc_41234_new_n4193_));
OAI21X1 OAI21X1_1085 ( .A(_abc_41234_new_n3279_), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n515__bF_buf4), .Y(_abc_41234_new_n4194_));
OAI21X1 OAI21X1_1086 ( .A(_abc_41234_new_n4190_), .B(_abc_41234_new_n4191_), .C(_abc_41234_new_n4195_), .Y(_abc_41234_new_n4196_));
OAI21X1 OAI21X1_1087 ( .A(_abc_41234_new_n1408_), .B(_abc_41234_new_n4146_), .C(_abc_41234_new_n3279_), .Y(_abc_41234_new_n4197_));
OAI21X1 OAI21X1_1088 ( .A(_abc_41234_new_n1637_), .B(_abc_41234_new_n1639__bF_buf2), .C(_abc_41234_new_n3619_), .Y(_abc_41234_new_n4199_));
OAI21X1 OAI21X1_1089 ( .A(sp_13_), .B(_abc_41234_new_n3914__bF_buf3), .C(_abc_41234_new_n660__bF_buf5), .Y(_abc_41234_new_n4204_));
OAI21X1 OAI21X1_109 ( .A(_abc_41234_new_n1119_), .B(_abc_41234_new_n1120_), .C(_abc_41234_new_n1118_), .Y(_abc_41234_new_n1121_));
OAI21X1 OAI21X1_1090 ( .A(_abc_41234_new_n895_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n4206_), .Y(_abc_41234_new_n4207_));
OAI21X1 OAI21X1_1091 ( .A(sp_14_), .B(_abc_41234_new_n4190_), .C(_abc_41234_new_n3936_), .Y(_abc_41234_new_n4212_));
OAI21X1 OAI21X1_1092 ( .A(sp_0_bF_buf3_), .B(_abc_41234_new_n3618_), .C(sp_14_), .Y(_abc_41234_new_n4214_));
OAI21X1 OAI21X1_1093 ( .A(sp_0_bF_buf2_), .B(_abc_41234_new_n4213_), .C(_abc_41234_new_n4214_), .Y(_abc_41234_new_n4215_));
OAI21X1 OAI21X1_1094 ( .A(_abc_41234_new_n1524_), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n515__bF_buf3), .Y(_abc_41234_new_n4216_));
OAI21X1 OAI21X1_1095 ( .A(_abc_41234_new_n4211_), .B(_abc_41234_new_n4212_), .C(_abc_41234_new_n4217_), .Y(_abc_41234_new_n4218_));
OAI21X1 OAI21X1_1096 ( .A(_abc_41234_new_n3639_), .B(_abc_41234_new_n3638_), .C(_abc_41234_new_n2463_), .Y(_abc_41234_new_n4221_));
OAI21X1 OAI21X1_1097 ( .A(sp_14_), .B(_abc_41234_new_n3914__bF_buf2), .C(_abc_41234_new_n660__bF_buf4), .Y(_abc_41234_new_n4226_));
OAI21X1 OAI21X1_1098 ( .A(_abc_41234_new_n3639_), .B(_abc_41234_new_n3638_), .C(_abc_41234_new_n3963_), .Y(_abc_41234_new_n4229_));
OAI21X1 OAI21X1_1099 ( .A(_abc_41234_new_n2947__bF_buf1), .B(_abc_41234_new_n4210_), .C(_abc_41234_new_n1569_), .Y(_abc_41234_new_n4235_));
OAI21X1 OAI21X1_11 ( .A(_abc_41234_new_n627_), .B(_abc_41234_new_n615_), .C(_abc_41234_new_n628_), .Y(_abc_41234_new_n629_));
OAI21X1 OAI21X1_110 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n899_), .C(_abc_41234_new_n1136_), .Y(_abc_41234_new_n1137_));
OAI21X1 OAI21X1_1100 ( .A(sp_0_bF_buf1_), .B(_abc_41234_new_n4213_), .C(_abc_41234_new_n1569_), .Y(_abc_41234_new_n4237_));
OAI21X1 OAI21X1_1101 ( .A(_abc_41234_new_n1524_), .B(_abc_41234_new_n4189_), .C(_abc_41234_new_n1569_), .Y(_abc_41234_new_n4242_));
OAI21X1 OAI21X1_1102 ( .A(_abc_41234_new_n1569_), .B(_abc_41234_new_n3927_), .C(_abc_41234_new_n4246_), .Y(_abc_41234_new_n4247_));
OAI21X1 OAI21X1_1103 ( .A(sp_15_), .B(_abc_41234_new_n3914__bF_buf1), .C(_abc_41234_new_n660__bF_buf3), .Y(_abc_41234_new_n4249_));
OAI21X1 OAI21X1_1104 ( .A(_abc_41234_new_n585_), .B(_abc_41234_new_n4257_), .C(_abc_41234_new_n4258_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_0_));
OAI21X1 OAI21X1_1105 ( .A(_abc_41234_new_n739_), .B(_abc_41234_new_n4257_), .C(_abc_41234_new_n4260_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_1_));
OAI21X1 OAI21X1_1106 ( .A(_abc_41234_new_n766_), .B(_abc_41234_new_n4257_), .C(_abc_41234_new_n4262_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_2_));
OAI21X1 OAI21X1_1107 ( .A(_abc_41234_new_n805_), .B(_abc_41234_new_n4257_), .C(_abc_41234_new_n4264_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_3_));
OAI21X1 OAI21X1_1108 ( .A(_abc_41234_new_n866_), .B(_abc_41234_new_n4257_), .C(_abc_41234_new_n4266_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_4_));
OAI21X1 OAI21X1_1109 ( .A(_abc_41234_new_n914_), .B(_abc_41234_new_n4257_), .C(_abc_41234_new_n4268_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_5_));
OAI21X1 OAI21X1_111 ( .A(regfil_5__5_), .B(regfil_3__5_), .C(_abc_41234_new_n1137_), .Y(_abc_41234_new_n1138_));
OAI21X1 OAI21X1_1110 ( .A(_abc_41234_new_n944_), .B(_abc_41234_new_n4257_), .C(_abc_41234_new_n4270_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_6_));
OAI21X1 OAI21X1_1111 ( .A(_abc_41234_new_n983_), .B(_abc_41234_new_n4257_), .C(_abc_41234_new_n4272_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_7_));
OAI21X1 OAI21X1_1112 ( .A(_abc_41234_new_n2353_), .B(_abc_41234_new_n606_), .C(_abc_41234_new_n3910_), .Y(_abc_41234_new_n4274_));
OAI21X1 OAI21X1_1113 ( .A(_abc_41234_new_n548_), .B(_abc_41234_new_n1105__bF_buf3), .C(_abc_41234_new_n1856_), .Y(_abc_41234_new_n4278_));
OAI21X1 OAI21X1_1114 ( .A(_abc_41234_new_n555_), .B(_abc_41234_new_n3916_), .C(_abc_41234_new_n538_), .Y(_abc_41234_new_n4279_));
OAI21X1 OAI21X1_1115 ( .A(_abc_41234_new_n1684_), .B(_abc_41234_new_n1051_), .C(_abc_41234_new_n4281_), .Y(_abc_41234_new_n4282_));
OAI21X1 OAI21X1_1116 ( .A(opcode_4_bF_buf1_), .B(_abc_41234_new_n536__bF_buf0), .C(_abc_41234_new_n528_), .Y(_abc_41234_new_n4283_));
OAI21X1 OAI21X1_1117 ( .A(_abc_41234_new_n2933_), .B(_abc_41234_new_n2935_), .C(_abc_41234_new_n4283_), .Y(_abc_41234_new_n4284_));
OAI21X1 OAI21X1_1118 ( .A(_abc_41234_new_n530_), .B(_abc_41234_new_n537__bF_buf3), .C(_abc_41234_new_n1628_), .Y(_abc_41234_new_n4286_));
OAI21X1 OAI21X1_1119 ( .A(_abc_41234_new_n1105__bF_buf2), .B(_abc_41234_new_n1051_), .C(_abc_41234_new_n3935_), .Y(_abc_41234_new_n4292_));
OAI21X1 OAI21X1_112 ( .A(_abc_41234_new_n1131_), .B(_abc_41234_new_n1138_), .C(_abc_41234_new_n1139_), .Y(_abc_41234_new_n1140_));
OAI21X1 OAI21X1_1120 ( .A(_abc_41234_new_n2915_), .B(_abc_41234_new_n4295_), .C(_abc_41234_new_n1647_), .Y(_abc_41234_new_n4296_));
OAI21X1 OAI21X1_1121 ( .A(_abc_41234_new_n665__bF_buf0), .B(_abc_41234_new_n4297__bF_buf3), .C(pc_0_), .Y(_abc_41234_new_n4298_));
OAI21X1 OAI21X1_1122 ( .A(opcode_4_bF_buf0_), .B(_abc_41234_new_n1038_), .C(_abc_41234_new_n4287_), .Y(_abc_41234_new_n4303_));
OAI21X1 OAI21X1_1123 ( .A(_abc_41234_new_n555_), .B(_abc_41234_new_n3916_), .C(_abc_41234_new_n4010_), .Y(_abc_41234_new_n4306_));
OAI21X1 OAI21X1_1124 ( .A(opcode_2_), .B(_abc_41234_new_n620__bF_buf5), .C(_abc_41234_new_n1626_), .Y(_abc_41234_new_n4309_));
OAI21X1 OAI21X1_1125 ( .A(_abc_41234_new_n4301_), .B(_abc_41234_new_n4312_), .C(pc_0_), .Y(_abc_41234_new_n4313_));
OAI21X1 OAI21X1_1126 ( .A(_abc_41234_new_n4309_), .B(_abc_41234_new_n4308_), .C(_abc_41234_new_n1647_), .Y(_abc_41234_new_n4314_));
OAI21X1 OAI21X1_1127 ( .A(pc_0_), .B(_abc_41234_new_n3914__bF_buf0), .C(_abc_41234_new_n4316_), .Y(_abc_41234_new_n4317_));
OAI21X1 OAI21X1_1128 ( .A(_abc_41234_new_n4294_), .B(_abc_41234_new_n4291_), .C(_abc_41234_new_n2707_), .Y(_abc_41234_new_n4320_));
OAI21X1 OAI21X1_1129 ( .A(_abc_41234_new_n2707_), .B(_abc_41234_new_n2916_), .C(_abc_41234_new_n4320_), .Y(_abc_41234_new_n4321_));
OAI21X1 OAI21X1_113 ( .A(_abc_41234_new_n1158_), .B(_abc_41234_new_n1159_), .C(_abc_41234_new_n1157_), .Y(_abc_41234_new_n1160_));
OAI21X1 OAI21X1_1130 ( .A(pc_1_), .B(_abc_41234_new_n2185__bF_buf4), .C(_abc_41234_new_n4322_), .Y(_abc_41234_new_n4323_));
OAI21X1 OAI21X1_1131 ( .A(_abc_41234_new_n4323_), .B(_abc_41234_new_n4321_), .C(_abc_41234_new_n515__bF_buf1), .Y(_abc_41234_new_n4324_));
OAI21X1 OAI21X1_1132 ( .A(_abc_41234_new_n2706_), .B(_abc_41234_new_n4328_), .C(_abc_41234_new_n4331_), .Y(_abc_41234_new_n4332_));
OAI21X1 OAI21X1_1133 ( .A(_abc_41234_new_n4332_), .B(_abc_41234_new_n4327_), .C(_abc_41234_new_n1046__bF_buf6), .Y(_abc_41234_new_n4333_));
OAI21X1 OAI21X1_1134 ( .A(_abc_41234_new_n3914__bF_buf3), .B(_abc_41234_new_n2706_), .C(_abc_41234_new_n4333_), .Y(_abc_41234_new_n4334_));
OAI21X1 OAI21X1_1135 ( .A(_abc_41234_new_n4325_), .B(_abc_41234_new_n4334_), .C(_abc_41234_new_n660__bF_buf0), .Y(_abc_41234_new_n4335_));
OAI21X1 OAI21X1_1136 ( .A(_abc_41234_new_n2739_), .B(_abc_41234_new_n2916_), .C(_abc_41234_new_n4339_), .Y(_abc_41234_new_n4340_));
OAI21X1 OAI21X1_1137 ( .A(pc_2_), .B(_abc_41234_new_n4322_), .C(_abc_41234_new_n515__bF_buf0), .Y(_abc_41234_new_n4342_));
OAI21X1 OAI21X1_1138 ( .A(_abc_41234_new_n2995_), .B(_abc_41234_new_n4328_), .C(_abc_41234_new_n4346_), .Y(_abc_41234_new_n4347_));
OAI21X1 OAI21X1_1139 ( .A(_abc_41234_new_n4347_), .B(_abc_41234_new_n4344_), .C(_abc_41234_new_n1046__bF_buf5), .Y(_abc_41234_new_n4348_));
OAI21X1 OAI21X1_114 ( .A(_abc_41234_new_n1193_), .B(_abc_41234_new_n1196_), .C(_abc_41234_new_n1200_), .Y(_abc_41234_new_n1201_));
OAI21X1 OAI21X1_1140 ( .A(_abc_41234_new_n3914__bF_buf2), .B(_abc_41234_new_n2995_), .C(_abc_41234_new_n4348_), .Y(_abc_41234_new_n4349_));
OAI21X1 OAI21X1_1141 ( .A(_abc_41234_new_n4343_), .B(_abc_41234_new_n4349_), .C(_abc_41234_new_n660__bF_buf7), .Y(_abc_41234_new_n4350_));
OAI21X1 OAI21X1_1142 ( .A(_abc_41234_new_n1614_), .B(_abc_41234_new_n1646_), .C(_abc_41234_new_n1613_), .Y(_abc_41234_new_n4354_));
OAI21X1 OAI21X1_1143 ( .A(_abc_41234_new_n2185__bF_buf3), .B(_abc_41234_new_n4355_), .C(_abc_41234_new_n4356_), .Y(_abc_41234_new_n4357_));
OAI21X1 OAI21X1_1144 ( .A(_abc_41234_new_n4297__bF_buf2), .B(_abc_41234_new_n4357_), .C(_abc_41234_new_n4358_), .Y(_abc_41234_new_n4359_));
OAI21X1 OAI21X1_1145 ( .A(_abc_41234_new_n2564_), .B(_abc_41234_new_n4355_), .C(_abc_41234_new_n4362_), .Y(_abc_41234_new_n4363_));
OAI21X1 OAI21X1_1146 ( .A(_abc_41234_new_n1613_), .B(_abc_41234_new_n4326_), .C(_abc_41234_new_n4364_), .Y(_abc_41234_new_n4365_));
OAI21X1 OAI21X1_1147 ( .A(_abc_41234_new_n4361_), .B(_abc_41234_new_n4365_), .C(_abc_41234_new_n1046__bF_buf4), .Y(_abc_41234_new_n4366_));
OAI21X1 OAI21X1_1148 ( .A(_abc_41234_new_n3914__bF_buf1), .B(_abc_41234_new_n2774_), .C(_abc_41234_new_n4366_), .Y(_abc_41234_new_n4367_));
OAI21X1 OAI21X1_1149 ( .A(_abc_41234_new_n4367_), .B(_abc_41234_new_n4360_), .C(_abc_41234_new_n660__bF_buf6), .Y(_abc_41234_new_n4368_));
OAI21X1 OAI21X1_115 ( .A(_abc_41234_new_n1198_), .B(_abc_41234_new_n1201_), .C(_abc_41234_new_n1156_), .Y(_abc_41234_new_n1202_));
OAI21X1 OAI21X1_1150 ( .A(_abc_41234_new_n2185__bF_buf2), .B(_abc_41234_new_n4371_), .C(_abc_41234_new_n4372_), .Y(_abc_41234_new_n4373_));
OAI21X1 OAI21X1_1151 ( .A(_abc_41234_new_n4297__bF_buf1), .B(_abc_41234_new_n4373_), .C(_abc_41234_new_n515__bF_buf6), .Y(_abc_41234_new_n4374_));
OAI21X1 OAI21X1_1152 ( .A(_abc_41234_new_n4376_), .B(_abc_41234_new_n4375_), .C(_abc_41234_new_n660__bF_buf5), .Y(_abc_41234_new_n4377_));
OAI21X1 OAI21X1_1153 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n1645_), .C(_abc_41234_new_n4379_), .Y(_abc_41234_new_n4380_));
OAI21X1 OAI21X1_1154 ( .A(_abc_41234_new_n2806_), .B(_abc_41234_new_n4326_), .C(_abc_41234_new_n4381_), .Y(_abc_41234_new_n4382_));
OAI21X1 OAI21X1_1155 ( .A(_abc_41234_new_n2656_), .B(_abc_41234_new_n4383_), .C(_abc_41234_new_n4384_), .Y(_abc_41234_new_n4385_));
OAI21X1 OAI21X1_1156 ( .A(_abc_41234_new_n4294_), .B(_abc_41234_new_n4291_), .C(_abc_41234_new_n4388_), .Y(_abc_41234_new_n4389_));
OAI21X1 OAI21X1_1157 ( .A(_abc_41234_new_n2806_), .B(_abc_41234_new_n4353_), .C(_abc_41234_new_n2831_), .Y(_abc_41234_new_n4390_));
OAI21X1 OAI21X1_1158 ( .A(_abc_41234_new_n1617_), .B(_abc_41234_new_n4353_), .C(_abc_41234_new_n4390_), .Y(_abc_41234_new_n4391_));
OAI21X1 OAI21X1_1159 ( .A(pc_5_), .B(_abc_41234_new_n4322_), .C(_abc_41234_new_n515__bF_buf5), .Y(_abc_41234_new_n4394_));
OAI21X1 OAI21X1_116 ( .A(_abc_41234_new_n1202_), .B(_abc_41234_new_n1154_), .C(_abc_41234_new_n1203_), .Y(_abc_41234_new_n1204_));
OAI21X1 OAI21X1_1160 ( .A(_abc_41234_new_n2835_), .B(_abc_41234_new_n4329_), .C(_abc_41234_new_n4398_), .Y(_abc_41234_new_n4399_));
OAI21X1 OAI21X1_1161 ( .A(_abc_41234_new_n2833_), .B(_abc_41234_new_n4328_), .C(_abc_41234_new_n4400_), .Y(_abc_41234_new_n4401_));
OAI21X1 OAI21X1_1162 ( .A(_abc_41234_new_n4401_), .B(_abc_41234_new_n4396_), .C(_abc_41234_new_n1046__bF_buf3), .Y(_abc_41234_new_n4402_));
OAI21X1 OAI21X1_1163 ( .A(_abc_41234_new_n3914__bF_buf3), .B(_abc_41234_new_n2833_), .C(_abc_41234_new_n4402_), .Y(_abc_41234_new_n4403_));
OAI21X1 OAI21X1_1164 ( .A(_abc_41234_new_n4395_), .B(_abc_41234_new_n4403_), .C(_abc_41234_new_n660__bF_buf4), .Y(_abc_41234_new_n4404_));
OAI21X1 OAI21X1_1165 ( .A(_abc_41234_new_n1617_), .B(_abc_41234_new_n4353_), .C(_abc_41234_new_n2865_), .Y(_abc_41234_new_n4409_));
OAI21X1 OAI21X1_1166 ( .A(_abc_41234_new_n2456_), .B(_abc_41234_new_n2931_), .C(_abc_41234_new_n4411_), .Y(_abc_41234_new_n4412_));
OAI21X1 OAI21X1_1167 ( .A(pc_6_), .B(_abc_41234_new_n4322_), .C(_abc_41234_new_n515__bF_buf4), .Y(_abc_41234_new_n4414_));
OAI21X1 OAI21X1_1168 ( .A(_abc_41234_new_n2469_), .B(_abc_41234_new_n1627_), .C(_abc_41234_new_n2858_), .Y(_abc_41234_new_n4416_));
OAI21X1 OAI21X1_1169 ( .A(_abc_41234_new_n2865_), .B(_abc_41234_new_n4326_), .C(_abc_41234_new_n4419_), .Y(_abc_41234_new_n4420_));
OAI21X1 OAI21X1_117 ( .A(_abc_41234_new_n1227_), .B(_abc_41234_new_n1225_), .C(_abc_41234_new_n1144_), .Y(_abc_41234_new_n1228_));
OAI21X1 OAI21X1_1170 ( .A(_abc_41234_new_n3914__bF_buf2), .B(_abc_41234_new_n2855_), .C(_abc_41234_new_n4421_), .Y(_abc_41234_new_n4422_));
OAI21X1 OAI21X1_1171 ( .A(_abc_41234_new_n4415_), .B(_abc_41234_new_n4422_), .C(_abc_41234_new_n660__bF_buf3), .Y(_abc_41234_new_n4423_));
OAI21X1 OAI21X1_1172 ( .A(_abc_41234_new_n2889_), .B(_abc_41234_new_n4328_), .C(_abc_41234_new_n4431_), .Y(_abc_41234_new_n4432_));
OAI21X1 OAI21X1_1173 ( .A(_abc_41234_new_n2882_), .B(_abc_41234_new_n4326_), .C(_abc_41234_new_n4433_), .Y(_abc_41234_new_n4434_));
OAI21X1 OAI21X1_1174 ( .A(_abc_41234_new_n2884_), .B(_abc_41234_new_n2916_), .C(_abc_41234_new_n4437_), .Y(_abc_41234_new_n4438_));
OAI21X1 OAI21X1_1175 ( .A(pc_7_), .B(_abc_41234_new_n4322_), .C(_abc_41234_new_n515__bF_buf3), .Y(_abc_41234_new_n4440_));
OAI21X1 OAI21X1_1176 ( .A(_abc_41234_new_n4439_), .B(_abc_41234_new_n4440_), .C(_abc_41234_new_n4435_), .Y(_abc_41234_new_n4441_));
OAI21X1 OAI21X1_1177 ( .A(_abc_41234_new_n4426_), .B(_abc_41234_new_n4441_), .C(_abc_41234_new_n660__bF_buf2), .Y(_abc_41234_new_n4442_));
OAI21X1 OAI21X1_1178 ( .A(_abc_41234_new_n2882_), .B(_abc_41234_new_n4408_), .C(_abc_41234_new_n1622_), .Y(_abc_41234_new_n4445_));
OAI21X1 OAI21X1_1179 ( .A(_abc_41234_new_n2185__bF_buf0), .B(_abc_41234_new_n4447_), .C(_abc_41234_new_n4449_), .Y(_abc_41234_new_n4450_));
OAI21X1 OAI21X1_118 ( .A(_abc_41234_new_n1065_), .B(_abc_41234_new_n1234_), .C(_abc_41234_new_n1064_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_0_));
OAI21X1 OAI21X1_1180 ( .A(_abc_41234_new_n4297__bF_buf1), .B(_abc_41234_new_n4450_), .C(_abc_41234_new_n515__bF_buf2), .Y(_abc_41234_new_n4451_));
OAI21X1 OAI21X1_1181 ( .A(_abc_41234_new_n2469_), .B(_abc_41234_new_n1627_), .C(_abc_41234_new_n1624_), .Y(_abc_41234_new_n4453_));
OAI21X1 OAI21X1_1182 ( .A(_abc_41234_new_n2564_), .B(_abc_41234_new_n4447_), .C(_abc_41234_new_n4453_), .Y(_abc_41234_new_n4454_));
OAI21X1 OAI21X1_1183 ( .A(_abc_41234_new_n1622_), .B(_abc_41234_new_n4326_), .C(_abc_41234_new_n4456_), .Y(_abc_41234_new_n4457_));
OAI21X1 OAI21X1_1184 ( .A(_abc_41234_new_n3914__bF_buf0), .B(_abc_41234_new_n1653_), .C(_abc_41234_new_n4458_), .Y(_abc_41234_new_n4459_));
OAI21X1 OAI21X1_1185 ( .A(_abc_41234_new_n4452_), .B(_abc_41234_new_n4459_), .C(_abc_41234_new_n660__bF_buf1), .Y(_abc_41234_new_n4460_));
OAI21X1 OAI21X1_1186 ( .A(_abc_41234_new_n1670_), .B(_abc_41234_new_n4326_), .C(_abc_41234_new_n4469_), .Y(_abc_41234_new_n4470_));
OAI21X1 OAI21X1_1187 ( .A(_abc_41234_new_n4464_), .B(_abc_41234_new_n4470_), .C(_abc_41234_new_n1046__bF_buf7), .Y(_abc_41234_new_n4471_));
OAI21X1 OAI21X1_1188 ( .A(_abc_41234_new_n2185__bF_buf5), .B(_abc_41234_new_n4467_), .C(_abc_41234_new_n4472_), .Y(_abc_41234_new_n4473_));
OAI21X1 OAI21X1_1189 ( .A(_abc_41234_new_n4297__bF_buf2), .B(_abc_41234_new_n4473_), .C(_abc_41234_new_n4474_), .Y(_abc_41234_new_n4475_));
OAI21X1 OAI21X1_119 ( .A(_abc_41234_new_n720_), .B(_abc_41234_new_n1060_), .C(_abc_41234_new_n1236_), .Y(_abc_41234_new_n1237_));
OAI21X1 OAI21X1_1190 ( .A(_abc_41234_new_n534__bF_buf4), .B(_abc_41234_new_n4475_), .C(_abc_41234_new_n4471_), .Y(_abc_41234_new_n4476_));
OAI21X1 OAI21X1_1191 ( .A(_abc_41234_new_n4463_), .B(_abc_41234_new_n4476_), .C(_abc_41234_new_n660__bF_buf0), .Y(_abc_41234_new_n4477_));
OAI21X1 OAI21X1_1192 ( .A(_abc_41234_new_n1670_), .B(_abc_41234_new_n4446_), .C(_abc_41234_new_n1705_), .Y(_abc_41234_new_n4482_));
OAI21X1 OAI21X1_1193 ( .A(_abc_41234_new_n2916_), .B(_abc_41234_new_n1709_), .C(_abc_41234_new_n4322_), .Y(_abc_41234_new_n4485_));
OAI21X1 OAI21X1_1194 ( .A(pc_10_), .B(_abc_41234_new_n4322_), .C(_abc_41234_new_n515__bF_buf1), .Y(_abc_41234_new_n4487_));
OAI21X1 OAI21X1_1195 ( .A(_abc_41234_new_n1709_), .B(_abc_41234_new_n4329_), .C(_abc_41234_new_n4490_), .Y(_abc_41234_new_n4491_));
OAI21X1 OAI21X1_1196 ( .A(_abc_41234_new_n4489_), .B(_abc_41234_new_n4492_), .C(_abc_41234_new_n1046__bF_buf6), .Y(_abc_41234_new_n4493_));
OAI21X1 OAI21X1_1197 ( .A(_abc_41234_new_n4488_), .B(_abc_41234_new_n4495_), .C(_abc_41234_new_n660__bF_buf7), .Y(_abc_41234_new_n4496_));
OAI21X1 OAI21X1_1198 ( .A(_abc_41234_new_n1705_), .B(_abc_41234_new_n4465_), .C(_abc_41234_new_n1727_), .Y(_abc_41234_new_n4501_));
OAI21X1 OAI21X1_1199 ( .A(_abc_41234_new_n2185__bF_buf4), .B(_abc_41234_new_n4502_), .C(_abc_41234_new_n4503_), .Y(_abc_41234_new_n4504_));
OAI21X1 OAI21X1_12 ( .A(_abc_41234_new_n606_), .B(_abc_41234_new_n609_), .C(_abc_41234_new_n632_), .Y(_abc_41234_new_n633_));
OAI21X1 OAI21X1_120 ( .A(regfil_2__1_), .B(_abc_41234_new_n1049__bF_buf1), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1239_));
OAI21X1 OAI21X1_1200 ( .A(_abc_41234_new_n4505_), .B(_abc_41234_new_n4504_), .C(_abc_41234_new_n515__bF_buf0), .Y(_abc_41234_new_n4506_));
OAI21X1 OAI21X1_1201 ( .A(_abc_41234_new_n1047__bF_buf2), .B(_abc_41234_new_n4328_), .C(_abc_41234_new_n3914__bF_buf3), .Y(_abc_41234_new_n4507_));
OAI21X1 OAI21X1_1202 ( .A(_abc_41234_new_n2564_), .B(_abc_41234_new_n4502_), .C(_abc_41234_new_n4510_), .Y(_abc_41234_new_n4511_));
OAI21X1 OAI21X1_1203 ( .A(_abc_41234_new_n4509_), .B(_abc_41234_new_n4511_), .C(_abc_41234_new_n1046__bF_buf5), .Y(_abc_41234_new_n4512_));
OAI21X1 OAI21X1_1204 ( .A(_abc_41234_new_n1727_), .B(_abc_41234_new_n4481_), .C(_abc_41234_new_n1750_), .Y(_abc_41234_new_n4517_));
OAI21X1 OAI21X1_1205 ( .A(_abc_41234_new_n2185__bF_buf3), .B(_abc_41234_new_n4519_), .C(_abc_41234_new_n4520_), .Y(_abc_41234_new_n4521_));
OAI21X1 OAI21X1_1206 ( .A(pc_12_), .B(_abc_41234_new_n4322_), .C(_abc_41234_new_n515__bF_buf6), .Y(_abc_41234_new_n4523_));
OAI21X1 OAI21X1_1207 ( .A(_abc_41234_new_n2937_), .B(_abc_41234_new_n4528_), .C(_abc_41234_new_n1756_), .Y(_abc_41234_new_n4529_));
OAI21X1 OAI21X1_1208 ( .A(_abc_41234_new_n4524_), .B(_abc_41234_new_n4533_), .C(_abc_41234_new_n660__bF_buf5), .Y(_abc_41234_new_n4534_));
OAI21X1 OAI21X1_1209 ( .A(_abc_41234_new_n1750_), .B(_abc_41234_new_n4500_), .C(_abc_41234_new_n1775_), .Y(_abc_41234_new_n4538_));
OAI21X1 OAI21X1_121 ( .A(regfil_4__0_), .B(_abc_41234_new_n1214_), .C(regfil_4__1_bF_buf1_), .Y(_abc_41234_new_n1242_));
OAI21X1 OAI21X1_1210 ( .A(_abc_41234_new_n2185__bF_buf2), .B(_abc_41234_new_n4539_), .C(_abc_41234_new_n4540_), .Y(_abc_41234_new_n4541_));
OAI21X1 OAI21X1_1211 ( .A(_abc_41234_new_n4297__bF_buf3), .B(_abc_41234_new_n4541_), .C(_abc_41234_new_n4542_), .Y(_abc_41234_new_n4543_));
OAI21X1 OAI21X1_1212 ( .A(_abc_41234_new_n2937_), .B(_abc_41234_new_n4528_), .C(_abc_41234_new_n1780_), .Y(_abc_41234_new_n4547_));
OAI21X1 OAI21X1_1213 ( .A(_abc_41234_new_n4545_), .B(_abc_41234_new_n4549_), .C(_abc_41234_new_n1046__bF_buf4), .Y(_abc_41234_new_n4550_));
OAI21X1 OAI21X1_1214 ( .A(_abc_41234_new_n3914__bF_buf1), .B(_abc_41234_new_n3273_), .C(_abc_41234_new_n4550_), .Y(_abc_41234_new_n4551_));
OAI21X1 OAI21X1_1215 ( .A(_abc_41234_new_n4544_), .B(_abc_41234_new_n4551_), .C(_abc_41234_new_n660__bF_buf4), .Y(_abc_41234_new_n4552_));
OAI21X1 OAI21X1_1216 ( .A(_abc_41234_new_n1775_), .B(_abc_41234_new_n4518_), .C(_abc_41234_new_n1798_), .Y(_abc_41234_new_n4557_));
OAI21X1 OAI21X1_1217 ( .A(_abc_41234_new_n4559_), .B(_abc_41234_new_n4562_), .C(_abc_41234_new_n4563_), .Y(_abc_41234_new_n4564_));
OAI21X1 OAI21X1_1218 ( .A(_abc_41234_new_n4566_), .B(_abc_41234_new_n4570_), .C(_abc_41234_new_n1046__bF_buf3), .Y(_abc_41234_new_n4571_));
OAI21X1 OAI21X1_1219 ( .A(_abc_41234_new_n3914__bF_buf0), .B(_abc_41234_new_n1804_), .C(_abc_41234_new_n4571_), .Y(_abc_41234_new_n4572_));
OAI21X1 OAI21X1_122 ( .A(_abc_41234_new_n1219_), .B(_abc_41234_new_n1243_), .C(_abc_41234_new_n1049__bF_buf0), .Y(_abc_41234_new_n1244_));
OAI21X1 OAI21X1_1220 ( .A(_abc_41234_new_n4565_), .B(_abc_41234_new_n4572_), .C(_abc_41234_new_n660__bF_buf3), .Y(_abc_41234_new_n4573_));
OAI21X1 OAI21X1_1221 ( .A(_abc_41234_new_n1798_), .B(_abc_41234_new_n1824_), .C(_abc_41234_new_n1828_), .Y(_abc_41234_new_n4576_));
OAI21X1 OAI21X1_1222 ( .A(_abc_41234_new_n1798_), .B(_abc_41234_new_n4537_), .C(_abc_41234_new_n1828_), .Y(_abc_41234_new_n4579_));
OAI21X1 OAI21X1_1223 ( .A(_abc_41234_new_n1798_), .B(_abc_41234_new_n1779_), .C(_abc_41234_new_n1828_), .Y(_abc_41234_new_n4582_));
OAI21X1 OAI21X1_1224 ( .A(_abc_41234_new_n4586_), .B(_abc_41234_new_n4585_), .C(_abc_41234_new_n515__bF_buf5), .Y(_abc_41234_new_n4587_));
OAI21X1 OAI21X1_1225 ( .A(_abc_41234_new_n4588_), .B(_abc_41234_new_n4592_), .C(_abc_41234_new_n1046__bF_buf2), .Y(_abc_41234_new_n4593_));
OAI21X1 OAI21X1_1226 ( .A(waitr), .B(_abc_41234_new_n4601_), .C(_auto_iopadmap_cc_368_execute_45653), .Y(_abc_41234_new_n4602_));
OAI21X1 OAI21X1_1227 ( .A(reset_bF_buf5), .B(_abc_41234_new_n4602_), .C(_abc_41234_new_n4599_), .Y(_0writemem_0_0_));
OAI21X1 OAI21X1_1228 ( .A(_abc_41234_new_n607_), .B(_abc_41234_new_n3959_), .C(_abc_41234_new_n2428_), .Y(_abc_41234_new_n4604_));
OAI21X1 OAI21X1_1229 ( .A(_abc_41234_new_n607_), .B(_abc_41234_new_n698_), .C(_abc_41234_new_n4605_), .Y(_abc_41234_new_n4606_));
OAI21X1 OAI21X1_123 ( .A(_abc_41234_new_n720_), .B(_abc_41234_new_n1231_), .C(_abc_41234_new_n1219_), .Y(_abc_41234_new_n1248_));
OAI21X1 OAI21X1_1230 ( .A(_auto_iopadmap_cc_368_execute_45649), .B(_abc_41234_new_n4608_), .C(_abc_41234_new_n516__bF_buf3), .Y(_abc_41234_new_n4609_));
OAI21X1 OAI21X1_1231 ( .A(_abc_41234_new_n607_), .B(_abc_41234_new_n1850_), .C(_abc_41234_new_n4612_), .Y(_abc_41234_new_n4613_));
OAI21X1 OAI21X1_1232 ( .A(_abc_41234_new_n4613_), .B(_abc_41234_new_n4606_), .C(_abc_41234_new_n516__bF_buf2), .Y(_abc_41234_new_n4614_));
OAI21X1 OAI21X1_1233 ( .A(reset_bF_buf4), .B(_abc_41234_new_n2671_), .C(_abc_41234_new_n4614_), .Y(_abc_41234_new_n4615_));
OAI21X1 OAI21X1_1234 ( .A(_abc_41234_new_n2910_), .B(_abc_41234_new_n2959__bF_buf3), .C(_abc_41234_new_n4616_), .Y(_abc_41234_new_n4617_));
OAI21X1 OAI21X1_1235 ( .A(_abc_41234_new_n2965_), .B(_abc_41234_new_n2959__bF_buf2), .C(_abc_41234_new_n4621_), .Y(_abc_41234_new_n4622_));
OAI21X1 OAI21X1_1236 ( .A(_abc_41234_new_n3003_), .B(_abc_41234_new_n2959__bF_buf1), .C(_abc_41234_new_n4626_), .Y(_abc_41234_new_n4627_));
OAI21X1 OAI21X1_1237 ( .A(_abc_41234_new_n3023_), .B(_abc_41234_new_n2959__bF_buf0), .C(_abc_41234_new_n4631_), .Y(_abc_41234_new_n4632_));
OAI21X1 OAI21X1_1238 ( .A(_abc_41234_new_n3049_), .B(_abc_41234_new_n2959__bF_buf3), .C(_abc_41234_new_n4636_), .Y(_abc_41234_new_n4637_));
OAI21X1 OAI21X1_1239 ( .A(_abc_41234_new_n3074_), .B(_abc_41234_new_n2959__bF_buf2), .C(_abc_41234_new_n4641_), .Y(_abc_41234_new_n4642_));
OAI21X1 OAI21X1_124 ( .A(_abc_41234_new_n1247_), .B(_abc_41234_new_n1248_), .C(_abc_41234_new_n1043_), .Y(_abc_41234_new_n1249_));
OAI21X1 OAI21X1_1240 ( .A(_abc_41234_new_n3101_), .B(_abc_41234_new_n2959__bF_buf1), .C(_abc_41234_new_n4646_), .Y(_abc_41234_new_n4647_));
OAI21X1 OAI21X1_1241 ( .A(_abc_41234_new_n3125_), .B(_abc_41234_new_n2959__bF_buf0), .C(_abc_41234_new_n4651_), .Y(_abc_41234_new_n4652_));
OAI21X1 OAI21X1_1242 ( .A(_abc_41234_new_n4659_), .B(_abc_41234_new_n4615_), .C(_abc_41234_new_n4664_), .Y(_0addr_15_0__9_));
OAI21X1 OAI21X1_1243 ( .A(_abc_41234_new_n4666_), .B(_abc_41234_new_n4615_), .C(_abc_41234_new_n4669_), .Y(_0addr_15_0__10_));
OAI21X1 OAI21X1_1244 ( .A(_abc_41234_new_n4671_), .B(_abc_41234_new_n4615_), .C(_abc_41234_new_n4674_), .Y(_0addr_15_0__11_));
OAI21X1 OAI21X1_1245 ( .A(_abc_41234_new_n4684_), .B(_abc_41234_new_n4615_), .C(_abc_41234_new_n4687_), .Y(_0addr_15_0__14_));
OAI21X1 OAI21X1_1246 ( .A(waitr), .B(_abc_41234_new_n755_), .C(_auto_iopadmap_cc_368_execute_45647), .Y(_abc_41234_new_n4693_));
OAI21X1 OAI21X1_1247 ( .A(_abc_41234_new_n4699_), .B(_abc_41234_new_n4605_), .C(_abc_41234_new_n4698_), .Y(_abc_41234_new_n4700_));
OAI21X1 OAI21X1_1248 ( .A(_abc_41234_new_n4700_), .B(_abc_41234_new_n4697_), .C(_abc_41234_new_n516__bF_buf4), .Y(_abc_41234_new_n4701_));
OAI21X1 OAI21X1_1249 ( .A(_abc_41234_new_n4706_), .B(_abc_41234_new_n4705_), .C(_abc_41234_new_n4703_), .Y(_0writeio_0_0_));
OAI21X1 OAI21X1_125 ( .A(_abc_41234_new_n1254_), .B(_abc_41234_new_n1103_), .C(_abc_41234_new_n1258_), .Y(_abc_41234_new_n1259_));
OAI21X1 OAI21X1_1250 ( .A(_abc_41234_new_n4708_), .B(_abc_41234_new_n4710_), .C(_abc_41234_new_n2604_), .Y(_abc_41234_new_n4711_));
OAI21X1 OAI21X1_1251 ( .A(_abc_41234_new_n4712_), .B(_abc_41234_new_n4714_), .C(_abc_41234_new_n4716_), .Y(_abc_41234_new_n4717_));
OAI21X1 OAI21X1_1252 ( .A(_abc_41234_new_n4717_), .B(_abc_41234_new_n4711_), .C(_abc_41234_new_n2639_), .Y(_abc_41234_new_n4718_));
OAI21X1 OAI21X1_1253 ( .A(statesel_2_), .B(_abc_41234_new_n2588_), .C(_abc_41234_new_n2557_), .Y(_abc_41234_new_n4721_));
OAI21X1 OAI21X1_1254 ( .A(statesel_2_), .B(_abc_41234_new_n4712_), .C(_abc_41234_new_n2604_), .Y(_abc_41234_new_n4723_));
OAI21X1 OAI21X1_1255 ( .A(_abc_41234_new_n4722_), .B(_abc_41234_new_n4723_), .C(_abc_41234_new_n4720_), .Y(_abc_41234_new_n4724_));
OAI21X1 OAI21X1_1256 ( .A(_abc_41234_new_n4713_), .B(_abc_41234_new_n4709_), .C(_abc_41234_new_n4727_), .Y(_abc_41234_new_n4728_));
OAI21X1 OAI21X1_1257 ( .A(_abc_41234_new_n2601_), .B(_abc_41234_new_n4709_), .C(_abc_41234_new_n4731_), .Y(_abc_41234_new_n4732_));
OAI21X1 OAI21X1_1258 ( .A(_abc_41234_new_n4726_), .B(_abc_41234_new_n4728_), .C(_abc_41234_new_n4732_), .Y(_abc_41234_new_n4733_));
OAI21X1 OAI21X1_1259 ( .A(_abc_41234_new_n2996_), .B(_abc_41234_new_n2917_), .C(_abc_41234_new_n4736_), .Y(_abc_41234_new_n4737_));
OAI21X1 OAI21X1_126 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1255_), .C(_abc_41234_new_n1253_), .Y(_abc_41234_new_n1261_));
OAI21X1 OAI21X1_1260 ( .A(_abc_41234_new_n546__bF_buf5), .B(_abc_41234_new_n721_), .C(_abc_41234_new_n616_), .Y(_abc_41234_new_n4740_));
OAI21X1 OAI21X1_1261 ( .A(_abc_41234_new_n529_), .B(opcode_3_bF_buf0_), .C(_abc_41234_new_n4741_), .Y(_abc_41234_new_n4742_));
OAI21X1 OAI21X1_1262 ( .A(_abc_41234_new_n4741_), .B(_abc_41234_new_n4743_), .C(_abc_41234_new_n4742_), .Y(_abc_41234_new_n4744_));
OAI21X1 OAI21X1_1263 ( .A(_abc_41234_new_n555_), .B(zero), .C(_abc_41234_new_n531_), .Y(_abc_41234_new_n4745_));
OAI21X1 OAI21X1_1264 ( .A(_abc_41234_new_n4748_), .B(_abc_41234_new_n4739_), .C(_abc_41234_new_n2450_), .Y(_abc_41234_new_n4749_));
OAI21X1 OAI21X1_1265 ( .A(opcode_3_bF_buf3_), .B(_abc_41234_new_n1105__bF_buf1), .C(_abc_41234_new_n516__bF_buf2), .Y(_abc_41234_new_n4750_));
OAI21X1 OAI21X1_1266 ( .A(parity), .B(_abc_41234_new_n2342_), .C(_abc_41234_new_n4751_), .Y(_abc_41234_new_n4752_));
OAI21X1 OAI21X1_1267 ( .A(_abc_41234_new_n4708_), .B(_abc_41234_new_n4710_), .C(_abc_41234_new_n4762_), .Y(_abc_41234_new_n4763_));
OAI21X1 OAI21X1_1268 ( .A(reset_bF_buf8), .B(_abc_41234_new_n4759_), .C(_abc_41234_new_n4764_), .Y(_abc_41234_new_n4765_));
OAI21X1 OAI21X1_1269 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n2428_), .C(_abc_41234_new_n4776_), .Y(_abc_41234_new_n4777_));
OAI21X1 OAI21X1_127 ( .A(_abc_41234_new_n1261_), .B(_abc_41234_new_n1260_), .C(_abc_41234_new_n1108_), .Y(_abc_41234_new_n1262_));
OAI21X1 OAI21X1_1270 ( .A(opcode_5_bF_buf2_), .B(_abc_41234_new_n1610_), .C(_abc_41234_new_n4280_), .Y(_abc_41234_new_n4785_));
OAI21X1 OAI21X1_1271 ( .A(_abc_41234_new_n4791_), .B(_abc_41234_new_n4780_), .C(_abc_41234_new_n4719_), .Y(_abc_41234_new_n4792_));
OAI21X1 OAI21X1_1272 ( .A(_abc_41234_new_n4714_), .B(_abc_41234_new_n4712_), .C(_abc_41234_new_n4721_), .Y(_abc_41234_new_n4793_));
OAI21X1 OAI21X1_1273 ( .A(_abc_41234_new_n2556_), .B(_abc_41234_new_n4710_), .C(_abc_41234_new_n4716_), .Y(_abc_41234_new_n4794_));
OAI21X1 OAI21X1_1274 ( .A(_abc_41234_new_n4790_), .B(_abc_41234_new_n4792_), .C(_abc_41234_new_n4795_), .Y(_abc_41234_new_n4796_));
OAI21X1 OAI21X1_1275 ( .A(_abc_41234_new_n2449_), .B(_abc_41234_new_n2481_), .C(_abc_41234_new_n4797_), .Y(_abc_41234_new_n4798_));
OAI21X1 OAI21X1_1276 ( .A(_abc_41234_new_n2533_), .B(_abc_41234_new_n2525_), .C(_abc_41234_new_n4801_), .Y(_abc_41234_new_n4802_));
OAI21X1 OAI21X1_1277 ( .A(_abc_41234_new_n4716_), .B(_abc_41234_new_n4802_), .C(_abc_41234_new_n4807_), .Y(_abc_41234_new_n4808_));
OAI21X1 OAI21X1_1278 ( .A(_abc_41234_new_n2640_), .B(_abc_41234_new_n4809_), .C(_abc_41234_new_n4810_), .Y(_abc_41234_new_n4811_));
OAI21X1 OAI21X1_1279 ( .A(_abc_41234_new_n4822_), .B(_abc_41234_new_n4821_), .C(_abc_41234_new_n4824_), .Y(_abc_41234_new_n4825_));
OAI21X1 OAI21X1_128 ( .A(_abc_41234_new_n1145_), .B(_abc_41234_new_n1148_), .C(_abc_41234_new_n1266_), .Y(_abc_41234_new_n1268_));
OAI21X1 OAI21X1_1280 ( .A(_abc_41234_new_n4827_), .B(_abc_41234_new_n4761_), .C(_abc_41234_new_n2639_), .Y(_abc_41234_new_n4828_));
OAI21X1 OAI21X1_1281 ( .A(reset_bF_buf4), .B(_abc_41234_new_n4841_), .C(_abc_41234_new_n4842_), .Y(_abc_41234_new_n4843_));
OAI21X1 OAI21X1_1282 ( .A(_abc_41234_new_n4827_), .B(_abc_41234_new_n2622_), .C(_abc_41234_new_n4729_), .Y(_abc_41234_new_n4848_));
OAI21X1 OAI21X1_1283 ( .A(_abc_41234_new_n2640_), .B(_abc_41234_new_n4847_), .C(_abc_41234_new_n4848_), .Y(_abc_41234_new_n4849_));
OAI21X1 OAI21X1_1284 ( .A(_abc_41234_new_n4849_), .B(_abc_41234_new_n4850_), .C(_abc_41234_new_n2535_), .Y(_abc_41234_new_n4851_));
OAI21X1 OAI21X1_1285 ( .A(_abc_41234_new_n4821_), .B(_abc_41234_new_n4845_), .C(_abc_41234_new_n4853_), .Y(_abc_41234_new_n4854_));
OAI21X1 OAI21X1_1286 ( .A(_abc_41234_new_n4845_), .B(_abc_41234_new_n4802_), .C(_abc_41234_new_n4834_), .Y(_abc_41234_new_n4862_));
OAI21X1 OAI21X1_1287 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n4704_), .C(_abc_41234_new_n4851_), .Y(_abc_41234_new_n4863_));
OAI21X1 OAI21X1_1288 ( .A(_abc_41234_new_n609_), .B(_abc_41234_new_n698_), .C(_abc_41234_new_n4832_), .Y(_abc_41234_new_n4872_));
OAI21X1 OAI21X1_1289 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n4601_), .C(_abc_41234_new_n4873_), .Y(_abc_41234_new_n4874_));
OAI21X1 OAI21X1_129 ( .A(_abc_41234_new_n1194_), .B(_abc_41234_new_n1192_), .C(_abc_41234_new_n1274_), .Y(_abc_41234_new_n1275_));
OAI21X1 OAI21X1_1290 ( .A(_abc_41234_new_n4716_), .B(_abc_41234_new_n4821_), .C(_abc_41234_new_n4852_), .Y(_abc_41234_new_n4879_));
OAI21X1 OAI21X1_1291 ( .A(_abc_41234_new_n4708_), .B(_abc_41234_new_n4710_), .C(_abc_41234_new_n4822_), .Y(_abc_41234_new_n4884_));
OAI21X1 OAI21X1_1292 ( .A(_abc_41234_new_n4766_), .B(_abc_41234_new_n4884_), .C(_abc_41234_new_n4760_), .Y(_abc_41234_new_n4885_));
OAI21X1 OAI21X1_1293 ( .A(_abc_41234_new_n4768_), .B(_abc_41234_new_n4780_), .C(_abc_41234_new_n4760_), .Y(_abc_41234_new_n4886_));
OAI21X1 OAI21X1_1294 ( .A(_abc_41234_new_n4605_), .B(_abc_41234_new_n4889_), .C(_abc_41234_new_n4892_), .Y(_0ei_0_0_));
OAI21X1 OAI21X1_1295 ( .A(alu__abc_40887_new_n45_), .B(alu__abc_40887_new_n44_), .C(alu__abc_40887_new_n43_), .Y(alu__abc_40887_new_n46_));
OAI21X1 OAI21X1_1296 ( .A(alu__abc_40887_new_n56_), .B(alu__abc_40887_new_n59_), .C(alu__abc_40887_new_n60_), .Y(alu__abc_40887_new_n65_));
OAI21X1 OAI21X1_1297 ( .A(alu__abc_40887_new_n65_), .B(alu__abc_40887_new_n64_), .C(alu__abc_40887_new_n42_), .Y(alu__abc_40887_new_n66_));
OAI21X1 OAI21X1_1298 ( .A(alu__abc_40887_new_n63_), .B(alu__abc_40887_new_n78_), .C(alu__abc_40887_new_n79_), .Y(alu__abc_40887_new_n80_));
OAI21X1 OAI21X1_1299 ( .A(alu__abc_40887_new_n47_), .B(alu__abc_40887_new_n82_), .C(alu__abc_40887_new_n84_), .Y(alu__abc_40887_new_n85_));
OAI21X1 OAI21X1_13 ( .A(_abc_41234_new_n640_), .B(_abc_41234_new_n636_), .C(regfil_0__0_), .Y(_abc_41234_new_n643_));
OAI21X1 OAI21X1_130 ( .A(_abc_41234_new_n1192_), .B(_abc_41234_new_n1277_), .C(_abc_41234_new_n1278_), .Y(_abc_41234_new_n1279_));
OAI21X1 OAI21X1_1300 ( .A(alu__abc_40887_new_n33_), .B(alu__abc_40887_new_n35_), .C(alu__abc_40887_new_n105_), .Y(alu__abc_40887_new_n106_));
OAI21X1 OAI21X1_1301 ( .A(alu__abc_40887_new_n97_), .B(alu__abc_40887_new_n78_), .C(alu__abc_40887_new_n77_), .Y(alu__abc_40887_new_n109_));
OAI21X1 OAI21X1_1302 ( .A(alu__abc_40887_new_n123_), .B(alu__abc_40887_new_n52_), .C(alu__abc_40887_new_n121_), .Y(alu__abc_40887_new_n124_));
OAI21X1 OAI21X1_1303 ( .A(alu__abc_40887_new_n44_), .B(alu__abc_40887_new_n127_), .C(alu__abc_40887_new_n129_), .Y(alu__abc_40887_new_n130_));
OAI21X1 OAI21X1_1304 ( .A(alu__abc_40887_new_n59_), .B(alu__abc_40887_new_n61_), .C(alu__abc_40887_new_n97_), .Y(alu__abc_40887_new_n133_));
OAI21X1 OAI21X1_1305 ( .A(alu__abc_40887_new_n124_), .B(alu__abc_40887_new_n132_), .C(alu__abc_40887_new_n134_), .Y(alu__abc_40887_new_n135_));
OAI21X1 OAI21X1_1306 ( .A(alu__abc_40887_new_n59_), .B(alu__abc_40887_new_n61_), .C(alu__abc_40887_new_n138_), .Y(alu__abc_40887_new_n139_));
OAI21X1 OAI21X1_1307 ( .A(alu_oprb_5_), .B(alu__abc_40887_new_n136_), .C(alu__abc_40887_new_n139_), .Y(alu__abc_40887_new_n140_));
OAI21X1 OAI21X1_1308 ( .A(alu__abc_40887_new_n144_), .B(alu__abc_40887_new_n142_), .C(alu__abc_40887_new_n37_), .Y(alu__abc_40887_new_n145_));
OAI21X1 OAI21X1_1309 ( .A(alu__abc_40887_new_n148_), .B(alu__abc_40887_new_n149_), .C(alu__abc_40887_new_n152_), .Y(alu__abc_40887_new_n153_));
OAI21X1 OAI21X1_131 ( .A(_abc_41234_new_n1276_), .B(_abc_41234_new_n1279_), .C(_abc_41234_new_n1156_), .Y(_abc_41234_new_n1280_));
OAI21X1 OAI21X1_1310 ( .A(alu__abc_40887_new_n140_), .B(alu__abc_40887_new_n154_), .C(alu__abc_40887_new_n41_), .Y(alu__abc_40887_new_n155_));
OAI21X1 OAI21X1_1311 ( .A(alu__abc_40887_new_n146_), .B(alu__abc_40887_new_n160_), .C(alu__abc_40887_new_n84_), .Y(alu__abc_40887_new_n161_));
OAI21X1 OAI21X1_1312 ( .A(alu__abc_40887_new_n148_), .B(alu__abc_40887_new_n149_), .C(alu__abc_40887_new_n162_), .Y(alu__abc_40887_new_n163_));
OAI21X1 OAI21X1_1313 ( .A(alu__abc_40887_new_n124_), .B(alu__abc_40887_new_n132_), .C(alu__abc_40887_new_n97_), .Y(alu__abc_40887_new_n175_));
OAI21X1 OAI21X1_1314 ( .A(alu__abc_40887_new_n58_), .B(alu__abc_40887_new_n177_), .C(alu__abc_40887_new_n179_), .Y(alu__abc_40887_new_n180_));
OAI21X1 OAI21X1_1315 ( .A(alu__abc_40887_new_n133_), .B(alu__abc_40887_new_n177_), .C(alu__abc_40887_new_n139_), .Y(alu__abc_40887_new_n188_));
OAI21X1 OAI21X1_1316 ( .A(alu__abc_40887_new_n149_), .B(alu__abc_40887_new_n192_), .C(alu__abc_40887_new_n168_), .Y(alu__abc_40887_new_n193_));
OAI21X1 OAI21X1_1317 ( .A(alu__abc_40887_new_n186_), .B(alu__abc_40887_new_n197_), .C(alu__abc_40887_new_n118_), .Y(alu__abc_40887_new_n198_));
OAI21X1 OAI21X1_1318 ( .A(alu_sel_2_), .B(alu__abc_40887_new_n203_), .C(alu__abc_40887_new_n204_), .Y(alu__abc_40887_new_n205_));
OAI21X1 OAI21X1_1319 ( .A(alu__abc_40887_new_n110_), .B(alu__abc_40887_new_n111_), .C(alu__abc_40887_new_n74_), .Y(alu__abc_40887_new_n220_));
OAI21X1 OAI21X1_132 ( .A(_abc_41234_new_n1270_), .B(_abc_41234_new_n1280_), .C(_abc_41234_new_n1281_), .Y(_abc_41234_new_n1282_));
OAI21X1 OAI21X1_1320 ( .A(alu__abc_40887_new_n189_), .B(alu__abc_40887_new_n195_), .C(alu__abc_40887_new_n159_), .Y(alu__abc_40887_new_n223_));
OAI21X1 OAI21X1_1321 ( .A(alu__abc_40887_new_n172_), .B(alu__abc_40887_new_n237_), .C(alu__abc_40887_new_n118_), .Y(alu__abc_40887_new_n238_));
OAI21X1 OAI21X1_1322 ( .A(alu__abc_40887_new_n167_), .B(alu__abc_40887_new_n239_), .C(alu__abc_40887_new_n235_), .Y(alu__abc_40887_new_n240_));
OAI21X1 OAI21X1_1323 ( .A(alu__abc_40887_new_n115_), .B(alu__abc_40887_new_n127_), .C(alu__abc_40887_new_n199_), .Y(alu__abc_40887_new_n244_));
OAI21X1 OAI21X1_1324 ( .A(alu__abc_40887_new_n44_), .B(alu__abc_40887_new_n208_), .C(alu__abc_40887_new_n244_), .Y(alu__abc_40887_new_n245_));
OAI21X1 OAI21X1_1325 ( .A(alu__abc_40887_new_n236_), .B(alu__abc_40887_new_n243_), .C(alu__abc_40887_new_n246_), .Y(alu__abc_40887_new_n247_));
OAI21X1 OAI21X1_1326 ( .A(alu__abc_40887_new_n104_), .B(alu__abc_40887_new_n118_), .C(alu__abc_40887_new_n92_), .Y(alu__abc_40887_new_n252_));
OAI21X1 OAI21X1_1327 ( .A(alu_oprb_0_), .B(alu_opra_0_), .C(alu__abc_40887_new_n209_), .Y(alu__abc_40887_new_n254_));
OAI21X1 OAI21X1_1328 ( .A(alu__abc_40887_new_n45_), .B(alu__abc_40887_new_n211_), .C(alu__abc_40887_new_n254_), .Y(alu__abc_40887_new_n255_));
OAI21X1 OAI21X1_1329 ( .A(alu__abc_40887_new_n174_), .B(alu__abc_40887_new_n259_), .C(alu__abc_40887_new_n118_), .Y(alu__abc_40887_new_n260_));
OAI21X1 OAI21X1_133 ( .A(_abc_41234_new_n1259_), .B(_abc_41234_new_n1262_), .C(_abc_41234_new_n1283_), .Y(_abc_41234_new_n1284_));
OAI21X1 OAI21X1_1330 ( .A(alu__abc_40887_new_n271_), .B(alu__abc_40887_new_n193_), .C(alu__abc_40887_new_n287_), .Y(alu__abc_40887_new_n288_));
OAI21X1 OAI21X1_1331 ( .A(alu__abc_40887_new_n194_), .B(alu__abc_40887_new_n294_), .C(alu__abc_40887_new_n118_), .Y(alu__abc_40887_new_n295_));
OAI21X1 OAI21X1_1332 ( .A(alu__abc_40887_new_n289_), .B(alu__abc_40887_new_n293_), .C(alu__abc_40887_new_n298_), .Y(alu__abc_40887_new_n299_));
OAI21X1 OAI21X1_1333 ( .A(alu__abc_40887_new_n302_), .B(alu__abc_40887_new_n303_), .C(alu__abc_40887_new_n301_), .Y(alu__abc_40887_new_n304_));
OAI21X1 OAI21X1_1334 ( .A(alu__abc_40887_new_n306_), .B(alu__abc_40887_new_n290_), .C(alu__abc_40887_new_n110_), .Y(alu__abc_40887_new_n307_));
OAI21X1 OAI21X1_1335 ( .A(alu__abc_40887_new_n154_), .B(alu__abc_40887_new_n309_), .C(alu__abc_40887_new_n195_), .Y(alu__abc_40887_new_n310_));
OAI21X1 OAI21X1_1336 ( .A(alu__abc_40887_new_n60_), .B(alu__abc_40887_new_n211_), .C(alu__abc_40887_new_n314_), .Y(alu__abc_40887_new_n315_));
OAI21X1 OAI21X1_1337 ( .A(alu__abc_40887_new_n290_), .B(alu__abc_40887_new_n306_), .C(alu__abc_40887_new_n320_), .Y(alu__abc_40887_new_n321_));
OAI21X1 OAI21X1_1338 ( .A(alu__abc_40887_new_n322_), .B(alu__abc_40887_new_n323_), .C(alu__abc_40887_new_n118_), .Y(alu__abc_40887_new_n324_));
OAI21X1 OAI21X1_1339 ( .A(alu_oprb_4_), .B(alu_opra_4_), .C(alu__abc_40887_new_n209_), .Y(alu__abc_40887_new_n325_));
OAI21X1 OAI21X1_134 ( .A(_abc_41234_new_n1239_), .B(_abc_41234_new_n1285_), .C(_abc_41234_new_n1238_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_1_));
OAI21X1 OAI21X1_1340 ( .A(alu__abc_40887_new_n97_), .B(alu__abc_40887_new_n210_), .C(alu__abc_40887_new_n325_), .Y(alu__abc_40887_new_n326_));
OAI21X1 OAI21X1_1341 ( .A(alu__abc_40887_new_n243_), .B(alu__abc_40887_new_n190_), .C(alu__abc_40887_new_n328_), .Y(alu__abc_40887_new_n329_));
OAI21X1 OAI21X1_1342 ( .A(alu__abc_40887_new_n81_), .B(alu__abc_40887_new_n314_), .C(alu__abc_40887_new_n318_), .Y(alu__abc_40887_new_n333_));
OAI21X1 OAI21X1_1343 ( .A(alu__abc_40887_new_n302_), .B(alu__abc_40887_new_n303_), .C(alu__abc_40887_new_n258_), .Y(alu__abc_40887_new_n338_));
OAI21X1 OAI21X1_1344 ( .A(alu__abc_40887_new_n251_), .B(alu__abc_40887_new_n256_), .C(alu__abc_40887_new_n204_), .Y(alu__abc_40887_new_n354_));
OAI21X1 OAI21X1_1345 ( .A(alu__abc_40887_new_n128_), .B(alu__abc_40887_new_n204_), .C(alu__abc_40887_new_n354_), .Y(alu_res_0_));
OAI21X1 OAI21X1_1346 ( .A(alu__abc_40887_new_n125_), .B(alu__abc_40887_new_n204_), .C(alu__abc_40887_new_n356_), .Y(alu_res_1_));
OAI21X1 OAI21X1_1347 ( .A(alu__abc_40887_new_n150_), .B(alu__abc_40887_new_n204_), .C(alu__abc_40887_new_n358_), .Y(alu_res_2_));
OAI21X1 OAI21X1_1348 ( .A(alu__abc_40887_new_n289_), .B(alu__abc_40887_new_n293_), .C(alu__abc_40887_new_n204_), .Y(alu__abc_40887_new_n360_));
OAI21X1 OAI21X1_1349 ( .A(alu__abc_40887_new_n119_), .B(alu__abc_40887_new_n204_), .C(alu__abc_40887_new_n360_), .Y(alu_res_3_));
OAI21X1 OAI21X1_135 ( .A(_abc_41234_new_n1058_), .B(_abc_41234_new_n1059_), .C(regfil_4__2_bF_buf2_), .Y(_abc_41234_new_n1287_));
OAI21X1 OAI21X1_1350 ( .A(alu__abc_40887_new_n137_), .B(alu__abc_40887_new_n204_), .C(alu__abc_40887_new_n362_), .Y(alu_res_4_));
OAI21X1 OAI21X1_1351 ( .A(alu__abc_40887_new_n143_), .B(alu__abc_40887_new_n204_), .C(alu__abc_40887_new_n365_), .Y(alu_res_6_));
OAI21X1 OAI21X1_1352 ( .A(alu__abc_40887_new_n367_), .B(alu__abc_40887_new_n204_), .C(alu__abc_40887_new_n368_), .Y(alu_res_7_));
OAI21X1 OAI21X1_1353 ( .A(alu_oprb_7_), .B(alu__abc_40887_new_n367_), .C(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n371_));
OAI21X1 OAI21X1_1354 ( .A(alu__abc_40887_new_n270_), .B(alu__abc_40887_new_n370_), .C(alu__abc_40887_new_n371_), .Y(alu__abc_40887_new_n372_));
OAI21X1 OAI21X1_1355 ( .A(alu__abc_40887_new_n118_), .B(alu__abc_40887_new_n205_), .C(alu__abc_40887_new_n372_), .Y(alu__abc_40887_new_n373_));
OAI21X1 OAI21X1_1356 ( .A(alu__abc_40887_new_n33_), .B(alu__abc_40887_new_n375_), .C(alu__abc_40887_new_n34_), .Y(alu__abc_40887_new_n376_));
OAI21X1 OAI21X1_1357 ( .A(alu__abc_40887_new_n104_), .B(alu__abc_40887_new_n201_), .C(alu__abc_40887_new_n376_), .Y(alu__abc_40887_new_n377_));
OAI21X1 OAI21X1_136 ( .A(_abc_41234_new_n1061_), .B(_abc_41234_new_n790_), .C(_abc_41234_new_n1287_), .Y(_abc_41234_new_n1288_));
OAI21X1 OAI21X1_137 ( .A(regfil_2__2_), .B(_abc_41234_new_n1049__bF_buf4), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1290_));
OAI21X1 OAI21X1_138 ( .A(regfil_4__2_bF_buf0_), .B(_abc_41234_new_n1241_), .C(_abc_41234_new_n1291_), .Y(_abc_41234_new_n1292_));
OAI21X1 OAI21X1_139 ( .A(_abc_41234_new_n720_), .B(_abc_41234_new_n1231_), .C(_abc_41234_new_n773_), .Y(_abc_41234_new_n1293_));
OAI21X1 OAI21X1_14 ( .A(_abc_41234_new_n613_), .B(_abc_41234_new_n650_), .C(_abc_41234_new_n649_), .Y(_abc_41234_new_n651_));
OAI21X1 OAI21X1_140 ( .A(_abc_41234_new_n1254_), .B(_abc_41234_new_n1103_), .C(_abc_41234_new_n1296_), .Y(_abc_41234_new_n1297_));
OAI21X1 OAI21X1_141 ( .A(regfil_2__1_), .B(regfil_4__1_bF_buf3_), .C(_abc_41234_new_n1145_), .Y(_abc_41234_new_n1312_));
OAI21X1 OAI21X1_142 ( .A(_abc_41234_new_n731_), .B(_abc_41234_new_n720_), .C(_abc_41234_new_n1312_), .Y(_abc_41234_new_n1313_));
OAI21X1 OAI21X1_143 ( .A(_abc_41234_new_n1313_), .B(_abc_41234_new_n1311_), .C(_abc_41234_new_n1317_), .Y(_abc_41234_new_n1318_));
OAI21X1 OAI21X1_144 ( .A(_abc_41234_new_n1314_), .B(_abc_41234_new_n1315_), .C(_abc_41234_new_n1319_), .Y(_abc_41234_new_n1320_));
OAI21X1 OAI21X1_145 ( .A(_abc_41234_new_n1271_), .B(_abc_41234_new_n1274_), .C(_abc_41234_new_n1326_), .Y(_abc_41234_new_n1327_));
OAI21X1 OAI21X1_146 ( .A(_abc_41234_new_n1277_), .B(_abc_41234_new_n1192_), .C(_abc_41234_new_n1328_), .Y(_abc_41234_new_n1329_));
OAI21X1 OAI21X1_147 ( .A(_abc_41234_new_n1290_), .B(_abc_41234_new_n1341_), .C(_abc_41234_new_n1289_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_2_));
OAI21X1 OAI21X1_148 ( .A(regfil_2__3_), .B(_abc_41234_new_n1049__bF_buf3), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1347_));
OAI21X1 OAI21X1_149 ( .A(regfil_4__2_bF_buf1_), .B(_abc_41234_new_n1241_), .C(regfil_4__3_), .Y(_abc_41234_new_n1351_));
OAI21X1 OAI21X1_15 ( .A(opcode_5_bF_buf1_), .B(_abc_41234_new_n615_), .C(_abc_41234_new_n651_), .Y(_abc_41234_new_n652_));
OAI21X1 OAI21X1_150 ( .A(_abc_41234_new_n1355_), .B(_abc_41234_new_n1354_), .C(_abc_41234_new_n1219_), .Y(_abc_41234_new_n1356_));
OAI21X1 OAI21X1_151 ( .A(_abc_41234_new_n1218_), .B(_abc_41234_new_n1206_), .C(_abc_41234_new_n1356_), .Y(_abc_41234_new_n1357_));
OAI21X1 OAI21X1_152 ( .A(_abc_41234_new_n1252_), .B(_abc_41234_new_n1259_), .C(_abc_41234_new_n1301_), .Y(_abc_41234_new_n1359_));
OAI21X1 OAI21X1_153 ( .A(_abc_41234_new_n773_), .B(_abc_41234_new_n1358_), .C(_abc_41234_new_n1359_), .Y(_abc_41234_new_n1360_));
OAI21X1 OAI21X1_154 ( .A(_abc_41234_new_n769_), .B(_abc_41234_new_n773_), .C(_abc_41234_new_n1318_), .Y(_abc_41234_new_n1370_));
OAI21X1 OAI21X1_155 ( .A(_abc_41234_new_n1370_), .B(_abc_41234_new_n1371_), .C(_abc_41234_new_n1372_), .Y(_abc_41234_new_n1373_));
OAI21X1 OAI21X1_156 ( .A(_abc_41234_new_n1378_), .B(_abc_41234_new_n1374_), .C(_abc_41234_new_n1200_), .Y(_abc_41234_new_n1380_));
OAI21X1 OAI21X1_157 ( .A(_abc_41234_new_n1379_), .B(_abc_41234_new_n1380_), .C(_abc_41234_new_n1152_), .Y(_abc_41234_new_n1381_));
OAI21X1 OAI21X1_158 ( .A(_abc_41234_new_n1347_), .B(_abc_41234_new_n1384_), .C(_abc_41234_new_n1346_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_3_));
OAI21X1 OAI21X1_159 ( .A(regfil_2__4_), .B(_abc_41234_new_n1049__bF_buf2), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1390_));
OAI21X1 OAI21X1_16 ( .A(opcode_4_bF_buf1_), .B(opcode_3_bF_buf2_), .C(opcode_5_bF_buf0_), .Y(_abc_41234_new_n666_));
OAI21X1 OAI21X1_160 ( .A(_abc_41234_new_n1393_), .B(_abc_41234_new_n1392_), .C(_abc_41234_new_n1218_), .Y(_abc_41234_new_n1394_));
OAI21X1 OAI21X1_161 ( .A(_abc_41234_new_n525__bF_buf0), .B(_abc_41234_new_n1217_), .C(_abc_41234_new_n1397_), .Y(_abc_41234_new_n1398_));
OAI21X1 OAI21X1_162 ( .A(_abc_41234_new_n1396_), .B(_abc_41234_new_n1398_), .C(_abc_41234_new_n1043_), .Y(_abc_41234_new_n1399_));
OAI21X1 OAI21X1_163 ( .A(regfil_4__3_), .B(sp_11_), .C(_abc_41234_new_n1300_), .Y(_abc_41234_new_n1403_));
OAI21X1 OAI21X1_164 ( .A(_abc_41234_new_n819_), .B(_abc_41234_new_n1362_), .C(_abc_41234_new_n1403_), .Y(_abc_41234_new_n1404_));
OAI21X1 OAI21X1_165 ( .A(_abc_41234_new_n1401_), .B(_abc_41234_new_n1103_), .C(_abc_41234_new_n1405_), .Y(_abc_41234_new_n1406_));
OAI21X1 OAI21X1_166 ( .A(_abc_41234_new_n1410_), .B(_abc_41234_new_n1406_), .C(_abc_41234_new_n1108_), .Y(_abc_41234_new_n1412_));
OAI21X1 OAI21X1_167 ( .A(regfil_2__3_), .B(regfil_4__3_), .C(_abc_41234_new_n1315_), .Y(_abc_41234_new_n1415_));
OAI21X1 OAI21X1_168 ( .A(_abc_41234_new_n815_), .B(_abc_41234_new_n819_), .C(_abc_41234_new_n1415_), .Y(_abc_41234_new_n1416_));
OAI21X1 OAI21X1_169 ( .A(_abc_41234_new_n1414_), .B(_abc_41234_new_n1141_), .C(_abc_41234_new_n1417_), .Y(_abc_41234_new_n1418_));
OAI21X1 OAI21X1_17 ( .A(_abc_41234_new_n555_), .B(_abc_41234_new_n536__bF_buf3), .C(_abc_41234_new_n667_), .Y(_abc_41234_new_n668_));
OAI21X1 OAI21X1_170 ( .A(_abc_41234_new_n1421_), .B(_abc_41234_new_n1418_), .C(_abc_41234_new_n1151_), .Y(_abc_41234_new_n1422_));
OAI21X1 OAI21X1_171 ( .A(_abc_41234_new_n1331_), .B(_abc_41234_new_n1376_), .C(_abc_41234_new_n1375_), .Y(_abc_41234_new_n1428_));
OAI21X1 OAI21X1_172 ( .A(_abc_41234_new_n1432_), .B(_abc_41234_new_n1192_), .C(_abc_41234_new_n1431_), .Y(_abc_41234_new_n1433_));
OAI21X1 OAI21X1_173 ( .A(_abc_41234_new_n1427_), .B(_abc_41234_new_n1433_), .C(_abc_41234_new_n1200_), .Y(_abc_41234_new_n1435_));
OAI21X1 OAI21X1_174 ( .A(_abc_41234_new_n1434_), .B(_abc_41234_new_n1435_), .C(_abc_41234_new_n1156_), .Y(_abc_41234_new_n1436_));
OAI21X1 OAI21X1_175 ( .A(_abc_41234_new_n1436_), .B(_abc_41234_new_n1423_), .C(_abc_41234_new_n1437_), .Y(_abc_41234_new_n1438_));
OAI21X1 OAI21X1_176 ( .A(_abc_41234_new_n1411_), .B(_abc_41234_new_n1412_), .C(_abc_41234_new_n1439_), .Y(_abc_41234_new_n1440_));
OAI21X1 OAI21X1_177 ( .A(_abc_41234_new_n1390_), .B(_abc_41234_new_n1441_), .C(_abc_41234_new_n1389_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_4_));
OAI21X1 OAI21X1_178 ( .A(regfil_2__5_), .B(_abc_41234_new_n1049__bF_buf0), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1447_));
OAI21X1 OAI21X1_179 ( .A(_abc_41234_new_n1448_), .B(_abc_41234_new_n1449_), .C(_abc_41234_new_n1218_), .Y(_abc_41234_new_n1450_));
OAI21X1 OAI21X1_18 ( .A(_abc_41234_new_n613_), .B(_abc_41234_new_n650_), .C(_abc_41234_new_n673_), .Y(_abc_41234_new_n674_));
OAI21X1 OAI21X1_180 ( .A(_abc_41234_new_n904_), .B(_abc_41234_new_n1397_), .C(_abc_41234_new_n1219_), .Y(_abc_41234_new_n1454_));
OAI21X1 OAI21X1_181 ( .A(_abc_41234_new_n1453_), .B(_abc_41234_new_n1454_), .C(_abc_41234_new_n1043_), .Y(_abc_41234_new_n1455_));
OAI21X1 OAI21X1_182 ( .A(_abc_41234_new_n849_), .B(_abc_41234_new_n1408_), .C(_abc_41234_new_n1459_), .Y(_abc_41234_new_n1460_));
OAI21X1 OAI21X1_183 ( .A(_abc_41234_new_n1411_), .B(_abc_41234_new_n1460_), .C(_abc_41234_new_n1467_), .Y(_abc_41234_new_n1468_));
OAI21X1 OAI21X1_184 ( .A(_abc_41234_new_n1471_), .B(_abc_41234_new_n1473_), .C(_abc_41234_new_n1425_), .Y(_abc_41234_new_n1474_));
OAI21X1 OAI21X1_185 ( .A(_abc_41234_new_n1483_), .B(_abc_41234_new_n1484_), .C(_abc_41234_new_n1482_), .Y(_abc_41234_new_n1485_));
OAI21X1 OAI21X1_186 ( .A(_abc_41234_new_n1140_), .B(_abc_41234_new_n1492_), .C(_abc_41234_new_n1494_), .Y(_abc_41234_new_n1495_));
OAI21X1 OAI21X1_187 ( .A(_abc_41234_new_n1447_), .B(_abc_41234_new_n1505_), .C(_abc_41234_new_n1446_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_5_));
OAI21X1 OAI21X1_188 ( .A(regfil_2__6_), .B(_abc_41234_new_n1049__bF_buf3), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1512_));
OAI21X1 OAI21X1_189 ( .A(regfil_4__5_), .B(_abc_41234_new_n1391_), .C(regfil_4__6_), .Y(_abc_41234_new_n1514_));
OAI21X1 OAI21X1_19 ( .A(opcode_3_bF_buf1_), .B(_abc_41234_new_n615_), .C(_abc_41234_new_n674_), .Y(_abc_41234_new_n675_));
OAI21X1 OAI21X1_190 ( .A(_abc_41234_new_n1219_), .B(_abc_41234_new_n1515_), .C(_abc_41234_new_n1049__bF_buf2), .Y(_abc_41234_new_n1516_));
OAI21X1 OAI21X1_191 ( .A(regfil_4__6_), .B(_abc_41234_new_n1517_), .C(_abc_41234_new_n1518_), .Y(_abc_41234_new_n1519_));
OAI21X1 OAI21X1_192 ( .A(_abc_41234_new_n1218_), .B(_abc_41234_new_n1206_), .C(_abc_41234_new_n1519_), .Y(_abc_41234_new_n1520_));
OAI21X1 OAI21X1_193 ( .A(_abc_41234_new_n1523_), .B(_abc_41234_new_n1525_), .C(_abc_41234_new_n1522_), .Y(_abc_41234_new_n1526_));
OAI21X1 OAI21X1_194 ( .A(_abc_41234_new_n900_), .B(_abc_41234_new_n904_), .C(_abc_41234_new_n1500_), .Y(_abc_41234_new_n1532_));
OAI21X1 OAI21X1_195 ( .A(_abc_41234_new_n1425_), .B(_abc_41234_new_n1471_), .C(_abc_41234_new_n1472_), .Y(_abc_41234_new_n1542_));
OAI21X1 OAI21X1_196 ( .A(_abc_41234_new_n1550_), .B(_abc_41234_new_n1549_), .C(_abc_41234_new_n1200_), .Y(_abc_41234_new_n1551_));
OAI21X1 OAI21X1_197 ( .A(_abc_41234_new_n1551_), .B(_abc_41234_new_n1548_), .C(_abc_41234_new_n1156_), .Y(_abc_41234_new_n1552_));
OAI21X1 OAI21X1_198 ( .A(_abc_41234_new_n1541_), .B(_abc_41234_new_n1552_), .C(_abc_41234_new_n1553_), .Y(_abc_41234_new_n1554_));
OAI21X1 OAI21X1_199 ( .A(_abc_41234_new_n1512_), .B(_abc_41234_new_n1556_), .C(_abc_41234_new_n1511_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_6_));
OAI21X1 OAI21X1_2 ( .A(regfil_7__2_), .B(regfil_7__1_), .C(regfil_7__3_), .Y(_abc_41234_new_n542_));
OAI21X1 OAI21X1_20 ( .A(regfil_7__6_), .B(regfil_7__5_), .C(regfil_7__7_), .Y(_abc_41234_new_n689_));
OAI21X1 OAI21X1_200 ( .A(_abc_41234_new_n1058_), .B(_abc_41234_new_n1059_), .C(regfil_4__7_), .Y(_abc_41234_new_n1559_));
OAI21X1 OAI21X1_201 ( .A(_abc_41234_new_n1061_), .B(_abc_41234_new_n1558_), .C(_abc_41234_new_n1559_), .Y(_abc_41234_new_n1560_));
OAI21X1 OAI21X1_202 ( .A(regfil_2__7_), .B(_abc_41234_new_n1049__bF_buf1), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1562_));
OAI21X1 OAI21X1_203 ( .A(_abc_41234_new_n1563_), .B(_abc_41234_new_n1564_), .C(_abc_41234_new_n1218_), .Y(_abc_41234_new_n1565_));
OAI21X1 OAI21X1_204 ( .A(_abc_41234_new_n1528_), .B(_abc_41234_new_n1522_), .C(_abc_41234_new_n1566_), .Y(_abc_41234_new_n1567_));
OAI21X1 OAI21X1_205 ( .A(_abc_41234_new_n1550_), .B(_abc_41234_new_n1549_), .C(_abc_41234_new_n1582_), .Y(_abc_41234_new_n1583_));
OAI21X1 OAI21X1_206 ( .A(_abc_41234_new_n1532_), .B(_abc_41234_new_n1498_), .C(_abc_41234_new_n1537_), .Y(_abc_41234_new_n1588_));
OAI21X1 OAI21X1_207 ( .A(_abc_41234_new_n1538_), .B(_abc_41234_new_n1533_), .C(_abc_41234_new_n1587_), .Y(_abc_41234_new_n1594_));
OAI21X1 OAI21X1_208 ( .A(_abc_41234_new_n1591_), .B(_abc_41234_new_n1594_), .C(_abc_41234_new_n1151_), .Y(_abc_41234_new_n1595_));
OAI21X1 OAI21X1_209 ( .A(_abc_41234_new_n1593_), .B(_abc_41234_new_n1595_), .C(_abc_41234_new_n1586_), .Y(_abc_41234_new_n1596_));
OAI21X1 OAI21X1_21 ( .A(carry), .B(_abc_41234_new_n690_), .C(_abc_41234_new_n701_), .Y(_abc_41234_new_n702_));
OAI21X1 OAI21X1_210 ( .A(_abc_41234_new_n1562_), .B(_abc_41234_new_n1603_), .C(_abc_41234_new_n1561_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_7_));
OAI21X1 OAI21X1_211 ( .A(_abc_41234_new_n544__bF_buf3), .B(_abc_41234_new_n1610_), .C(wdatahold2_0_), .Y(_abc_41234_new_n1611_));
OAI21X1 OAI21X1_212 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n1611_), .Y(_abc_41234_new_n1612_));
OAI21X1 OAI21X1_213 ( .A(pc_1_), .B(pc_0_), .C(_abc_41234_new_n1615_), .Y(_abc_41234_new_n1616_));
OAI21X1 OAI21X1_214 ( .A(_abc_41234_new_n1619_), .B(_abc_41234_new_n1616_), .C(_abc_41234_new_n1622_), .Y(_abc_41234_new_n1623_));
OAI21X1 OAI21X1_215 ( .A(_abc_41234_new_n1625_), .B(_abc_41234_new_n547_), .C(_abc_41234_new_n618_), .Y(_abc_41234_new_n1626_));
OAI21X1 OAI21X1_216 ( .A(_abc_41234_new_n1627_), .B(_abc_41234_new_n1632_), .C(_abc_41234_new_n1624_), .Y(_abc_41234_new_n1633_));
OAI21X1 OAI21X1_217 ( .A(_abc_41234_new_n528_), .B(_abc_41234_new_n1634_), .C(_abc_41234_new_n544__bF_buf2), .Y(_abc_41234_new_n1635_));
OAI21X1 OAI21X1_218 ( .A(_abc_41234_new_n536__bF_buf2), .B(_abc_41234_new_n548_), .C(_abc_41234_new_n1635_), .Y(_abc_41234_new_n1636_));
OAI21X1 OAI21X1_219 ( .A(_abc_41234_new_n1322_), .B(_abc_41234_new_n1629_), .C(_abc_41234_new_n1640_), .Y(_abc_41234_new_n1641_));
OAI21X1 OAI21X1_22 ( .A(_abc_41234_new_n646_), .B(_abc_41234_new_n679_), .C(_abc_41234_new_n712_), .Y(_abc_41234_new_n713_));
OAI21X1 OAI21X1_220 ( .A(_abc_41234_new_n1619_), .B(_abc_41234_new_n1649_), .C(_abc_41234_new_n1622_), .Y(_abc_41234_new_n1650_));
OAI21X1 OAI21X1_221 ( .A(opcode_4_bF_buf3_), .B(regfil_0__0_), .C(_abc_41234_new_n1655_), .Y(_abc_41234_new_n1656_));
OAI21X1 OAI21X1_222 ( .A(_abc_41234_new_n1657_), .B(_abc_41234_new_n1654_), .C(_abc_41234_new_n1639__bF_buf2), .Y(_abc_41234_new_n1658_));
OAI21X1 OAI21X1_223 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1040__bF_buf2), .C(_abc_41234_new_n1658_), .Y(_abc_41234_new_n1659_));
OAI21X1 OAI21X1_224 ( .A(_abc_41234_new_n1653_), .B(_abc_41234_new_n1645_), .C(_abc_41234_new_n1660_), .Y(_abc_41234_new_n1661_));
OAI21X1 OAI21X1_225 ( .A(_abc_41234_new_n544__bF_buf0), .B(_abc_41234_new_n1610_), .C(wdatahold2_1_), .Y(_abc_41234_new_n1667_));
OAI21X1 OAI21X1_226 ( .A(_abc_41234_new_n720_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n1667_), .Y(_abc_41234_new_n1668_));
OAI21X1 OAI21X1_227 ( .A(_abc_41234_new_n1622_), .B(_abc_41234_new_n1671_), .C(_abc_41234_new_n1670_), .Y(_abc_41234_new_n1672_));
OAI21X1 OAI21X1_228 ( .A(_abc_41234_new_n1627_), .B(_abc_41234_new_n1675_), .C(_abc_41234_new_n1674_), .Y(_abc_41234_new_n1676_));
OAI21X1 OAI21X1_229 ( .A(_abc_41234_new_n1622_), .B(_abc_41234_new_n1677_), .C(_abc_41234_new_n1670_), .Y(_abc_41234_new_n1678_));
OAI21X1 OAI21X1_23 ( .A(_abc_41234_new_n570_), .B(_abc_41234_new_n722__bF_buf2), .C(_abc_41234_new_n728_), .Y(_abc_41234_new_n729_));
OAI21X1 OAI21X1_230 ( .A(_abc_41234_new_n539_), .B(_abc_41234_new_n1636_), .C(_abc_41234_new_n1680_), .Y(_abc_41234_new_n1681_));
OAI21X1 OAI21X1_231 ( .A(opcode_4_bF_buf1_), .B(regfil_0__1_), .C(_abc_41234_new_n1685_), .Y(_abc_41234_new_n1686_));
OAI21X1 OAI21X1_232 ( .A(_abc_41234_new_n1640_), .B(_abc_41234_new_n1688_), .C(_abc_41234_new_n1689_), .Y(_abc_41234_new_n1690_));
OAI21X1 OAI21X1_233 ( .A(_abc_41234_new_n544__bF_buf2), .B(_abc_41234_new_n1610_), .C(wdatahold2_2_), .Y(_abc_41234_new_n1698_));
OAI21X1 OAI21X1_234 ( .A(_abc_41234_new_n773_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n1698_), .Y(_abc_41234_new_n1699_));
OAI21X1 OAI21X1_235 ( .A(opcode_4_bF_buf6_), .B(regfil_0__2_), .C(_abc_41234_new_n1700_), .Y(_abc_41234_new_n1701_));
OAI21X1 OAI21X1_236 ( .A(_abc_41234_new_n751_), .B(_abc_41234_new_n1105__bF_buf0), .C(_abc_41234_new_n1368_), .Y(_abc_41234_new_n1703_));
OAI21X1 OAI21X1_237 ( .A(_abc_41234_new_n1702_), .B(_abc_41234_new_n1703_), .C(_abc_41234_new_n1639__bF_buf1), .Y(_abc_41234_new_n1704_));
OAI21X1 OAI21X1_238 ( .A(_abc_41234_new_n1670_), .B(_abc_41234_new_n1621_), .C(_abc_41234_new_n1705_), .Y(_abc_41234_new_n1708_));
OAI21X1 OAI21X1_239 ( .A(intcyc_bF_buf2), .B(_abc_41234_new_n1710_), .C(_abc_41234_new_n1711_), .Y(_abc_41234_new_n1712_));
OAI21X1 OAI21X1_24 ( .A(_abc_41234_new_n732_), .B(_abc_41234_new_n729_), .C(_abc_41234_new_n546__bF_buf0), .Y(_abc_41234_new_n733_));
OAI21X1 OAI21X1_240 ( .A(_abc_41234_new_n773_), .B(_abc_41234_new_n1040__bF_buf1), .C(_abc_41234_new_n1712_), .Y(_abc_41234_new_n1713_));
OAI21X1 OAI21X1_241 ( .A(_abc_41234_new_n1670_), .B(_abc_41234_new_n1652_), .C(_abc_41234_new_n1705_), .Y(_abc_41234_new_n1714_));
OAI21X1 OAI21X1_242 ( .A(_abc_41234_new_n539_), .B(_abc_41234_new_n1636_), .C(_abc_41234_new_n1716_), .Y(_abc_41234_new_n1717_));
OAI21X1 OAI21X1_243 ( .A(_abc_41234_new_n1626_), .B(_abc_41234_new_n1709_), .C(_abc_41234_new_n1717_), .Y(_abc_41234_new_n1718_));
OAI21X1 OAI21X1_244 ( .A(_abc_41234_new_n544__bF_buf1), .B(_abc_41234_new_n1610_), .C(wdatahold2_3_), .Y(_abc_41234_new_n1725_));
OAI21X1 OAI21X1_245 ( .A(_abc_41234_new_n819_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n1725_), .Y(_abc_41234_new_n1726_));
OAI21X1 OAI21X1_246 ( .A(_abc_41234_new_n1729_), .B(pc_11_), .C(_abc_41234_new_n1630_), .Y(_abc_41234_new_n1730_));
OAI21X1 OAI21X1_247 ( .A(_abc_41234_new_n1627_), .B(_abc_41234_new_n1731_), .C(_abc_41234_new_n1728_), .Y(_abc_41234_new_n1732_));
OAI21X1 OAI21X1_248 ( .A(_abc_41234_new_n1639__bF_buf0), .B(_abc_41234_new_n581_), .C(_abc_41234_new_n537__bF_buf1), .Y(_abc_41234_new_n1735_));
OAI21X1 OAI21X1_249 ( .A(opcode_4_bF_buf4_), .B(regfil_0__3_), .C(_abc_41234_new_n1736_), .Y(_abc_41234_new_n1737_));
OAI21X1 OAI21X1_25 ( .A(_abc_41234_new_n546__bF_buf5), .B(_abc_41234_new_n727_), .C(_abc_41234_new_n733_), .Y(_abc_41234_new_n734_));
OAI21X1 OAI21X1_250 ( .A(_abc_41234_new_n819_), .B(_abc_41234_new_n1735_), .C(_abc_41234_new_n1739_), .Y(_abc_41234_new_n1740_));
OAI21X1 OAI21X1_251 ( .A(_abc_41234_new_n544__bF_buf0), .B(_abc_41234_new_n1610_), .C(wdatahold2_4_), .Y(_abc_41234_new_n1747_));
OAI21X1 OAI21X1_252 ( .A(_abc_41234_new_n849_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n1747_), .Y(_abc_41234_new_n1748_));
OAI21X1 OAI21X1_253 ( .A(_abc_41234_new_n1727_), .B(_abc_41234_new_n1707_), .C(_abc_41234_new_n1750_), .Y(_abc_41234_new_n1751_));
OAI21X1 OAI21X1_254 ( .A(_abc_41234_new_n1727_), .B(_abc_41234_new_n1715_), .C(_abc_41234_new_n1750_), .Y(_abc_41234_new_n1753_));
OAI21X1 OAI21X1_255 ( .A(intcyc_bF_buf2), .B(_abc_41234_new_n1752_), .C(_abc_41234_new_n1758_), .Y(_abc_41234_new_n1759_));
OAI21X1 OAI21X1_256 ( .A(opcode_4_bF_buf2_), .B(regfil_0__4_), .C(_abc_41234_new_n1760_), .Y(_abc_41234_new_n1761_));
OAI21X1 OAI21X1_257 ( .A(_abc_41234_new_n851_), .B(_abc_41234_new_n1105__bF_buf2), .C(_abc_41234_new_n1469_), .Y(_abc_41234_new_n1763_));
OAI21X1 OAI21X1_258 ( .A(_abc_41234_new_n1762_), .B(_abc_41234_new_n1763_), .C(_abc_41234_new_n1639__bF_buf2), .Y(_abc_41234_new_n1764_));
OAI21X1 OAI21X1_259 ( .A(_abc_41234_new_n849_), .B(_abc_41234_new_n1040__bF_buf0), .C(_abc_41234_new_n1764_), .Y(_abc_41234_new_n1765_));
OAI21X1 OAI21X1_26 ( .A(_abc_41234_new_n615_), .B(_abc_41234_new_n735_), .C(_abc_41234_new_n736_), .Y(_abc_41234_new_n737_));
OAI21X1 OAI21X1_260 ( .A(_abc_41234_new_n544__bF_buf3), .B(_abc_41234_new_n1610_), .C(wdatahold2_5_), .Y(_abc_41234_new_n1772_));
OAI21X1 OAI21X1_261 ( .A(_abc_41234_new_n904_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n1772_), .Y(_abc_41234_new_n1773_));
OAI21X1 OAI21X1_262 ( .A(_abc_41234_new_n1627_), .B(_abc_41234_new_n1776_), .C(_abc_41234_new_n1774_), .Y(_abc_41234_new_n1777_));
OAI21X1 OAI21X1_263 ( .A(opcode_4_bF_buf0_), .B(regfil_0__5_), .C(_abc_41234_new_n1782_), .Y(_abc_41234_new_n1783_));
OAI21X1 OAI21X1_264 ( .A(_abc_41234_new_n904_), .B(_abc_41234_new_n1735_), .C(_abc_41234_new_n1786_), .Y(_abc_41234_new_n1787_));
OAI21X1 OAI21X1_265 ( .A(_abc_41234_new_n544__bF_buf2), .B(_abc_41234_new_n1610_), .C(wdatahold2_6_), .Y(_abc_41234_new_n1794_));
OAI21X1 OAI21X1_266 ( .A(_abc_41234_new_n1509_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n1794_), .Y(_abc_41234_new_n1795_));
OAI21X1 OAI21X1_267 ( .A(_abc_41234_new_n1775_), .B(_abc_41234_new_n1749_), .C(_abc_41234_new_n1798_), .Y(_abc_41234_new_n1799_));
OAI21X1 OAI21X1_268 ( .A(_abc_41234_new_n1775_), .B(_abc_41234_new_n1754_), .C(_abc_41234_new_n1798_), .Y(_abc_41234_new_n1801_));
OAI21X1 OAI21X1_269 ( .A(intcyc_bF_buf2), .B(_abc_41234_new_n1800_), .C(_abc_41234_new_n1807_), .Y(_abc_41234_new_n1808_));
OAI21X1 OAI21X1_27 ( .A(_abc_41234_new_n738_), .B(_abc_41234_new_n741_), .C(_abc_41234_new_n600_), .Y(_abc_41234_new_n742_));
OAI21X1 OAI21X1_270 ( .A(opcode_4_bF_buf5_), .B(regfil_0__6_), .C(_abc_41234_new_n1811_), .Y(_abc_41234_new_n1812_));
OAI21X1 OAI21X1_271 ( .A(_abc_41234_new_n1810_), .B(_abc_41234_new_n1813_), .C(_abc_41234_new_n1639__bF_buf0), .Y(_abc_41234_new_n1814_));
OAI21X1 OAI21X1_272 ( .A(_abc_41234_new_n1509_), .B(_abc_41234_new_n1040__bF_buf4), .C(_abc_41234_new_n1814_), .Y(_abc_41234_new_n1815_));
OAI21X1 OAI21X1_273 ( .A(_abc_41234_new_n544__bF_buf0), .B(_abc_41234_new_n1610_), .C(wdatahold2_7_), .Y(_abc_41234_new_n1822_));
OAI21X1 OAI21X1_274 ( .A(_abc_41234_new_n997_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n1822_), .Y(_abc_41234_new_n1823_));
OAI21X1 OAI21X1_275 ( .A(_abc_41234_new_n1798_), .B(_abc_41234_new_n1824_), .C(pc_15_), .Y(_abc_41234_new_n1825_));
OAI21X1 OAI21X1_276 ( .A(_abc_41234_new_n1627_), .B(_abc_41234_new_n1829_), .C(_abc_41234_new_n1827_), .Y(_abc_41234_new_n1830_));
OAI21X1 OAI21X1_277 ( .A(_abc_41234_new_n1798_), .B(_abc_41234_new_n1779_), .C(pc_15_), .Y(_abc_41234_new_n1831_));
OAI21X1 OAI21X1_278 ( .A(opcode_4_bF_buf3_), .B(regfil_0__7_), .C(_abc_41234_new_n1835_), .Y(_abc_41234_new_n1836_));
OAI21X1 OAI21X1_279 ( .A(_abc_41234_new_n997_), .B(_abc_41234_new_n1735_), .C(_abc_41234_new_n1839_), .Y(_abc_41234_new_n1840_));
OAI21X1 OAI21X1_28 ( .A(_abc_41234_new_n718_), .B(_abc_41234_new_n632_), .C(_abc_41234_new_n747_), .Y(_abc_41234_new_n748_));
OAI21X1 OAI21X1_280 ( .A(_abc_41234_new_n518_), .B(_abc_41234_new_n1850_), .C(_abc_41234_new_n1854_), .Y(_abc_41234_new_n1855_));
OAI21X1 OAI21X1_281 ( .A(_abc_41234_new_n598_), .B(_abc_41234_new_n581_), .C(_abc_41234_new_n530_), .Y(_abc_41234_new_n1856_));
OAI21X1 OAI21X1_282 ( .A(_abc_41234_new_n646_), .B(_abc_41234_new_n1847_), .C(_abc_41234_new_n1860_), .Y(_abc_41234_new_n1861_));
OAI21X1 OAI21X1_283 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold2_0_), .Y(_abc_41234_new_n1863_));
OAI21X1 OAI21X1_284 ( .A(regfil_3__0_), .B(_abc_41234_new_n1864_), .C(_abc_41234_new_n1049__bF_buf4), .Y(_abc_41234_new_n1865_));
OAI21X1 OAI21X1_285 ( .A(regfil_5__0_), .B(_abc_41234_new_n1049__bF_buf3), .C(_abc_41234_new_n1865_), .Y(_abc_41234_new_n1866_));
OAI21X1 OAI21X1_286 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n748_), .C(_abc_41234_new_n1868_), .Y(_abc_41234_new_n1869_));
OAI21X1 OAI21X1_287 ( .A(_abc_41234_new_n1872_), .B(_abc_41234_new_n1874_), .C(_abc_41234_new_n1876_), .Y(_abc_41234_new_n1877_));
OAI21X1 OAI21X1_288 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n791_), .C(_abc_41234_new_n1884_), .Y(_abc_41234_new_n1885_));
OAI21X1 OAI21X1_289 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold2_2_), .Y(_abc_41234_new_n1886_));
OAI21X1 OAI21X1_29 ( .A(regfil_7__1_), .B(_abc_41234_new_n678_), .C(_abc_41234_new_n710_), .Y(_abc_41234_new_n750_));
OAI21X1 OAI21X1_290 ( .A(regfil_3__0_), .B(regfil_3__1_), .C(regfil_3__2_), .Y(_abc_41234_new_n1889_));
OAI21X1 OAI21X1_291 ( .A(_abc_41234_new_n1848_), .B(_abc_41234_new_n730_), .C(_abc_41234_new_n768_), .Y(_abc_41234_new_n1891_));
OAI21X1 OAI21X1_292 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n829_), .C(_abc_41234_new_n1897_), .Y(_abc_41234_new_n1898_));
OAI21X1 OAI21X1_293 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold2_3_), .Y(_abc_41234_new_n1899_));
OAI21X1 OAI21X1_294 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n879_), .C(_abc_41234_new_n1908_), .Y(_abc_41234_new_n1909_));
OAI21X1 OAI21X1_295 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold2_4_), .Y(_abc_41234_new_n1910_));
OAI21X1 OAI21X1_296 ( .A(_abc_41234_new_n1913_), .B(_abc_41234_new_n1914_), .C(_abc_41234_new_n1873_), .Y(_abc_41234_new_n1915_));
OAI21X1 OAI21X1_297 ( .A(_abc_41234_new_n814_), .B(_abc_41234_new_n1892_), .C(_abc_41234_new_n858_), .Y(_abc_41234_new_n1916_));
OAI21X1 OAI21X1_298 ( .A(_abc_41234_new_n1918_), .B(_abc_41234_new_n1887_), .C(_abc_41234_new_n1915_), .Y(_abc_41234_new_n1919_));
OAI21X1 OAI21X1_299 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n924_), .C(_abc_41234_new_n1922_), .Y(_abc_41234_new_n1923_));
OAI21X1 OAI21X1_3 ( .A(auxcar), .B(_abc_41234_new_n543_), .C(_abc_41234_new_n551_), .Y(_abc_41234_new_n552_));
OAI21X1 OAI21X1_30 ( .A(_abc_41234_new_n525__bF_buf1), .B(_abc_41234_new_n538_), .C(_abc_41234_new_n552_), .Y(_abc_41234_new_n752_));
OAI21X1 OAI21X1_300 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold2_5_), .Y(_abc_41234_new_n1924_));
OAI21X1 OAI21X1_301 ( .A(_abc_41234_new_n1926_), .B(_abc_41234_new_n1927_), .C(_abc_41234_new_n1873_), .Y(_abc_41234_new_n1928_));
OAI21X1 OAI21X1_302 ( .A(_abc_41234_new_n858_), .B(_abc_41234_new_n1903_), .C(_abc_41234_new_n899_), .Y(_abc_41234_new_n1931_));
OAI21X1 OAI21X1_303 ( .A(_abc_41234_new_n1932_), .B(_abc_41234_new_n1887_), .C(_abc_41234_new_n1928_), .Y(_abc_41234_new_n1933_));
OAI21X1 OAI21X1_304 ( .A(_abc_41234_new_n1847_), .B(_abc_41234_new_n963_), .C(_abc_41234_new_n1937_), .Y(_abc_41234_new_n1938_));
OAI21X1 OAI21X1_305 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold2_6_), .Y(_abc_41234_new_n1939_));
OAI21X1 OAI21X1_306 ( .A(_abc_41234_new_n1940_), .B(_abc_41234_new_n1941_), .C(_abc_41234_new_n1873_), .Y(_abc_41234_new_n1942_));
OAI21X1 OAI21X1_307 ( .A(regfil_3__6_), .B(_abc_41234_new_n1929_), .C(_abc_41234_new_n1875_), .Y(_abc_41234_new_n1945_));
OAI21X1 OAI21X1_308 ( .A(_abc_41234_new_n1944_), .B(_abc_41234_new_n1945_), .C(_abc_41234_new_n1942_), .Y(_abc_41234_new_n1946_));
OAI21X1 OAI21X1_309 ( .A(_abc_41234_new_n1010_), .B(_abc_41234_new_n1847_), .C(_abc_41234_new_n1949_), .Y(_abc_41234_new_n1950_));
OAI21X1 OAI21X1_31 ( .A(_abc_41234_new_n751_), .B(_abc_41234_new_n688_), .C(_abc_41234_new_n753_), .Y(_abc_41234_new_n754_));
OAI21X1 OAI21X1_310 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold2_7_), .Y(_abc_41234_new_n1951_));
OAI21X1 OAI21X1_311 ( .A(regfil_3__6_), .B(_abc_41234_new_n1925_), .C(regfil_3__7_), .Y(_abc_41234_new_n1957_));
OAI21X1 OAI21X1_312 ( .A(_abc_41234_new_n1958_), .B(_abc_41234_new_n1956_), .C(_abc_41234_new_n1955_), .Y(_abc_41234_new_n1959_));
OAI21X1 OAI21X1_313 ( .A(regfil_3__7_), .B(_abc_41234_new_n1944_), .C(_abc_41234_new_n1961_), .Y(_abc_41234_new_n1962_));
OAI21X1 OAI21X1_314 ( .A(_abc_41234_new_n1953_), .B(_abc_41234_new_n1962_), .C(_abc_41234_new_n1959_), .Y(_abc_41234_new_n1963_));
OAI21X1 OAI21X1_315 ( .A(_abc_41234_new_n1066__bF_buf0), .B(_abc_41234_new_n1963_), .C(_abc_41234_new_n1952_), .Y(_abc_41234_new_n1964_));
OAI21X1 OAI21X1_316 ( .A(_abc_41234_new_n652_), .B(_abc_41234_new_n648_), .C(_abc_41234_new_n1057_), .Y(_abc_41234_new_n1966_));
OAI21X1 OAI21X1_317 ( .A(_abc_41234_new_n646_), .B(_abc_41234_new_n1967_), .C(_abc_41234_new_n1968_), .Y(_abc_41234_new_n1969_));
OAI21X1 OAI21X1_318 ( .A(_abc_41234_new_n1967_), .B(_abc_41234_new_n748_), .C(_abc_41234_new_n1973_), .Y(_abc_41234_new_n1974_));
OAI21X1 OAI21X1_319 ( .A(_abc_41234_new_n583_), .B(_abc_41234_new_n1977_), .C(_abc_41234_new_n1978_), .Y(_abc_41234_new_n1979_));
OAI21X1 OAI21X1_32 ( .A(_abc_41234_new_n718_), .B(_abc_41234_new_n512_), .C(_abc_41234_new_n759_), .Y(_abc_41234_new_n760_));
OAI21X1 OAI21X1_320 ( .A(_abc_41234_new_n1967_), .B(_abc_41234_new_n791_), .C(_abc_41234_new_n1982_), .Y(_abc_41234_new_n1983_));
OAI21X1 OAI21X1_321 ( .A(regfil_1__0_), .B(regfil_1__1_), .C(regfil_1__2_), .Y(_abc_41234_new_n1984_));
OAI21X1 OAI21X1_322 ( .A(_abc_41234_new_n569_), .B(_abc_41234_new_n570_), .C(_abc_41234_new_n634_), .Y(_abc_41234_new_n1986_));
OAI21X1 OAI21X1_323 ( .A(_abc_41234_new_n1967_), .B(_abc_41234_new_n829_), .C(_abc_41234_new_n1991_), .Y(_abc_41234_new_n1992_));
OAI21X1 OAI21X1_324 ( .A(regfil_1__2_), .B(_abc_41234_new_n1976_), .C(regfil_1__3_), .Y(_abc_41234_new_n1993_));
OAI21X1 OAI21X1_325 ( .A(_abc_41234_new_n634_), .B(_abc_41234_new_n1975_), .C(_abc_41234_new_n568_), .Y(_abc_41234_new_n1996_));
OAI21X1 OAI21X1_326 ( .A(_abc_41234_new_n648_), .B(_abc_41234_new_n2001_), .C(_abc_41234_new_n2006_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_4_));
OAI21X1 OAI21X1_327 ( .A(regfil_1__4_), .B(_abc_41234_new_n636_), .C(regfil_1__5_), .Y(_abc_41234_new_n2010_));
OAI21X1 OAI21X1_328 ( .A(_abc_41234_new_n855_), .B(_abc_41234_new_n1995_), .C(_abc_41234_new_n896_), .Y(_abc_41234_new_n2012_));
OAI21X1 OAI21X1_329 ( .A(_abc_41234_new_n1995_), .B(_abc_41234_new_n574_), .C(_abc_41234_new_n2012_), .Y(_abc_41234_new_n2013_));
OAI21X1 OAI21X1_33 ( .A(_abc_41234_new_n514_), .B(_abc_41234_new_n702_), .C(_abc_41234_new_n761_), .Y(_abc_41234_new_n762_));
OAI21X1 OAI21X1_330 ( .A(_abc_41234_new_n648_), .B(_abc_41234_new_n2008_), .C(_abc_41234_new_n2015_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_5_));
OAI21X1 OAI21X1_331 ( .A(_abc_41234_new_n638_), .B(_abc_41234_new_n2021_), .C(_abc_41234_new_n583_), .Y(_abc_41234_new_n2022_));
OAI21X1 OAI21X1_332 ( .A(_abc_41234_new_n648_), .B(_abc_41234_new_n2017_), .C(_abc_41234_new_n2024_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_6_));
OAI21X1 OAI21X1_333 ( .A(regfil_1__6_), .B(_abc_41234_new_n2009_), .C(regfil_1__7_), .Y(_abc_41234_new_n2027_));
OAI21X1 OAI21X1_334 ( .A(_abc_41234_new_n641_), .B(_abc_41234_new_n2028_), .C(_abc_41234_new_n631_), .Y(_abc_41234_new_n2029_));
OAI21X1 OAI21X1_335 ( .A(_abc_41234_new_n2030_), .B(_abc_41234_new_n2031_), .C(_abc_41234_new_n2029_), .Y(_abc_41234_new_n2032_));
OAI21X1 OAI21X1_336 ( .A(_abc_41234_new_n648_), .B(_abc_41234_new_n2026_), .C(_abc_41234_new_n2033_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_7_));
OAI21X1 OAI21X1_337 ( .A(_abc_41234_new_n725_), .B(_abc_41234_new_n2035_), .C(_abc_41234_new_n2038_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_1_));
OAI21X1 OAI21X1_338 ( .A(_abc_41234_new_n775_), .B(_abc_41234_new_n2035_), .C(_abc_41234_new_n2040_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_2_));
OAI21X1 OAI21X1_339 ( .A(_abc_41234_new_n822_), .B(_abc_41234_new_n2035_), .C(_abc_41234_new_n2042_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_3_));
OAI21X1 OAI21X1_34 ( .A(_abc_41234_new_n750_), .B(_abc_41234_new_n749_), .C(_abc_41234_new_n763_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_1_));
OAI21X1 OAI21X1_340 ( .A(_abc_41234_new_n852_), .B(_abc_41234_new_n2035_), .C(_abc_41234_new_n2044_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_4_));
OAI21X1 OAI21X1_341 ( .A(_abc_41234_new_n907_), .B(_abc_41234_new_n2035_), .C(_abc_41234_new_n2046_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_5_));
OAI21X1 OAI21X1_342 ( .A(_abc_41234_new_n2048_), .B(_abc_41234_new_n2035_), .C(_abc_41234_new_n2049_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_6_));
OAI21X1 OAI21X1_343 ( .A(_abc_41234_new_n999_), .B(_abc_41234_new_n2035_), .C(_abc_41234_new_n2051_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_7_));
OAI21X1 OAI21X1_344 ( .A(_abc_41234_new_n646_), .B(_abc_41234_new_n2053_), .C(_abc_41234_new_n2054_), .Y(_abc_41234_new_n2055_));
OAI21X1 OAI21X1_345 ( .A(_abc_41234_new_n2057_), .B(_abc_41234_new_n2058_), .C(_abc_41234_new_n1873_), .Y(_abc_41234_new_n2059_));
OAI21X1 OAI21X1_346 ( .A(regfil_2__0_), .B(_abc_41234_new_n1953_), .C(_abc_41234_new_n2062_), .Y(_abc_41234_new_n2063_));
OAI21X1 OAI21X1_347 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1049__bF_buf2), .C(_abc_41234_new_n2064_), .Y(_abc_41234_new_n2065_));
OAI21X1 OAI21X1_348 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n748_), .C(_abc_41234_new_n2068_), .Y(_abc_41234_new_n2069_));
OAI21X1 OAI21X1_349 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold_1_), .Y(_abc_41234_new_n2070_));
OAI21X1 OAI21X1_35 ( .A(_abc_41234_new_n770_), .B(_abc_41234_new_n767_), .C(_abc_41234_new_n546__bF_buf4), .Y(_abc_41234_new_n771_));
OAI21X1 OAI21X1_350 ( .A(regfil_2__0_), .B(_abc_41234_new_n2056_), .C(regfil_2__1_), .Y(_abc_41234_new_n2073_));
OAI21X1 OAI21X1_351 ( .A(_abc_41234_new_n731_), .B(_abc_41234_new_n2060_), .C(_abc_41234_new_n1875_), .Y(_abc_41234_new_n2076_));
OAI21X1 OAI21X1_352 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n791_), .C(_abc_41234_new_n2080_), .Y(_abc_41234_new_n2081_));
OAI21X1 OAI21X1_353 ( .A(_abc_41234_new_n2083_), .B(_abc_41234_new_n2082_), .C(_abc_41234_new_n1873_), .Y(_abc_41234_new_n2084_));
OAI21X1 OAI21X1_354 ( .A(_abc_41234_new_n731_), .B(_abc_41234_new_n2060_), .C(_abc_41234_new_n769_), .Y(_abc_41234_new_n2085_));
OAI21X1 OAI21X1_355 ( .A(_abc_41234_new_n773_), .B(_abc_41234_new_n1049__bF_buf1), .C(_abc_41234_new_n2088_), .Y(_abc_41234_new_n2089_));
OAI21X1 OAI21X1_356 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n829_), .C(_abc_41234_new_n2092_), .Y(_abc_41234_new_n2093_));
OAI21X1 OAI21X1_357 ( .A(regfil_2__3_), .B(_abc_41234_new_n2095_), .C(_abc_41234_new_n1875_), .Y(_abc_41234_new_n2096_));
OAI21X1 OAI21X1_358 ( .A(_abc_41234_new_n2098_), .B(_abc_41234_new_n2099_), .C(_abc_41234_new_n1873_), .Y(_abc_41234_new_n2100_));
OAI21X1 OAI21X1_359 ( .A(_abc_41234_new_n2094_), .B(_abc_41234_new_n2096_), .C(_abc_41234_new_n2101_), .Y(_abc_41234_new_n2102_));
OAI21X1 OAI21X1_36 ( .A(_abc_41234_new_n776_), .B(_abc_41234_new_n774_), .C(opcode_2_), .Y(_abc_41234_new_n777_));
OAI21X1 OAI21X1_360 ( .A(regfil_2__4_), .B(_abc_41234_new_n2094_), .C(_abc_41234_new_n1875_), .Y(_abc_41234_new_n2109_));
OAI21X1 OAI21X1_361 ( .A(_abc_41234_new_n2097_), .B(_abc_41234_new_n2056_), .C(regfil_2__4_), .Y(_abc_41234_new_n2111_));
OAI21X1 OAI21X1_362 ( .A(_abc_41234_new_n2108_), .B(_abc_41234_new_n2109_), .C(_abc_41234_new_n2113_), .Y(_abc_41234_new_n2114_));
OAI21X1 OAI21X1_363 ( .A(_abc_41234_new_n1859_), .B(_abc_41234_new_n2106_), .C(_abc_41234_new_n2116_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_4_));
OAI21X1 OAI21X1_364 ( .A(regfil_2__5_), .B(_abc_41234_new_n2108_), .C(_abc_41234_new_n1875_), .Y(_abc_41234_new_n2120_));
OAI21X1 OAI21X1_365 ( .A(_abc_41234_new_n2119_), .B(_abc_41234_new_n2120_), .C(_abc_41234_new_n2125_), .Y(_abc_41234_new_n2126_));
OAI21X1 OAI21X1_366 ( .A(_abc_41234_new_n1859_), .B(_abc_41234_new_n2118_), .C(_abc_41234_new_n2128_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_5_));
OAI21X1 OAI21X1_367 ( .A(_abc_41234_new_n2053_), .B(_abc_41234_new_n963_), .C(_abc_41234_new_n2130_), .Y(_abc_41234_new_n2131_));
OAI21X1 OAI21X1_368 ( .A(_abc_41234_new_n2147_), .B(_abc_41234_new_n2146_), .C(regfil_2__6_), .Y(_abc_41234_new_n2148_));
OAI21X1 OAI21X1_369 ( .A(_abc_41234_new_n2151_), .B(_abc_41234_new_n2150_), .C(_abc_41234_new_n2137_), .Y(_abc_41234_new_n2152_));
OAI21X1 OAI21X1_37 ( .A(_abc_41234_new_n782_), .B(_abc_41234_new_n784_), .C(_abc_41234_new_n600_), .Y(_abc_41234_new_n785_));
OAI21X1 OAI21X1_370 ( .A(_abc_41234_new_n2137_), .B(_abc_41234_new_n2149_), .C(_abc_41234_new_n2152_), .Y(_abc_41234_new_n2153_));
OAI21X1 OAI21X1_371 ( .A(_abc_41234_new_n2133_), .B(_abc_41234_new_n2154_), .C(_abc_41234_new_n2155_), .Y(_abc_41234_new_n2156_));
OAI21X1 OAI21X1_372 ( .A(_abc_41234_new_n1010_), .B(_abc_41234_new_n2053_), .C(_abc_41234_new_n2159_), .Y(_abc_41234_new_n2160_));
OAI21X1 OAI21X1_373 ( .A(_abc_41234_new_n1862_), .B(_abc_41234_new_n1853_), .C(rdatahold_7_), .Y(_abc_41234_new_n2161_));
OAI21X1 OAI21X1_374 ( .A(regfil_2__7_), .B(_abc_41234_new_n2163_), .C(_abc_41234_new_n1955_), .Y(_abc_41234_new_n2165_));
OAI21X1 OAI21X1_375 ( .A(_abc_41234_new_n1535_), .B(_abc_41234_new_n2166_), .C(_abc_41234_new_n993_), .Y(_abc_41234_new_n2169_));
OAI21X1 OAI21X1_376 ( .A(_abc_41234_new_n2164_), .B(_abc_41234_new_n2165_), .C(_abc_41234_new_n2170_), .Y(_abc_41234_new_n2171_));
OAI21X1 OAI21X1_377 ( .A(_abc_41234_new_n1066__bF_buf0), .B(_abc_41234_new_n2171_), .C(_abc_41234_new_n2162_), .Y(_abc_41234_new_n2172_));
OAI21X1 OAI21X1_378 ( .A(_abc_41234_new_n661_), .B(opcode_7_), .C(_abc_41234_new_n524_), .Y(_abc_41234_new_n2175_));
OAI21X1 OAI21X1_379 ( .A(_abc_41234_new_n534__bF_buf3), .B(_abc_41234_new_n2174_), .C(_abc_41234_new_n2176_), .Y(_abc_41234_new_n2177_));
OAI21X1 OAI21X1_38 ( .A(regfil_7__2_), .B(_abc_41234_new_n678_), .C(_abc_41234_new_n710_), .Y(_abc_41234_new_n793_));
OAI21X1 OAI21X1_380 ( .A(_abc_41234_new_n546__bF_buf2), .B(_abc_41234_new_n620__bF_buf2), .C(_abc_41234_new_n1046__bF_buf3), .Y(_abc_41234_new_n2178_));
OAI21X1 OAI21X1_381 ( .A(_abc_41234_new_n2179_), .B(_abc_41234_new_n2177_), .C(alu_sel_0_), .Y(_abc_41234_new_n2180_));
OAI21X1 OAI21X1_382 ( .A(_abc_41234_new_n661_), .B(_abc_41234_new_n665__bF_buf2), .C(opcode_7_), .Y(_abc_41234_new_n2181_));
OAI21X1 OAI21X1_383 ( .A(_abc_41234_new_n2181_), .B(_abc_41234_new_n2182_), .C(_abc_41234_new_n2180_), .Y(_0alusel_2_0__0_));
OAI21X1 OAI21X1_384 ( .A(alu_sel_1_), .B(_abc_41234_new_n665__bF_buf0), .C(_abc_41234_new_n1046__bF_buf2), .Y(_abc_41234_new_n2187_));
OAI21X1 OAI21X1_385 ( .A(alu_sel_1_), .B(_abc_41234_new_n2174_), .C(_abc_41234_new_n1626_), .Y(_abc_41234_new_n2191_));
OAI21X1 OAI21X1_386 ( .A(_abc_41234_new_n2192_), .B(_abc_41234_new_n2188_), .C(_abc_41234_new_n524_), .Y(_abc_41234_new_n2193_));
OAI21X1 OAI21X1_387 ( .A(_abc_41234_new_n2184_), .B(_abc_41234_new_n2176_), .C(_abc_41234_new_n2193_), .Y(_0alusel_2_0__1_));
OAI21X1 OAI21X1_388 ( .A(_abc_41234_new_n546__bF_buf1), .B(_abc_41234_new_n620__bF_buf1), .C(_abc_41234_new_n2196_), .Y(_abc_41234_new_n2197_));
OAI21X1 OAI21X1_389 ( .A(opcode_5_bF_buf4_), .B(_abc_41234_new_n2185__bF_buf4), .C(_abc_41234_new_n524_), .Y(_abc_41234_new_n2199_));
OAI21X1 OAI21X1_39 ( .A(_abc_41234_new_n751_), .B(_abc_41234_new_n702_), .C(_abc_41234_new_n801_), .Y(_abc_41234_new_n802_));
OAI21X1 OAI21X1_390 ( .A(_abc_41234_new_n2198_), .B(_abc_41234_new_n2199_), .C(_abc_41234_new_n2195_), .Y(_0alusel_2_0__2_));
OAI21X1 OAI21X1_391 ( .A(_abc_41234_new_n523__bF_buf0), .B(_abc_41234_new_n2181_), .C(alu_cin), .Y(_abc_41234_new_n2203_));
OAI21X1 OAI21X1_392 ( .A(_abc_41234_new_n1013_), .B(_abc_41234_new_n2202_), .C(_abc_41234_new_n2203_), .Y(_0alucin_0_0_));
OAI21X1 OAI21X1_393 ( .A(_abc_41234_new_n2206_), .B(_abc_41234_new_n2189__bF_buf3), .C(_abc_41234_new_n2209_), .Y(_abc_41234_new_n2210_));
OAI21X1 OAI21X1_394 ( .A(_abc_41234_new_n705_), .B(_abc_41234_new_n2213_), .C(_abc_41234_new_n692_), .Y(_abc_41234_new_n2214_));
OAI21X1 OAI21X1_395 ( .A(_abc_41234_new_n660__bF_buf3), .B(_abc_41234_new_n2215_), .C(_abc_41234_new_n516__bF_buf5), .Y(_abc_41234_new_n2216_));
OAI21X1 OAI21X1_396 ( .A(_abc_41234_new_n523__bF_buf4), .B(_abc_41234_new_n2211_), .C(_abc_41234_new_n2218_), .Y(_0aluoprb_7_0__0_));
OAI21X1 OAI21X1_397 ( .A(opcode_7_), .B(_abc_41234_new_n2174_), .C(_abc_41234_new_n661_), .Y(_abc_41234_new_n2221_));
OAI21X1 OAI21X1_398 ( .A(_abc_41234_new_n2220_), .B(_abc_41234_new_n2222_), .C(_abc_41234_new_n2225_), .Y(_0aluoprb_7_0__1_));
OAI21X1 OAI21X1_399 ( .A(_abc_41234_new_n2227_), .B(_abc_41234_new_n2222_), .C(_abc_41234_new_n2228_), .Y(_0aluoprb_7_0__2_));
OAI21X1 OAI21X1_4 ( .A(opcode_4_bF_buf2_), .B(_abc_41234_new_n560_), .C(_abc_41234_new_n561_), .Y(_abc_41234_new_n562_));
OAI21X1 OAI21X1_40 ( .A(_abc_41234_new_n793_), .B(_abc_41234_new_n792_), .C(_abc_41234_new_n803_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_2_));
OAI21X1 OAI21X1_400 ( .A(_abc_41234_new_n523__bF_buf2), .B(_abc_41234_new_n2230_), .C(_abc_41234_new_n2231_), .Y(_0aluoprb_7_0__3_));
OAI21X1 OAI21X1_401 ( .A(_abc_41234_new_n2233_), .B(_abc_41234_new_n2222_), .C(_abc_41234_new_n2234_), .Y(_0aluoprb_7_0__4_));
OAI21X1 OAI21X1_402 ( .A(_abc_41234_new_n2236_), .B(_abc_41234_new_n2222_), .C(_abc_41234_new_n2237_), .Y(_0aluoprb_7_0__5_));
OAI21X1 OAI21X1_403 ( .A(_abc_41234_new_n523__bF_buf1), .B(_abc_41234_new_n2239_), .C(_abc_41234_new_n2240_), .Y(_0aluoprb_7_0__6_));
OAI21X1 OAI21X1_404 ( .A(_abc_41234_new_n2242_), .B(_abc_41234_new_n2222_), .C(_abc_41234_new_n2243_), .Y(_0aluoprb_7_0__7_));
OAI21X1 OAI21X1_405 ( .A(_abc_41234_new_n569_), .B(_abc_41234_new_n2253_), .C(_abc_41234_new_n536__bF_buf5), .Y(_abc_41234_new_n2254_));
OAI21X1 OAI21X1_406 ( .A(_abc_41234_new_n1848_), .B(_abc_41234_new_n2255_), .C(_abc_41234_new_n2256_), .Y(_abc_41234_new_n2257_));
OAI21X1 OAI21X1_407 ( .A(_abc_41234_new_n2254_), .B(_abc_41234_new_n2257_), .C(_abc_41234_new_n2208_), .Y(_abc_41234_new_n2258_));
OAI21X1 OAI21X1_408 ( .A(reset_bF_buf5), .B(_abc_41234_new_n2262_), .C(_abc_41234_new_n523__bF_buf0), .Y(_abc_41234_new_n2264_));
OAI21X1 OAI21X1_409 ( .A(_abc_41234_new_n1045_), .B(_abc_41234_new_n2185__bF_buf3), .C(_abc_41234_new_n2221_), .Y(_abc_41234_new_n2265_));
OAI21X1 OAI21X1_41 ( .A(_abc_41234_new_n808_), .B(_abc_41234_new_n807_), .C(_abc_41234_new_n631_), .Y(_abc_41234_new_n809_));
OAI21X1 OAI21X1_410 ( .A(_abc_41234_new_n523__bF_buf4), .B(_abc_41234_new_n2265_), .C(_abc_41234_new_n2264_), .Y(_abc_41234_new_n2266_));
OAI21X1 OAI21X1_411 ( .A(_abc_41234_new_n2175_), .B(_abc_41234_new_n2260_), .C(_abc_41234_new_n2267_), .Y(_0aluopra_7_0__0_));
OAI21X1 OAI21X1_412 ( .A(_abc_41234_new_n570_), .B(_abc_41234_new_n2253_), .C(_abc_41234_new_n536__bF_buf3), .Y(_abc_41234_new_n2273_));
OAI21X1 OAI21X1_413 ( .A(_abc_41234_new_n730_), .B(_abc_41234_new_n2255_), .C(_abc_41234_new_n2274_), .Y(_abc_41234_new_n2275_));
OAI21X1 OAI21X1_414 ( .A(_abc_41234_new_n2273_), .B(_abc_41234_new_n2275_), .C(_abc_41234_new_n2208_), .Y(_abc_41234_new_n2276_));
OAI21X1 OAI21X1_415 ( .A(_abc_41234_new_n2175_), .B(_abc_41234_new_n2278_), .C(_abc_41234_new_n2279_), .Y(_0aluopra_7_0__1_));
OAI21X1 OAI21X1_416 ( .A(_abc_41234_new_n634_), .B(_abc_41234_new_n2253_), .C(_abc_41234_new_n536__bF_buf1), .Y(_abc_41234_new_n2285_));
OAI21X1 OAI21X1_417 ( .A(_abc_41234_new_n768_), .B(_abc_41234_new_n2255_), .C(_abc_41234_new_n2286_), .Y(_abc_41234_new_n2287_));
OAI21X1 OAI21X1_418 ( .A(_abc_41234_new_n2285_), .B(_abc_41234_new_n2287_), .C(_abc_41234_new_n2208_), .Y(_abc_41234_new_n2288_));
OAI21X1 OAI21X1_419 ( .A(_abc_41234_new_n2175_), .B(_abc_41234_new_n2290_), .C(_abc_41234_new_n2291_), .Y(_0aluopra_7_0__2_));
OAI21X1 OAI21X1_42 ( .A(regfil_0__3_), .B(_abc_41234_new_n784_), .C(_abc_41234_new_n810_), .Y(_abc_41234_new_n811_));
OAI21X1 OAI21X1_420 ( .A(_abc_41234_new_n568_), .B(_abc_41234_new_n2253_), .C(_abc_41234_new_n536__bF_buf5), .Y(_abc_41234_new_n2297_));
OAI21X1 OAI21X1_421 ( .A(_abc_41234_new_n814_), .B(_abc_41234_new_n2255_), .C(_abc_41234_new_n2298_), .Y(_abc_41234_new_n2299_));
OAI21X1 OAI21X1_422 ( .A(_abc_41234_new_n2297_), .B(_abc_41234_new_n2299_), .C(_abc_41234_new_n2208_), .Y(_abc_41234_new_n2300_));
OAI21X1 OAI21X1_423 ( .A(_abc_41234_new_n2175_), .B(_abc_41234_new_n2302_), .C(_abc_41234_new_n2303_), .Y(_0aluopra_7_0__3_));
OAI21X1 OAI21X1_424 ( .A(_abc_41234_new_n855_), .B(_abc_41234_new_n2253_), .C(_abc_41234_new_n536__bF_buf3), .Y(_abc_41234_new_n2309_));
OAI21X1 OAI21X1_425 ( .A(_abc_41234_new_n858_), .B(_abc_41234_new_n2255_), .C(_abc_41234_new_n2310_), .Y(_abc_41234_new_n2311_));
OAI21X1 OAI21X1_426 ( .A(_abc_41234_new_n2309_), .B(_abc_41234_new_n2311_), .C(_abc_41234_new_n2208_), .Y(_abc_41234_new_n2312_));
OAI21X1 OAI21X1_427 ( .A(_abc_41234_new_n2175_), .B(_abc_41234_new_n2314_), .C(_abc_41234_new_n2315_), .Y(_0aluopra_7_0__4_));
OAI21X1 OAI21X1_428 ( .A(_abc_41234_new_n896_), .B(_abc_41234_new_n2253_), .C(_abc_41234_new_n536__bF_buf2), .Y(_abc_41234_new_n2317_));
OAI21X1 OAI21X1_429 ( .A(_abc_41234_new_n899_), .B(_abc_41234_new_n2255_), .C(_abc_41234_new_n2318_), .Y(_abc_41234_new_n2319_));
OAI21X1 OAI21X1_43 ( .A(_abc_41234_new_n568_), .B(_abc_41234_new_n722__bF_buf3), .C(_abc_41234_new_n812_), .Y(_abc_41234_new_n813_));
OAI21X1 OAI21X1_430 ( .A(_abc_41234_new_n906_), .B(_abc_41234_new_n2255_), .C(opcode_5_bF_buf3_), .Y(_abc_41234_new_n2321_));
OAI21X1 OAI21X1_431 ( .A(_abc_41234_new_n907_), .B(_abc_41234_new_n2322_), .C(_abc_41234_new_n2323_), .Y(_abc_41234_new_n2324_));
OAI21X1 OAI21X1_432 ( .A(_abc_41234_new_n2321_), .B(_abc_41234_new_n2324_), .C(_abc_41234_new_n2208_), .Y(_abc_41234_new_n2325_));
OAI21X1 OAI21X1_433 ( .A(_abc_41234_new_n2175_), .B(_abc_41234_new_n2327_), .C(_abc_41234_new_n2328_), .Y(_0aluopra_7_0__5_));
OAI21X1 OAI21X1_434 ( .A(_abc_41234_new_n638_), .B(_abc_41234_new_n2253_), .C(_abc_41234_new_n536__bF_buf1), .Y(_abc_41234_new_n2330_));
OAI21X1 OAI21X1_435 ( .A(_abc_41234_new_n1936_), .B(_abc_41234_new_n2255_), .C(_abc_41234_new_n2331_), .Y(_abc_41234_new_n2332_));
OAI21X1 OAI21X1_436 ( .A(_abc_41234_new_n967_), .B(_abc_41234_new_n2255_), .C(opcode_5_bF_buf2_), .Y(_abc_41234_new_n2334_));
OAI21X1 OAI21X1_437 ( .A(_abc_41234_new_n2048_), .B(_abc_41234_new_n2322_), .C(_abc_41234_new_n2335_), .Y(_abc_41234_new_n2336_));
OAI21X1 OAI21X1_438 ( .A(_abc_41234_new_n2334_), .B(_abc_41234_new_n2336_), .C(_abc_41234_new_n2208_), .Y(_abc_41234_new_n2337_));
OAI21X1 OAI21X1_439 ( .A(_abc_41234_new_n2175_), .B(_abc_41234_new_n2339_), .C(_abc_41234_new_n2340_), .Y(_0aluopra_7_0__6_));
OAI21X1 OAI21X1_44 ( .A(_abc_41234_new_n816_), .B(_abc_41234_new_n813_), .C(_abc_41234_new_n546__bF_buf3), .Y(_abc_41234_new_n817_));
OAI21X1 OAI21X1_440 ( .A(_abc_41234_new_n2344_), .B(_abc_41234_new_n2343_), .C(_abc_41234_new_n536__bF_buf0), .Y(_abc_41234_new_n2345_));
OAI21X1 OAI21X1_441 ( .A(_abc_41234_new_n2346_), .B(_abc_41234_new_n2347_), .C(opcode_5_bF_buf1_), .Y(_abc_41234_new_n2348_));
OAI21X1 OAI21X1_442 ( .A(_abc_41234_new_n2175_), .B(_abc_41234_new_n2350_), .C(_abc_41234_new_n2351_), .Y(_0aluopra_7_0__7_));
OAI21X1 OAI21X1_443 ( .A(intcyc_bF_buf3), .B(_abc_41234_new_n2358_), .C(_abc_41234_new_n516__bF_buf3), .Y(_abc_41234_new_n2359_));
OAI21X1 OAI21X1_444 ( .A(state_4_), .B(_abc_41234_new_n612_), .C(_abc_41234_new_n706_), .Y(_abc_41234_new_n2362_));
OAI21X1 OAI21X1_445 ( .A(_abc_41234_new_n509_), .B(_abc_41234_new_n2362_), .C(_abc_41234_new_n516__bF_buf2), .Y(_abc_41234_new_n2363_));
OAI21X1 OAI21X1_446 ( .A(_abc_41234_new_n1878_), .B(_abc_41234_new_n1851_), .C(parity), .Y(_abc_41234_new_n2366_));
OAI21X1 OAI21X1_447 ( .A(_abc_41234_new_n2365_), .B(_abc_41234_new_n510_), .C(_abc_41234_new_n2366_), .Y(_abc_41234_new_n2367_));
OAI21X1 OAI21X1_448 ( .A(_abc_41234_new_n1878_), .B(_abc_41234_new_n1851_), .C(zero), .Y(_abc_41234_new_n2372_));
OAI21X1 OAI21X1_449 ( .A(_abc_41234_new_n2371_), .B(_abc_41234_new_n510_), .C(_abc_41234_new_n2372_), .Y(_abc_41234_new_n2373_));
OAI21X1 OAI21X1_45 ( .A(_abc_41234_new_n823_), .B(_abc_41234_new_n820_), .C(opcode_2_), .Y(_abc_41234_new_n824_));
OAI21X1 OAI21X1_450 ( .A(reset_bF_buf3), .B(_abc_41234_new_n2374_), .C(_abc_41234_new_n2370_), .Y(_0zero_0_0_));
OAI21X1 OAI21X1_451 ( .A(_abc_41234_new_n2379_), .B(_abc_41234_new_n706_), .C(_abc_41234_new_n2380_), .Y(_abc_41234_new_n2381_));
OAI21X1 OAI21X1_452 ( .A(_abc_41234_new_n550_), .B(_abc_41234_new_n2384_), .C(_abc_41234_new_n2385_), .Y(_abc_41234_new_n2386_));
OAI21X1 OAI21X1_453 ( .A(_abc_41234_new_n508_), .B(_abc_41234_new_n2387_), .C(_abc_41234_new_n2388_), .Y(_abc_41234_new_n2389_));
OAI21X1 OAI21X1_454 ( .A(reset_bF_buf1), .B(_abc_41234_new_n2390_), .C(_abc_41234_new_n2391_), .Y(_0auxcar_0_0_));
OAI21X1 OAI21X1_455 ( .A(_abc_41234_new_n504_), .B(_abc_41234_new_n659_), .C(_abc_41234_new_n706_), .Y(_abc_41234_new_n2393_));
OAI21X1 OAI21X1_456 ( .A(_abc_41234_new_n509_), .B(_abc_41234_new_n2393_), .C(_abc_41234_new_n516__bF_buf1), .Y(_abc_41234_new_n2394_));
OAI21X1 OAI21X1_457 ( .A(_abc_41234_new_n1545_), .B(_abc_41234_new_n1549_), .C(_abc_41234_new_n2396_), .Y(_abc_41234_new_n2397_));
OAI21X1 OAI21X1_458 ( .A(_abc_41234_new_n1579_), .B(_abc_41234_new_n2397_), .C(_abc_41234_new_n2399_), .Y(_abc_41234_new_n2400_));
OAI21X1 OAI21X1_459 ( .A(_abc_41234_new_n2402_), .B(_abc_41234_new_n1533_), .C(_abc_41234_new_n2401_), .Y(_abc_41234_new_n2403_));
OAI21X1 OAI21X1_46 ( .A(regfil_7__3_), .B(_abc_41234_new_n678_), .C(_abc_41234_new_n710_), .Y(_abc_41234_new_n831_));
OAI21X1 OAI21X1_460 ( .A(_abc_41234_new_n680_), .B(_abc_41234_new_n532_), .C(_abc_41234_new_n2404_), .Y(_abc_41234_new_n2405_));
OAI21X1 OAI21X1_461 ( .A(_abc_41234_new_n997_), .B(_abc_41234_new_n1575_), .C(_abc_41234_new_n2406_), .Y(_abc_41234_new_n2407_));
OAI21X1 OAI21X1_462 ( .A(_abc_41234_new_n1570_), .B(_abc_41234_new_n1567_), .C(_abc_41234_new_n2409_), .Y(_abc_41234_new_n2410_));
OAI21X1 OAI21X1_463 ( .A(_abc_41234_new_n2414_), .B(_abc_41234_new_n2411_), .C(_abc_41234_new_n2416_), .Y(_abc_41234_new_n2417_));
OAI21X1 OAI21X1_464 ( .A(_abc_41234_new_n2418_), .B(_abc_41234_new_n706_), .C(_abc_41234_new_n2419_), .Y(_abc_41234_new_n2420_));
OAI21X1 OAI21X1_465 ( .A(_abc_41234_new_n1878_), .B(_abc_41234_new_n1851_), .C(carry), .Y(_abc_41234_new_n2422_));
OAI21X1 OAI21X1_466 ( .A(_abc_41234_new_n2421_), .B(_abc_41234_new_n510_), .C(_abc_41234_new_n2422_), .Y(_abc_41234_new_n2423_));
OAI21X1 OAI21X1_467 ( .A(reset_bF_buf0), .B(_abc_41234_new_n2425_), .C(_abc_41234_new_n2395_), .Y(_0carry_0_0_));
OAI21X1 OAI21X1_468 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n2428_), .C(opcode_1_), .Y(_abc_41234_new_n2433_));
OAI21X1 OAI21X1_469 ( .A(_abc_41234_new_n2432_), .B(_abc_41234_new_n2430_), .C(_abc_41234_new_n2433_), .Y(_0opcode_7_0__1_));
OAI21X1 OAI21X1_47 ( .A(_abc_41234_new_n821_), .B(_abc_41234_new_n834_), .C(_abc_41234_new_n795_), .Y(_abc_41234_new_n835_));
OAI21X1 OAI21X1_470 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n2428_), .C(opcode_3_bF_buf0_), .Y(_abc_41234_new_n2438_));
OAI21X1 OAI21X1_471 ( .A(_abc_41234_new_n2437_), .B(_abc_41234_new_n2430_), .C(_abc_41234_new_n2438_), .Y(_0opcode_7_0__3_));
OAI21X1 OAI21X1_472 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n2428_), .C(opcode_6_), .Y(_abc_41234_new_n2444_));
OAI21X1 OAI21X1_473 ( .A(_abc_41234_new_n2443_), .B(_abc_41234_new_n2430_), .C(_abc_41234_new_n2444_), .Y(_0opcode_7_0__6_));
OAI21X1 OAI21X1_474 ( .A(_abc_41234_new_n757_), .B(_abc_41234_new_n2428_), .C(opcode_7_), .Y(_abc_41234_new_n2446_));
OAI21X1 OAI21X1_475 ( .A(_abc_41234_new_n1016_), .B(_abc_41234_new_n2430_), .C(_abc_41234_new_n2446_), .Y(_0opcode_7_0__7_));
OAI21X1 OAI21X1_476 ( .A(_abc_41234_new_n2353_), .B(_abc_41234_new_n2212_), .C(eienb), .Y(_abc_41234_new_n2448_));
OAI21X1 OAI21X1_477 ( .A(_abc_41234_new_n1322_), .B(_abc_41234_new_n1051_), .C(_abc_41234_new_n2456_), .Y(_abc_41234_new_n2457_));
OAI21X1 OAI21X1_478 ( .A(_abc_41234_new_n556_), .B(_abc_41234_new_n722__bF_buf3), .C(_abc_41234_new_n1645_), .Y(_abc_41234_new_n2463_));
OAI21X1 OAI21X1_479 ( .A(_abc_41234_new_n546__bF_buf4), .B(_abc_41234_new_n620__bF_buf0), .C(_abc_41234_new_n1040__bF_buf3), .Y(_abc_41234_new_n2465_));
OAI21X1 OAI21X1_48 ( .A(regfil_7__3_), .B(_abc_41234_new_n540_), .C(_abc_41234_new_n835_), .Y(_abc_41234_new_n836_));
OAI21X1 OAI21X1_480 ( .A(_abc_41234_new_n530_), .B(_abc_41234_new_n531_), .C(_abc_41234_new_n2466_), .Y(_abc_41234_new_n2467_));
OAI21X1 OAI21X1_481 ( .A(_abc_41234_new_n2322_), .B(_abc_41234_new_n2471_), .C(_abc_41234_new_n2470_), .Y(_abc_41234_new_n2472_));
OAI21X1 OAI21X1_482 ( .A(_abc_41234_new_n580_), .B(_abc_41234_new_n722__bF_buf2), .C(_abc_41234_new_n2481_), .Y(_abc_41234_new_n2482_));
OAI21X1 OAI21X1_483 ( .A(_abc_41234_new_n2455_), .B(_abc_41234_new_n2480_), .C(_abc_41234_new_n2484_), .Y(_abc_41234_new_n2485_));
OAI21X1 OAI21X1_484 ( .A(_abc_41234_new_n537__bF_buf0), .B(_abc_41234_new_n1684_), .C(_abc_41234_new_n2469_), .Y(_abc_41234_new_n2486_));
OAI21X1 OAI21X1_485 ( .A(_abc_41234_new_n721_), .B(_abc_41234_new_n616_), .C(opcode_2_), .Y(_abc_41234_new_n2489_));
OAI21X1 OAI21X1_486 ( .A(_abc_41234_new_n536__bF_buf3), .B(_abc_41234_new_n2488_), .C(_abc_41234_new_n2489_), .Y(_abc_41234_new_n2490_));
OAI21X1 OAI21X1_487 ( .A(_abc_41234_new_n2174_), .B(_abc_41234_new_n2493_), .C(_abc_41234_new_n515__bF_buf6), .Y(_abc_41234_new_n2494_));
OAI21X1 OAI21X1_488 ( .A(_abc_41234_new_n668__bF_buf4), .B(_abc_41234_new_n2493_), .C(statesel_0_), .Y(_abc_41234_new_n2495_));
OAI21X1 OAI21X1_489 ( .A(_abc_41234_new_n2342_), .B(_abc_41234_new_n2471_), .C(_abc_41234_new_n2496_), .Y(_abc_41234_new_n2497_));
OAI21X1 OAI21X1_49 ( .A(regfil_7__2_), .B(_abc_41234_new_n839_), .C(_abc_41234_new_n688_), .Y(_abc_41234_new_n840_));
OAI21X1 OAI21X1_490 ( .A(opcode_3_bF_buf3_), .B(_abc_41234_new_n1105__bF_buf3), .C(_abc_41234_new_n665__bF_buf3), .Y(_abc_41234_new_n2499_));
OAI21X1 OAI21X1_491 ( .A(_abc_41234_new_n546__bF_buf3), .B(_abc_41234_new_n620__bF_buf3), .C(_abc_41234_new_n2189__bF_buf5), .Y(_abc_41234_new_n2501_));
OAI21X1 OAI21X1_492 ( .A(_abc_41234_new_n2185__bF_buf1), .B(_abc_41234_new_n669__bF_buf2), .C(_abc_41234_new_n662_), .Y(_abc_41234_new_n2502_));
OAI21X1 OAI21X1_493 ( .A(_abc_41234_new_n546__bF_buf2), .B(_abc_41234_new_n620__bF_buf2), .C(_abc_41234_new_n669__bF_buf1), .Y(_abc_41234_new_n2504_));
OAI21X1 OAI21X1_494 ( .A(statesel_0_), .B(_abc_41234_new_n2505_), .C(_abc_41234_new_n2503_), .Y(_abc_41234_new_n2506_));
OAI21X1 OAI21X1_495 ( .A(_abc_41234_new_n2455_), .B(_abc_41234_new_n2501_), .C(_abc_41234_new_n2506_), .Y(_abc_41234_new_n2507_));
OAI21X1 OAI21X1_496 ( .A(_abc_41234_new_n2494_), .B(_abc_41234_new_n2495_), .C(_abc_41234_new_n2508_), .Y(_abc_41234_new_n2509_));
OAI21X1 OAI21X1_497 ( .A(_abc_41234_new_n607_), .B(_abc_41234_new_n2212_), .C(_abc_41234_new_n2515_), .Y(_abc_41234_new_n2516_));
OAI21X1 OAI21X1_498 ( .A(_abc_41234_new_n693_), .B(_abc_41234_new_n612_), .C(_abc_41234_new_n2519_), .Y(_abc_41234_new_n2520_));
OAI21X1 OAI21X1_499 ( .A(_abc_41234_new_n659_), .B(_abc_41234_new_n604_), .C(_abc_41234_new_n2521_), .Y(_abc_41234_new_n2522_));
OAI21X1 OAI21X1_5 ( .A(_abc_41234_new_n513_), .B(_abc_41234_new_n564_), .C(_abc_41234_new_n566_), .Y(_abc_41234_new_n567_));
OAI21X1 OAI21X1_50 ( .A(_abc_41234_new_n840_), .B(_abc_41234_new_n838_), .C(_abc_41234_new_n841_), .Y(_abc_41234_new_n842_));
OAI21X1 OAI21X1_500 ( .A(_abc_41234_new_n504_), .B(_abc_41234_new_n659_), .C(_abc_41234_new_n2526_), .Y(_abc_41234_new_n2527_));
OAI21X1 OAI21X1_501 ( .A(_abc_41234_new_n2527_), .B(_abc_41234_new_n2525_), .C(_abc_41234_new_n516__bF_buf4), .Y(_abc_41234_new_n2528_));
OAI21X1 OAI21X1_502 ( .A(reset_bF_buf9), .B(_abc_41234_new_n2531_), .C(_abc_41234_new_n2529_), .Y(_abc_41234_new_n2532_));
OAI21X1 OAI21X1_503 ( .A(_abc_41234_new_n2533_), .B(_abc_41234_new_n2525_), .C(_abc_41234_new_n516__bF_buf3), .Y(_abc_41234_new_n2534_));
OAI21X1 OAI21X1_504 ( .A(_abc_41234_new_n523__bF_buf2), .B(_abc_41234_new_n2510_), .C(_abc_41234_new_n2536_), .Y(_0statesel_5_0__0_));
OAI21X1 OAI21X1_505 ( .A(_abc_41234_new_n580_), .B(_abc_41234_new_n722__bF_buf1), .C(_abc_41234_new_n2476_), .Y(_abc_41234_new_n2539_));
OAI21X1 OAI21X1_506 ( .A(_abc_41234_new_n2541_), .B(_abc_41234_new_n2493_), .C(statesel_1_), .Y(_abc_41234_new_n2542_));
OAI21X1 OAI21X1_507 ( .A(_abc_41234_new_n2466_), .B(_abc_41234_new_n1608_), .C(_abc_41234_new_n537__bF_buf3), .Y(_abc_41234_new_n2543_));
OAI21X1 OAI21X1_508 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n2488_), .C(_abc_41234_new_n2499_), .Y(_abc_41234_new_n2545_));
OAI21X1 OAI21X1_509 ( .A(statesel_1_), .B(_abc_41234_new_n665__bF_buf2), .C(_abc_41234_new_n2189__bF_buf4), .Y(_abc_41234_new_n2549_));
OAI21X1 OAI21X1_51 ( .A(_abc_41234_new_n821_), .B(_abc_41234_new_n702_), .C(_abc_41234_new_n843_), .Y(_abc_41234_new_n844_));
OAI21X1 OAI21X1_510 ( .A(_abc_41234_new_n665__bF_buf0), .B(_abc_41234_new_n668__bF_buf2), .C(_abc_41234_new_n662_), .Y(_abc_41234_new_n2551_));
OAI21X1 OAI21X1_511 ( .A(_abc_41234_new_n2551_), .B(_abc_41234_new_n2550_), .C(_abc_41234_new_n2549_), .Y(_abc_41234_new_n2552_));
OAI21X1 OAI21X1_512 ( .A(_abc_41234_new_n1047__bF_buf1), .B(_abc_41234_new_n2540_), .C(_abc_41234_new_n2553_), .Y(_abc_41234_new_n2554_));
OAI21X1 OAI21X1_513 ( .A(reset_bF_buf8), .B(_abc_41234_new_n2555_), .C(_abc_41234_new_n2561_), .Y(_0statesel_5_0__1_));
OAI21X1 OAI21X1_514 ( .A(_abc_41234_new_n2502_), .B(_abc_41234_new_n2505_), .C(_abc_41234_new_n2501_), .Y(_abc_41234_new_n2567_));
OAI21X1 OAI21X1_515 ( .A(opcode_5_bF_buf0_), .B(_abc_41234_new_n2488_), .C(_abc_41234_new_n2185__bF_buf0), .Y(_abc_41234_new_n2569_));
OAI21X1 OAI21X1_516 ( .A(statesel_2_), .B(_abc_41234_new_n2571_), .C(_abc_41234_new_n515__bF_buf3), .Y(_abc_41234_new_n2572_));
OAI21X1 OAI21X1_517 ( .A(_abc_41234_new_n1047__bF_buf0), .B(_abc_41234_new_n2566_), .C(_abc_41234_new_n2574_), .Y(_abc_41234_new_n2575_));
OAI21X1 OAI21X1_518 ( .A(_abc_41234_new_n2581_), .B(_abc_41234_new_n2582_), .C(_abc_41234_new_n2533_), .Y(_abc_41234_new_n2583_));
OAI21X1 OAI21X1_519 ( .A(_abc_41234_new_n2580_), .B(_abc_41234_new_n2577_), .C(_abc_41234_new_n2583_), .Y(_abc_41234_new_n2584_));
OAI21X1 OAI21X1_52 ( .A(_abc_41234_new_n831_), .B(_abc_41234_new_n830_), .C(_abc_41234_new_n845_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_3_));
OAI21X1 OAI21X1_520 ( .A(reset_bF_buf6), .B(_abc_41234_new_n2576_), .C(_abc_41234_new_n2586_), .Y(_0statesel_5_0__2_));
OAI21X1 OAI21X1_521 ( .A(_abc_41234_new_n536__bF_buf1), .B(_abc_41234_new_n2488_), .C(_abc_41234_new_n2185__bF_buf5), .Y(_abc_41234_new_n2591_));
OAI21X1 OAI21X1_522 ( .A(statesel_3_), .B(_abc_41234_new_n2571_), .C(_abc_41234_new_n515__bF_buf2), .Y(_abc_41234_new_n2594_));
OAI21X1 OAI21X1_523 ( .A(_abc_41234_new_n2190__bF_buf1), .B(_abc_41234_new_n2185__bF_buf4), .C(_abc_41234_new_n2588_), .Y(_abc_41234_new_n2596_));
OAI21X1 OAI21X1_524 ( .A(_abc_41234_new_n2502_), .B(_abc_41234_new_n2505_), .C(_abc_41234_new_n2190__bF_buf0), .Y(_abc_41234_new_n2597_));
OAI21X1 OAI21X1_525 ( .A(_abc_41234_new_n1047__bF_buf4), .B(_abc_41234_new_n2590_), .C(_abc_41234_new_n2598_), .Y(_abc_41234_new_n2599_));
OAI21X1 OAI21X1_526 ( .A(_abc_41234_new_n2526_), .B(_abc_41234_new_n2580_), .C(_abc_41234_new_n2531_), .Y(_abc_41234_new_n2606_));
OAI21X1 OAI21X1_527 ( .A(_abc_41234_new_n2606_), .B(_abc_41234_new_n2605_), .C(statesel_3_), .Y(_abc_41234_new_n2607_));
OAI21X1 OAI21X1_528 ( .A(_abc_41234_new_n2600_), .B(_abc_41234_new_n2604_), .C(_abc_41234_new_n2607_), .Y(_abc_41234_new_n2608_));
OAI21X1 OAI21X1_529 ( .A(_abc_41234_new_n668__bF_buf1), .B(_abc_41234_new_n2207__bF_buf1), .C(_abc_41234_new_n2486_), .Y(_abc_41234_new_n2615_));
OAI21X1 OAI21X1_53 ( .A(_abc_41234_new_n855_), .B(_abc_41234_new_n722__bF_buf0), .C(_abc_41234_new_n856_), .Y(_abc_41234_new_n857_));
OAI21X1 OAI21X1_530 ( .A(_abc_41234_new_n2185__bF_buf3), .B(_abc_41234_new_n2190__bF_buf3), .C(_abc_41234_new_n2616_), .Y(_abc_41234_new_n2617_));
OAI21X1 OAI21X1_531 ( .A(_abc_41234_new_n1047__bF_buf3), .B(_abc_41234_new_n2612_), .C(_abc_41234_new_n2618_), .Y(_abc_41234_new_n2619_));
OAI21X1 OAI21X1_532 ( .A(_abc_41234_new_n2533_), .B(_abc_41234_new_n2525_), .C(_abc_41234_new_n2624_), .Y(_abc_41234_new_n2625_));
OAI21X1 OAI21X1_533 ( .A(statesel_5_), .B(_abc_41234_new_n2480_), .C(_abc_41234_new_n1046__bF_buf6), .Y(_abc_41234_new_n2629_));
OAI21X1 OAI21X1_534 ( .A(waitr), .B(_abc_41234_new_n2624_), .C(_abc_41234_new_n2634_), .Y(_abc_41234_new_n2635_));
OAI21X1 OAI21X1_535 ( .A(_abc_41234_new_n2633_), .B(_abc_41234_new_n2577_), .C(_abc_41234_new_n2635_), .Y(_abc_41234_new_n2636_));
OAI21X1 OAI21X1_536 ( .A(reset_bF_buf3), .B(_abc_41234_new_n2637_), .C(_abc_41234_new_n2642_), .Y(_0statesel_5_0__5_));
OAI21X1 OAI21X1_537 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n2644_), .C(_abc_41234_new_n2645_), .Y(_0popdes_1_0__0_));
OAI21X1 OAI21X1_538 ( .A(_abc_41234_new_n536__bF_buf0), .B(_abc_41234_new_n2644_), .C(_abc_41234_new_n2647_), .Y(_0popdes_1_0__1_));
OAI21X1 OAI21X1_539 ( .A(_abc_41234_new_n504_), .B(_abc_41234_new_n659_), .C(_abc_41234_new_n2671_), .Y(_abc_41234_new_n2672_));
OAI21X1 OAI21X1_54 ( .A(_abc_41234_new_n860_), .B(_abc_41234_new_n857_), .C(_abc_41234_new_n546__bF_buf2), .Y(_abc_41234_new_n861_));
OAI21X1 OAI21X1_540 ( .A(_abc_41234_new_n693_), .B(_abc_41234_new_n612_), .C(_abc_41234_new_n2515_), .Y(_abc_41234_new_n2673_));
OAI21X1 OAI21X1_541 ( .A(_abc_41234_new_n661_), .B(_abc_41234_new_n1644_), .C(opcode_7_), .Y(_abc_41234_new_n2676_));
OAI21X1 OAI21X1_542 ( .A(_abc_41234_new_n680_), .B(_abc_41234_new_n537__bF_buf2), .C(_abc_41234_new_n1608_), .Y(_abc_41234_new_n2678_));
OAI21X1 OAI21X1_543 ( .A(_abc_41234_new_n2677_), .B(_abc_41234_new_n2678_), .C(_abc_41234_new_n2679_), .Y(_abc_41234_new_n2680_));
OAI21X1 OAI21X1_544 ( .A(wdatahold_0_), .B(_abc_41234_new_n2505_), .C(_abc_41234_new_n662_), .Y(_abc_41234_new_n2682_));
OAI21X1 OAI21X1_545 ( .A(_abc_41234_new_n2682_), .B(_abc_41234_new_n2681_), .C(_abc_41234_new_n2680_), .Y(_abc_41234_new_n2683_));
OAI21X1 OAI21X1_546 ( .A(_abc_41234_new_n1013_), .B(_abc_41234_new_n1105__bF_buf2), .C(_abc_41234_new_n2686_), .Y(_abc_41234_new_n2687_));
OAI21X1 OAI21X1_547 ( .A(regfil_1__0_), .B(_abc_41234_new_n1322_), .C(_abc_41234_new_n1639__bF_buf1), .Y(_abc_41234_new_n2688_));
OAI21X1 OAI21X1_548 ( .A(_abc_41234_new_n1221_), .B(_abc_41234_new_n1040__bF_buf1), .C(_abc_41234_new_n2688_), .Y(_abc_41234_new_n2689_));
OAI21X1 OAI21X1_549 ( .A(pc_0_), .B(_abc_41234_new_n1638_), .C(_abc_41234_new_n2690_), .Y(_abc_41234_new_n2691_));
OAI21X1 OAI21X1_55 ( .A(_abc_41234_new_n546__bF_buf1), .B(_abc_41234_new_n854_), .C(_abc_41234_new_n861_), .Y(_abc_41234_new_n862_));
OAI21X1 OAI21X1_550 ( .A(_abc_41234_new_n2670_), .B(_abc_41234_new_n2676_), .C(_abc_41234_new_n2692_), .Y(_abc_41234_new_n2693_));
OAI21X1 OAI21X1_551 ( .A(_abc_41234_new_n565_), .B(_abc_41234_new_n2515_), .C(_abc_41234_new_n2697_), .Y(_abc_41234_new_n2698_));
OAI21X1 OAI21X1_552 ( .A(opcode_6_), .B(_abc_41234_new_n1608_), .C(_abc_41234_new_n2551_), .Y(_abc_41234_new_n2703_));
OAI21X1 OAI21X1_553 ( .A(_abc_41234_new_n2703_), .B(_abc_41234_new_n2702_), .C(wdatahold_1_), .Y(_abc_41234_new_n2704_));
OAI21X1 OAI21X1_554 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n730_), .C(_abc_41234_new_n1105__bF_buf1), .Y(_abc_41234_new_n2712_));
OAI21X1 OAI21X1_555 ( .A(_abc_41234_new_n2712_), .B(_abc_41234_new_n2711_), .C(_abc_41234_new_n1639__bF_buf0), .Y(_abc_41234_new_n2713_));
OAI21X1 OAI21X1_556 ( .A(_abc_41234_new_n536__bF_buf4), .B(_abc_41234_new_n719_), .C(_abc_41234_new_n2713_), .Y(_abc_41234_new_n2714_));
OAI21X1 OAI21X1_557 ( .A(_abc_41234_new_n2710_), .B(_abc_41234_new_n1639__bF_buf3), .C(_abc_41234_new_n2714_), .Y(_abc_41234_new_n2715_));
OAI21X1 OAI21X1_558 ( .A(_abc_41234_new_n1645_), .B(_abc_41234_new_n2706_), .C(_abc_41234_new_n2716_), .Y(_abc_41234_new_n2717_));
OAI21X1 OAI21X1_559 ( .A(opcode_4_bF_buf3_), .B(_abc_41234_new_n536__bF_buf3), .C(_abc_41234_new_n1608_), .Y(_abc_41234_new_n2719_));
OAI21X1 OAI21X1_56 ( .A(_abc_41234_new_n615_), .B(_abc_41234_new_n863_), .C(_abc_41234_new_n864_), .Y(_abc_41234_new_n865_));
OAI21X1 OAI21X1_560 ( .A(_abc_41234_new_n735_), .B(_abc_41234_new_n2721_), .C(_abc_41234_new_n2190__bF_buf1), .Y(_abc_41234_new_n2722_));
OAI21X1 OAI21X1_561 ( .A(_abc_41234_new_n1646_), .B(_abc_41234_new_n1647_), .C(_abc_41234_new_n1614_), .Y(_abc_41234_new_n2734_));
OAI21X1 OAI21X1_562 ( .A(pc_1_), .B(pc_0_), .C(pc_2_), .Y(_abc_41234_new_n2736_));
OAI21X1 OAI21X1_563 ( .A(pc_0_), .B(_abc_41234_new_n2738_), .C(_abc_41234_new_n2736_), .Y(_abc_41234_new_n2739_));
OAI21X1 OAI21X1_564 ( .A(_abc_41234_new_n2361_), .B(_abc_41234_new_n1105__bF_buf0), .C(_abc_41234_new_n2741_), .Y(_abc_41234_new_n2742_));
OAI21X1 OAI21X1_565 ( .A(regfil_1__2_), .B(_abc_41234_new_n1322_), .C(_abc_41234_new_n2742_), .Y(_abc_41234_new_n2743_));
OAI21X1 OAI21X1_566 ( .A(pc_2_), .B(_abc_41234_new_n1729_), .C(_abc_41234_new_n2746_), .Y(_abc_41234_new_n2747_));
OAI21X1 OAI21X1_567 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n1040__bF_buf0), .C(_abc_41234_new_n2747_), .Y(_abc_41234_new_n2748_));
OAI21X1 OAI21X1_568 ( .A(_abc_41234_new_n751_), .B(_abc_41234_new_n537__bF_buf3), .C(_abc_41234_new_n2752_), .Y(_abc_41234_new_n2753_));
OAI21X1 OAI21X1_569 ( .A(_abc_41234_new_n1610_), .B(_abc_41234_new_n2753_), .C(_abc_41234_new_n2754_), .Y(_abc_41234_new_n2755_));
OAI21X1 OAI21X1_57 ( .A(_abc_41234_new_n847_), .B(_abc_41234_new_n632_), .C(_abc_41234_new_n878_), .Y(_abc_41234_new_n879_));
OAI21X1 OAI21X1_570 ( .A(opcode_6_), .B(_abc_41234_new_n1045_), .C(_abc_41234_new_n2551_), .Y(_abc_41234_new_n2756_));
OAI21X1 OAI21X1_571 ( .A(_abc_41234_new_n2758_), .B(_abc_41234_new_n2750_), .C(_abc_41234_new_n660__bF_buf2), .Y(_abc_41234_new_n2759_));
OAI21X1 OAI21X1_572 ( .A(_abc_41234_new_n821_), .B(_abc_41234_new_n537__bF_buf2), .C(_abc_41234_new_n1608_), .Y(_abc_41234_new_n2766_));
OAI21X1 OAI21X1_573 ( .A(_abc_41234_new_n2504_), .B(_abc_41234_new_n825_), .C(_abc_41234_new_n2768_), .Y(_abc_41234_new_n2769_));
OAI21X1 OAI21X1_574 ( .A(_abc_41234_new_n534__bF_buf3), .B(_abc_41234_new_n2767_), .C(_abc_41234_new_n2769_), .Y(_abc_41234_new_n2770_));
OAI21X1 OAI21X1_575 ( .A(_abc_41234_new_n1647_), .B(_abc_41234_new_n2771_), .C(_abc_41234_new_n1613_), .Y(_abc_41234_new_n2772_));
OAI21X1 OAI21X1_576 ( .A(_abc_41234_new_n1614_), .B(_abc_41234_new_n2705_), .C(_abc_41234_new_n1613_), .Y(_abc_41234_new_n2775_));
OAI21X1 OAI21X1_577 ( .A(_abc_41234_new_n1613_), .B(_abc_41234_new_n1729_), .C(_abc_41234_new_n2777_), .Y(_abc_41234_new_n2778_));
OAI21X1 OAI21X1_578 ( .A(regfil_1__3_), .B(_abc_41234_new_n1322_), .C(_abc_41234_new_n1639__bF_buf2), .Y(_abc_41234_new_n2781_));
OAI21X1 OAI21X1_579 ( .A(_abc_41234_new_n2780_), .B(_abc_41234_new_n2781_), .C(_abc_41234_new_n2782_), .Y(_abc_41234_new_n2783_));
OAI21X1 OAI21X1_58 ( .A(regfil_7__4_), .B(_abc_41234_new_n678_), .C(_abc_41234_new_n710_), .Y(_abc_41234_new_n881_));
OAI21X1 OAI21X1_580 ( .A(_abc_41234_new_n2774_), .B(_abc_41234_new_n1645_), .C(_abc_41234_new_n2784_), .Y(_abc_41234_new_n2785_));
OAI21X1 OAI21X1_581 ( .A(_abc_41234_new_n2764_), .B(_abc_41234_new_n2676_), .C(_abc_41234_new_n2786_), .Y(_abc_41234_new_n2787_));
OAI21X1 OAI21X1_582 ( .A(_abc_41234_new_n832_), .B(_abc_41234_new_n2515_), .C(_abc_41234_new_n2788_), .Y(_abc_41234_new_n2789_));
OAI21X1 OAI21X1_583 ( .A(_abc_41234_new_n2189__bF_buf2), .B(_abc_41234_new_n2702_), .C(wdatahold_4_), .Y(_abc_41234_new_n2793_));
OAI21X1 OAI21X1_584 ( .A(_abc_41234_new_n851_), .B(_abc_41234_new_n537__bF_buf0), .C(_abc_41234_new_n2794_), .Y(_abc_41234_new_n2795_));
OAI21X1 OAI21X1_585 ( .A(_abc_41234_new_n620__bF_buf1), .B(_abc_41234_new_n580_), .C(_abc_41234_new_n2792_), .Y(_abc_41234_new_n2796_));
OAI21X1 OAI21X1_586 ( .A(_abc_41234_new_n2795_), .B(_abc_41234_new_n1610_), .C(_abc_41234_new_n2796_), .Y(_abc_41234_new_n2797_));
OAI21X1 OAI21X1_587 ( .A(_abc_41234_new_n2504_), .B(_abc_41234_new_n862_), .C(_abc_41234_new_n2798_), .Y(_abc_41234_new_n2799_));
OAI21X1 OAI21X1_588 ( .A(_abc_41234_new_n534__bF_buf2), .B(_abc_41234_new_n2797_), .C(_abc_41234_new_n2799_), .Y(_abc_41234_new_n2800_));
OAI21X1 OAI21X1_589 ( .A(intcyc_bF_buf0), .B(_abc_41234_new_n2805_), .C(_abc_41234_new_n2807_), .Y(_abc_41234_new_n2808_));
OAI21X1 OAI21X1_59 ( .A(regfil_7__4_), .B(_abc_41234_new_n835_), .C(_abc_41234_new_n839_), .Y(_abc_41234_new_n885_));
OAI21X1 OAI21X1_590 ( .A(_abc_41234_new_n2809_), .B(_abc_41234_new_n1105__bF_buf3), .C(_abc_41234_new_n2794_), .Y(_abc_41234_new_n2810_));
OAI21X1 OAI21X1_591 ( .A(regfil_1__4_), .B(_abc_41234_new_n1322_), .C(_abc_41234_new_n1639__bF_buf1), .Y(_abc_41234_new_n2813_));
OAI21X1 OAI21X1_592 ( .A(_abc_41234_new_n1645_), .B(_abc_41234_new_n2802_), .C(_abc_41234_new_n2816_), .Y(_abc_41234_new_n2817_));
OAI21X1 OAI21X1_593 ( .A(_abc_41234_new_n847_), .B(_abc_41234_new_n2515_), .C(_abc_41234_new_n2820_), .Y(_abc_41234_new_n2821_));
OAI21X1 OAI21X1_594 ( .A(_abc_41234_new_n2821_), .B(_abc_41234_new_n2819_), .C(_abc_41234_new_n516__bF_buf2), .Y(_abc_41234_new_n2822_));
OAI21X1 OAI21X1_595 ( .A(_abc_41234_new_n2792_), .B(_abc_41234_new_n2675_), .C(_abc_41234_new_n2822_), .Y(_0wdatahold_7_0__4_));
OAI21X1 OAI21X1_596 ( .A(_abc_41234_new_n906_), .B(_abc_41234_new_n537__bF_buf3), .C(_abc_41234_new_n1608_), .Y(_abc_41234_new_n2826_));
OAI21X1 OAI21X1_597 ( .A(_abc_41234_new_n2504_), .B(_abc_41234_new_n910_), .C(_abc_41234_new_n2828_), .Y(_abc_41234_new_n2829_));
OAI21X1 OAI21X1_598 ( .A(_abc_41234_new_n534__bF_buf1), .B(_abc_41234_new_n2827_), .C(_abc_41234_new_n2829_), .Y(_abc_41234_new_n2830_));
OAI21X1 OAI21X1_599 ( .A(_abc_41234_new_n2806_), .B(_abc_41234_new_n1649_), .C(_abc_41234_new_n2831_), .Y(_abc_41234_new_n2832_));
OAI21X1 OAI21X1_6 ( .A(regfil_0__0_), .B(_abc_41234_new_n578_), .C(_abc_41234_new_n587_), .Y(_abc_41234_new_n588_));
OAI21X1 OAI21X1_60 ( .A(_abc_41234_new_n890_), .B(_abc_41234_new_n683_), .C(_abc_41234_new_n891_), .Y(_abc_41234_new_n892_));
OAI21X1 OAI21X1_600 ( .A(_abc_41234_new_n1617_), .B(_abc_41234_new_n1649_), .C(_abc_41234_new_n2832_), .Y(_abc_41234_new_n2833_));
OAI21X1 OAI21X1_601 ( .A(_abc_41234_new_n2806_), .B(_abc_41234_new_n1616_), .C(_abc_41234_new_n2831_), .Y(_abc_41234_new_n2834_));
OAI21X1 OAI21X1_602 ( .A(_abc_41234_new_n1616_), .B(_abc_41234_new_n1617_), .C(_abc_41234_new_n2834_), .Y(_abc_41234_new_n2835_));
OAI21X1 OAI21X1_603 ( .A(pc_5_), .B(_abc_41234_new_n1729_), .C(_abc_41234_new_n1630_), .Y(_abc_41234_new_n2836_));
OAI21X1 OAI21X1_604 ( .A(_abc_41234_new_n1729_), .B(_abc_41234_new_n2836_), .C(_abc_41234_new_n2835_), .Y(_abc_41234_new_n2837_));
OAI21X1 OAI21X1_605 ( .A(_abc_41234_new_n546__bF_buf1), .B(_abc_41234_new_n723_), .C(_abc_41234_new_n2836_), .Y(_abc_41234_new_n2838_));
OAI21X1 OAI21X1_606 ( .A(regfil_1__5_), .B(_abc_41234_new_n1322_), .C(_abc_41234_new_n1639__bF_buf0), .Y(_abc_41234_new_n2841_));
OAI21X1 OAI21X1_607 ( .A(_abc_41234_new_n1645_), .B(_abc_41234_new_n2833_), .C(_abc_41234_new_n2843_), .Y(_abc_41234_new_n2844_));
OAI21X1 OAI21X1_608 ( .A(_abc_41234_new_n2824_), .B(_abc_41234_new_n2676_), .C(_abc_41234_new_n2845_), .Y(_abc_41234_new_n2846_));
OAI21X1 OAI21X1_609 ( .A(_abc_41234_new_n895_), .B(_abc_41234_new_n2515_), .C(_abc_41234_new_n2847_), .Y(_abc_41234_new_n2848_));
OAI21X1 OAI21X1_61 ( .A(_abc_41234_new_n881_), .B(_abc_41234_new_n880_), .C(_abc_41234_new_n893_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_4_));
OAI21X1 OAI21X1_610 ( .A(_abc_41234_new_n2756_), .B(_abc_41234_new_n2702_), .C(wdatahold_6_), .Y(_abc_41234_new_n2852_));
OAI21X1 OAI21X1_611 ( .A(intcyc_bF_buf3), .B(_abc_41234_new_n1631_), .C(_abc_41234_new_n1626_), .Y(_abc_41234_new_n2859_));
OAI21X1 OAI21X1_612 ( .A(regfil_3__6_), .B(_abc_41234_new_n529_), .C(_abc_41234_new_n536__bF_buf4), .Y(_abc_41234_new_n2862_));
OAI21X1 OAI21X1_613 ( .A(regfil_1__6_), .B(_abc_41234_new_n1322_), .C(_abc_41234_new_n2863_), .Y(_abc_41234_new_n2864_));
OAI21X1 OAI21X1_614 ( .A(_abc_41234_new_n1640_), .B(_abc_41234_new_n2864_), .C(_abc_41234_new_n2867_), .Y(_abc_41234_new_n2868_));
OAI21X1 OAI21X1_615 ( .A(_abc_41234_new_n1645_), .B(_abc_41234_new_n2855_), .C(_abc_41234_new_n2869_), .Y(_abc_41234_new_n2870_));
OAI21X1 OAI21X1_616 ( .A(_abc_41234_new_n967_), .B(_abc_41234_new_n537__bF_buf1), .C(_abc_41234_new_n2861_), .Y(_abc_41234_new_n2871_));
OAI21X1 OAI21X1_617 ( .A(_abc_41234_new_n1610_), .B(_abc_41234_new_n2871_), .C(_abc_41234_new_n2872_), .Y(_abc_41234_new_n2873_));
OAI21X1 OAI21X1_618 ( .A(_abc_41234_new_n2721_), .B(_abc_41234_new_n950_), .C(_abc_41234_new_n2873_), .Y(_abc_41234_new_n2874_));
OAI21X1 OAI21X1_619 ( .A(_abc_41234_new_n940_), .B(_abc_41234_new_n2515_), .C(_abc_41234_new_n2877_), .Y(_abc_41234_new_n2878_));
OAI21X1 OAI21X1_62 ( .A(_abc_41234_new_n896_), .B(_abc_41234_new_n722__bF_buf3), .C(_abc_41234_new_n897_), .Y(_abc_41234_new_n898_));
OAI21X1 OAI21X1_620 ( .A(_abc_41234_new_n2865_), .B(_abc_41234_new_n2857_), .C(_abc_41234_new_n2882_), .Y(_abc_41234_new_n2883_));
OAI21X1 OAI21X1_621 ( .A(_abc_41234_new_n1616_), .B(_abc_41234_new_n1619_), .C(_abc_41234_new_n2883_), .Y(_abc_41234_new_n2884_));
OAI21X1 OAI21X1_622 ( .A(pc_7_), .B(_abc_41234_new_n1729_), .C(_abc_41234_new_n1630_), .Y(_abc_41234_new_n2885_));
OAI21X1 OAI21X1_623 ( .A(_abc_41234_new_n2865_), .B(_abc_41234_new_n2853_), .C(_abc_41234_new_n2882_), .Y(_abc_41234_new_n2888_));
OAI21X1 OAI21X1_624 ( .A(_abc_41234_new_n1618_), .B(_abc_41234_new_n2853_), .C(_abc_41234_new_n2888_), .Y(_abc_41234_new_n2889_));
OAI21X1 OAI21X1_625 ( .A(_abc_41234_new_n2376_), .B(_abc_41234_new_n1105__bF_buf2), .C(_abc_41234_new_n2891_), .Y(_abc_41234_new_n2892_));
OAI21X1 OAI21X1_626 ( .A(regfil_1__7_), .B(_abc_41234_new_n1322_), .C(_abc_41234_new_n2892_), .Y(_abc_41234_new_n2893_));
OAI21X1 OAI21X1_627 ( .A(_abc_41234_new_n2881_), .B(_abc_41234_new_n1643__bF_buf3), .C(_abc_41234_new_n2895_), .Y(_abc_41234_new_n2896_));
OAI21X1 OAI21X1_628 ( .A(_abc_41234_new_n2886_), .B(_abc_41234_new_n2896_), .C(_abc_41234_new_n1046__bF_buf7), .Y(_abc_41234_new_n2897_));
OAI21X1 OAI21X1_629 ( .A(_abc_41234_new_n2899_), .B(_abc_41234_new_n2898_), .C(_abc_41234_new_n515__bF_buf0), .Y(_abc_41234_new_n2900_));
OAI21X1 OAI21X1_63 ( .A(_abc_41234_new_n908_), .B(_abc_41234_new_n905_), .C(opcode_2_), .Y(_abc_41234_new_n909_));
OAI21X1 OAI21X1_630 ( .A(wdatahold_7_), .B(_abc_41234_new_n2505_), .C(_abc_41234_new_n662_), .Y(_abc_41234_new_n2902_));
OAI21X1 OAI21X1_631 ( .A(_abc_41234_new_n2901_), .B(_abc_41234_new_n2902_), .C(_abc_41234_new_n2900_), .Y(_abc_41234_new_n2903_));
OAI21X1 OAI21X1_632 ( .A(_abc_41234_new_n691_), .B(_abc_41234_new_n2380_), .C(_abc_41234_new_n2906_), .Y(_abc_41234_new_n2907_));
OAI21X1 OAI21X1_633 ( .A(_abc_41234_new_n693_), .B(_abc_41234_new_n2512_), .C(_abc_41234_new_n2415__bF_buf0), .Y(_abc_41234_new_n2912_));
OAI21X1 OAI21X1_634 ( .A(_abc_41234_new_n2911_), .B(_abc_41234_new_n2912_), .C(_abc_41234_new_n516__bF_buf1), .Y(_abc_41234_new_n2913_));
OAI21X1 OAI21X1_635 ( .A(_abc_41234_new_n580_), .B(_abc_41234_new_n722__bF_buf0), .C(_abc_41234_new_n2486_), .Y(_abc_41234_new_n2915_));
OAI21X1 OAI21X1_636 ( .A(_abc_41234_new_n546__bF_buf0), .B(_abc_41234_new_n620__bF_buf0), .C(_abc_41234_new_n2916_), .Y(_abc_41234_new_n2917_));
OAI21X1 OAI21X1_637 ( .A(opcode_4_bF_buf4_), .B(regfil_1__0_), .C(_abc_41234_new_n2685_), .Y(_abc_41234_new_n2921_));
OAI21X1 OAI21X1_638 ( .A(raddrhold_0_), .B(_abc_41234_new_n669__bF_buf1), .C(_abc_41234_new_n2923_), .Y(_abc_41234_new_n2924_));
OAI21X1 OAI21X1_639 ( .A(_abc_41234_new_n2467_), .B(_abc_41234_new_n2921_), .C(_abc_41234_new_n2924_), .Y(_abc_41234_new_n2925_));
OAI21X1 OAI21X1_64 ( .A(opcode_2_), .B(_abc_41234_new_n902_), .C(_abc_41234_new_n909_), .Y(_abc_41234_new_n910_));
OAI21X1 OAI21X1_640 ( .A(pc_0_), .B(_abc_41234_new_n2918_), .C(_abc_41234_new_n2926_), .Y(_abc_41234_new_n2927_));
OAI21X1 OAI21X1_641 ( .A(raddrhold_0_), .B(_abc_41234_new_n2919__bF_buf2), .C(_abc_41234_new_n2927_), .Y(_abc_41234_new_n2928_));
OAI21X1 OAI21X1_642 ( .A(_abc_41234_new_n546__bF_buf5), .B(_abc_41234_new_n620__bF_buf5), .C(raddrhold_0_), .Y(_abc_41234_new_n2929_));
OAI21X1 OAI21X1_643 ( .A(_abc_41234_new_n1221_), .B(_abc_41234_new_n2185__bF_buf1), .C(_abc_41234_new_n2929_), .Y(_abc_41234_new_n2930_));
OAI21X1 OAI21X1_644 ( .A(_abc_41234_new_n2456_), .B(_abc_41234_new_n2931_), .C(_abc_41234_new_n1040__bF_buf1), .Y(_abc_41234_new_n2932_));
OAI21X1 OAI21X1_645 ( .A(opcode_5_bF_buf3_), .B(_abc_41234_new_n2245_), .C(_abc_41234_new_n2934_), .Y(_abc_41234_new_n2935_));
OAI21X1 OAI21X1_646 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n555_), .C(_abc_41234_new_n2939_), .Y(_abc_41234_new_n2940_));
OAI21X1 OAI21X1_647 ( .A(_abc_41234_new_n2948_), .B(_abc_41234_new_n2946_), .C(_abc_41234_new_n1046__bF_buf6), .Y(_abc_41234_new_n2949_));
OAI21X1 OAI21X1_648 ( .A(raddrhold_0_), .B(_abc_41234_new_n2953_), .C(_abc_41234_new_n662_), .Y(_abc_41234_new_n2954_));
OAI21X1 OAI21X1_649 ( .A(_abc_41234_new_n2952_), .B(_abc_41234_new_n2954_), .C(_abc_41234_new_n2949_), .Y(_abc_41234_new_n2955_));
OAI21X1 OAI21X1_65 ( .A(_abc_41234_new_n615_), .B(_abc_41234_new_n911_), .C(_abc_41234_new_n912_), .Y(_abc_41234_new_n913_));
OAI21X1 OAI21X1_650 ( .A(_abc_41234_new_n534__bF_buf5), .B(_abc_41234_new_n2928_), .C(_abc_41234_new_n2956_), .Y(_abc_41234_new_n2957_));
OAI21X1 OAI21X1_651 ( .A(opcode_4_bF_buf2_), .B(regfil_1__1_), .C(_abc_41234_new_n2963_), .Y(_abc_41234_new_n2964_));
OAI21X1 OAI21X1_652 ( .A(regfil_5__1_), .B(_abc_41234_new_n668__bF_buf2), .C(_abc_41234_new_n2966_), .Y(_abc_41234_new_n2967_));
OAI21X1 OAI21X1_653 ( .A(_abc_41234_new_n2467_), .B(_abc_41234_new_n2964_), .C(_abc_41234_new_n2967_), .Y(_abc_41234_new_n2968_));
OAI21X1 OAI21X1_654 ( .A(_abc_41234_new_n2706_), .B(_abc_41234_new_n2918_), .C(_abc_41234_new_n2969_), .Y(_abc_41234_new_n2970_));
OAI21X1 OAI21X1_655 ( .A(raddrhold_1_), .B(_abc_41234_new_n2919__bF_buf1), .C(_abc_41234_new_n2970_), .Y(_abc_41234_new_n2971_));
OAI21X1 OAI21X1_656 ( .A(_abc_41234_new_n2974_), .B(_abc_41234_new_n2972_), .C(_abc_41234_new_n1046__bF_buf5), .Y(_abc_41234_new_n2975_));
OAI21X1 OAI21X1_657 ( .A(_abc_41234_new_n668__bF_buf1), .B(_abc_41234_new_n2185__bF_buf0), .C(_abc_41234_new_n662_), .Y(_abc_41234_new_n2976_));
OAI21X1 OAI21X1_658 ( .A(_abc_41234_new_n546__bF_buf4), .B(_abc_41234_new_n620__bF_buf4), .C(_abc_41234_new_n2965_), .Y(_abc_41234_new_n2978_));
OAI21X1 OAI21X1_659 ( .A(regfil_5__1_), .B(_abc_41234_new_n2185__bF_buf5), .C(_abc_41234_new_n2978_), .Y(_abc_41234_new_n2979_));
OAI21X1 OAI21X1_66 ( .A(_abc_41234_new_n866_), .B(_abc_41234_new_n870_), .C(regfil_0__5_), .Y(_abc_41234_new_n916_));
OAI21X1 OAI21X1_660 ( .A(_abc_41234_new_n534__bF_buf4), .B(_abc_41234_new_n2971_), .C(_abc_41234_new_n2983_), .Y(_abc_41234_new_n2984_));
OAI21X1 OAI21X1_661 ( .A(reset_bF_buf3), .B(_abc_41234_new_n2985_), .C(_abc_41234_new_n2991_), .Y(_0raddrhold_15_0__1_));
OAI21X1 OAI21X1_662 ( .A(_abc_41234_new_n2207__bF_buf1), .B(_abc_41234_new_n2993_), .C(_abc_41234_new_n2919__bF_buf0), .Y(_abc_41234_new_n2994_));
OAI21X1 OAI21X1_663 ( .A(opcode_4_bF_buf1_), .B(regfil_1__2_), .C(_abc_41234_new_n2740_), .Y(_abc_41234_new_n2998_));
OAI21X1 OAI21X1_664 ( .A(_abc_41234_new_n2995_), .B(_abc_41234_new_n2918_), .C(_abc_41234_new_n3000_), .Y(_abc_41234_new_n3001_));
OAI21X1 OAI21X1_665 ( .A(_abc_41234_new_n546__bF_buf3), .B(_abc_41234_new_n620__bF_buf3), .C(_abc_41234_new_n3003_), .Y(_abc_41234_new_n3004_));
OAI21X1 OAI21X1_666 ( .A(regfil_5__2_), .B(_abc_41234_new_n2185__bF_buf4), .C(_abc_41234_new_n3004_), .Y(_abc_41234_new_n3005_));
OAI21X1 OAI21X1_667 ( .A(_abc_41234_new_n2951__bF_buf0), .B(_abc_41234_new_n3006_), .C(_abc_41234_new_n3007_), .Y(_abc_41234_new_n3008_));
OAI21X1 OAI21X1_668 ( .A(_abc_41234_new_n534__bF_buf3), .B(_abc_41234_new_n3002_), .C(_abc_41234_new_n3008_), .Y(_abc_41234_new_n3009_));
OAI21X1 OAI21X1_669 ( .A(_abc_41234_new_n3011_), .B(_abc_41234_new_n3010_), .C(_abc_41234_new_n1046__bF_buf4), .Y(_abc_41234_new_n3012_));
OAI21X1 OAI21X1_67 ( .A(regfil_0__4_), .B(_abc_41234_new_n806_), .C(regfil_0__5_), .Y(_abc_41234_new_n920_));
OAI21X1 OAI21X1_670 ( .A(_abc_41234_new_n2190__bF_buf3), .B(_abc_41234_new_n3005_), .C(_abc_41234_new_n3012_), .Y(_abc_41234_new_n3013_));
OAI21X1 OAI21X1_671 ( .A(_abc_41234_new_n3009_), .B(_abc_41234_new_n3013_), .C(_abc_41234_new_n660__bF_buf3), .Y(_abc_41234_new_n3014_));
OAI21X1 OAI21X1_672 ( .A(reset_bF_buf2), .B(_abc_41234_new_n3016_), .C(_abc_41234_new_n3021_), .Y(_0raddrhold_15_0__2_));
OAI21X1 OAI21X1_673 ( .A(raddrhold_3_), .B(_abc_41234_new_n3019_), .C(_abc_41234_new_n2911_), .Y(_abc_41234_new_n3025_));
OAI21X1 OAI21X1_674 ( .A(_abc_41234_new_n2207__bF_buf3), .B(_abc_41234_new_n3027_), .C(_abc_41234_new_n2919__bF_buf3), .Y(_abc_41234_new_n3028_));
OAI21X1 OAI21X1_675 ( .A(opcode_4_bF_buf0_), .B(regfil_1__3_), .C(_abc_41234_new_n2779_), .Y(_abc_41234_new_n3030_));
OAI21X1 OAI21X1_676 ( .A(_abc_41234_new_n2774_), .B(_abc_41234_new_n2918_), .C(_abc_41234_new_n3032_), .Y(_abc_41234_new_n3033_));
OAI21X1 OAI21X1_677 ( .A(_abc_41234_new_n546__bF_buf2), .B(_abc_41234_new_n620__bF_buf2), .C(_abc_41234_new_n3023_), .Y(_abc_41234_new_n3035_));
OAI21X1 OAI21X1_678 ( .A(regfil_5__3_bF_buf3_), .B(_abc_41234_new_n2185__bF_buf3), .C(_abc_41234_new_n3035_), .Y(_abc_41234_new_n3036_));
OAI21X1 OAI21X1_679 ( .A(_abc_41234_new_n2951__bF_buf2), .B(_abc_41234_new_n3037_), .C(_abc_41234_new_n3038_), .Y(_abc_41234_new_n3039_));
OAI21X1 OAI21X1_68 ( .A(_abc_41234_new_n895_), .B(_abc_41234_new_n632_), .C(_abc_41234_new_n923_), .Y(_abc_41234_new_n924_));
OAI21X1 OAI21X1_680 ( .A(_abc_41234_new_n534__bF_buf2), .B(_abc_41234_new_n3034_), .C(_abc_41234_new_n3039_), .Y(_abc_41234_new_n3040_));
OAI21X1 OAI21X1_681 ( .A(_abc_41234_new_n3042_), .B(_abc_41234_new_n3041_), .C(_abc_41234_new_n1046__bF_buf3), .Y(_abc_41234_new_n3043_));
OAI21X1 OAI21X1_682 ( .A(_abc_41234_new_n2190__bF_buf2), .B(_abc_41234_new_n3036_), .C(_abc_41234_new_n3043_), .Y(_abc_41234_new_n3044_));
OAI21X1 OAI21X1_683 ( .A(_abc_41234_new_n3040_), .B(_abc_41234_new_n3044_), .C(_abc_41234_new_n660__bF_buf2), .Y(_abc_41234_new_n3045_));
OAI21X1 OAI21X1_684 ( .A(_abc_41234_new_n2654_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3045_), .Y(_abc_41234_new_n3046_));
OAI21X1 OAI21X1_685 ( .A(_abc_41234_new_n3026_), .B(_abc_41234_new_n3046_), .C(_abc_41234_new_n516__bF_buf5), .Y(_abc_41234_new_n3047_));
OAI21X1 OAI21X1_686 ( .A(_abc_41234_new_n3023_), .B(_abc_41234_new_n2914_), .C(_abc_41234_new_n3047_), .Y(_0raddrhold_15_0__3_));
OAI21X1 OAI21X1_687 ( .A(raddrhold_4_), .B(_abc_41234_new_n3024_), .C(_abc_41234_new_n2911_), .Y(_abc_41234_new_n3050_));
OAI21X1 OAI21X1_688 ( .A(_abc_41234_new_n2207__bF_buf1), .B(_abc_41234_new_n3052_), .C(_abc_41234_new_n2919__bF_buf2), .Y(_abc_41234_new_n3053_));
OAI21X1 OAI21X1_689 ( .A(opcode_4_bF_buf6_), .B(regfil_1__4_), .C(_abc_41234_new_n2811_), .Y(_abc_41234_new_n3055_));
OAI21X1 OAI21X1_69 ( .A(regfil_7__5_), .B(_abc_41234_new_n678_), .C(_abc_41234_new_n710_), .Y(_abc_41234_new_n926_));
OAI21X1 OAI21X1_690 ( .A(_abc_41234_new_n2802_), .B(_abc_41234_new_n2918_), .C(_abc_41234_new_n3057_), .Y(_abc_41234_new_n3058_));
OAI21X1 OAI21X1_691 ( .A(_abc_41234_new_n546__bF_buf1), .B(_abc_41234_new_n620__bF_buf1), .C(_abc_41234_new_n3049_), .Y(_abc_41234_new_n3060_));
OAI21X1 OAI21X1_692 ( .A(regfil_5__4_), .B(_abc_41234_new_n2185__bF_buf2), .C(_abc_41234_new_n3060_), .Y(_abc_41234_new_n3061_));
OAI21X1 OAI21X1_693 ( .A(_abc_41234_new_n2951__bF_buf0), .B(_abc_41234_new_n3062_), .C(_abc_41234_new_n3063_), .Y(_abc_41234_new_n3064_));
OAI21X1 OAI21X1_694 ( .A(_abc_41234_new_n534__bF_buf1), .B(_abc_41234_new_n3059_), .C(_abc_41234_new_n3064_), .Y(_abc_41234_new_n3065_));
OAI21X1 OAI21X1_695 ( .A(_abc_41234_new_n3067_), .B(_abc_41234_new_n3066_), .C(_abc_41234_new_n1046__bF_buf2), .Y(_abc_41234_new_n3068_));
OAI21X1 OAI21X1_696 ( .A(_abc_41234_new_n2190__bF_buf1), .B(_abc_41234_new_n3061_), .C(_abc_41234_new_n3068_), .Y(_abc_41234_new_n3069_));
OAI21X1 OAI21X1_697 ( .A(_abc_41234_new_n3065_), .B(_abc_41234_new_n3069_), .C(_abc_41234_new_n660__bF_buf1), .Y(_abc_41234_new_n3070_));
OAI21X1 OAI21X1_698 ( .A(_abc_41234_new_n2656_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3070_), .Y(_abc_41234_new_n3071_));
OAI21X1 OAI21X1_699 ( .A(_abc_41234_new_n3051_), .B(_abc_41234_new_n3071_), .C(_abc_41234_new_n516__bF_buf4), .Y(_abc_41234_new_n3072_));
OAI21X1 OAI21X1_7 ( .A(_abc_41234_new_n518_), .B(_abc_41234_new_n592_), .C(_abc_41234_new_n595_), .Y(_abc_41234_new_n596_));
OAI21X1 OAI21X1_70 ( .A(regfil_7__4_), .B(_abc_41234_new_n839_), .C(_abc_41234_new_n688_), .Y(_abc_41234_new_n929_));
OAI21X1 OAI21X1_700 ( .A(_abc_41234_new_n3049_), .B(_abc_41234_new_n2914_), .C(_abc_41234_new_n3072_), .Y(_0raddrhold_15_0__4_));
OAI21X1 OAI21X1_701 ( .A(_abc_41234_new_n2207__bF_buf3), .B(_abc_41234_new_n3079_), .C(_abc_41234_new_n2919__bF_buf1), .Y(_abc_41234_new_n3080_));
OAI21X1 OAI21X1_702 ( .A(opcode_4_bF_buf5_), .B(regfil_1__5_), .C(_abc_41234_new_n2839_), .Y(_abc_41234_new_n3082_));
OAI21X1 OAI21X1_703 ( .A(_abc_41234_new_n2833_), .B(_abc_41234_new_n2918_), .C(_abc_41234_new_n3084_), .Y(_abc_41234_new_n3085_));
OAI21X1 OAI21X1_704 ( .A(_abc_41234_new_n546__bF_buf0), .B(_abc_41234_new_n620__bF_buf0), .C(_abc_41234_new_n3074_), .Y(_abc_41234_new_n3087_));
OAI21X1 OAI21X1_705 ( .A(regfil_5__5_), .B(_abc_41234_new_n2185__bF_buf1), .C(_abc_41234_new_n3087_), .Y(_abc_41234_new_n3088_));
OAI21X1 OAI21X1_706 ( .A(_abc_41234_new_n2951__bF_buf2), .B(_abc_41234_new_n3089_), .C(_abc_41234_new_n3090_), .Y(_abc_41234_new_n3091_));
OAI21X1 OAI21X1_707 ( .A(_abc_41234_new_n534__bF_buf0), .B(_abc_41234_new_n3086_), .C(_abc_41234_new_n3091_), .Y(_abc_41234_new_n3092_));
OAI21X1 OAI21X1_708 ( .A(_abc_41234_new_n3094_), .B(_abc_41234_new_n3093_), .C(_abc_41234_new_n1046__bF_buf1), .Y(_abc_41234_new_n3095_));
OAI21X1 OAI21X1_709 ( .A(_abc_41234_new_n2190__bF_buf0), .B(_abc_41234_new_n3088_), .C(_abc_41234_new_n3095_), .Y(_abc_41234_new_n3096_));
OAI21X1 OAI21X1_71 ( .A(_abc_41234_new_n929_), .B(_abc_41234_new_n934_), .C(_abc_41234_new_n928_), .Y(_abc_41234_new_n935_));
OAI21X1 OAI21X1_710 ( .A(_abc_41234_new_n3092_), .B(_abc_41234_new_n3096_), .C(_abc_41234_new_n660__bF_buf0), .Y(_abc_41234_new_n3097_));
OAI21X1 OAI21X1_711 ( .A(_abc_41234_new_n2658_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3097_), .Y(_abc_41234_new_n3098_));
OAI21X1 OAI21X1_712 ( .A(regfil_5__6_bF_buf2_), .B(_abc_41234_new_n668__bF_buf1), .C(_abc_41234_new_n3102_), .Y(_abc_41234_new_n3103_));
OAI21X1 OAI21X1_713 ( .A(opcode_4_bF_buf3_), .B(regfil_1__6_), .C(_abc_41234_new_n3104_), .Y(_abc_41234_new_n3105_));
OAI21X1 OAI21X1_714 ( .A(raddrhold_6_), .B(_abc_41234_new_n2919__bF_buf3), .C(_abc_41234_new_n3108_), .Y(_abc_41234_new_n3109_));
OAI21X1 OAI21X1_715 ( .A(_abc_41234_new_n3111_), .B(_abc_41234_new_n3110_), .C(_abc_41234_new_n1046__bF_buf0), .Y(_abc_41234_new_n3112_));
OAI21X1 OAI21X1_716 ( .A(_abc_41234_new_n546__bF_buf5), .B(_abc_41234_new_n620__bF_buf5), .C(_abc_41234_new_n3101_), .Y(_abc_41234_new_n3113_));
OAI21X1 OAI21X1_717 ( .A(regfil_5__6_bF_buf1_), .B(_abc_41234_new_n2185__bF_buf0), .C(_abc_41234_new_n3113_), .Y(_abc_41234_new_n3114_));
OAI21X1 OAI21X1_718 ( .A(_abc_41234_new_n534__bF_buf5), .B(_abc_41234_new_n3109_), .C(_abc_41234_new_n3118_), .Y(_abc_41234_new_n3119_));
OAI21X1 OAI21X1_719 ( .A(_abc_41234_new_n3101_), .B(_abc_41234_new_n3076_), .C(_abc_41234_new_n3120_), .Y(_abc_41234_new_n3121_));
OAI21X1 OAI21X1_72 ( .A(regfil_7__5_), .B(_abc_41234_new_n702_), .C(_abc_41234_new_n936_), .Y(_abc_41234_new_n937_));
OAI21X1 OAI21X1_720 ( .A(_abc_41234_new_n2371_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3121_), .Y(_abc_41234_new_n3122_));
OAI21X1 OAI21X1_721 ( .A(opcode_4_bF_buf2_), .B(regfil_1__7_), .C(_abc_41234_new_n2890_), .Y(_abc_41234_new_n3126_));
OAI21X1 OAI21X1_722 ( .A(raddrhold_7_), .B(_abc_41234_new_n669__bF_buf0), .C(_abc_41234_new_n3128_), .Y(_abc_41234_new_n3129_));
OAI21X1 OAI21X1_723 ( .A(_abc_41234_new_n2467_), .B(_abc_41234_new_n3126_), .C(_abc_41234_new_n3129_), .Y(_abc_41234_new_n3130_));
OAI21X1 OAI21X1_724 ( .A(_abc_41234_new_n2889_), .B(_abc_41234_new_n2918_), .C(_abc_41234_new_n3131_), .Y(_abc_41234_new_n3132_));
OAI21X1 OAI21X1_725 ( .A(raddrhold_7_), .B(_abc_41234_new_n2919__bF_buf2), .C(_abc_41234_new_n3132_), .Y(_abc_41234_new_n3133_));
OAI21X1 OAI21X1_726 ( .A(_abc_41234_new_n3135_), .B(_abc_41234_new_n3134_), .C(_abc_41234_new_n1046__bF_buf7), .Y(_abc_41234_new_n3136_));
OAI21X1 OAI21X1_727 ( .A(_abc_41234_new_n546__bF_buf4), .B(_abc_41234_new_n620__bF_buf4), .C(raddrhold_7_), .Y(_abc_41234_new_n3137_));
OAI21X1 OAI21X1_728 ( .A(_abc_41234_new_n996_), .B(_abc_41234_new_n2185__bF_buf5), .C(_abc_41234_new_n3137_), .Y(_abc_41234_new_n3138_));
OAI21X1 OAI21X1_729 ( .A(_abc_41234_new_n3125_), .B(_abc_41234_new_n2953_), .C(_abc_41234_new_n3139_), .Y(_abc_41234_new_n3140_));
OAI21X1 OAI21X1_73 ( .A(_abc_41234_new_n926_), .B(_abc_41234_new_n925_), .C(_abc_41234_new_n938_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_5_));
OAI21X1 OAI21X1_730 ( .A(_abc_41234_new_n534__bF_buf4), .B(_abc_41234_new_n3133_), .C(_abc_41234_new_n3142_), .Y(_abc_41234_new_n3143_));
OAI21X1 OAI21X1_731 ( .A(_abc_41234_new_n3101_), .B(_abc_41234_new_n3076_), .C(_abc_41234_new_n3125_), .Y(_abc_41234_new_n3146_));
OAI21X1 OAI21X1_732 ( .A(_abc_41234_new_n2377_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3147_), .Y(_abc_41234_new_n3148_));
OAI21X1 OAI21X1_733 ( .A(raddrhold_8_), .B(_abc_41234_new_n669__bF_buf3), .C(_abc_41234_new_n3153_), .Y(_abc_41234_new_n3154_));
OAI21X1 OAI21X1_734 ( .A(_abc_41234_new_n1656_), .B(_abc_41234_new_n2467_), .C(_abc_41234_new_n3154_), .Y(_abc_41234_new_n3155_));
OAI21X1 OAI21X1_735 ( .A(_abc_41234_new_n1653_), .B(_abc_41234_new_n2918_), .C(_abc_41234_new_n3156_), .Y(_abc_41234_new_n3157_));
OAI21X1 OAI21X1_736 ( .A(raddrhold_8_), .B(_abc_41234_new_n2919__bF_buf1), .C(_abc_41234_new_n3157_), .Y(_abc_41234_new_n3158_));
OAI21X1 OAI21X1_737 ( .A(_abc_41234_new_n3160_), .B(_abc_41234_new_n3159_), .C(_abc_41234_new_n1046__bF_buf6), .Y(_abc_41234_new_n3161_));
OAI21X1 OAI21X1_738 ( .A(_abc_41234_new_n546__bF_buf3), .B(_abc_41234_new_n620__bF_buf3), .C(raddrhold_8_), .Y(_abc_41234_new_n3162_));
OAI21X1 OAI21X1_739 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n2185__bF_buf4), .C(_abc_41234_new_n3162_), .Y(_abc_41234_new_n3163_));
OAI21X1 OAI21X1_74 ( .A(_abc_41234_new_n945_), .B(_abc_41234_new_n947_), .C(_abc_41234_new_n546__bF_buf0), .Y(_abc_41234_new_n948_));
OAI21X1 OAI21X1_740 ( .A(_abc_41234_new_n3151_), .B(_abc_41234_new_n2953_), .C(_abc_41234_new_n3164_), .Y(_abc_41234_new_n3165_));
OAI21X1 OAI21X1_741 ( .A(_abc_41234_new_n534__bF_buf3), .B(_abc_41234_new_n3158_), .C(_abc_41234_new_n3167_), .Y(_abc_41234_new_n3168_));
OAI21X1 OAI21X1_742 ( .A(_abc_41234_new_n3125_), .B(_abc_41234_new_n3144_), .C(_abc_41234_new_n3151_), .Y(_abc_41234_new_n3170_));
OAI21X1 OAI21X1_743 ( .A(_abc_41234_new_n565_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3171_), .Y(_abc_41234_new_n3172_));
OAI21X1 OAI21X1_744 ( .A(_abc_41234_new_n3151_), .B(_abc_41234_new_n3145_), .C(_abc_41234_new_n3175_), .Y(_abc_41234_new_n3176_));
OAI21X1 OAI21X1_745 ( .A(raddrhold_9_), .B(_abc_41234_new_n669__bF_buf2), .C(_abc_41234_new_n3180_), .Y(_abc_41234_new_n3181_));
OAI21X1 OAI21X1_746 ( .A(raddrhold_9_), .B(_abc_41234_new_n2919__bF_buf3), .C(_abc_41234_new_n3183_), .Y(_abc_41234_new_n3184_));
OAI21X1 OAI21X1_747 ( .A(_abc_41234_new_n546__bF_buf2), .B(_abc_41234_new_n620__bF_buf2), .C(_abc_41234_new_n3175_), .Y(_abc_41234_new_n3185_));
OAI21X1 OAI21X1_748 ( .A(regfil_4__1_bF_buf1_), .B(_abc_41234_new_n2185__bF_buf3), .C(_abc_41234_new_n3185_), .Y(_abc_41234_new_n3186_));
OAI21X1 OAI21X1_749 ( .A(_abc_41234_new_n2951__bF_buf0), .B(_abc_41234_new_n3187_), .C(_abc_41234_new_n3188_), .Y(_abc_41234_new_n3189_));
OAI21X1 OAI21X1_75 ( .A(_abc_41234_new_n546__bF_buf5), .B(_abc_41234_new_n943_), .C(_abc_41234_new_n948_), .Y(_abc_41234_new_n949_));
OAI21X1 OAI21X1_750 ( .A(_abc_41234_new_n534__bF_buf2), .B(_abc_41234_new_n3184_), .C(_abc_41234_new_n3189_), .Y(_abc_41234_new_n3190_));
OAI21X1 OAI21X1_751 ( .A(_abc_41234_new_n2473_), .B(_abc_41234_new_n2943_), .C(_abc_41234_new_n1680_), .Y(_abc_41234_new_n3192_));
OAI21X1 OAI21X1_752 ( .A(_abc_41234_new_n1251_), .B(_abc_41234_new_n2942__bF_buf1), .C(_abc_41234_new_n3192_), .Y(_abc_41234_new_n3193_));
OAI21X1 OAI21X1_753 ( .A(_abc_41234_new_n3193_), .B(_abc_41234_new_n3191_), .C(_abc_41234_new_n1046__bF_buf5), .Y(_abc_41234_new_n3194_));
OAI21X1 OAI21X1_754 ( .A(_abc_41234_new_n2190__bF_buf2), .B(_abc_41234_new_n3186_), .C(_abc_41234_new_n3194_), .Y(_abc_41234_new_n3195_));
OAI21X1 OAI21X1_755 ( .A(_abc_41234_new_n3190_), .B(_abc_41234_new_n3195_), .C(_abc_41234_new_n660__bF_buf4), .Y(_abc_41234_new_n3196_));
OAI21X1 OAI21X1_756 ( .A(_abc_41234_new_n718_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3196_), .Y(_abc_41234_new_n3197_));
OAI21X1 OAI21X1_757 ( .A(_abc_41234_new_n2473_), .B(_abc_41234_new_n2943_), .C(_abc_41234_new_n1716_), .Y(_abc_41234_new_n3202_));
OAI21X1 OAI21X1_758 ( .A(_abc_41234_new_n1358_), .B(_abc_41234_new_n2942__bF_buf0), .C(_abc_41234_new_n3202_), .Y(_abc_41234_new_n3203_));
OAI21X1 OAI21X1_759 ( .A(_abc_41234_new_n3203_), .B(_abc_41234_new_n3201_), .C(_abc_41234_new_n1046__bF_buf4), .Y(_abc_41234_new_n3204_));
OAI21X1 OAI21X1_76 ( .A(_abc_41234_new_n615_), .B(_abc_41234_new_n950_), .C(_abc_41234_new_n951_), .Y(_abc_41234_new_n952_));
OAI21X1 OAI21X1_760 ( .A(raddrhold_10_), .B(_abc_41234_new_n669__bF_buf1), .C(_abc_41234_new_n3206_), .Y(_abc_41234_new_n3207_));
OAI21X1 OAI21X1_761 ( .A(_abc_41234_new_n546__bF_buf1), .B(_abc_41234_new_n620__bF_buf1), .C(_abc_41234_new_n3200_), .Y(_abc_41234_new_n3212_));
OAI21X1 OAI21X1_762 ( .A(regfil_4__2_bF_buf1_), .B(_abc_41234_new_n2185__bF_buf2), .C(_abc_41234_new_n3212_), .Y(_abc_41234_new_n3213_));
OAI21X1 OAI21X1_763 ( .A(_abc_41234_new_n2976_), .B(_abc_41234_new_n3213_), .C(_abc_41234_new_n3215_), .Y(_abc_41234_new_n3216_));
OAI21X1 OAI21X1_764 ( .A(raddrhold_11_), .B(_abc_41234_new_n669__bF_buf0), .C(_abc_41234_new_n2174_), .Y(_abc_41234_new_n3227_));
OAI21X1 OAI21X1_765 ( .A(_abc_41234_new_n3226_), .B(_abc_41234_new_n3227_), .C(_abc_41234_new_n3229_), .Y(_abc_41234_new_n3230_));
OAI21X1 OAI21X1_766 ( .A(_abc_41234_new_n546__bF_buf0), .B(_abc_41234_new_n620__bF_buf0), .C(raddrhold_11_), .Y(_abc_41234_new_n3232_));
OAI21X1 OAI21X1_767 ( .A(_abc_41234_new_n819_), .B(_abc_41234_new_n2185__bF_buf1), .C(_abc_41234_new_n3232_), .Y(_abc_41234_new_n3233_));
OAI21X1 OAI21X1_768 ( .A(opcode_6_), .B(_abc_41234_new_n1045_), .C(_abc_41234_new_n2976_), .Y(_abc_41234_new_n3234_));
OAI21X1 OAI21X1_769 ( .A(_abc_41234_new_n2473_), .B(_abc_41234_new_n2943_), .C(_abc_41234_new_n1734_), .Y(_abc_41234_new_n3236_));
OAI21X1 OAI21X1_77 ( .A(_abc_41234_new_n953_), .B(_abc_41234_new_n870_), .C(regfil_0__6_), .Y(_abc_41234_new_n956_));
OAI21X1 OAI21X1_770 ( .A(_abc_41234_new_n1362_), .B(_abc_41234_new_n2942__bF_buf3), .C(_abc_41234_new_n3236_), .Y(_abc_41234_new_n3237_));
OAI21X1 OAI21X1_771 ( .A(_abc_41234_new_n534__bF_buf5), .B(_abc_41234_new_n2919__bF_buf1), .C(_abc_41234_new_n2953_), .Y(_abc_41234_new_n3240_));
OAI21X1 OAI21X1_772 ( .A(_abc_41234_new_n3240_), .B(_abc_41234_new_n3239_), .C(raddrhold_11_), .Y(_abc_41234_new_n3241_));
OAI21X1 OAI21X1_773 ( .A(_abc_41234_new_n3225_), .B(_abc_41234_new_n3220_), .C(_abc_41234_new_n2911_), .Y(_abc_41234_new_n3244_));
OAI21X1 OAI21X1_774 ( .A(_abc_41234_new_n2918_), .B(_abc_41234_new_n1755_), .C(_abc_41234_new_n3252_), .Y(_abc_41234_new_n3253_));
OAI21X1 OAI21X1_775 ( .A(_abc_41234_new_n3254_), .B(_abc_41234_new_n3253_), .C(_abc_41234_new_n515__bF_buf6), .Y(_abc_41234_new_n3255_));
OAI21X1 OAI21X1_776 ( .A(_abc_41234_new_n546__bF_buf5), .B(_abc_41234_new_n620__bF_buf5), .C(raddrhold_12_), .Y(_abc_41234_new_n3258_));
OAI21X1 OAI21X1_777 ( .A(_abc_41234_new_n849_), .B(_abc_41234_new_n2185__bF_buf0), .C(_abc_41234_new_n3258_), .Y(_abc_41234_new_n3259_));
OAI21X1 OAI21X1_778 ( .A(_abc_41234_new_n1047__bF_buf4), .B(_abc_41234_new_n2945_), .C(_abc_41234_new_n2953_), .Y(_abc_41234_new_n3260_));
OAI21X1 OAI21X1_779 ( .A(raddrhold_13_), .B(_abc_41234_new_n669__bF_buf2), .C(_abc_41234_new_n2174_), .Y(_abc_41234_new_n3276_));
OAI21X1 OAI21X1_78 ( .A(_abc_41234_new_n940_), .B(_abc_41234_new_n632_), .C(_abc_41234_new_n962_), .Y(_abc_41234_new_n963_));
OAI21X1 OAI21X1_780 ( .A(_abc_41234_new_n3277_), .B(_abc_41234_new_n3274_), .C(_abc_41234_new_n3231_), .Y(_abc_41234_new_n3278_));
OAI21X1 OAI21X1_781 ( .A(_abc_41234_new_n546__bF_buf4), .B(_abc_41234_new_n620__bF_buf4), .C(_abc_41234_new_n3272_), .Y(_abc_41234_new_n3284_));
OAI21X1 OAI21X1_782 ( .A(regfil_4__5_), .B(_abc_41234_new_n2185__bF_buf5), .C(_abc_41234_new_n3284_), .Y(_abc_41234_new_n3285_));
OAI21X1 OAI21X1_783 ( .A(raddrhold_14_), .B(_abc_41234_new_n669__bF_buf1), .C(_abc_41234_new_n2174_), .Y(_abc_41234_new_n3296_));
OAI21X1 OAI21X1_784 ( .A(_abc_41234_new_n2918_), .B(_abc_41234_new_n1804_), .C(_abc_41234_new_n3298_), .Y(_abc_41234_new_n3299_));
OAI21X1 OAI21X1_785 ( .A(_abc_41234_new_n3303_), .B(_abc_41234_new_n3302_), .C(_abc_41234_new_n1046__bF_buf0), .Y(_abc_41234_new_n3304_));
OAI21X1 OAI21X1_786 ( .A(_abc_41234_new_n546__bF_buf3), .B(_abc_41234_new_n620__bF_buf3), .C(raddrhold_14_), .Y(_abc_41234_new_n3305_));
OAI21X1 OAI21X1_787 ( .A(_abc_41234_new_n1509_), .B(_abc_41234_new_n2185__bF_buf4), .C(_abc_41234_new_n3305_), .Y(_abc_41234_new_n3306_));
OAI21X1 OAI21X1_788 ( .A(_abc_41234_new_n3310_), .B(_abc_41234_new_n3311_), .C(_abc_41234_new_n2911_), .Y(_abc_41234_new_n3312_));
OAI21X1 OAI21X1_789 ( .A(_abc_41234_new_n940_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3312_), .Y(_abc_41234_new_n3313_));
OAI21X1 OAI21X1_79 ( .A(regfil_7__6_), .B(_abc_41234_new_n678_), .C(_abc_41234_new_n710_), .Y(_abc_41234_new_n965_));
OAI21X1 OAI21X1_790 ( .A(raddrhold_15_), .B(_abc_41234_new_n669__bF_buf0), .C(_abc_41234_new_n3319_), .Y(_abc_41234_new_n3320_));
OAI21X1 OAI21X1_791 ( .A(_abc_41234_new_n1836_), .B(_abc_41234_new_n2467_), .C(_abc_41234_new_n3320_), .Y(_abc_41234_new_n3321_));
OAI21X1 OAI21X1_792 ( .A(_abc_41234_new_n3322_), .B(_abc_41234_new_n3317_), .C(_abc_41234_new_n3323_), .Y(_abc_41234_new_n3324_));
OAI21X1 OAI21X1_793 ( .A(_abc_41234_new_n3326_), .B(_abc_41234_new_n3325_), .C(_abc_41234_new_n1046__bF_buf7), .Y(_abc_41234_new_n3327_));
OAI21X1 OAI21X1_794 ( .A(_abc_41234_new_n546__bF_buf2), .B(_abc_41234_new_n620__bF_buf2), .C(raddrhold_15_), .Y(_abc_41234_new_n3328_));
OAI21X1 OAI21X1_795 ( .A(_abc_41234_new_n997_), .B(_abc_41234_new_n2185__bF_buf3), .C(_abc_41234_new_n3328_), .Y(_abc_41234_new_n3329_));
OAI21X1 OAI21X1_796 ( .A(_abc_41234_new_n2672_), .B(_abc_41234_new_n2520_), .C(_abc_41234_new_n516__bF_buf3), .Y(_abc_41234_new_n3338_));
OAI21X1 OAI21X1_797 ( .A(waddrhold_0_), .B(_abc_41234_new_n1643__bF_buf1), .C(_abc_41234_new_n3340_), .Y(_abc_41234_new_n3341_));
OAI21X1 OAI21X1_798 ( .A(_abc_41234_new_n546__bF_buf1), .B(_abc_41234_new_n620__bF_buf1), .C(_abc_41234_new_n515__bF_buf5), .Y(_abc_41234_new_n3342_));
OAI21X1 OAI21X1_799 ( .A(_abc_41234_new_n3342_), .B(_abc_41234_new_n2497_), .C(_abc_41234_new_n2950_), .Y(_abc_41234_new_n3343_));
OAI21X1 OAI21X1_8 ( .A(_abc_41234_new_n525__bF_buf3), .B(_abc_41234_new_n582_), .C(_abc_41234_new_n600_), .Y(_abc_41234_new_n601_));
OAI21X1 OAI21X1_80 ( .A(_abc_41234_new_n906_), .B(_abc_41234_new_n839_), .C(_abc_41234_new_n972_), .Y(_abc_41234_new_n973_));
OAI21X1 OAI21X1_800 ( .A(_abc_41234_new_n546__bF_buf0), .B(_abc_41234_new_n620__bF_buf0), .C(_abc_41234_new_n662_), .Y(_abc_41234_new_n3346_));
OAI21X1 OAI21X1_801 ( .A(_abc_41234_new_n534__bF_buf0), .B(_abc_41234_new_n2185__bF_buf2), .C(_abc_41234_new_n3346_), .Y(_abc_41234_new_n3347_));
OAI21X1 OAI21X1_802 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3344_), .C(_abc_41234_new_n3348_), .Y(_abc_41234_new_n3349_));
OAI21X1 OAI21X1_803 ( .A(_abc_41234_new_n1047__bF_buf2), .B(_abc_41234_new_n3341_), .C(_abc_41234_new_n3350_), .Y(_abc_41234_new_n3351_));
OAI21X1 OAI21X1_804 ( .A(_abc_41234_new_n1221_), .B(_abc_41234_new_n2694_), .C(_abc_41234_new_n3354_), .Y(_abc_41234_new_n3355_));
OAI21X1 OAI21X1_805 ( .A(_abc_41234_new_n2973_), .B(_abc_41234_new_n1040__bF_buf0), .C(_abc_41234_new_n3360_), .Y(_abc_41234_new_n3361_));
OAI21X1 OAI21X1_806 ( .A(_abc_41234_new_n3362_), .B(_abc_41234_new_n3361_), .C(_abc_41234_new_n1046__bF_buf6), .Y(_abc_41234_new_n3363_));
OAI21X1 OAI21X1_807 ( .A(opcode_3_bF_buf1_), .B(_abc_41234_new_n1105__bF_buf1), .C(_abc_41234_new_n3358_), .Y(_abc_41234_new_n3367_));
OAI21X1 OAI21X1_808 ( .A(regfil_5__1_), .B(_abc_41234_new_n668__bF_buf2), .C(_abc_41234_new_n3367_), .Y(_abc_41234_new_n3368_));
OAI21X1 OAI21X1_809 ( .A(_abc_41234_new_n3368_), .B(_abc_41234_new_n3366_), .C(_abc_41234_new_n2190__bF_buf0), .Y(_abc_41234_new_n3369_));
OAI21X1 OAI21X1_81 ( .A(_abc_41234_new_n560_), .B(_abc_41234_new_n688_), .C(_abc_41234_new_n512_), .Y(_abc_41234_new_n974_));
OAI21X1 OAI21X1_810 ( .A(_abc_41234_new_n719_), .B(_abc_41234_new_n2694_), .C(_abc_41234_new_n3377_), .Y(_abc_41234_new_n3378_));
OAI21X1 OAI21X1_811 ( .A(_abc_41234_new_n1071_), .B(_abc_41234_new_n1040__bF_buf4), .C(_abc_41234_new_n1643__bF_buf5), .Y(_abc_41234_new_n3386_));
OAI21X1 OAI21X1_812 ( .A(waddrhold_2_), .B(_abc_41234_new_n1643__bF_buf4), .C(_abc_41234_new_n1046__bF_buf5), .Y(_abc_41234_new_n3388_));
OAI21X1 OAI21X1_813 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3389_), .C(_abc_41234_new_n3391_), .Y(_abc_41234_new_n3392_));
OAI21X1 OAI21X1_814 ( .A(_abc_41234_new_n3388_), .B(_abc_41234_new_n3387_), .C(_abc_41234_new_n3393_), .Y(_abc_41234_new_n3394_));
OAI21X1 OAI21X1_815 ( .A(_abc_41234_new_n3337_), .B(_abc_41234_new_n3358_), .C(_abc_41234_new_n3381_), .Y(_abc_41234_new_n3396_));
OAI21X1 OAI21X1_816 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n2694_), .C(_abc_41234_new_n3399_), .Y(_abc_41234_new_n3400_));
OAI21X1 OAI21X1_817 ( .A(_abc_41234_new_n1067_), .B(_abc_41234_new_n1040__bF_buf3), .C(_abc_41234_new_n1643__bF_buf3), .Y(_abc_41234_new_n3405_));
OAI21X1 OAI21X1_818 ( .A(waddrhold_3_), .B(_abc_41234_new_n1643__bF_buf2), .C(_abc_41234_new_n1046__bF_buf4), .Y(_abc_41234_new_n3407_));
OAI21X1 OAI21X1_819 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3408_), .C(_abc_41234_new_n3410_), .Y(_abc_41234_new_n3411_));
OAI21X1 OAI21X1_82 ( .A(_abc_41234_new_n974_), .B(_abc_41234_new_n973_), .C(_abc_41234_new_n966_), .Y(_abc_41234_new_n975_));
OAI21X1 OAI21X1_820 ( .A(_abc_41234_new_n3407_), .B(_abc_41234_new_n3406_), .C(_abc_41234_new_n3412_), .Y(_abc_41234_new_n3413_));
OAI21X1 OAI21X1_821 ( .A(_abc_41234_new_n818_), .B(_abc_41234_new_n2694_), .C(_abc_41234_new_n3418_), .Y(_abc_41234_new_n3419_));
OAI21X1 OAI21X1_822 ( .A(_abc_41234_new_n1090_), .B(_abc_41234_new_n1040__bF_buf2), .C(_abc_41234_new_n1643__bF_buf1), .Y(_abc_41234_new_n3428_));
OAI21X1 OAI21X1_823 ( .A(waddrhold_4_), .B(_abc_41234_new_n1643__bF_buf0), .C(_abc_41234_new_n1046__bF_buf3), .Y(_abc_41234_new_n3430_));
OAI21X1 OAI21X1_824 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3431_), .C(_abc_41234_new_n3433_), .Y(_abc_41234_new_n3434_));
OAI21X1 OAI21X1_825 ( .A(_abc_41234_new_n3430_), .B(_abc_41234_new_n3429_), .C(_abc_41234_new_n3435_), .Y(_abc_41234_new_n3436_));
OAI21X1 OAI21X1_826 ( .A(waddrhold_4_), .B(_abc_41234_new_n3415_), .C(_abc_41234_new_n2696__bF_buf4), .Y(_abc_41234_new_n3441_));
OAI21X1 OAI21X1_827 ( .A(_abc_41234_new_n3441_), .B(_abc_41234_new_n3440_), .C(_abc_41234_new_n3438_), .Y(_abc_41234_new_n3442_));
OAI21X1 OAI21X1_828 ( .A(sp_4_), .B(_abc_41234_new_n3423_), .C(sp_5_), .Y(_abc_41234_new_n3446_));
OAI21X1 OAI21X1_829 ( .A(_abc_41234_new_n1094_), .B(_abc_41234_new_n1040__bF_buf1), .C(_abc_41234_new_n1643__bF_buf5), .Y(_abc_41234_new_n3450_));
OAI21X1 OAI21X1_83 ( .A(_abc_41234_new_n976_), .B(_abc_41234_new_n977_), .C(_abc_41234_new_n703_), .Y(_abc_41234_new_n978_));
OAI21X1 OAI21X1_830 ( .A(waddrhold_5_), .B(_abc_41234_new_n1643__bF_buf4), .C(_abc_41234_new_n1046__bF_buf2), .Y(_abc_41234_new_n3452_));
OAI21X1 OAI21X1_831 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3453_), .C(_abc_41234_new_n3455_), .Y(_abc_41234_new_n3456_));
OAI21X1 OAI21X1_832 ( .A(_abc_41234_new_n3452_), .B(_abc_41234_new_n3451_), .C(_abc_41234_new_n3457_), .Y(_abc_41234_new_n3458_));
OAI21X1 OAI21X1_833 ( .A(waddrhold_5_), .B(_abc_41234_new_n3440_), .C(_abc_41234_new_n2696__bF_buf3), .Y(_abc_41234_new_n3462_));
OAI21X1 OAI21X1_834 ( .A(_abc_41234_new_n3461_), .B(_abc_41234_new_n3462_), .C(_abc_41234_new_n3460_), .Y(_abc_41234_new_n3463_));
OAI21X1 OAI21X1_835 ( .A(sp_5_), .B(_abc_41234_new_n3425_), .C(sp_6_), .Y(_abc_41234_new_n3468_));
OAI21X1 OAI21X1_836 ( .A(_abc_41234_new_n1085_), .B(_abc_41234_new_n1040__bF_buf0), .C(_abc_41234_new_n1643__bF_buf3), .Y(_abc_41234_new_n3470_));
OAI21X1 OAI21X1_837 ( .A(waddrhold_6_), .B(_abc_41234_new_n1643__bF_buf2), .C(_abc_41234_new_n1046__bF_buf1), .Y(_abc_41234_new_n3472_));
OAI21X1 OAI21X1_838 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3473_), .C(_abc_41234_new_n3475_), .Y(_abc_41234_new_n3476_));
OAI21X1 OAI21X1_839 ( .A(_abc_41234_new_n3472_), .B(_abc_41234_new_n3471_), .C(_abc_41234_new_n3477_), .Y(_abc_41234_new_n3478_));
OAI21X1 OAI21X1_84 ( .A(_abc_41234_new_n965_), .B(_abc_41234_new_n964_), .C(_abc_41234_new_n981_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_6_));
OAI21X1 OAI21X1_840 ( .A(waddrhold_6_), .B(_abc_41234_new_n3461_), .C(_abc_41234_new_n2696__bF_buf2), .Y(_abc_41234_new_n3483_));
OAI21X1 OAI21X1_841 ( .A(_abc_41234_new_n3483_), .B(_abc_41234_new_n3482_), .C(_abc_41234_new_n3480_), .Y(_abc_41234_new_n3484_));
OAI21X1 OAI21X1_842 ( .A(sp_6_), .B(_abc_41234_new_n3448_), .C(sp_7_), .Y(_abc_41234_new_n3488_));
OAI21X1 OAI21X1_843 ( .A(_abc_41234_new_n1080_), .B(_abc_41234_new_n1040__bF_buf4), .C(_abc_41234_new_n1643__bF_buf1), .Y(_abc_41234_new_n3491_));
OAI21X1 OAI21X1_844 ( .A(waddrhold_7_), .B(_abc_41234_new_n1643__bF_buf0), .C(_abc_41234_new_n1046__bF_buf0), .Y(_abc_41234_new_n3493_));
OAI21X1 OAI21X1_845 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3494_), .C(_abc_41234_new_n3496_), .Y(_abc_41234_new_n3497_));
OAI21X1 OAI21X1_846 ( .A(_abc_41234_new_n3493_), .B(_abc_41234_new_n3492_), .C(_abc_41234_new_n3498_), .Y(_abc_41234_new_n3499_));
OAI21X1 OAI21X1_847 ( .A(waddrhold_7_), .B(_abc_41234_new_n3482_), .C(_abc_41234_new_n2696__bF_buf1), .Y(_abc_41234_new_n3503_));
OAI21X1 OAI21X1_848 ( .A(_abc_41234_new_n3502_), .B(_abc_41234_new_n3503_), .C(_abc_41234_new_n3501_), .Y(_abc_41234_new_n3504_));
OAI21X1 OAI21X1_849 ( .A(_abc_41234_new_n1255_), .B(_abc_41234_new_n1040__bF_buf3), .C(_abc_41234_new_n1643__bF_buf5), .Y(_abc_41234_new_n3509_));
OAI21X1 OAI21X1_85 ( .A(_abc_41234_new_n944_), .B(_abc_41234_new_n954_), .C(_abc_41234_new_n983_), .Y(_abc_41234_new_n984_));
OAI21X1 OAI21X1_850 ( .A(waddrhold_8_), .B(_abc_41234_new_n1643__bF_buf4), .C(_abc_41234_new_n1046__bF_buf7), .Y(_abc_41234_new_n3511_));
OAI21X1 OAI21X1_851 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3512_), .C(_abc_41234_new_n3514_), .Y(_abc_41234_new_n3515_));
OAI21X1 OAI21X1_852 ( .A(_abc_41234_new_n3511_), .B(_abc_41234_new_n3510_), .C(_abc_41234_new_n3516_), .Y(_abc_41234_new_n3517_));
OAI21X1 OAI21X1_853 ( .A(waddrhold_8_), .B(_abc_41234_new_n3502_), .C(_abc_41234_new_n2696__bF_buf0), .Y(_abc_41234_new_n3522_));
OAI21X1 OAI21X1_854 ( .A(_abc_41234_new_n3522_), .B(_abc_41234_new_n3521_), .C(_abc_41234_new_n3519_), .Y(_abc_41234_new_n3523_));
OAI21X1 OAI21X1_855 ( .A(sp_8_), .B(_abc_41234_new_n3489_), .C(sp_9_), .Y(_abc_41234_new_n3527_));
OAI21X1 OAI21X1_856 ( .A(_abc_41234_new_n3489_), .B(_abc_41234_new_n3529_), .C(_abc_41234_new_n3527_), .Y(_abc_41234_new_n3530_));
OAI21X1 OAI21X1_857 ( .A(_abc_41234_new_n1251_), .B(_abc_41234_new_n1040__bF_buf2), .C(_abc_41234_new_n1643__bF_buf3), .Y(_abc_41234_new_n3531_));
OAI21X1 OAI21X1_858 ( .A(waddrhold_9_), .B(_abc_41234_new_n1643__bF_buf2), .C(_abc_41234_new_n1046__bF_buf6), .Y(_abc_41234_new_n3533_));
OAI21X1 OAI21X1_859 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3534_), .C(_abc_41234_new_n3536_), .Y(_abc_41234_new_n3537_));
OAI21X1 OAI21X1_86 ( .A(regfil_0__6_), .B(_abc_41234_new_n919_), .C(_abc_41234_new_n983_), .Y(_abc_41234_new_n989_));
OAI21X1 OAI21X1_860 ( .A(_abc_41234_new_n3533_), .B(_abc_41234_new_n3532_), .C(_abc_41234_new_n3538_), .Y(_abc_41234_new_n3539_));
OAI21X1 OAI21X1_861 ( .A(waddrhold_9_), .B(_abc_41234_new_n3521_), .C(_abc_41234_new_n2696__bF_buf4), .Y(_abc_41234_new_n3543_));
OAI21X1 OAI21X1_862 ( .A(_abc_41234_new_n3542_), .B(_abc_41234_new_n3543_), .C(_abc_41234_new_n3541_), .Y(_abc_41234_new_n3544_));
OAI21X1 OAI21X1_863 ( .A(_abc_41234_new_n3529_), .B(_abc_41234_new_n3489_), .C(sp_10_), .Y(_abc_41234_new_n3550_));
OAI21X1 OAI21X1_864 ( .A(_abc_41234_new_n1358_), .B(_abc_41234_new_n1040__bF_buf1), .C(_abc_41234_new_n1643__bF_buf1), .Y(_abc_41234_new_n3552_));
OAI21X1 OAI21X1_865 ( .A(waddrhold_10_), .B(_abc_41234_new_n1643__bF_buf0), .C(_abc_41234_new_n1046__bF_buf5), .Y(_abc_41234_new_n3554_));
OAI21X1 OAI21X1_866 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3555_), .C(_abc_41234_new_n3557_), .Y(_abc_41234_new_n3558_));
OAI21X1 OAI21X1_867 ( .A(_abc_41234_new_n3554_), .B(_abc_41234_new_n3553_), .C(_abc_41234_new_n3559_), .Y(_abc_41234_new_n3560_));
OAI21X1 OAI21X1_868 ( .A(waddrhold_10_), .B(_abc_41234_new_n3542_), .C(_abc_41234_new_n2696__bF_buf3), .Y(_abc_41234_new_n3565_));
OAI21X1 OAI21X1_869 ( .A(_abc_41234_new_n3565_), .B(_abc_41234_new_n3564_), .C(_abc_41234_new_n3562_), .Y(_abc_41234_new_n3566_));
OAI21X1 OAI21X1_87 ( .A(_abc_41234_new_n994_), .B(_abc_41234_new_n991_), .C(_abc_41234_new_n546__bF_buf4), .Y(_abc_41234_new_n995_));
OAI21X1 OAI21X1_870 ( .A(sp_10_), .B(_abc_41234_new_n3570_), .C(sp_11_), .Y(_abc_41234_new_n3571_));
OAI21X1 OAI21X1_871 ( .A(_abc_41234_new_n3489_), .B(_abc_41234_new_n3572_), .C(_abc_41234_new_n3571_), .Y(_abc_41234_new_n3573_));
OAI21X1 OAI21X1_872 ( .A(_abc_41234_new_n1362_), .B(_abc_41234_new_n1040__bF_buf0), .C(_abc_41234_new_n1643__bF_buf5), .Y(_abc_41234_new_n3574_));
OAI21X1 OAI21X1_873 ( .A(waddrhold_11_), .B(_abc_41234_new_n1643__bF_buf4), .C(_abc_41234_new_n1046__bF_buf4), .Y(_abc_41234_new_n3576_));
OAI21X1 OAI21X1_874 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3577_), .C(_abc_41234_new_n3579_), .Y(_abc_41234_new_n3580_));
OAI21X1 OAI21X1_875 ( .A(_abc_41234_new_n3576_), .B(_abc_41234_new_n3575_), .C(_abc_41234_new_n3581_), .Y(_abc_41234_new_n3582_));
OAI21X1 OAI21X1_876 ( .A(waddrhold_11_), .B(_abc_41234_new_n3564_), .C(_abc_41234_new_n2696__bF_buf2), .Y(_abc_41234_new_n3587_));
OAI21X1 OAI21X1_877 ( .A(_abc_41234_new_n3586_), .B(_abc_41234_new_n3587_), .C(_abc_41234_new_n3584_), .Y(_abc_41234_new_n3588_));
OAI21X1 OAI21X1_878 ( .A(_abc_41234_new_n3572_), .B(_abc_41234_new_n3489_), .C(sp_12_), .Y(_abc_41234_new_n3594_));
OAI21X1 OAI21X1_879 ( .A(_abc_41234_new_n1408_), .B(_abc_41234_new_n1040__bF_buf4), .C(_abc_41234_new_n1643__bF_buf3), .Y(_abc_41234_new_n3596_));
OAI21X1 OAI21X1_88 ( .A(_abc_41234_new_n1000_), .B(_abc_41234_new_n998_), .C(opcode_2_), .Y(_abc_41234_new_n1001_));
OAI21X1 OAI21X1_880 ( .A(waddrhold_12_), .B(_abc_41234_new_n1643__bF_buf2), .C(_abc_41234_new_n1046__bF_buf3), .Y(_abc_41234_new_n3598_));
OAI21X1 OAI21X1_881 ( .A(waddrhold_12_), .B(_abc_41234_new_n669__bF_buf3), .C(_abc_41234_new_n3250_), .Y(_abc_41234_new_n3599_));
OAI21X1 OAI21X1_882 ( .A(_abc_41234_new_n3366_), .B(_abc_41234_new_n3599_), .C(_abc_41234_new_n3601_), .Y(_abc_41234_new_n3602_));
OAI21X1 OAI21X1_883 ( .A(_abc_41234_new_n3598_), .B(_abc_41234_new_n3597_), .C(_abc_41234_new_n3603_), .Y(_abc_41234_new_n3604_));
OAI21X1 OAI21X1_884 ( .A(reset_bF_buf7), .B(_abc_41234_new_n3607_), .C(_abc_41234_new_n3612_), .Y(_0waddrhold_15_0__12_));
OAI21X1 OAI21X1_885 ( .A(sp_12_), .B(_abc_41234_new_n3615_), .C(sp_13_), .Y(_abc_41234_new_n3616_));
OAI21X1 OAI21X1_886 ( .A(_abc_41234_new_n3279_), .B(_abc_41234_new_n1040__bF_buf3), .C(_abc_41234_new_n1643__bF_buf1), .Y(_abc_41234_new_n3620_));
OAI21X1 OAI21X1_887 ( .A(waddrhold_13_), .B(_abc_41234_new_n1643__bF_buf0), .C(_abc_41234_new_n1046__bF_buf2), .Y(_abc_41234_new_n3622_));
OAI21X1 OAI21X1_888 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3623_), .C(_abc_41234_new_n3626_), .Y(_abc_41234_new_n3627_));
OAI21X1 OAI21X1_889 ( .A(_abc_41234_new_n3622_), .B(_abc_41234_new_n3621_), .C(_abc_41234_new_n3628_), .Y(_abc_41234_new_n3629_));
OAI21X1 OAI21X1_89 ( .A(regfil_7__7_), .B(_abc_41234_new_n678_), .C(_abc_41234_new_n710_), .Y(_abc_41234_new_n1012_));
OAI21X1 OAI21X1_890 ( .A(waddrhold_13_), .B(_abc_41234_new_n3632_), .C(_abc_41234_new_n3634_), .Y(_abc_41234_new_n3635_));
OAI21X1 OAI21X1_891 ( .A(reset_bF_buf6), .B(_abc_41234_new_n3631_), .C(_abc_41234_new_n3635_), .Y(_0waddrhold_15_0__13_));
OAI21X1 OAI21X1_892 ( .A(_abc_41234_new_n3639_), .B(_abc_41234_new_n3638_), .C(_abc_41234_new_n3359_), .Y(_abc_41234_new_n3640_));
OAI21X1 OAI21X1_893 ( .A(_abc_41234_new_n1524_), .B(_abc_41234_new_n1040__bF_buf2), .C(_abc_41234_new_n3640_), .Y(_abc_41234_new_n3641_));
OAI21X1 OAI21X1_894 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3643_), .C(_abc_41234_new_n3646_), .Y(_abc_41234_new_n3647_));
OAI21X1 OAI21X1_895 ( .A(_abc_41234_new_n1047__bF_buf1), .B(_abc_41234_new_n3642_), .C(_abc_41234_new_n3648_), .Y(_abc_41234_new_n3649_));
OAI21X1 OAI21X1_896 ( .A(sp_14_), .B(_abc_41234_new_n3618_), .C(sp_15_), .Y(_abc_41234_new_n3657_));
OAI21X1 OAI21X1_897 ( .A(_abc_41234_new_n1569_), .B(_abc_41234_new_n1040__bF_buf1), .C(_abc_41234_new_n1643__bF_buf5), .Y(_abc_41234_new_n3660_));
OAI21X1 OAI21X1_898 ( .A(_abc_41234_new_n3660_), .B(_abc_41234_new_n3659_), .C(_abc_41234_new_n3662_), .Y(_abc_41234_new_n3663_));
OAI21X1 OAI21X1_899 ( .A(_abc_41234_new_n2498_), .B(_abc_41234_new_n3664_), .C(_abc_41234_new_n3666_), .Y(_abc_41234_new_n3667_));
OAI21X1 OAI21X1_9 ( .A(_abc_41234_new_n606_), .B(_abc_41234_new_n609_), .C(_abc_41234_new_n614_), .Y(_abc_41234_new_n615_));
OAI21X1 OAI21X1_90 ( .A(_abc_41234_new_n1016_), .B(_abc_41234_new_n683_), .C(_abc_41234_new_n1017_), .Y(_abc_41234_new_n1018_));
OAI21X1 OAI21X1_900 ( .A(waddrhold_15_), .B(_abc_41234_new_n2190__bF_buf3), .C(_abc_41234_new_n660__bF_buf5), .Y(_abc_41234_new_n3669_));
OAI21X1 OAI21X1_901 ( .A(_abc_41234_new_n3656_), .B(_abc_41234_new_n3670_), .C(_abc_41234_new_n516__bF_buf2), .Y(_abc_41234_new_n3671_));
OAI21X1 OAI21X1_902 ( .A(_abc_41234_new_n3661_), .B(_abc_41234_new_n3653_), .C(_abc_41234_new_n3672_), .Y(_abc_41234_new_n3673_));
OAI21X1 OAI21X1_903 ( .A(_abc_41234_new_n609_), .B(_abc_41234_new_n1850_), .C(_abc_41234_new_n3610_), .Y(_abc_41234_new_n3676_));
OAI21X1 OAI21X1_904 ( .A(_abc_41234_new_n714_), .B(_abc_41234_new_n3676_), .C(_abc_41234_new_n3678_), .Y(_0datao_7_0__0_));
OAI21X1 OAI21X1_905 ( .A(_abc_41234_new_n2432_), .B(_abc_41234_new_n3676_), .C(_abc_41234_new_n3680_), .Y(_0datao_7_0__1_));
OAI21X1 OAI21X1_906 ( .A(_abc_41234_new_n2435_), .B(_abc_41234_new_n3676_), .C(_abc_41234_new_n3682_), .Y(_0datao_7_0__2_));
OAI21X1 OAI21X1_907 ( .A(_abc_41234_new_n2437_), .B(_abc_41234_new_n3676_), .C(_abc_41234_new_n3684_), .Y(_0datao_7_0__3_));
OAI21X1 OAI21X1_908 ( .A(_abc_41234_new_n890_), .B(_abc_41234_new_n3676_), .C(_abc_41234_new_n3686_), .Y(_0datao_7_0__4_));
OAI21X1 OAI21X1_909 ( .A(_abc_41234_new_n2441_), .B(_abc_41234_new_n3676_), .C(_abc_41234_new_n3688_), .Y(_0datao_7_0__5_));
OAI21X1 OAI21X1_91 ( .A(_abc_41234_new_n1013_), .B(_abc_41234_new_n1020_), .C(_abc_41234_new_n1019_), .Y(_abc_41234_new_n1021_));
OAI21X1 OAI21X1_910 ( .A(_abc_41234_new_n2443_), .B(_abc_41234_new_n3676_), .C(_abc_41234_new_n3690_), .Y(_0datao_7_0__6_));
OAI21X1 OAI21X1_911 ( .A(_abc_41234_new_n1016_), .B(_abc_41234_new_n3676_), .C(_abc_41234_new_n3692_), .Y(_0datao_7_0__7_));
OAI21X1 OAI21X1_912 ( .A(opcode_7_), .B(_abc_41234_new_n523__bF_buf1), .C(regd_0_), .Y(_abc_41234_new_n3694_));
OAI21X1 OAI21X1_913 ( .A(_abc_41234_new_n2185__bF_buf1), .B(_abc_41234_new_n2951__bF_buf0), .C(_abc_41234_new_n673_), .Y(_abc_41234_new_n3695_));
OAI21X1 OAI21X1_914 ( .A(_abc_41234_new_n555_), .B(_abc_41234_new_n663_), .C(_abc_41234_new_n2502_), .Y(_abc_41234_new_n3696_));
OAI21X1 OAI21X1_915 ( .A(_abc_41234_new_n523__bF_buf0), .B(_abc_41234_new_n3700_), .C(_abc_41234_new_n3694_), .Y(_0regd_2_0__0_));
OAI21X1 OAI21X1_916 ( .A(opcode_7_), .B(_abc_41234_new_n523__bF_buf4), .C(regd_1_), .Y(_abc_41234_new_n3702_));
OAI21X1 OAI21X1_917 ( .A(_abc_41234_new_n2185__bF_buf0), .B(_abc_41234_new_n2951__bF_buf3), .C(_abc_41234_new_n654_), .Y(_abc_41234_new_n3703_));
OAI21X1 OAI21X1_918 ( .A(_abc_41234_new_n523__bF_buf3), .B(_abc_41234_new_n3706_), .C(_abc_41234_new_n3702_), .Y(_0regd_2_0__1_));
OAI21X1 OAI21X1_919 ( .A(opcode_7_), .B(_abc_41234_new_n523__bF_buf2), .C(regd_2_), .Y(_abc_41234_new_n3708_));
OAI21X1 OAI21X1_92 ( .A(_abc_41234_new_n967_), .B(_abc_41234_new_n968_), .C(_abc_41234_new_n553_), .Y(_abc_41234_new_n1022_));
OAI21X1 OAI21X1_920 ( .A(_abc_41234_new_n2185__bF_buf5), .B(_abc_41234_new_n2951__bF_buf2), .C(_abc_41234_new_n649_), .Y(_abc_41234_new_n3709_));
OAI21X1 OAI21X1_921 ( .A(_abc_41234_new_n523__bF_buf1), .B(_abc_41234_new_n3712_), .C(_abc_41234_new_n3708_), .Y(_0regd_2_0__2_));
OAI21X1 OAI21X1_922 ( .A(regfil_5__0_), .B(_abc_41234_new_n3716_), .C(_abc_41234_new_n1055_), .Y(_abc_41234_new_n3717_));
OAI21X1 OAI21X1_923 ( .A(_abc_41234_new_n3715_), .B(_abc_41234_new_n3717_), .C(_abc_41234_new_n3728_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_0_));
OAI21X1 OAI21X1_924 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n748_), .C(_abc_41234_new_n3730_), .Y(_abc_41234_new_n3731_));
OAI21X1 OAI21X1_925 ( .A(_abc_41234_new_n3732_), .B(_abc_41234_new_n1219_), .C(_abc_41234_new_n1049__bF_buf4), .Y(_abc_41234_new_n3733_));
OAI21X1 OAI21X1_926 ( .A(_abc_41234_new_n3736_), .B(_abc_41234_new_n1109_), .C(_abc_41234_new_n1263_), .Y(_abc_41234_new_n3737_));
OAI21X1 OAI21X1_927 ( .A(_abc_41234_new_n1158_), .B(_abc_41234_new_n3740_), .C(_abc_41234_new_n1325_), .Y(_abc_41234_new_n3741_));
OAI21X1 OAI21X1_928 ( .A(_abc_41234_new_n3722_), .B(_abc_41234_new_n3739_), .C(_abc_41234_new_n1308_), .Y(_abc_41234_new_n3742_));
OAI21X1 OAI21X1_929 ( .A(_abc_41234_new_n1221_), .B(_abc_41234_new_n1304_), .C(_abc_41234_new_n3748_), .Y(_abc_41234_new_n3749_));
OAI21X1 OAI21X1_93 ( .A(_abc_41234_new_n969_), .B(_abc_41234_new_n552_), .C(regfil_7__7_), .Y(_abc_41234_new_n1024_));
OAI21X1 OAI21X1_930 ( .A(_abc_41234_new_n3732_), .B(_abc_41234_new_n1263_), .C(_abc_41234_new_n1219_), .Y(_abc_41234_new_n3751_));
OAI21X1 OAI21X1_931 ( .A(_abc_41234_new_n2651_), .B(_abc_41234_new_n1044_), .C(_abc_41234_new_n3754_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_1_));
OAI21X1 OAI21X1_932 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n791_), .C(_abc_41234_new_n1055_), .Y(_abc_41234_new_n3757_));
OAI21X1 OAI21X1_933 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n1207_), .C(_abc_41234_new_n1218_), .Y(_abc_41234_new_n3759_));
OAI21X1 OAI21X1_934 ( .A(_abc_41234_new_n1224_), .B(_abc_41234_new_n3761_), .C(_abc_41234_new_n1206_), .Y(_abc_41234_new_n3762_));
OAI21X1 OAI21X1_935 ( .A(_abc_41234_new_n3772_), .B(_abc_41234_new_n1308_), .C(_abc_41234_new_n1304_), .Y(_abc_41234_new_n3773_));
OAI21X1 OAI21X1_936 ( .A(_abc_41234_new_n1043_), .B(_abc_41234_new_n3775_), .C(_abc_41234_new_n3762_), .Y(_abc_41234_new_n3776_));
OAI21X1 OAI21X1_937 ( .A(_abc_41234_new_n3760_), .B(_abc_41234_new_n3776_), .C(_abc_41234_new_n1049__bF_buf2), .Y(_abc_41234_new_n3777_));
OAI21X1 OAI21X1_938 ( .A(_abc_41234_new_n3756_), .B(_abc_41234_new_n3757_), .C(_abc_41234_new_n3778_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_2_));
OAI21X1 OAI21X1_939 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n829_), .C(_abc_41234_new_n1055_), .Y(_abc_41234_new_n3780_));
OAI21X1 OAI21X1_94 ( .A(_abc_41234_new_n541_), .B(_abc_41234_new_n553_), .C(_abc_41234_new_n1024_), .Y(_abc_41234_new_n1025_));
OAI21X1 OAI21X1_940 ( .A(_abc_41234_new_n3785_), .B(_abc_41234_new_n1109_), .C(_abc_41234_new_n1263_), .Y(_abc_41234_new_n3786_));
OAI21X1 OAI21X1_941 ( .A(_abc_41234_new_n634_), .B(_abc_41234_new_n772_), .C(_abc_41234_new_n3767_), .Y(_abc_41234_new_n3787_));
OAI21X1 OAI21X1_942 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n768_), .C(_abc_41234_new_n3770_), .Y(_abc_41234_new_n3791_));
OAI21X1 OAI21X1_943 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n1304_), .C(_abc_41234_new_n3793_), .Y(_abc_41234_new_n3794_));
OAI21X1 OAI21X1_944 ( .A(_abc_41234_new_n3795_), .B(_abc_41234_new_n3796_), .C(_abc_41234_new_n1206_), .Y(_abc_41234_new_n3797_));
OAI21X1 OAI21X1_945 ( .A(_abc_41234_new_n3786_), .B(_abc_41234_new_n3794_), .C(_abc_41234_new_n3797_), .Y(_abc_41234_new_n3798_));
OAI21X1 OAI21X1_946 ( .A(regfil_3__3_), .B(_abc_41234_new_n1049__bF_buf1), .C(_abc_41234_new_n3799_), .Y(_abc_41234_new_n3800_));
OAI21X1 OAI21X1_947 ( .A(_abc_41234_new_n2654_), .B(_abc_41234_new_n1044_), .C(_abc_41234_new_n3800_), .Y(_abc_41234_new_n3801_));
OAI21X1 OAI21X1_948 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n879_), .C(_abc_41234_new_n1055_), .Y(_abc_41234_new_n3803_));
OAI21X1 OAI21X1_949 ( .A(_abc_41234_new_n1211_), .B(_abc_41234_new_n3805_), .C(_abc_41234_new_n1218_), .Y(_abc_41234_new_n3806_));
OAI21X1 OAI21X1_95 ( .A(_abc_41234_new_n1025_), .B(_abc_41234_new_n1023_), .C(_abc_41234_new_n1026_), .Y(_abc_41234_new_n1027_));
OAI21X1 OAI21X1_950 ( .A(_abc_41234_new_n818_), .B(_abc_41234_new_n1223_), .C(_abc_41234_new_n848_), .Y(_abc_41234_new_n3808_));
OAI21X1 OAI21X1_951 ( .A(regfil_5__3_bF_buf0_), .B(_abc_41234_new_n1304_), .C(_abc_41234_new_n3819_), .Y(_abc_41234_new_n3820_));
OAI21X1 OAI21X1_952 ( .A(_abc_41234_new_n2656_), .B(_abc_41234_new_n1044_), .C(_abc_41234_new_n3824_), .Y(_abc_41234_new_n3825_));
OAI21X1 OAI21X1_953 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n924_), .C(_abc_41234_new_n3827_), .Y(_abc_41234_new_n3828_));
OAI21X1 OAI21X1_954 ( .A(_abc_41234_new_n3830_), .B(_abc_41234_new_n1219_), .C(_abc_41234_new_n1049__bF_buf3), .Y(_abc_41234_new_n3831_));
OAI21X1 OAI21X1_955 ( .A(_abc_41234_new_n1109_), .B(_abc_41234_new_n3833_), .C(_abc_41234_new_n1263_), .Y(_abc_41234_new_n3834_));
OAI21X1 OAI21X1_956 ( .A(_abc_41234_new_n3811_), .B(_abc_41234_new_n3810_), .C(_abc_41234_new_n1136_), .Y(_abc_41234_new_n3835_));
OAI21X1 OAI21X1_957 ( .A(_abc_41234_new_n855_), .B(_abc_41234_new_n848_), .C(_abc_41234_new_n3816_), .Y(_abc_41234_new_n3837_));
OAI21X1 OAI21X1_958 ( .A(_abc_41234_new_n3838_), .B(_abc_41234_new_n3840_), .C(_abc_41234_new_n1308_), .Y(_abc_41234_new_n3841_));
OAI21X1 OAI21X1_959 ( .A(_abc_41234_new_n1308_), .B(_abc_41234_new_n3836_), .C(_abc_41234_new_n3841_), .Y(_abc_41234_new_n3842_));
OAI21X1 OAI21X1_96 ( .A(opcode_4_bF_buf6_), .B(_abc_41234_new_n680_), .C(_abc_41234_new_n533_), .Y(_abc_41234_new_n1028_));
OAI21X1 OAI21X1_960 ( .A(_abc_41234_new_n848_), .B(_abc_41234_new_n1304_), .C(_abc_41234_new_n3842_), .Y(_abc_41234_new_n3843_));
OAI21X1 OAI21X1_961 ( .A(_abc_41234_new_n3845_), .B(_abc_41234_new_n3846_), .C(_abc_41234_new_n1206_), .Y(_abc_41234_new_n3847_));
OAI21X1 OAI21X1_962 ( .A(_abc_41234_new_n525__bF_buf1), .B(_abc_41234_new_n1217_), .C(_abc_41234_new_n3847_), .Y(_abc_41234_new_n3848_));
OAI21X1 OAI21X1_963 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n963_), .C(_abc_41234_new_n3852_), .Y(_abc_41234_new_n3853_));
OAI21X1 OAI21X1_964 ( .A(_abc_41234_new_n1219_), .B(_abc_41234_new_n3855_), .C(_abc_41234_new_n1049__bF_buf1), .Y(_abc_41234_new_n3856_));
OAI21X1 OAI21X1_965 ( .A(_abc_41234_new_n3857_), .B(_abc_41234_new_n3858_), .C(_abc_41234_new_n1130_), .Y(_abc_41234_new_n3859_));
OAI21X1 OAI21X1_966 ( .A(_abc_41234_new_n1128_), .B(_abc_41234_new_n1129_), .C(_abc_41234_new_n3860_), .Y(_abc_41234_new_n3861_));
OAI21X1 OAI21X1_967 ( .A(_abc_41234_new_n3864_), .B(_abc_41234_new_n3866_), .C(_abc_41234_new_n1325_), .Y(_abc_41234_new_n3868_));
OAI21X1 OAI21X1_968 ( .A(_abc_41234_new_n3867_), .B(_abc_41234_new_n3868_), .C(_abc_41234_new_n1304_), .Y(_abc_41234_new_n3869_));
OAI21X1 OAI21X1_969 ( .A(_abc_41234_new_n1098_), .B(_abc_41234_new_n3871_), .C(_abc_41234_new_n1101_), .Y(_abc_41234_new_n3872_));
OAI21X1 OAI21X1_97 ( .A(_abc_41234_new_n1012_), .B(_abc_41234_new_n1011_), .C(_abc_41234_new_n1029_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_7_));
OAI21X1 OAI21X1_970 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n1229_), .C(_abc_41234_new_n1084_), .Y(_abc_41234_new_n3876_));
OAI21X1 OAI21X1_971 ( .A(_abc_41234_new_n1058_), .B(_abc_41234_new_n677_), .C(regfil_5__7_), .Y(_abc_41234_new_n3881_));
OAI21X1 OAI21X1_972 ( .A(_abc_41234_new_n3714_), .B(_abc_41234_new_n1558_), .C(_abc_41234_new_n3881_), .Y(_abc_41234_new_n3882_));
OAI21X1 OAI21X1_973 ( .A(regfil_3__7_), .B(_abc_41234_new_n1049__bF_buf4), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n3884_));
OAI21X1 OAI21X1_974 ( .A(regfil_5__6_bF_buf3_), .B(_abc_41234_new_n1212_), .C(regfil_5__7_), .Y(_abc_41234_new_n3885_));
OAI21X1 OAI21X1_975 ( .A(_abc_41234_new_n1219_), .B(_abc_41234_new_n3886_), .C(_abc_41234_new_n1049__bF_buf3), .Y(_abc_41234_new_n3887_));
OAI21X1 OAI21X1_976 ( .A(_abc_41234_new_n996_), .B(_abc_41234_new_n3875_), .C(_abc_41234_new_n1219_), .Y(_abc_41234_new_n3889_));
OAI21X1 OAI21X1_977 ( .A(_abc_41234_new_n3888_), .B(_abc_41234_new_n3889_), .C(_abc_41234_new_n1043_), .Y(_abc_41234_new_n3890_));
OAI21X1 OAI21X1_978 ( .A(_abc_41234_new_n1171_), .B(_abc_41234_new_n1172_), .C(_abc_41234_new_n3892_), .Y(_abc_41234_new_n3893_));
OAI21X1 OAI21X1_979 ( .A(_abc_41234_new_n1174_), .B(_abc_41234_new_n3891_), .C(_abc_41234_new_n1173_), .Y(_abc_41234_new_n3894_));
OAI21X1 OAI21X1_98 ( .A(_abc_41234_new_n1032_), .B(_abc_41234_new_n508_), .C(_abc_41234_new_n1034_), .Y(_abc_41234_new_n1035_));
OAI21X1 OAI21X1_980 ( .A(_abc_41234_new_n1084_), .B(_abc_41234_new_n1936_), .C(_abc_41234_new_n3859_), .Y(_abc_41234_new_n3896_));
OAI21X1 OAI21X1_981 ( .A(_abc_41234_new_n1152_), .B(_abc_41234_new_n3897_), .C(_abc_41234_new_n3895_), .Y(_abc_41234_new_n3898_));
OAI21X1 OAI21X1_982 ( .A(_abc_41234_new_n525__bF_buf0), .B(_abc_41234_new_n3899_), .C(_abc_41234_new_n1109_), .Y(_abc_41234_new_n3900_));
OAI21X1 OAI21X1_983 ( .A(_abc_41234_new_n1084_), .B(_abc_41234_new_n1085_), .C(_abc_41234_new_n3902_), .Y(_abc_41234_new_n3903_));
OAI21X1 OAI21X1_984 ( .A(_abc_41234_new_n3901_), .B(_abc_41234_new_n3903_), .C(_abc_41234_new_n3904_), .Y(_abc_41234_new_n3905_));
OAI21X1 OAI21X1_985 ( .A(_abc_41234_new_n3900_), .B(_abc_41234_new_n3898_), .C(_abc_41234_new_n3905_), .Y(_abc_41234_new_n3906_));
OAI21X1 OAI21X1_986 ( .A(_abc_41234_new_n525__bF_buf3), .B(_abc_41234_new_n1040__bF_buf0), .C(_abc_41234_new_n3906_), .Y(_abc_41234_new_n3907_));
OAI21X1 OAI21X1_987 ( .A(_abc_41234_new_n3884_), .B(_abc_41234_new_n3908_), .C(_abc_41234_new_n3883_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_7_));
OAI21X1 OAI21X1_988 ( .A(_abc_41234_new_n522_), .B(_abc_41234_new_n2427_), .C(_abc_41234_new_n692_), .Y(_abc_41234_new_n3910_));
OAI21X1 OAI21X1_989 ( .A(_abc_41234_new_n3911_), .B(_abc_41234_new_n522_), .C(_abc_41234_new_n517_), .Y(_abc_41234_new_n3912_));
OAI21X1 OAI21X1_99 ( .A(reset_bF_buf1), .B(_abc_41234_new_n1031_), .C(_abc_41234_new_n1036_), .Y(_abc_41234_new_n1037_));
OAI21X1 OAI21X1_990 ( .A(sp_0_bF_buf1_), .B(_abc_41234_new_n3914__bF_buf3), .C(_abc_41234_new_n660__bF_buf4), .Y(_abc_41234_new_n3915_));
OAI21X1 OAI21X1_991 ( .A(_abc_41234_new_n2947__bF_buf0), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n515__bF_buf0), .Y(_abc_41234_new_n3918_));
OAI21X1 OAI21X1_992 ( .A(_abc_41234_new_n2947__bF_buf2), .B(_abc_41234_new_n1106_), .C(_abc_41234_new_n3921_), .Y(_abc_41234_new_n3922_));
OAI21X1 OAI21X1_993 ( .A(_abc_41234_new_n1105__bF_buf0), .B(_abc_41234_new_n1051_), .C(_abc_41234_new_n2464_), .Y(_abc_41234_new_n3927_));
OAI21X1 OAI21X1_994 ( .A(_abc_41234_new_n719_), .B(_abc_41234_new_n1107_), .C(_abc_41234_new_n1046__bF_buf1), .Y(_abc_41234_new_n3928_));
OAI21X1 OAI21X1_995 ( .A(_abc_41234_new_n2973_), .B(_abc_41234_new_n3927_), .C(_abc_41234_new_n3929_), .Y(_abc_41234_new_n3930_));
OAI21X1 OAI21X1_996 ( .A(_abc_41234_new_n3931_), .B(_abc_41234_new_n3932_), .C(_abc_41234_new_n2452_), .Y(_abc_41234_new_n3933_));
OAI21X1 OAI21X1_997 ( .A(_abc_41234_new_n2973_), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n515__bF_buf6), .Y(_abc_41234_new_n3937_));
OAI21X1 OAI21X1_998 ( .A(sp_1_), .B(_abc_41234_new_n3914__bF_buf2), .C(_abc_41234_new_n660__bF_buf3), .Y(_abc_41234_new_n3939_));
OAI21X1 OAI21X1_999 ( .A(_abc_41234_new_n1639__bF_buf3), .B(_abc_41234_new_n1637_), .C(_abc_41234_new_n3385_), .Y(_abc_41234_new_n3944_));
OAI22X1 OAI22X1_1 ( .A(_abc_41234_new_n714_), .B(_abc_41234_new_n683_), .C(_abc_41234_new_n680_), .D(_abc_41234_new_n702_), .Y(_abc_41234_new_n715_));
OAI22X1 OAI22X1_10 ( .A(_abc_41234_new_n818_), .B(_abc_41234_new_n722__bF_buf2), .C(_abc_41234_new_n819_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n820_));
OAI22X1 OAI22X1_100 ( .A(_abc_41234_new_n3248_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf4), .D(_abc_41234_new_n3270_), .Y(_0raddrhold_15_0__12_));
OAI22X1 OAI22X1_101 ( .A(_abc_41234_new_n1783_), .B(_abc_41234_new_n2467_), .C(_abc_41234_new_n3275_), .D(_abc_41234_new_n3276_), .Y(_abc_41234_new_n3277_));
OAI22X1 OAI22X1_102 ( .A(_abc_41234_new_n3279_), .B(_abc_41234_new_n2942__bF_buf1), .C(_abc_41234_new_n2944_), .D(_abc_41234_new_n3273_), .Y(_abc_41234_new_n3280_));
OAI22X1 OAI22X1_103 ( .A(_abc_41234_new_n534__bF_buf4), .B(_abc_41234_new_n2919__bF_buf3), .C(_abc_41234_new_n1047__bF_buf3), .D(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3282_));
OAI22X1 OAI22X1_104 ( .A(_abc_41234_new_n3272_), .B(_abc_41234_new_n2953_), .C(_abc_41234_new_n3285_), .D(_abc_41234_new_n3283_), .Y(_abc_41234_new_n3286_));
OAI22X1 OAI22X1_105 ( .A(_abc_41234_new_n895_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n2959__bF_buf2), .D(_abc_41234_new_n3290_), .Y(_abc_41234_new_n3291_));
OAI22X1 OAI22X1_106 ( .A(_abc_41234_new_n3272_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf3), .D(_abc_41234_new_n3292_), .Y(_0raddrhold_15_0__13_));
OAI22X1 OAI22X1_107 ( .A(_abc_41234_new_n1812_), .B(_abc_41234_new_n2467_), .C(_abc_41234_new_n3295_), .D(_abc_41234_new_n3296_), .Y(_abc_41234_new_n3297_));
OAI22X1 OAI22X1_108 ( .A(_abc_41234_new_n1524_), .B(_abc_41234_new_n2942__bF_buf0), .C(_abc_41234_new_n3294_), .D(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3303_));
OAI22X1 OAI22X1_109 ( .A(_abc_41234_new_n3294_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf2), .D(_abc_41234_new_n3314_), .Y(_0raddrhold_15_0__14_));
OAI22X1 OAI22X1_11 ( .A(_abc_41234_new_n821_), .B(_abc_41234_new_n526__bF_buf1), .C(_abc_41234_new_n822_), .D(_abc_41234_new_n620__bF_buf4), .Y(_abc_41234_new_n823_));
OAI22X1 OAI22X1_110 ( .A(_abc_41234_new_n1569_), .B(_abc_41234_new_n2942__bF_buf3), .C(_abc_41234_new_n3316_), .D(_abc_41234_new_n2945_), .Y(_abc_41234_new_n3326_));
OAI22X1 OAI22X1_111 ( .A(_abc_41234_new_n1005_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n2959__bF_buf1), .D(_abc_41234_new_n3333_), .Y(_abc_41234_new_n3334_));
OAI22X1 OAI22X1_112 ( .A(_abc_41234_new_n3316_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf1), .D(_abc_41234_new_n3335_), .Y(_0raddrhold_15_0__15_));
OAI22X1 OAI22X1_113 ( .A(_abc_41234_new_n3337_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf0), .D(_abc_41234_new_n3356_), .Y(_0waddrhold_15_0__0_));
OAI22X1 OAI22X1_114 ( .A(_abc_41234_new_n3358_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf9), .D(_abc_41234_new_n3379_), .Y(_0waddrhold_15_0__1_));
OAI22X1 OAI22X1_115 ( .A(_abc_41234_new_n3381_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf8), .D(_abc_41234_new_n3401_), .Y(_0waddrhold_15_0__2_));
OAI22X1 OAI22X1_116 ( .A(_abc_41234_new_n3403_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf7), .D(_abc_41234_new_n3420_), .Y(_0waddrhold_15_0__3_));
OAI22X1 OAI22X1_117 ( .A(_abc_41234_new_n3422_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf6), .D(_abc_41234_new_n3443_), .Y(_0waddrhold_15_0__4_));
OAI22X1 OAI22X1_118 ( .A(_abc_41234_new_n3445_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf5), .D(_abc_41234_new_n3464_), .Y(_0waddrhold_15_0__5_));
OAI22X1 OAI22X1_119 ( .A(_abc_41234_new_n3466_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf4), .D(_abc_41234_new_n3485_), .Y(_0waddrhold_15_0__6_));
OAI22X1 OAI22X1_12 ( .A(_abc_41234_new_n848_), .B(_abc_41234_new_n722__bF_buf1), .C(_abc_41234_new_n849_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n850_));
OAI22X1 OAI22X1_120 ( .A(_abc_41234_new_n3487_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf3), .D(_abc_41234_new_n3505_), .Y(_0waddrhold_15_0__7_));
OAI22X1 OAI22X1_121 ( .A(_abc_41234_new_n3507_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf2), .D(_abc_41234_new_n3524_), .Y(_0waddrhold_15_0__8_));
OAI22X1 OAI22X1_122 ( .A(_abc_41234_new_n3526_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf1), .D(_abc_41234_new_n3545_), .Y(_0waddrhold_15_0__9_));
OAI22X1 OAI22X1_123 ( .A(_abc_41234_new_n3547_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf0), .D(_abc_41234_new_n3567_), .Y(_0waddrhold_15_0__10_));
OAI22X1 OAI22X1_124 ( .A(_abc_41234_new_n3569_), .B(_abc_41234_new_n3339_), .C(reset_bF_buf9), .D(_abc_41234_new_n3589_), .Y(_0waddrhold_15_0__11_));
OAI22X1 OAI22X1_125 ( .A(_abc_41234_new_n847_), .B(_abc_41234_new_n2519_), .C(_abc_41234_new_n849_), .D(_abc_41234_new_n2694_), .Y(_abc_41234_new_n3591_));
OAI22X1 OAI22X1_126 ( .A(_abc_41234_new_n895_), .B(_abc_41234_new_n2519_), .C(_abc_41234_new_n904_), .D(_abc_41234_new_n2694_), .Y(_abc_41234_new_n3614_));
OAI22X1 OAI22X1_127 ( .A(_abc_41234_new_n3624_), .B(_abc_41234_new_n3339_), .C(_abc_41234_new_n3610_), .D(_abc_41234_new_n3633_), .Y(_abc_41234_new_n3634_));
OAI22X1 OAI22X1_128 ( .A(_abc_41234_new_n940_), .B(_abc_41234_new_n2519_), .C(_abc_41234_new_n1509_), .D(_abc_41234_new_n2694_), .Y(_abc_41234_new_n3637_));
OAI22X1 OAI22X1_129 ( .A(_abc_41234_new_n3652_), .B(_abc_41234_new_n3654_), .C(reset_bF_buf5), .D(_abc_41234_new_n3651_), .Y(_0waddrhold_15_0__14_));
OAI22X1 OAI22X1_13 ( .A(_abc_41234_new_n851_), .B(_abc_41234_new_n526__bF_buf0), .C(_abc_41234_new_n852_), .D(_abc_41234_new_n620__bF_buf3), .Y(_abc_41234_new_n853_));
OAI22X1 OAI22X1_130 ( .A(_abc_41234_new_n1005_), .B(_abc_41234_new_n2519_), .C(_abc_41234_new_n997_), .D(_abc_41234_new_n2694_), .Y(_abc_41234_new_n3656_));
OAI22X1 OAI22X1_131 ( .A(regfil_3__1_), .B(_abc_41234_new_n1049__bF_buf3), .C(_abc_41234_new_n3733_), .D(_abc_41234_new_n3752_), .Y(_abc_41234_new_n3753_));
OAI22X1 OAI22X1_132 ( .A(regfil_5__1_), .B(_abc_41234_new_n1304_), .C(_abc_41234_new_n3769_), .D(_abc_41234_new_n3773_), .Y(_abc_41234_new_n3774_));
OAI22X1 OAI22X1_133 ( .A(regfil_3__4_), .B(_abc_41234_new_n1049__bF_buf4), .C(_abc_41234_new_n3807_), .D(_abc_41234_new_n3823_), .Y(_abc_41234_new_n3824_));
OAI22X1 OAI22X1_134 ( .A(regfil_3__5_), .B(_abc_41234_new_n1049__bF_buf2), .C(_abc_41234_new_n3831_), .D(_abc_41234_new_n3849_), .Y(_abc_41234_new_n3850_));
OAI22X1 OAI22X1_135 ( .A(regfil_5__5_), .B(_abc_41234_new_n1304_), .C(_abc_41234_new_n3869_), .D(_abc_41234_new_n3863_), .Y(_abc_41234_new_n3870_));
OAI22X1 OAI22X1_136 ( .A(regfil_3__6_), .B(_abc_41234_new_n1049__bF_buf0), .C(_abc_41234_new_n3856_), .D(_abc_41234_new_n3878_), .Y(_abc_41234_new_n3879_));
OAI22X1 OAI22X1_137 ( .A(_abc_41234_new_n2421_), .B(_abc_41234_new_n3923_), .C(_abc_41234_new_n2947__bF_buf1), .D(_abc_41234_new_n3910_), .Y(_abc_41234_new_n3924_));
OAI22X1 OAI22X1_138 ( .A(_abc_41234_new_n2947__bF_buf0), .B(_abc_41234_new_n3913_), .C(reset_bF_buf3), .D(_abc_41234_new_n3925_), .Y(_0sp_15_0__0_));
OAI22X1 OAI22X1_139 ( .A(_abc_41234_new_n2651_), .B(_abc_41234_new_n3923_), .C(sp_1_), .D(_abc_41234_new_n3910_), .Y(_abc_41234_new_n3941_));
OAI22X1 OAI22X1_14 ( .A(_abc_41234_new_n858_), .B(_abc_41234_new_n526__bF_buf3), .C(_abc_41234_new_n859_), .D(_abc_41234_new_n620__bF_buf2), .Y(_abc_41234_new_n860_));
OAI22X1 OAI22X1_140 ( .A(_abc_41234_new_n2973_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf2), .D(_abc_41234_new_n3942_), .Y(_0sp_15_0__1_));
OAI22X1 OAI22X1_141 ( .A(_abc_41234_new_n1071_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf1), .D(_abc_41234_new_n3967_), .Y(_0sp_15_0__2_));
OAI22X1 OAI22X1_142 ( .A(_abc_41234_new_n1067_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf0), .D(_abc_41234_new_n3988_), .Y(_0sp_15_0__3_));
OAI22X1 OAI22X1_143 ( .A(_abc_41234_new_n848_), .B(_abc_41234_new_n1107_), .C(_abc_41234_new_n2488_), .D(_abc_41234_new_n3990_), .Y(_abc_41234_new_n3991_));
OAI22X1 OAI22X1_144 ( .A(_abc_41234_new_n1090_), .B(_abc_41234_new_n3917_), .C(_abc_41234_new_n3935_), .D(_abc_41234_new_n3996_), .Y(_abc_41234_new_n3997_));
OAI22X1 OAI22X1_145 ( .A(_abc_41234_new_n1090_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf9), .D(_abc_41234_new_n4007_), .Y(_0sp_15_0__4_));
OAI22X1 OAI22X1_146 ( .A(_abc_41234_new_n1080_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf8), .D(_abc_41234_new_n4077_), .Y(_0sp_15_0__7_));
OAI22X1 OAI22X1_147 ( .A(_abc_41234_new_n1255_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf7), .D(_abc_41234_new_n4099_), .Y(_0sp_15_0__8_));
OAI22X1 OAI22X1_148 ( .A(_abc_41234_new_n1251_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf6), .D(_abc_41234_new_n4121_), .Y(_0sp_15_0__9_));
OAI22X1 OAI22X1_149 ( .A(_abc_41234_new_n1362_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf5), .D(_abc_41234_new_n4167_), .Y(_0sp_15_0__11_));
OAI22X1 OAI22X1_15 ( .A(_abc_41234_new_n821_), .B(_abc_41234_new_n839_), .C(_abc_41234_new_n885_), .D(_abc_41234_new_n884_), .Y(_abc_41234_new_n886_));
OAI22X1 OAI22X1_150 ( .A(_abc_41234_new_n3279_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf4), .D(_abc_41234_new_n4208_), .Y(_0sp_15_0__13_));
OAI22X1 OAI22X1_151 ( .A(_abc_41234_new_n1524_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf3), .D(_abc_41234_new_n4232_), .Y(_0sp_15_0__14_));
OAI22X1 OAI22X1_152 ( .A(_abc_41234_new_n1569_), .B(_abc_41234_new_n3913_), .C(reset_bF_buf2), .D(_abc_41234_new_n4255_), .Y(_0sp_15_0__15_));
OAI22X1 OAI22X1_153 ( .A(_abc_41234_new_n719_), .B(_abc_41234_new_n1575_), .C(_abc_41234_new_n2707_), .D(_abc_41234_new_n4329_), .Y(_abc_41234_new_n4330_));
OAI22X1 OAI22X1_154 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n1575_), .C(_abc_41234_new_n2739_), .D(_abc_41234_new_n4329_), .Y(_abc_41234_new_n4345_));
OAI22X1 OAI22X1_155 ( .A(_abc_41234_new_n1051_), .B(_abc_41234_new_n2794_), .C(_abc_41234_new_n2564_), .D(_abc_41234_new_n4371_), .Y(_abc_41234_new_n4378_));
OAI22X1 OAI22X1_156 ( .A(_abc_41234_new_n2185__bF_buf1), .B(_abc_41234_new_n4391_), .C(_abc_41234_new_n2835_), .D(_abc_41234_new_n2916_), .Y(_abc_41234_new_n4392_));
OAI22X1 OAI22X1_157 ( .A(_abc_41234_new_n1144_), .B(_abc_41234_new_n1575_), .C(_abc_41234_new_n1653_), .D(_abc_41234_new_n4328_), .Y(_abc_41234_new_n4455_));
OAI22X1 OAI22X1_158 ( .A(_abc_41234_new_n720_), .B(_abc_41234_new_n1575_), .C(_abc_41234_new_n2564_), .D(_abc_41234_new_n4467_), .Y(_abc_41234_new_n4468_));
OAI22X1 OAI22X1_159 ( .A(_abc_41234_new_n3914__bF_buf2), .B(_abc_41234_new_n1755_), .C(_abc_41234_new_n1047__bF_buf1), .D(_abc_41234_new_n4532_), .Y(_abc_41234_new_n4533_));
OAI22X1 OAI22X1_16 ( .A(_abc_41234_new_n899_), .B(_abc_41234_new_n526__bF_buf2), .C(_abc_41234_new_n900_), .D(_abc_41234_new_n620__bF_buf1), .Y(_abc_41234_new_n901_));
OAI22X1 OAI22X1_160 ( .A(_abc_41234_new_n4605_), .B(_abc_41234_new_n2356_), .C(intcyc_bF_buf2), .D(_abc_41234_new_n2959__bF_buf0), .Y(_abc_41234_new_n4608_));
OAI22X1 OAI22X1_161 ( .A(reset_bF_buf3), .B(_abc_41234_new_n4618_), .C(_abc_41234_new_n4611_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__0_));
OAI22X1 OAI22X1_162 ( .A(reset_bF_buf2), .B(_abc_41234_new_n4623_), .C(_abc_41234_new_n4620_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__1_));
OAI22X1 OAI22X1_163 ( .A(reset_bF_buf1), .B(_abc_41234_new_n4628_), .C(_abc_41234_new_n4625_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__2_));
OAI22X1 OAI22X1_164 ( .A(reset_bF_buf0), .B(_abc_41234_new_n4633_), .C(_abc_41234_new_n4630_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__3_));
OAI22X1 OAI22X1_165 ( .A(reset_bF_buf9), .B(_abc_41234_new_n4638_), .C(_abc_41234_new_n4635_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__4_));
OAI22X1 OAI22X1_166 ( .A(reset_bF_buf8), .B(_abc_41234_new_n4643_), .C(_abc_41234_new_n4640_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__5_));
OAI22X1 OAI22X1_167 ( .A(reset_bF_buf7), .B(_abc_41234_new_n4648_), .C(_abc_41234_new_n4645_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__6_));
OAI22X1 OAI22X1_168 ( .A(reset_bF_buf6), .B(_abc_41234_new_n4653_), .C(_abc_41234_new_n4650_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__7_));
OAI22X1 OAI22X1_169 ( .A(_abc_41234_new_n3507_), .B(_abc_41234_new_n2671_), .C(_abc_41234_new_n1622_), .D(_abc_41234_new_n4605_), .Y(_abc_41234_new_n4656_));
OAI22X1 OAI22X1_17 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n722__bF_buf2), .C(_abc_41234_new_n904_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n905_));
OAI22X1 OAI22X1_170 ( .A(reset_bF_buf5), .B(_abc_41234_new_n4657_), .C(_abc_41234_new_n4655_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__8_));
OAI22X1 OAI22X1_171 ( .A(_abc_41234_new_n1670_), .B(_abc_41234_new_n4661_), .C(_abc_41234_new_n4662_), .D(_abc_41234_new_n2959__bF_buf3), .Y(_abc_41234_new_n4663_));
OAI22X1 OAI22X1_172 ( .A(_abc_41234_new_n1705_), .B(_abc_41234_new_n4661_), .C(_abc_41234_new_n4667_), .D(_abc_41234_new_n2959__bF_buf2), .Y(_abc_41234_new_n4668_));
OAI22X1 OAI22X1_173 ( .A(_abc_41234_new_n1727_), .B(_abc_41234_new_n4661_), .C(_abc_41234_new_n4672_), .D(_abc_41234_new_n2959__bF_buf1), .Y(_abc_41234_new_n4673_));
OAI22X1 OAI22X1_174 ( .A(_abc_41234_new_n3605_), .B(_abc_41234_new_n2671_), .C(_abc_41234_new_n1750_), .D(_abc_41234_new_n4605_), .Y(_abc_41234_new_n4677_));
OAI22X1 OAI22X1_175 ( .A(reset_bF_buf4), .B(_abc_41234_new_n4678_), .C(_abc_41234_new_n4676_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__12_));
OAI22X1 OAI22X1_176 ( .A(_abc_41234_new_n3624_), .B(_abc_41234_new_n2671_), .C(_abc_41234_new_n1775_), .D(_abc_41234_new_n4605_), .Y(_abc_41234_new_n4681_));
OAI22X1 OAI22X1_177 ( .A(reset_bF_buf3), .B(_abc_41234_new_n4682_), .C(_abc_41234_new_n4680_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__13_));
OAI22X1 OAI22X1_178 ( .A(_abc_41234_new_n1798_), .B(_abc_41234_new_n4661_), .C(reset_bF_buf2), .D(_abc_41234_new_n4685_), .Y(_abc_41234_new_n4686_));
OAI22X1 OAI22X1_179 ( .A(_abc_41234_new_n3661_), .B(_abc_41234_new_n2671_), .C(_abc_41234_new_n1828_), .D(_abc_41234_new_n4605_), .Y(_abc_41234_new_n4690_));
OAI22X1 OAI22X1_18 ( .A(_abc_41234_new_n906_), .B(_abc_41234_new_n526__bF_buf1), .C(_abc_41234_new_n907_), .D(_abc_41234_new_n620__bF_buf0), .Y(_abc_41234_new_n908_));
OAI22X1 OAI22X1_180 ( .A(reset_bF_buf1), .B(_abc_41234_new_n4691_), .C(_abc_41234_new_n4689_), .D(_abc_41234_new_n4615_), .Y(_0addr_15_0__15_));
OAI22X1 OAI22X1_181 ( .A(_abc_41234_new_n2950_), .B(_abc_41234_new_n4750_), .C(_abc_41234_new_n4740_), .D(_abc_41234_new_n4753_), .Y(_abc_41234_new_n4754_));
OAI22X1 OAI22X1_182 ( .A(_abc_41234_new_n2604_), .B(_abc_41234_new_n4726_), .C(_abc_41234_new_n4778_), .D(_abc_41234_new_n2638_), .Y(_abc_41234_new_n4850_));
OAI22X1 OAI22X1_183 ( .A(alu__abc_40887_new_n67_), .B(alu__abc_40887_new_n69_), .C(alu__abc_40887_new_n74_), .D(alu__abc_40887_new_n100_), .Y(alu__abc_40887_new_n101_));
OAI22X1 OAI22X1_184 ( .A(alu__abc_40887_new_n51_), .B(alu__abc_40887_new_n50_), .C(alu__abc_40887_new_n47_), .D(alu__abc_40887_new_n48_), .Y(alu__abc_40887_new_n131_));
OAI22X1 OAI22X1_185 ( .A(alu__abc_40887_new_n34_), .B(alu__abc_40887_new_n211_), .C(alu__abc_40887_new_n210_), .D(alu__abc_40887_new_n37_), .Y(alu__abc_40887_new_n212_));
OAI22X1 OAI22X1_186 ( .A(alu__abc_40887_new_n38_), .B(alu__abc_40887_new_n211_), .C(alu__abc_40887_new_n39_), .D(alu__abc_40887_new_n208_), .Y(alu__abc_40887_new_n228_));
OAI22X1 OAI22X1_187 ( .A(alu__abc_40887_new_n90_), .B(alu__abc_40887_new_n92_), .C(alu__abc_40887_new_n274_), .D(alu__abc_40887_new_n82_), .Y(alu__abc_40887_new_n275_));
OAI22X1 OAI22X1_188 ( .A(alu__abc_40887_new_n86_), .B(alu__abc_40887_new_n211_), .C(alu__abc_40887_new_n162_), .D(alu__abc_40887_new_n210_), .Y(alu__abc_40887_new_n281_));
OAI22X1 OAI22X1_189 ( .A(alu__abc_40887_new_n59_), .B(alu__abc_40887_new_n208_), .C(alu__abc_40887_new_n210_), .D(alu__abc_40887_new_n178_), .Y(alu__abc_40887_new_n313_));
OAI22X1 OAI22X1_19 ( .A(regfil_7__5_), .B(_abc_41234_new_n540_), .C(_abc_41234_new_n931_), .D(_abc_41234_new_n686_), .Y(_abc_41234_new_n932_));
OAI22X1 OAI22X1_190 ( .A(alu__abc_40887_new_n344_), .B(alu__abc_40887_new_n345_), .C(alu__abc_40887_new_n346_), .D(alu__abc_40887_new_n347_), .Y(alu__abc_40887_new_n348_));
OAI22X1 OAI22X1_2 ( .A(_abc_41234_new_n719_), .B(_abc_41234_new_n722__bF_buf3), .C(_abc_41234_new_n720_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n724_));
OAI22X1 OAI22X1_20 ( .A(_abc_41234_new_n638_), .B(_abc_41234_new_n722__bF_buf1), .C(_abc_41234_new_n944_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n945_));
OAI22X1 OAI22X1_21 ( .A(regfil_7__6_), .B(_abc_41234_new_n540_), .C(_abc_41234_new_n969_), .D(_abc_41234_new_n686_), .Y(_abc_41234_new_n970_));
OAI22X1 OAI22X1_22 ( .A(_abc_41234_new_n637_), .B(_abc_41234_new_n722__bF_buf0), .C(_abc_41234_new_n983_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n991_));
OAI22X1 OAI22X1_23 ( .A(_abc_41234_new_n992_), .B(_abc_41234_new_n526__bF_buf0), .C(_abc_41234_new_n993_), .D(_abc_41234_new_n620__bF_buf5), .Y(_abc_41234_new_n994_));
OAI22X1 OAI22X1_24 ( .A(_abc_41234_new_n996_), .B(_abc_41234_new_n722__bF_buf3), .C(_abc_41234_new_n997_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n998_));
OAI22X1 OAI22X1_25 ( .A(_abc_41234_new_n560_), .B(_abc_41234_new_n526__bF_buf3), .C(_abc_41234_new_n999_), .D(_abc_41234_new_n620__bF_buf4), .Y(_abc_41234_new_n1000_));
OAI22X1 OAI22X1_26 ( .A(_abc_41234_new_n1475_), .B(_abc_41234_new_n1481_), .C(_abc_41234_new_n1486_), .D(_abc_41234_new_n1501_), .Y(_abc_41234_new_n1502_));
OAI22X1 OAI22X1_27 ( .A(_abc_41234_new_n680_), .B(_abc_41234_new_n1105__bF_buf2), .C(_abc_41234_new_n1144_), .D(_abc_41234_new_n544__bF_buf1), .Y(_abc_41234_new_n1654_));
OAI22X1 OAI22X1_28 ( .A(_abc_41234_new_n1605_), .B(_abc_41234_new_n1607_), .C(_abc_41234_new_n523__bF_buf4), .D(_abc_41234_new_n1664_), .Y(_0wdatahold2_7_0__0_));
OAI22X1 OAI22X1_29 ( .A(_abc_41234_new_n1666_), .B(_abc_41234_new_n1607_), .C(_abc_41234_new_n523__bF_buf3), .D(_abc_41234_new_n1695_), .Y(_0wdatahold2_7_0__1_));
OAI22X1 OAI22X1_3 ( .A(_abc_41234_new_n514_), .B(_abc_41234_new_n526__bF_buf2), .C(_abc_41234_new_n725_), .D(_abc_41234_new_n620__bF_buf3), .Y(_abc_41234_new_n726_));
OAI22X1 OAI22X1_30 ( .A(_abc_41234_new_n1697_), .B(_abc_41234_new_n1607_), .C(_abc_41234_new_n523__bF_buf2), .D(_abc_41234_new_n1722_), .Y(_0wdatahold2_7_0__2_));
OAI22X1 OAI22X1_31 ( .A(_abc_41234_new_n821_), .B(_abc_41234_new_n1105__bF_buf3), .C(opcode_5_bF_buf0_), .D(_abc_41234_new_n1737_), .Y(_abc_41234_new_n1738_));
OAI22X1 OAI22X1_32 ( .A(_abc_41234_new_n1724_), .B(_abc_41234_new_n1607_), .C(_abc_41234_new_n523__bF_buf1), .D(_abc_41234_new_n1744_), .Y(_0wdatahold2_7_0__3_));
OAI22X1 OAI22X1_33 ( .A(_abc_41234_new_n1746_), .B(_abc_41234_new_n1607_), .C(_abc_41234_new_n523__bF_buf0), .D(_abc_41234_new_n1769_), .Y(_0wdatahold2_7_0__4_));
OAI22X1 OAI22X1_34 ( .A(_abc_41234_new_n906_), .B(_abc_41234_new_n1105__bF_buf1), .C(opcode_5_bF_buf3_), .D(_abc_41234_new_n1783_), .Y(_abc_41234_new_n1784_));
OAI22X1 OAI22X1_35 ( .A(_abc_41234_new_n1771_), .B(_abc_41234_new_n1607_), .C(_abc_41234_new_n523__bF_buf4), .D(_abc_41234_new_n1791_), .Y(_0wdatahold2_7_0__5_));
OAI22X1 OAI22X1_36 ( .A(opcode_5_bF_buf2_), .B(_abc_41234_new_n1812_), .C(_abc_41234_new_n1509_), .D(_abc_41234_new_n544__bF_buf1), .Y(_abc_41234_new_n1813_));
OAI22X1 OAI22X1_37 ( .A(_abc_41234_new_n1793_), .B(_abc_41234_new_n1607_), .C(_abc_41234_new_n523__bF_buf3), .D(_abc_41234_new_n1819_), .Y(_0wdatahold2_7_0__6_));
OAI22X1 OAI22X1_38 ( .A(_abc_41234_new_n560_), .B(_abc_41234_new_n1105__bF_buf0), .C(opcode_5_bF_buf1_), .D(_abc_41234_new_n1836_), .Y(_abc_41234_new_n1837_));
OAI22X1 OAI22X1_39 ( .A(_abc_41234_new_n1821_), .B(_abc_41234_new_n1607_), .C(_abc_41234_new_n523__bF_buf2), .D(_abc_41234_new_n1844_), .Y(_0wdatahold2_7_0__7_));
OAI22X1 OAI22X1_4 ( .A(_abc_41234_new_n730_), .B(_abc_41234_new_n526__bF_buf1), .C(_abc_41234_new_n731_), .D(_abc_41234_new_n620__bF_buf2), .Y(_abc_41234_new_n732_));
OAI22X1 OAI22X1_40 ( .A(_abc_41234_new_n1890_), .B(_abc_41234_new_n1874_), .C(_abc_41234_new_n1887_), .D(_abc_41234_new_n1893_), .Y(_abc_41234_new_n1894_));
OAI22X1 OAI22X1_41 ( .A(_abc_41234_new_n1900_), .B(_abc_41234_new_n1874_), .C(_abc_41234_new_n1887_), .D(_abc_41234_new_n1904_), .Y(_abc_41234_new_n1905_));
OAI22X1 OAI22X1_42 ( .A(_abc_41234_new_n600_), .B(_abc_41234_new_n2003_), .C(_abc_41234_new_n2004_), .D(_abc_41234_new_n584_), .Y(_abc_41234_new_n2005_));
OAI22X1 OAI22X1_43 ( .A(_abc_41234_new_n600_), .B(_abc_41234_new_n2011_), .C(_abc_41234_new_n2013_), .D(_abc_41234_new_n584_), .Y(_abc_41234_new_n2014_));
OAI22X1 OAI22X1_44 ( .A(_abc_41234_new_n600_), .B(_abc_41234_new_n2018_), .C(_abc_41234_new_n2020_), .D(_abc_41234_new_n2022_), .Y(_abc_41234_new_n2023_));
OAI22X1 OAI22X1_45 ( .A(_abc_41234_new_n1874_), .B(_abc_41234_new_n2074_), .C(_abc_41234_new_n2076_), .D(_abc_41234_new_n2075_), .Y(_abc_41234_new_n2077_));
OAI22X1 OAI22X1_46 ( .A(_abc_41234_new_n529_), .B(_abc_41234_new_n2190__bF_buf3), .C(_abc_41234_new_n534__bF_buf2), .D(_abc_41234_new_n2191_), .Y(_abc_41234_new_n2192_));
OAI22X1 OAI22X1_47 ( .A(_abc_41234_new_n983_), .B(_abc_41234_new_n2342_), .C(_abc_41234_new_n992_), .D(_abc_41234_new_n2255_), .Y(_abc_41234_new_n2343_));
OAI22X1 OAI22X1_48 ( .A(_abc_41234_new_n993_), .B(_abc_41234_new_n2322_), .C(_abc_41234_new_n637_), .D(_abc_41234_new_n2253_), .Y(_abc_41234_new_n2344_));
OAI22X1 OAI22X1_49 ( .A(_abc_41234_new_n997_), .B(_abc_41234_new_n2342_), .C(_abc_41234_new_n996_), .D(_abc_41234_new_n2253_), .Y(_abc_41234_new_n2346_));
OAI22X1 OAI22X1_5 ( .A(_abc_41234_new_n634_), .B(_abc_41234_new_n722__bF_buf1), .C(_abc_41234_new_n766_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n767_));
OAI22X1 OAI22X1_50 ( .A(_abc_41234_new_n999_), .B(_abc_41234_new_n2322_), .C(_abc_41234_new_n560_), .D(_abc_41234_new_n2255_), .Y(_abc_41234_new_n2347_));
OAI22X1 OAI22X1_51 ( .A(reset_bF_buf4), .B(_abc_41234_new_n2368_), .C(_abc_41234_new_n2361_), .D(_abc_41234_new_n2364_), .Y(_0parity_0_0_));
OAI22X1 OAI22X1_52 ( .A(reset_bF_buf2), .B(_abc_41234_new_n2382_), .C(_abc_41234_new_n2376_), .D(_abc_41234_new_n2364_), .Y(_0sign_0_0_));
OAI22X1 OAI22X1_53 ( .A(statesel_2_), .B(_abc_41234_new_n669__bF_buf3), .C(_abc_41234_new_n2174_), .D(_abc_41234_new_n2493_), .Y(_abc_41234_new_n2568_));
OAI22X1 OAI22X1_54 ( .A(statesel_3_), .B(_abc_41234_new_n669__bF_buf2), .C(_abc_41234_new_n2174_), .D(_abc_41234_new_n2493_), .Y(_abc_41234_new_n2593_));
OAI22X1 OAI22X1_55 ( .A(_abc_41234_new_n2588_), .B(_abc_41234_new_n2529_), .C(reset_bF_buf5), .D(_abc_41234_new_n2609_), .Y(_0statesel_5_0__3_));
OAI22X1 OAI22X1_56 ( .A(_abc_41234_new_n2611_), .B(_abc_41234_new_n2531_), .C(_abc_41234_new_n2623_), .D(_abc_41234_new_n2625_), .Y(_abc_41234_new_n2626_));
OAI22X1 OAI22X1_57 ( .A(_abc_41234_new_n2611_), .B(_abc_41234_new_n2529_), .C(reset_bF_buf4), .D(_abc_41234_new_n2627_), .Y(_0statesel_5_0__4_));
OAI22X1 OAI22X1_58 ( .A(_abc_41234_new_n2185__bF_buf2), .B(_abc_41234_new_n2190__bF_buf2), .C(_abc_41234_new_n668__bF_buf0), .D(_abc_41234_new_n2209_), .Y(_abc_41234_new_n2630_));
OAI22X1 OAI22X1_59 ( .A(_abc_41234_new_n2670_), .B(_abc_41234_new_n2675_), .C(reset_bF_buf1), .D(_abc_41234_new_n2699_), .Y(_0wdatahold_7_0__0_));
OAI22X1 OAI22X1_6 ( .A(_abc_41234_new_n768_), .B(_abc_41234_new_n526__bF_buf0), .C(_abc_41234_new_n769_), .D(_abc_41234_new_n620__bF_buf1), .Y(_abc_41234_new_n770_));
OAI22X1 OAI22X1_60 ( .A(_abc_41234_new_n719_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n514_), .D(_abc_41234_new_n2719_), .Y(_abc_41234_new_n2720_));
OAI22X1 OAI22X1_61 ( .A(_abc_41234_new_n2701_), .B(_abc_41234_new_n2675_), .C(reset_bF_buf0), .D(_abc_41234_new_n2729_), .Y(_0wdatahold_7_0__1_));
OAI22X1 OAI22X1_62 ( .A(_abc_41234_new_n1626_), .B(_abc_41234_new_n2739_), .C(_abc_41234_new_n1640_), .D(_abc_41234_new_n2743_), .Y(_abc_41234_new_n2744_));
OAI22X1 OAI22X1_63 ( .A(_abc_41234_new_n794_), .B(_abc_41234_new_n2515_), .C(_abc_41234_new_n1697_), .D(_abc_41234_new_n2671_), .Y(_abc_41234_new_n2760_));
OAI22X1 OAI22X1_64 ( .A(_abc_41234_new_n2731_), .B(_abc_41234_new_n2675_), .C(reset_bF_buf9), .D(_abc_41234_new_n2762_), .Y(_0wdatahold_7_0__2_));
OAI22X1 OAI22X1_65 ( .A(wdatahold_3_), .B(_abc_41234_new_n1608_), .C(_abc_41234_new_n2765_), .D(_abc_41234_new_n2766_), .Y(_abc_41234_new_n2767_));
OAI22X1 OAI22X1_66 ( .A(_abc_41234_new_n2764_), .B(_abc_41234_new_n2675_), .C(reset_bF_buf8), .D(_abc_41234_new_n2790_), .Y(_0wdatahold_7_0__3_));
OAI22X1 OAI22X1_67 ( .A(_abc_41234_new_n848_), .B(_abc_41234_new_n1040__bF_buf4), .C(_abc_41234_new_n2813_), .D(_abc_41234_new_n2812_), .Y(_abc_41234_new_n2814_));
OAI22X1 OAI22X1_68 ( .A(wdatahold_5_), .B(_abc_41234_new_n1608_), .C(_abc_41234_new_n2825_), .D(_abc_41234_new_n2826_), .Y(_abc_41234_new_n2827_));
OAI22X1 OAI22X1_69 ( .A(_abc_41234_new_n903_), .B(_abc_41234_new_n1040__bF_buf3), .C(_abc_41234_new_n2841_), .D(_abc_41234_new_n2840_), .Y(_abc_41234_new_n2842_));
OAI22X1 OAI22X1_7 ( .A(_abc_41234_new_n772_), .B(_abc_41234_new_n722__bF_buf0), .C(_abc_41234_new_n773_), .D(_abc_41234_new_n723_), .Y(_abc_41234_new_n774_));
OAI22X1 OAI22X1_70 ( .A(_abc_41234_new_n2824_), .B(_abc_41234_new_n2675_), .C(reset_bF_buf7), .D(_abc_41234_new_n2849_), .Y(_0wdatahold_7_0__5_));
OAI22X1 OAI22X1_71 ( .A(_abc_41234_new_n2851_), .B(_abc_41234_new_n2675_), .C(reset_bF_buf6), .D(_abc_41234_new_n2879_), .Y(_0wdatahold_7_0__6_));
OAI22X1 OAI22X1_72 ( .A(_abc_41234_new_n996_), .B(_abc_41234_new_n1040__bF_buf2), .C(_abc_41234_new_n1626_), .D(_abc_41234_new_n2884_), .Y(_abc_41234_new_n2887_));
OAI22X1 OAI22X1_73 ( .A(_abc_41234_new_n1640_), .B(_abc_41234_new_n2893_), .C(_abc_41234_new_n2889_), .D(_abc_41234_new_n1645_), .Y(_abc_41234_new_n2894_));
OAI22X1 OAI22X1_74 ( .A(_abc_41234_new_n996_), .B(_abc_41234_new_n1609_), .C(_abc_41234_new_n560_), .D(_abc_41234_new_n2719_), .Y(_abc_41234_new_n2898_));
OAI22X1 OAI22X1_75 ( .A(_abc_41234_new_n2881_), .B(_abc_41234_new_n2675_), .C(reset_bF_buf5), .D(_abc_41234_new_n2908_), .Y(_0wdatahold_7_0__7_));
OAI22X1 OAI22X1_76 ( .A(_abc_41234_new_n2947__bF_buf3), .B(_abc_41234_new_n2942__bF_buf2), .C(pc_0_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n2948_));
OAI22X1 OAI22X1_77 ( .A(_abc_41234_new_n2421_), .B(_abc_41234_new_n2958_), .C(raddrhold_0_), .D(_abc_41234_new_n2959__bF_buf3), .Y(_abc_41234_new_n2960_));
OAI22X1 OAI22X1_78 ( .A(_abc_41234_new_n2910_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf4), .D(_abc_41234_new_n2961_), .Y(_0raddrhold_15_0__0_));
OAI22X1 OAI22X1_79 ( .A(_abc_41234_new_n2973_), .B(_abc_41234_new_n2942__bF_buf1), .C(_abc_41234_new_n2706_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n2974_));
OAI22X1 OAI22X1_8 ( .A(_abc_41234_new_n751_), .B(_abc_41234_new_n526__bF_buf3), .C(_abc_41234_new_n775_), .D(_abc_41234_new_n620__bF_buf0), .Y(_abc_41234_new_n776_));
OAI22X1 OAI22X1_80 ( .A(_abc_41234_new_n2190__bF_buf0), .B(_abc_41234_new_n2979_), .C(_abc_41234_new_n2965_), .D(_abc_41234_new_n2953_), .Y(_abc_41234_new_n2981_));
OAI22X1 OAI22X1_81 ( .A(_abc_41234_new_n1071_), .B(_abc_41234_new_n2942__bF_buf0), .C(_abc_41234_new_n2995_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n3011_));
OAI22X1 OAI22X1_82 ( .A(_abc_41234_new_n1067_), .B(_abc_41234_new_n2942__bF_buf3), .C(_abc_41234_new_n2774_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n3042_));
OAI22X1 OAI22X1_83 ( .A(_abc_41234_new_n1090_), .B(_abc_41234_new_n2942__bF_buf2), .C(_abc_41234_new_n2802_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n3067_));
OAI22X1 OAI22X1_84 ( .A(_abc_41234_new_n1094_), .B(_abc_41234_new_n2942__bF_buf1), .C(_abc_41234_new_n2833_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n3094_));
OAI22X1 OAI22X1_85 ( .A(_abc_41234_new_n3074_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf1), .D(_abc_41234_new_n3099_), .Y(_0raddrhold_15_0__5_));
OAI22X1 OAI22X1_86 ( .A(_abc_41234_new_n1085_), .B(_abc_41234_new_n2942__bF_buf0), .C(_abc_41234_new_n2855_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n3111_));
OAI22X1 OAI22X1_87 ( .A(_abc_41234_new_n2190__bF_buf3), .B(_abc_41234_new_n3114_), .C(_abc_41234_new_n3101_), .D(_abc_41234_new_n2953_), .Y(_abc_41234_new_n3116_));
OAI22X1 OAI22X1_88 ( .A(_abc_41234_new_n3101_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf0), .D(_abc_41234_new_n3123_), .Y(_0raddrhold_15_0__6_));
OAI22X1 OAI22X1_89 ( .A(_abc_41234_new_n1080_), .B(_abc_41234_new_n2942__bF_buf3), .C(_abc_41234_new_n2889_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n3135_));
OAI22X1 OAI22X1_9 ( .A(_abc_41234_new_n814_), .B(_abc_41234_new_n526__bF_buf2), .C(_abc_41234_new_n815_), .D(_abc_41234_new_n620__bF_buf5), .Y(_abc_41234_new_n816_));
OAI22X1 OAI22X1_90 ( .A(_abc_41234_new_n3125_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf9), .D(_abc_41234_new_n3149_), .Y(_0raddrhold_15_0__7_));
OAI22X1 OAI22X1_91 ( .A(_abc_41234_new_n1255_), .B(_abc_41234_new_n2942__bF_buf2), .C(_abc_41234_new_n1653_), .D(_abc_41234_new_n2944_), .Y(_abc_41234_new_n3160_));
OAI22X1 OAI22X1_92 ( .A(_abc_41234_new_n3151_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf8), .D(_abc_41234_new_n3173_), .Y(_0raddrhold_15_0__8_));
OAI22X1 OAI22X1_93 ( .A(_abc_41234_new_n3175_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf7), .D(_abc_41234_new_n3198_), .Y(_0raddrhold_15_0__9_));
OAI22X1 OAI22X1_94 ( .A(_abc_41234_new_n794_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3219_), .D(_abc_41234_new_n3221_), .Y(_abc_41234_new_n3222_));
OAI22X1 OAI22X1_95 ( .A(_abc_41234_new_n3200_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf6), .D(_abc_41234_new_n3223_), .Y(_0raddrhold_15_0__10_));
OAI22X1 OAI22X1_96 ( .A(_abc_41234_new_n832_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n3243_), .D(_abc_41234_new_n3244_), .Y(_abc_41234_new_n3245_));
OAI22X1 OAI22X1_97 ( .A(_abc_41234_new_n3225_), .B(_abc_41234_new_n2914_), .C(reset_bF_buf5), .D(_abc_41234_new_n3246_), .Y(_0raddrhold_15_0__11_));
OAI22X1 OAI22X1_98 ( .A(_abc_41234_new_n1408_), .B(_abc_41234_new_n2942__bF_buf2), .C(_abc_41234_new_n2944_), .D(_abc_41234_new_n1755_), .Y(_abc_41234_new_n3256_));
OAI22X1 OAI22X1_99 ( .A(_abc_41234_new_n847_), .B(_abc_41234_new_n2958_), .C(_abc_41234_new_n2959__bF_buf3), .D(_abc_41234_new_n3268_), .Y(_abc_41234_new_n3269_));
OR2X2 OR2X2_1 ( .A(_abc_41234_new_n525__bF_buf0), .B(_abc_41234_new_n599_), .Y(_abc_41234_new_n600_));
OR2X2 OR2X2_10 ( .A(_abc_41234_new_n1252_), .B(_abc_41234_new_n1250_), .Y(_abc_41234_new_n1253_));
OR2X2 OR2X2_11 ( .A(_abc_41234_new_n1253_), .B(_abc_41234_new_n1104_), .Y(_abc_41234_new_n1254_));
OR2X2 OR2X2_12 ( .A(_abc_41234_new_n1315_), .B(_abc_41234_new_n1314_), .Y(_abc_41234_new_n1316_));
OR2X2 OR2X2_13 ( .A(_abc_41234_new_n1329_), .B(_abc_41234_new_n1333_), .Y(_abc_41234_new_n1335_));
OR2X2 OR2X2_14 ( .A(_abc_41234_new_n1304_), .B(regfil_4__1_bF_buf2_), .Y(_abc_41234_new_n1338_));
OR2X2 OR2X2_15 ( .A(_abc_41234_new_n829_), .B(_abc_41234_new_n1061_), .Y(_abc_41234_new_n1343_));
OR2X2 OR2X2_16 ( .A(_abc_41234_new_n1360_), .B(_abc_41234_new_n1364_), .Y(_abc_41234_new_n1366_));
OR2X2 OR2X2_17 ( .A(_abc_41234_new_n1254_), .B(_abc_41234_new_n1400_), .Y(_abc_41234_new_n1401_));
OR2X2 OR2X2_18 ( .A(_abc_41234_new_n1458_), .B(_abc_41234_new_n1456_), .Y(_abc_41234_new_n1459_));
OR2X2 OR2X2_19 ( .A(_abc_41234_new_n1316_), .B(_abc_41234_new_n1371_), .Y(_abc_41234_new_n1493_));
OR2X2 OR2X2_2 ( .A(_abc_41234_new_n635_), .B(regfil_1__3_), .Y(_abc_41234_new_n636_));
OR2X2 OR2X2_20 ( .A(_abc_41234_new_n1465_), .B(_abc_41234_new_n1458_), .Y(_abc_41234_new_n1521_));
OR2X2 OR2X2_21 ( .A(_abc_41234_new_n1522_), .B(_abc_41234_new_n1528_), .Y(_abc_41234_new_n1529_));
OR2X2 OR2X2_22 ( .A(_abc_41234_new_n1567_), .B(_abc_41234_new_n1571_), .Y(_abc_41234_new_n1572_));
OR2X2 OR2X2_23 ( .A(_abc_41234_new_n1579_), .B(_abc_41234_new_n1577_), .Y(_abc_41234_new_n1580_));
OR2X2 OR2X2_24 ( .A(_abc_41234_new_n1617_), .B(_abc_41234_new_n1618_), .Y(_abc_41234_new_n1619_));
OR2X2 OR2X2_25 ( .A(_abc_41234_new_n1636_), .B(_abc_41234_new_n539_), .Y(_abc_41234_new_n1637_));
OR2X2 OR2X2_26 ( .A(_abc_41234_new_n1679_), .B(_abc_41234_new_n1705_), .Y(_abc_41234_new_n1715_));
OR2X2 OR2X2_27 ( .A(_abc_41234_new_n1754_), .B(_abc_41234_new_n1775_), .Y(_abc_41234_new_n1779_));
OR2X2 OR2X2_28 ( .A(_abc_41234_new_n1749_), .B(_abc_41234_new_n1775_), .Y(_abc_41234_new_n1824_));
OR2X2 OR2X2_29 ( .A(_abc_41234_new_n1797_), .B(pc_15_), .Y(_abc_41234_new_n1826_));
OR2X2 OR2X2_3 ( .A(_abc_41234_new_n685_), .B(_abc_41234_new_n684_), .Y(_abc_41234_new_n686_));
OR2X2 OR2X2_30 ( .A(_abc_41234_new_n1057_), .B(_abc_41234_new_n653_), .Y(_abc_41234_new_n1846_));
OR2X2 OR2X2_31 ( .A(_abc_41234_new_n1846_), .B(_abc_41234_new_n677_), .Y(_abc_41234_new_n1847_));
OR2X2 OR2X2_32 ( .A(_abc_41234_new_n677_), .B(_abc_41234_new_n1966_), .Y(_abc_41234_new_n1967_));
OR2X2 OR2X2_33 ( .A(_abc_41234_new_n1846_), .B(_abc_41234_new_n1059_), .Y(_abc_41234_new_n2053_));
OR2X2 OR2X2_34 ( .A(_abc_41234_new_n2468_), .B(_abc_41234_new_n2472_), .Y(_abc_41234_new_n2473_));
OR2X2 OR2X2_35 ( .A(_abc_41234_new_n2479_), .B(_abc_41234_new_n2461_), .Y(_abc_41234_new_n2480_));
OR2X2 OR2X2_36 ( .A(_abc_41234_new_n1648_), .B(_abc_41234_new_n2705_), .Y(_abc_41234_new_n2706_));
OR2X2 OR2X2_37 ( .A(_abc_41234_new_n1649_), .B(_abc_41234_new_n1617_), .Y(_abc_41234_new_n2853_));
OR2X2 OR2X2_38 ( .A(_abc_41234_new_n2932_), .B(_abc_41234_new_n2936_), .Y(_abc_41234_new_n2937_));
OR2X2 OR2X2_39 ( .A(_abc_41234_new_n3076_), .B(_abc_41234_new_n3101_), .Y(_abc_41234_new_n3144_));
OR2X2 OR2X2_4 ( .A(_abc_41234_new_n886_), .B(_abc_41234_new_n513_), .Y(_abc_41234_new_n887_));
OR2X2 OR2X2_40 ( .A(_abc_41234_new_n3144_), .B(_abc_41234_new_n3125_), .Y(_abc_41234_new_n3145_));
OR2X2 OR2X2_41 ( .A(_abc_41234_new_n3145_), .B(_abc_41234_new_n3151_), .Y(_abc_41234_new_n3169_));
OR2X2 OR2X2_42 ( .A(_abc_41234_new_n2920_), .B(_abc_41234_new_n3321_), .Y(_abc_41234_new_n3322_));
OR2X2 OR2X2_43 ( .A(_abc_41234_new_n2921_), .B(_abc_41234_new_n534__bF_buf1), .Y(_abc_41234_new_n3344_));
OR2X2 OR2X2_44 ( .A(_abc_41234_new_n3126_), .B(_abc_41234_new_n534__bF_buf4), .Y(_abc_41234_new_n3494_));
OR2X2 OR2X2_45 ( .A(_abc_41234_new_n1656_), .B(_abc_41234_new_n534__bF_buf3), .Y(_abc_41234_new_n3512_));
OR2X2 OR2X2_46 ( .A(_abc_41234_new_n3489_), .B(_abc_41234_new_n3572_), .Y(_abc_41234_new_n3615_));
OR2X2 OR2X2_47 ( .A(_abc_41234_new_n1783_), .B(_abc_41234_new_n534__bF_buf1), .Y(_abc_41234_new_n3623_));
OR2X2 OR2X2_48 ( .A(_abc_41234_new_n1812_), .B(_abc_41234_new_n534__bF_buf0), .Y(_abc_41234_new_n3643_));
OR2X2 OR2X2_49 ( .A(_abc_41234_new_n1836_), .B(_abc_41234_new_n534__bF_buf5), .Y(_abc_41234_new_n3664_));
OR2X2 OR2X2_5 ( .A(_abc_41234_new_n806_), .B(_abc_41234_new_n918_), .Y(_abc_41234_new_n919_));
OR2X2 OR2X2_50 ( .A(_abc_41234_new_n677_), .B(_abc_41234_new_n1058_), .Y(_abc_41234_new_n3714_));
OR2X2 OR2X2_51 ( .A(_abc_41234_new_n1077_), .B(_abc_41234_new_n1076_), .Y(_abc_41234_new_n3764_));
OR2X2 OR2X2_52 ( .A(_abc_41234_new_n1160_), .B(_abc_41234_new_n1166_), .Y(_abc_41234_new_n3766_));
OR2X2 OR2X2_53 ( .A(_abc_41234_new_n1122_), .B(_abc_41234_new_n1121_), .Y(_abc_41234_new_n3771_));
OR2X2 OR2X2_54 ( .A(_abc_41234_new_n3787_), .B(_abc_41234_new_n1163_), .Y(_abc_41234_new_n3788_));
OR2X2 OR2X2_55 ( .A(_abc_41234_new_n3781_), .B(_abc_41234_new_n3801_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_3_));
OR2X2 OR2X2_56 ( .A(_abc_41234_new_n1170_), .B(_abc_41234_new_n1180_), .Y(_abc_41234_new_n3817_));
OR2X2 OR2X2_57 ( .A(_abc_41234_new_n3804_), .B(_abc_41234_new_n3825_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_4_));
OR2X2 OR2X2_58 ( .A(_abc_41234_new_n3991_), .B(_abc_41234_new_n1047__bF_buf3), .Y(_abc_41234_new_n3992_));
OR2X2 OR2X2_59 ( .A(_abc_41234_new_n4148_), .B(_abc_41234_new_n2488_), .Y(_abc_41234_new_n4149_));
OR2X2 OR2X2_6 ( .A(_abc_41234_new_n870_), .B(_abc_41234_new_n953_), .Y(_abc_41234_new_n954_));
OR2X2 OR2X2_60 ( .A(_abc_41234_new_n4210_), .B(_abc_41234_new_n1569_), .Y(_abc_41234_new_n4243_));
OR2X2 OR2X2_61 ( .A(_abc_41234_new_n4291_), .B(_abc_41234_new_n4294_), .Y(_abc_41234_new_n4295_));
OR2X2 OR2X2_62 ( .A(_abc_41234_new_n4491_), .B(_abc_41234_new_n1369_), .Y(_abc_41234_new_n4492_));
OR2X2 OR2X2_63 ( .A(_abc_41234_new_n4825_), .B(_abc_41234_new_n4765_), .Y(_abc_41234_new_n4855_));
OR2X2 OR2X2_64 ( .A(alu_oprb_3_), .B(alu_opra_3_), .Y(alu__abc_40887_new_n54_));
OR2X2 OR2X2_65 ( .A(alu_oprb_4_), .B(alu_opra_4_), .Y(alu__abc_40887_new_n57_));
OR2X2 OR2X2_66 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_40887_new_n89_));
OR2X2 OR2X2_67 ( .A(alu_oprb_0_), .B(alu_opra_0_), .Y(alu__abc_40887_new_n91_));
OR2X2 OR2X2_68 ( .A(alu__abc_40887_new_n46_), .B(alu__abc_40887_new_n49_), .Y(alu__abc_40887_new_n94_));
OR2X2 OR2X2_69 ( .A(alu__abc_40887_new_n125_), .B(alu_oprb_1_), .Y(alu__abc_40887_new_n126_));
OR2X2 OR2X2_7 ( .A(_abc_41234_new_n954_), .B(regfil_0__6_), .Y(_abc_41234_new_n955_));
OR2X2 OR2X2_70 ( .A(alu__abc_40887_new_n103_), .B(alu__abc_40887_new_n115_), .Y(alu__abc_40887_new_n210_));
OR2X2 OR2X2_71 ( .A(alu__abc_40887_new_n253_), .B(alu__abc_40887_new_n255_), .Y(alu__abc_40887_new_n256_));
OR2X2 OR2X2_72 ( .A(alu__abc_40887_new_n313_), .B(alu__abc_40887_new_n315_), .Y(alu__abc_40887_new_n316_));
OR2X2 OR2X2_73 ( .A(alu__abc_40887_new_n113_), .B(alu__abc_40887_new_n241_), .Y(alu__abc_40887_new_n374_));
OR2X2 OR2X2_8 ( .A(_abc_41234_new_n659_), .B(_abc_41234_new_n604_), .Y(_abc_41234_new_n1031_));
OR2X2 OR2X2_9 ( .A(_abc_41234_new_n1225_), .B(_abc_41234_new_n1227_), .Y(_abc_41234_new_n1245_));
XNOR2X1 XNOR2X1_1 ( .A(_abc_41234_new_n796_), .B(_abc_41234_new_n751_), .Y(_abc_41234_new_n797_));
XNOR2X1 XNOR2X1_10 ( .A(_abc_41234_new_n573_), .B(regfil_1__4_), .Y(_abc_41234_new_n2004_));
XNOR2X1 XNOR2X1_11 ( .A(_abc_41234_new_n2009_), .B(_abc_41234_new_n638_), .Y(_abc_41234_new_n2018_));
XNOR2X1 XNOR2X1_12 ( .A(pc_0_), .B(intcyc_bF_buf2), .Y(_abc_41234_new_n2684_));
XNOR2X1 XNOR2X1_13 ( .A(_abc_41234_new_n1649_), .B(pc_4_), .Y(_abc_41234_new_n2801_));
XNOR2X1 XNOR2X1_14 ( .A(_abc_41234_new_n2803_), .B(pc_4_), .Y(_abc_41234_new_n2804_));
XNOR2X1 XNOR2X1_15 ( .A(_abc_41234_new_n2853_), .B(pc_6_), .Y(_abc_41234_new_n2854_));
XNOR2X1 XNOR2X1_16 ( .A(_abc_41234_new_n2857_), .B(pc_6_), .Y(_abc_41234_new_n2858_));
XNOR2X1 XNOR2X1_17 ( .A(_abc_41234_new_n3267_), .B(raddrhold_12_), .Y(_abc_41234_new_n3268_));
XNOR2X1 XNOR2X1_18 ( .A(_abc_41234_new_n3289_), .B(_abc_41234_new_n3272_), .Y(_abc_41234_new_n3290_));
XNOR2X1 XNOR2X1_19 ( .A(_abc_41234_new_n3332_), .B(raddrhold_15_), .Y(_abc_41234_new_n3333_));
XNOR2X1 XNOR2X1_2 ( .A(regfil_4__0_), .B(sp_8_), .Y(_abc_41234_new_n1104_));
XNOR2X1 XNOR2X1_20 ( .A(_abc_41234_new_n3382_), .B(_abc_41234_new_n1067_), .Y(_abc_41234_new_n3404_));
XNOR2X1 XNOR2X1_21 ( .A(_abc_41234_new_n3489_), .B(sp_8_), .Y(_abc_41234_new_n3508_));
XNOR2X1 XNOR2X1_22 ( .A(_abc_41234_new_n3735_), .B(_abc_41234_new_n1075_), .Y(_abc_41234_new_n3736_));
XNOR2X1 XNOR2X1_23 ( .A(_abc_41234_new_n3745_), .B(_abc_41234_new_n1119_), .Y(_abc_41234_new_n3746_));
XNOR2X1 XNOR2X1_24 ( .A(_abc_41234_new_n1208_), .B(regfil_5__3_bF_buf2_), .Y(_abc_41234_new_n3782_));
XNOR2X1 XNOR2X1_25 ( .A(_abc_41234_new_n1210_), .B(_abc_41234_new_n903_), .Y(_abc_41234_new_n3830_));
XNOR2X1 XNOR2X1_26 ( .A(_abc_41234_new_n1212_), .B(_abc_41234_new_n1084_), .Y(_abc_41234_new_n3855_));
XNOR2X1 XNOR2X1_27 ( .A(_abc_41234_new_n3896_), .B(_abc_41234_new_n1127_), .Y(_abc_41234_new_n3897_));
XNOR2X1 XNOR2X1_28 ( .A(_abc_41234_new_n3953_), .B(sp_3_), .Y(_abc_41234_new_n3977_));
XNOR2X1 XNOR2X1_29 ( .A(_abc_41234_new_n3969_), .B(_abc_41234_new_n1090_), .Y(_abc_41234_new_n3990_));
XNOR2X1 XNOR2X1_3 ( .A(regfil_2__3_), .B(regfil_4__3_), .Y(_abc_41234_new_n1371_));
XNOR2X1 XNOR2X1_30 ( .A(_abc_41234_new_n4189_), .B(sp_14_), .Y(_abc_41234_new_n4219_));
XNOR2X1 XNOR2X1_31 ( .A(_abc_41234_new_n4353_), .B(_abc_41234_new_n2806_), .Y(_abc_41234_new_n4371_));
XNOR2X1 XNOR2X1_32 ( .A(alu__abc_40887_new_n170_), .B(alu__abc_40887_new_n234_), .Y(alu__abc_40887_new_n235_));
XNOR2X1 XNOR2X1_33 ( .A(alu__abc_40887_new_n249_), .B(alu__abc_40887_new_n257_), .Y(alu__abc_40887_new_n301_));
XNOR2X1 XNOR2X1_4 ( .A(regfil_5__6_bF_buf3_), .B(regfil_3__6_), .Y(_abc_41234_new_n1489_));
XNOR2X1 XNOR2X1_5 ( .A(_abc_41234_new_n1706_), .B(_abc_41234_new_n1727_), .Y(_abc_41234_new_n1728_));
XNOR2X1 XNOR2X1_6 ( .A(_abc_41234_new_n1733_), .B(_abc_41234_new_n1727_), .Y(_abc_41234_new_n1734_));
XNOR2X1 XNOR2X1_7 ( .A(_abc_41234_new_n1749_), .B(pc_13_), .Y(_abc_41234_new_n1774_));
XNOR2X1 XNOR2X1_8 ( .A(_abc_41234_new_n1888_), .B(_abc_41234_new_n814_), .Y(_abc_41234_new_n1900_));
XNOR2X1 XNOR2X1_9 ( .A(_abc_41234_new_n2002_), .B(regfil_1__4_), .Y(_abc_41234_new_n2003_));
XOR2X1 XOR2X1_1 ( .A(regfil_5__2_), .B(sp_2_), .Y(_abc_41234_new_n1077_));
XOR2X1 XOR2X1_10 ( .A(_abc_41234_new_n3832_), .B(_abc_41234_new_n1097_), .Y(_abc_41234_new_n3833_));
XOR2X1 XOR2X1_11 ( .A(_abc_41234_new_n3835_), .B(_abc_41234_new_n1132_), .Y(_abc_41234_new_n3836_));
XOR2X1 XOR2X1_12 ( .A(_abc_41234_new_n3872_), .B(_abc_41234_new_n1088_), .Y(_abc_41234_new_n3873_));
XOR2X1 XOR2X1_13 ( .A(alu_sout), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n233_));
XOR2X1 XOR2X1_14 ( .A(alu__abc_40887_new_n249_), .B(alu__abc_40887_new_n257_), .Y(alu__abc_40887_new_n258_));
XOR2X1 XOR2X1_2 ( .A(regfil_5__2_), .B(regfil_3__2_), .Y(_abc_41234_new_n1122_));
XOR2X1 XOR2X1_3 ( .A(regfil_5__5_), .B(regfil_3__5_), .Y(_abc_41234_new_n1132_));
XOR2X1 XOR2X1_4 ( .A(regfil_5__4_), .B(regfil_3__4_), .Y(_abc_41234_new_n1133_));
XOR2X1 XOR2X1_5 ( .A(_abc_41234_new_n1297_), .B(_abc_41234_new_n1301_), .Y(_abc_41234_new_n1302_));
XOR2X1 XOR2X1_6 ( .A(regfil_3__0_), .B(regfil_5__0_), .Y(_abc_41234_new_n3721_));
XOR2X1 XOR2X1_7 ( .A(_abc_41234_new_n1078_), .B(_abc_41234_new_n3784_), .Y(_abc_41234_new_n3785_));
XOR2X1 XOR2X1_8 ( .A(_abc_41234_new_n3791_), .B(_abc_41234_new_n1117_), .Y(_abc_41234_new_n3792_));
XOR2X1 XOR2X1_9 ( .A(_abc_41234_new_n1079_), .B(_abc_41234_new_n1093_), .Y(_abc_41234_new_n3821_));


endmodule