module completogpio(\WAddress[0] , \WAddress[1] , \WAddress[2] , \WAddress[3] , \WAddress[4] , \WAddress[5] , \WAddress[6] , \WAddress[7] , \WAddress[8] , \WAddress[9] , \WAddress[10] , \WAddress[11] , \WAddress[12] , \WAddress[13] , \WAddress[14] , \WAddress[15] , \WAddress[16] , \WAddress[17] , \WAddress[18] , \WAddress[19] , \WAddress[20] , \WAddress[21] , \WAddress[22] , \WAddress[23] , \WAddress[24] , \WAddress[25] , \WAddress[26] , \WAddress[27] , \WAddress[28] , \WAddress[29] , \WAddress[30] , \WAddress[31] , \Wdata[0] , \Wdata[1] , \Wdata[2] , \Wdata[3] , \Wdata[4] , \Wdata[5] , \Wdata[6] , \Wdata[7] , \Wdata[8] , \Wdata[9] , \Wdata[10] , \Wdata[11] , \Wdata[12] , \Wdata[13] , \Wdata[14] , \Wdata[15] , \Wdata[16] , \Wdata[17] , \Wdata[18] , \Wdata[19] , \Wdata[20] , \Wdata[21] , \Wdata[22] , \Wdata[23] , \Wdata[24] , \Wdata[25] , \Wdata[26] , \Wdata[27] , \Wdata[28] , \Wdata[29] , \Wdata[30] , \Wdata[31] , AWvalid, \pindata[0] , \pindata[1] , \pindata[2] , \pindata[3] , \pindata[4] , \pindata[5] , \pindata[6] , \pindata[7] , \RAddress[0] , \RAddress[1] , \RAddress[2] , \RAddress[3] , \RAddress[4] , \RAddress[5] , \RAddress[6] , \RAddress[7] , \RAddress[8] , \RAddress[9] , \RAddress[10] , \RAddress[11] , \RAddress[12] , \RAddress[13] , \RAddress[14] , \RAddress[15] , \RAddress[16] , \RAddress[17] , \RAddress[18] , \RAddress[19] , \RAddress[20] , \RAddress[21] , \RAddress[22] , \RAddress[23] , \RAddress[24] , \RAddress[25] , \RAddress[26] , \RAddress[27] , \RAddress[28] , \RAddress[29] , \RAddress[30] , \RAddress[31] , Wvalid, clock, ARvalid, reset, Rready, Bready, ARready, Rvalid, AWready, Wready, Bvalid, \Rx[0] , \Rx[1] , \Rx[2] , \Rx[3] , \Rx[4] , \Rx[5] , \Rx[6] , \Rx[7] , \datanw[0] , \datanw[1] , \datanw[2] , \datanw[3] , \datanw[4] , \datanw[5] , \datanw[6] , \datanw[7] , \Tx[0] , \Tx[1] , \Tx[2] , \Tx[3] , \Tx[4] , \Tx[5] , \Tx[6] , \Tx[7] , \DSE[0] , \DSE[1] , \DSE[2] , \DSE[3] , \DSE[4] , \DSE[5] , \DSE[6] , \DSE[7] , \Rdata[0] , \Rdata[1] , \Rdata[2] , \Rdata[3] , \Rdata[4] , \Rdata[5] , \Rdata[6] , \Rdata[7] , \Rdata[8] , \Rdata[9] , \Rdata[10] , \Rdata[11] , \Rdata[12] , \Rdata[13] , \Rdata[14] , \Rdata[15] , \Rdata[16] , \Rdata[17] , \Rdata[18] , \Rdata[19] , \Rdata[20] , \Rdata[21] , \Rdata[22] , \Rdata[23] , \Rdata[24] , \Rdata[25] , \Rdata[26] , \Rdata[27] , \Rdata[28] , \Rdata[29] , \Rdata[30] , \Rdata[31] );

output ARready;
input ARvalid;
output AWready;
input AWvalid;
input Bready;
output Bvalid;
output \DSE[0] ;
output \DSE[1] ;
output \DSE[2] ;
output \DSE[3] ;
output \DSE[4] ;
output \DSE[5] ;
output \DSE[6] ;
output \DSE[7] ;
wire LRAddress_0_; 
wire LRAddress_1_; 
wire LRAddress_2_; 
wire LWAddress_0_; 
wire LWAddress_1_; 
wire LWAddress_2_; 
input \RAddress[0] ;
input \RAddress[10] ;
input \RAddress[11] ;
input \RAddress[12] ;
input \RAddress[13] ;
input \RAddress[14] ;
input \RAddress[15] ;
input \RAddress[16] ;
input \RAddress[17] ;
input \RAddress[18] ;
input \RAddress[19] ;
input \RAddress[1] ;
input \RAddress[20] ;
input \RAddress[21] ;
input \RAddress[22] ;
input \RAddress[23] ;
input \RAddress[24] ;
input \RAddress[25] ;
input \RAddress[26] ;
input \RAddress[27] ;
input \RAddress[28] ;
input \RAddress[29] ;
input \RAddress[2] ;
input \RAddress[30] ;
input \RAddress[31] ;
input \RAddress[3] ;
input \RAddress[4] ;
input \RAddress[5] ;
input \RAddress[6] ;
input \RAddress[7] ;
input \RAddress[8] ;
input \RAddress[9] ;
output \Rdata[0] ;
output \Rdata[10] ;
output \Rdata[11] ;
output \Rdata[12] ;
output \Rdata[13] ;
output \Rdata[14] ;
output \Rdata[15] ;
output \Rdata[16] ;
output \Rdata[17] ;
output \Rdata[18] ;
output \Rdata[19] ;
output \Rdata[1] ;
output \Rdata[20] ;
output \Rdata[21] ;
output \Rdata[22] ;
output \Rdata[23] ;
output \Rdata[24] ;
output \Rdata[25] ;
output \Rdata[26] ;
output \Rdata[27] ;
output \Rdata[28] ;
output \Rdata[29] ;
output \Rdata[2] ;
output \Rdata[30] ;
output \Rdata[31] ;
output \Rdata[3] ;
output \Rdata[4] ;
output \Rdata[5] ;
output \Rdata[6] ;
output \Rdata[7] ;
output \Rdata[8] ;
output \Rdata[9] ;
input Rready;
output Rvalid;
output \Rx[0] ;
output \Rx[1] ;
output \Rx[2] ;
output \Rx[3] ;
output \Rx[4] ;
output \Rx[5] ;
output \Rx[6] ;
output \Rx[7] ;
output \Tx[0] ;
output \Tx[1] ;
output \Tx[2] ;
output \Tx[3] ;
output \Tx[4] ;
output \Tx[5] ;
output \Tx[6] ;
output \Tx[7] ;
input \WAddress[0] ;
input \WAddress[10] ;
input \WAddress[11] ;
input \WAddress[12] ;
input \WAddress[13] ;
input \WAddress[14] ;
input \WAddress[15] ;
input \WAddress[16] ;
input \WAddress[17] ;
input \WAddress[18] ;
input \WAddress[19] ;
input \WAddress[1] ;
input \WAddress[20] ;
input \WAddress[21] ;
input \WAddress[22] ;
input \WAddress[23] ;
input \WAddress[24] ;
input \WAddress[25] ;
input \WAddress[26] ;
input \WAddress[27] ;
input \WAddress[28] ;
input \WAddress[29] ;
input \WAddress[2] ;
input \WAddress[30] ;
input \WAddress[31] ;
input \WAddress[3] ;
input \WAddress[4] ;
input \WAddress[5] ;
input \WAddress[6] ;
input \WAddress[7] ;
input \WAddress[8] ;
input \WAddress[9] ;
input \Wdata[0] ;
input \Wdata[10] ;
input \Wdata[11] ;
input \Wdata[12] ;
input \Wdata[13] ;
input \Wdata[14] ;
input \Wdata[15] ;
input \Wdata[16] ;
input \Wdata[17] ;
input \Wdata[18] ;
input \Wdata[19] ;
input \Wdata[1] ;
input \Wdata[20] ;
input \Wdata[21] ;
input \Wdata[22] ;
input \Wdata[23] ;
input \Wdata[24] ;
input \Wdata[25] ;
input \Wdata[26] ;
input \Wdata[27] ;
input \Wdata[28] ;
input \Wdata[29] ;
input \Wdata[2] ;
input \Wdata[30] ;
input \Wdata[31] ;
input \Wdata[3] ;
input \Wdata[4] ;
input \Wdata[5] ;
input \Wdata[6] ;
input \Wdata[7] ;
input \Wdata[8] ;
input \Wdata[9] ;
output Wready;
input Wvalid;
wire _0Rdata_0_0_; 
wire _0vel_0_0_; 
wire _abc_1210_new_n18_; 
wire _abc_1210_new_n19_; 
wire _abc_1210_new_n20_; 
wire _abc_1210_new_n21_; 
wire _abc_1210_new_n22_; 
wire _abc_1210_new_n24_; 
wire _abc_1210_new_n25_; 
wire _abc_1210_new_n26_; 
wire _abc_1210_new_n27_; 
wire _abc_1210_new_n28_; 
wire _abc_1210_new_n29_; 
wire _abc_1210_new_n30_; 
wire _abc_1210_new_n31_; 
wire _abc_1210_new_n32_; 
wire _abc_1210_new_n33_; 
wire _abc_1210_new_n34_; 
wire _abc_1210_new_n35_; 
wire _abc_1210_new_n36_; 
wire _abc_1210_new_n37_; 
wire _abc_1210_new_n38_; 
wire _abc_1210_new_n39_; 
wire _abc_1210_new_n40_; 
wire _abc_1210_new_n41_; 
wire _abc_1210_new_n42_; 
wire _abc_1210_new_n43_; 
wire _abc_1210_new_n44_; 
wire _abc_1210_new_n45_; 
wire _abc_1210_new_n46_; 
wire _abc_1210_new_n47_; 
wire _auto_iopadmap_cc_368_execute_1371; 
wire _auto_iopadmap_cc_368_execute_1373; 
wire _auto_iopadmap_cc_368_execute_1375; 
wire _auto_iopadmap_cc_368_execute_1386_0_; 
wire _auto_iopadmap_cc_368_execute_1419; 
wire _auto_iopadmap_cc_368_execute_1439; 
input clock;
wire clock_bF_buf0; 
wire clock_bF_buf1; 
wire clock_bF_buf2; 
wire clock_bF_buf3; 
wire clock_bF_buf4; 
wire clock_bF_buf5; 
wire clock_bF_buf6; 
output \datanw[0] ;
output \datanw[1] ;
output \datanw[2] ;
output \datanw[3] ;
output \datanw[4] ;
output \datanw[5] ;
output \datanw[6] ;
output \datanw[7] ;
wire decor__abc_1242_new_n13_; 
wire decor__abc_1242_new_n14_; 
wire decor__abc_1242_new_n15_; 
wire decor__abc_1242_new_n16_; 
wire decor__abc_1242_new_n17_; 
wire decor__abc_1242_new_n19_; 
wire decor__abc_1242_new_n21_; 
wire decor__abc_1242_new_n23_; 
wire decor__abc_1242_new_n25_; 
wire decow__abc_1242_new_n13_; 
wire decow__abc_1242_new_n14_; 
wire decow__abc_1242_new_n15_; 
wire decow__abc_1242_new_n16_; 
wire decow__abc_1242_new_n17_; 
wire decow__abc_1242_new_n19_; 
wire decow__abc_1242_new_n21_; 
wire decow__abc_1242_new_n23_; 
wire decow__abc_1242_new_n25_; 
wire flip1_R1; 
wire flip1_Rx; 
wire flip1_Tx; 
wire flip1_W1; 
wire flip1__0Rx_0_0_; 
wire flip1__0Tx_0_0_; 
wire flip1__abc_1260_new_n10_; 
wire flip1__abc_1260_new_n11_; 
wire flip1__abc_1260_new_n12_; 
wire flip1__abc_1260_new_n13_; 
wire flip1__abc_1260_new_n15_; 
wire flip1__abc_1260_new_n16_; 
wire flip1__abc_1260_new_n8_; 
wire flip1__abc_1260_new_n9_; 
wire flip2_R1; 
wire flip2_Rx; 
wire flip2_Tx; 
wire flip2_W1; 
wire flip2__0Rx_0_0_; 
wire flip2__0Tx_0_0_; 
wire flip2__abc_1260_new_n10_; 
wire flip2__abc_1260_new_n11_; 
wire flip2__abc_1260_new_n12_; 
wire flip2__abc_1260_new_n13_; 
wire flip2__abc_1260_new_n15_; 
wire flip2__abc_1260_new_n16_; 
wire flip2__abc_1260_new_n8_; 
wire flip2__abc_1260_new_n9_; 
wire flip3_R1; 
wire flip3_Rx; 
wire flip3_Tx; 
wire flip3_W1; 
wire flip3__0Rx_0_0_; 
wire flip3__0Tx_0_0_; 
wire flip3__abc_1260_new_n10_; 
wire flip3__abc_1260_new_n11_; 
wire flip3__abc_1260_new_n12_; 
wire flip3__abc_1260_new_n13_; 
wire flip3__abc_1260_new_n15_; 
wire flip3__abc_1260_new_n16_; 
wire flip3__abc_1260_new_n8_; 
wire flip3__abc_1260_new_n9_; 
wire flip4_R1; 
wire flip4_Rx; 
wire flip4_Tx; 
wire flip4_W1; 
wire flip4__0Rx_0_0_; 
wire flip4__0Tx_0_0_; 
wire flip4__abc_1260_new_n10_; 
wire flip4__abc_1260_new_n11_; 
wire flip4__abc_1260_new_n12_; 
wire flip4__abc_1260_new_n13_; 
wire flip4__abc_1260_new_n15_; 
wire flip4__abc_1260_new_n16_; 
wire flip4__abc_1260_new_n8_; 
wire flip4__abc_1260_new_n9_; 
wire flip5_R1; 
wire flip5_Rx; 
wire flip5_Tx; 
wire flip5_W1; 
wire flip5__0Rx_0_0_; 
wire flip5__0Tx_0_0_; 
wire flip5__abc_1260_new_n10_; 
wire flip5__abc_1260_new_n11_; 
wire flip5__abc_1260_new_n12_; 
wire flip5__abc_1260_new_n13_; 
wire flip5__abc_1260_new_n15_; 
wire flip5__abc_1260_new_n16_; 
wire flip5__abc_1260_new_n8_; 
wire flip5__abc_1260_new_n9_; 
wire flip6_R1; 
wire flip6_Rx; 
wire flip6_Tx; 
wire flip6_W1; 
wire flip6__0Rx_0_0_; 
wire flip6__0Tx_0_0_; 
wire flip6__abc_1260_new_n10_; 
wire flip6__abc_1260_new_n11_; 
wire flip6__abc_1260_new_n12_; 
wire flip6__abc_1260_new_n13_; 
wire flip6__abc_1260_new_n15_; 
wire flip6__abc_1260_new_n16_; 
wire flip6__abc_1260_new_n8_; 
wire flip6__abc_1260_new_n9_; 
wire flip7_R1; 
wire flip7_Rx; 
wire flip7_Tx; 
wire flip7_W1; 
wire flip7__0Rx_0_0_; 
wire flip7__0Tx_0_0_; 
wire flip7__abc_1260_new_n10_; 
wire flip7__abc_1260_new_n11_; 
wire flip7__abc_1260_new_n12_; 
wire flip7__abc_1260_new_n13_; 
wire flip7__abc_1260_new_n15_; 
wire flip7__abc_1260_new_n16_; 
wire flip7__abc_1260_new_n8_; 
wire flip7__abc_1260_new_n9_; 
wire flip8_R1; 
wire flip8_Rx; 
wire flip8_Tx; 
wire flip8_W1; 
wire flip8__0Rx_0_0_; 
wire flip8__0Tx_0_0_; 
wire flip8__abc_1260_new_n10_; 
wire flip8__abc_1260_new_n11_; 
wire flip8__abc_1260_new_n12_; 
wire flip8__abc_1260_new_n13_; 
wire flip8__abc_1260_new_n15_; 
wire flip8__abc_1260_new_n16_; 
wire flip8__abc_1260_new_n8_; 
wire flip8__abc_1260_new_n9_; 
wire flipw1_DS; 
wire flipw1__0DS_0_0_; 
wire flipw1__0outdata_0_0_; 
wire flipw1__abc_1271_new_n10_; 
wire flipw1__abc_1271_new_n11_; 
wire flipw1__abc_1271_new_n12_; 
wire flipw1__abc_1271_new_n14_; 
wire flipw1__abc_1271_new_n15_; 
wire flipw1__abc_1271_new_n16_; 
wire flipw1__abc_1271_new_n9_; 
wire flipw1_outdata; 
wire flipw2_DS; 
wire flipw2__0DS_0_0_; 
wire flipw2__0outdata_0_0_; 
wire flipw2__abc_1271_new_n10_; 
wire flipw2__abc_1271_new_n11_; 
wire flipw2__abc_1271_new_n12_; 
wire flipw2__abc_1271_new_n14_; 
wire flipw2__abc_1271_new_n15_; 
wire flipw2__abc_1271_new_n16_; 
wire flipw2__abc_1271_new_n9_; 
wire flipw2_outdata; 
wire flipw3_DS; 
wire flipw3__0DS_0_0_; 
wire flipw3__0outdata_0_0_; 
wire flipw3__abc_1271_new_n10_; 
wire flipw3__abc_1271_new_n11_; 
wire flipw3__abc_1271_new_n12_; 
wire flipw3__abc_1271_new_n14_; 
wire flipw3__abc_1271_new_n15_; 
wire flipw3__abc_1271_new_n16_; 
wire flipw3__abc_1271_new_n9_; 
wire flipw3_outdata; 
wire flipw4_DS; 
wire flipw4__0DS_0_0_; 
wire flipw4__0outdata_0_0_; 
wire flipw4__abc_1271_new_n10_; 
wire flipw4__abc_1271_new_n11_; 
wire flipw4__abc_1271_new_n12_; 
wire flipw4__abc_1271_new_n14_; 
wire flipw4__abc_1271_new_n15_; 
wire flipw4__abc_1271_new_n16_; 
wire flipw4__abc_1271_new_n9_; 
wire flipw4_outdata; 
wire flipw5_DS; 
wire flipw5__0DS_0_0_; 
wire flipw5__0outdata_0_0_; 
wire flipw5__abc_1271_new_n10_; 
wire flipw5__abc_1271_new_n11_; 
wire flipw5__abc_1271_new_n12_; 
wire flipw5__abc_1271_new_n14_; 
wire flipw5__abc_1271_new_n15_; 
wire flipw5__abc_1271_new_n16_; 
wire flipw5__abc_1271_new_n9_; 
wire flipw5_outdata; 
wire flipw6_DS; 
wire flipw6__0DS_0_0_; 
wire flipw6__0outdata_0_0_; 
wire flipw6__abc_1271_new_n10_; 
wire flipw6__abc_1271_new_n11_; 
wire flipw6__abc_1271_new_n12_; 
wire flipw6__abc_1271_new_n14_; 
wire flipw6__abc_1271_new_n15_; 
wire flipw6__abc_1271_new_n16_; 
wire flipw6__abc_1271_new_n9_; 
wire flipw6_outdata; 
wire flipw7_DS; 
wire flipw7__0DS_0_0_; 
wire flipw7__0outdata_0_0_; 
wire flipw7__abc_1271_new_n10_; 
wire flipw7__abc_1271_new_n11_; 
wire flipw7__abc_1271_new_n12_; 
wire flipw7__abc_1271_new_n14_; 
wire flipw7__abc_1271_new_n15_; 
wire flipw7__abc_1271_new_n16_; 
wire flipw7__abc_1271_new_n9_; 
wire flipw7_outdata; 
wire flipw8_DS; 
wire flipw8__0DS_0_0_; 
wire flipw8__0outdata_0_0_; 
wire flipw8__abc_1271_new_n10_; 
wire flipw8__abc_1271_new_n11_; 
wire flipw8__abc_1271_new_n12_; 
wire flipw8__abc_1271_new_n14_; 
wire flipw8__abc_1271_new_n15_; 
wire flipw8__abc_1271_new_n16_; 
wire flipw8__abc_1271_new_n9_; 
wire flipw8_outdata; 
wire latchR__0LWAddres_2_0__0_; 
wire latchR__0LWAddres_2_0__1_; 
wire latchR__0LWAddres_2_0__2_; 
wire latchR__abc_1281_new_n12_; 
wire latchR__abc_1281_new_n13_; 
wire latchR__abc_1281_new_n14_; 
wire latchR__abc_1281_new_n15_; 
wire latchR__abc_1281_new_n17_; 
wire latchR__abc_1281_new_n18_; 
wire latchR__abc_1281_new_n19_; 
wire latchR__abc_1281_new_n21_; 
wire latchR__abc_1281_new_n22_; 
wire latchR__abc_1281_new_n23_; 
wire latchW__0LWAddres_2_0__0_; 
wire latchW__0LWAddres_2_0__1_; 
wire latchW__0LWAddres_2_0__2_; 
wire latchW__abc_1281_new_n12_; 
wire latchW__abc_1281_new_n13_; 
wire latchW__abc_1281_new_n14_; 
wire latchW__abc_1281_new_n15_; 
wire latchW__abc_1281_new_n17_; 
wire latchW__abc_1281_new_n18_; 
wire latchW__abc_1281_new_n19_; 
wire latchW__abc_1281_new_n21_; 
wire latchW__abc_1281_new_n22_; 
wire latchW__abc_1281_new_n23_; 
wire maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_477; 
wire maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_490; 
wire maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_494; 
wire maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_498; 
wire maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_502; 
wire maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_506; 
wire maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_510; 
wire maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_0_; 
wire maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_10_; 
wire maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_2_; 
wire maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_9_; 
wire maquina__abc_1295_new_n101_; 
wire maquina__abc_1295_new_n102_; 
wire maquina__abc_1295_new_n35_; 
wire maquina__abc_1295_new_n36_; 
wire maquina__abc_1295_new_n37_; 
wire maquina__abc_1295_new_n38_; 
wire maquina__abc_1295_new_n39_; 
wire maquina__abc_1295_new_n40_; 
wire maquina__abc_1295_new_n41_; 
wire maquina__abc_1295_new_n42_; 
wire maquina__abc_1295_new_n43_; 
wire maquina__abc_1295_new_n44_; 
wire maquina__abc_1295_new_n46_; 
wire maquina__abc_1295_new_n47_; 
wire maquina__abc_1295_new_n48_; 
wire maquina__abc_1295_new_n49_; 
wire maquina__abc_1295_new_n50_; 
wire maquina__abc_1295_new_n52_; 
wire maquina__abc_1295_new_n53_; 
wire maquina__abc_1295_new_n54_; 
wire maquina__abc_1295_new_n55_; 
wire maquina__abc_1295_new_n56_; 
wire maquina__abc_1295_new_n57_; 
wire maquina__abc_1295_new_n58_; 
wire maquina__abc_1295_new_n60_; 
wire maquina__abc_1295_new_n61_; 
wire maquina__abc_1295_new_n62_; 
wire maquina__abc_1295_new_n63_; 
wire maquina__abc_1295_new_n64_; 
wire maquina__abc_1295_new_n65_; 
wire maquina__abc_1295_new_n67_; 
wire maquina__abc_1295_new_n68_; 
wire maquina__abc_1295_new_n69_; 
wire maquina__abc_1295_new_n70_; 
wire maquina__abc_1295_new_n71_; 
wire maquina__abc_1295_new_n72_; 
wire maquina__abc_1295_new_n73_; 
wire maquina__abc_1295_new_n74_; 
wire maquina__abc_1295_new_n75_; 
wire maquina__abc_1295_new_n76_; 
wire maquina__abc_1295_new_n77_; 
wire maquina__abc_1295_new_n79_; 
wire maquina__abc_1295_new_n80_; 
wire maquina__abc_1295_new_n81_; 
wire maquina__abc_1295_new_n83_; 
wire maquina__abc_1295_new_n84_; 
wire maquina__abc_1295_new_n85_; 
wire maquina__abc_1295_new_n87_; 
wire maquina__abc_1295_new_n88_; 
wire maquina__abc_1295_new_n89_; 
wire maquina__abc_1295_new_n90_; 
wire maquina__abc_1295_new_n91_; 
wire maquina__abc_1295_new_n92_; 
wire maquina__abc_1295_new_n93_; 
wire maquina__abc_1295_new_n94_; 
wire maquina__abc_1295_new_n95_; 
wire maquina__abc_1295_new_n97_; 
wire maquina__abc_1295_new_n98_; 
wire maquina__abc_1295_new_n99_; 
wire maquina_state_0_; 
wire maquina_state_10_; 
wire maquina_state_1_; 
wire maquina_state_2_; 
wire maquina_state_3_; 
wire maquina_state_4_; 
wire maquina_state_5_; 
wire maquina_state_6_; 
wire maquina_state_7_; 
wire maquina_state_8_; 
wire maquina_state_9_; 
wire maquina_vel; 
input \pindata[0] ;
input \pindata[1] ;
input \pindata[2] ;
input \pindata[3] ;
input \pindata[4] ;
input \pindata[5] ;
input \pindata[6] ;
input \pindata[7] ;
input reset;
wire reset_bF_buf0; 
wire reset_bF_buf1; 
wire reset_bF_buf2; 
wire reset_bF_buf3; 
wire reset_bF_buf4; 
wire reset_bF_buf5; 
wire reset_bF_buf6; 
AND2X2 AND2X2_1 ( .A(_abc_1210_new_n18_), .B(maquina_vel), .Y(_abc_1210_new_n19_));
AND2X2 AND2X2_10 ( .A(LRAddress_0_), .B(\pindata[1] ), .Y(_abc_1210_new_n41_));
AND2X2 AND2X2_100 ( .A(flipw5__abc_1271_new_n10_), .B(flipw5_outdata), .Y(flipw5__abc_1271_new_n11_));
AND2X2 AND2X2_101 ( .A(flipw5__abc_1271_new_n12_), .B(reset_bF_buf1), .Y(flipw5__0outdata_0_0_));
AND2X2 AND2X2_102 ( .A(flip5_W1), .B(\Wdata[1] ), .Y(flipw5__abc_1271_new_n14_));
AND2X2 AND2X2_103 ( .A(flipw5__abc_1271_new_n10_), .B(flipw5_DS), .Y(flipw5__abc_1271_new_n15_));
AND2X2 AND2X2_104 ( .A(flipw5__abc_1271_new_n16_), .B(reset_bF_buf0), .Y(flipw5__0DS_0_0_));
AND2X2 AND2X2_105 ( .A(\Wdata[0] ), .B(flip6_W1), .Y(flipw6__abc_1271_new_n9_));
AND2X2 AND2X2_106 ( .A(flipw6__abc_1271_new_n10_), .B(flipw6_outdata), .Y(flipw6__abc_1271_new_n11_));
AND2X2 AND2X2_107 ( .A(flipw6__abc_1271_new_n12_), .B(reset_bF_buf6), .Y(flipw6__0outdata_0_0_));
AND2X2 AND2X2_108 ( .A(flip6_W1), .B(\Wdata[1] ), .Y(flipw6__abc_1271_new_n14_));
AND2X2 AND2X2_109 ( .A(flipw6__abc_1271_new_n10_), .B(flipw6_DS), .Y(flipw6__abc_1271_new_n15_));
AND2X2 AND2X2_11 ( .A(_abc_1210_new_n27_), .B(\pindata[0] ), .Y(_abc_1210_new_n42_));
AND2X2 AND2X2_110 ( .A(flipw6__abc_1271_new_n16_), .B(reset_bF_buf5), .Y(flipw6__0DS_0_0_));
AND2X2 AND2X2_111 ( .A(\Wdata[0] ), .B(flip7_W1), .Y(flipw7__abc_1271_new_n9_));
AND2X2 AND2X2_112 ( .A(flipw7__abc_1271_new_n10_), .B(flipw7_outdata), .Y(flipw7__abc_1271_new_n11_));
AND2X2 AND2X2_113 ( .A(flipw7__abc_1271_new_n12_), .B(reset_bF_buf4), .Y(flipw7__0outdata_0_0_));
AND2X2 AND2X2_114 ( .A(flip7_W1), .B(\Wdata[1] ), .Y(flipw7__abc_1271_new_n14_));
AND2X2 AND2X2_115 ( .A(flipw7__abc_1271_new_n10_), .B(flipw7_DS), .Y(flipw7__abc_1271_new_n15_));
AND2X2 AND2X2_116 ( .A(flipw7__abc_1271_new_n16_), .B(reset_bF_buf3), .Y(flipw7__0DS_0_0_));
AND2X2 AND2X2_117 ( .A(\Wdata[0] ), .B(flip8_W1), .Y(flipw8__abc_1271_new_n9_));
AND2X2 AND2X2_118 ( .A(flipw8__abc_1271_new_n10_), .B(flipw8_outdata), .Y(flipw8__abc_1271_new_n11_));
AND2X2 AND2X2_119 ( .A(flipw8__abc_1271_new_n12_), .B(reset_bF_buf2), .Y(flipw8__0outdata_0_0_));
AND2X2 AND2X2_12 ( .A(_abc_1210_new_n40_), .B(_abc_1210_new_n44_), .Y(_abc_1210_new_n45_));
AND2X2 AND2X2_120 ( .A(flip8_W1), .B(\Wdata[1] ), .Y(flipw8__abc_1271_new_n14_));
AND2X2 AND2X2_121 ( .A(flipw8__abc_1271_new_n10_), .B(flipw8_DS), .Y(flipw8__abc_1271_new_n15_));
AND2X2 AND2X2_122 ( .A(flipw8__abc_1271_new_n16_), .B(reset_bF_buf1), .Y(flipw8__0DS_0_0_));
AND2X2 AND2X2_123 ( .A(\RAddress[0] ), .B(ARvalid), .Y(latchR__abc_1281_new_n12_));
AND2X2 AND2X2_124 ( .A(latchR__abc_1281_new_n13_), .B(LRAddress_0_), .Y(latchR__abc_1281_new_n14_));
AND2X2 AND2X2_125 ( .A(latchR__abc_1281_new_n15_), .B(reset_bF_buf0), .Y(latchR__0LWAddres_2_0__0_));
AND2X2 AND2X2_126 ( .A(ARvalid), .B(\RAddress[1] ), .Y(latchR__abc_1281_new_n17_));
AND2X2 AND2X2_127 ( .A(latchR__abc_1281_new_n13_), .B(LRAddress_1_), .Y(latchR__abc_1281_new_n18_));
AND2X2 AND2X2_128 ( .A(latchR__abc_1281_new_n19_), .B(reset_bF_buf6), .Y(latchR__0LWAddres_2_0__1_));
AND2X2 AND2X2_129 ( .A(ARvalid), .B(\RAddress[2] ), .Y(latchR__abc_1281_new_n21_));
AND2X2 AND2X2_13 ( .A(_abc_1210_new_n46_), .B(reset_bF_buf5), .Y(_abc_1210_new_n47_));
AND2X2 AND2X2_130 ( .A(latchR__abc_1281_new_n13_), .B(LRAddress_2_), .Y(latchR__abc_1281_new_n22_));
AND2X2 AND2X2_131 ( .A(latchR__abc_1281_new_n23_), .B(reset_bF_buf5), .Y(latchR__0LWAddres_2_0__2_));
AND2X2 AND2X2_132 ( .A(\WAddress[0] ), .B(AWvalid), .Y(latchW__abc_1281_new_n12_));
AND2X2 AND2X2_133 ( .A(latchW__abc_1281_new_n13_), .B(LWAddress_0_), .Y(latchW__abc_1281_new_n14_));
AND2X2 AND2X2_134 ( .A(latchW__abc_1281_new_n15_), .B(reset_bF_buf4), .Y(latchW__0LWAddres_2_0__0_));
AND2X2 AND2X2_135 ( .A(AWvalid), .B(\WAddress[1] ), .Y(latchW__abc_1281_new_n17_));
AND2X2 AND2X2_136 ( .A(latchW__abc_1281_new_n13_), .B(LWAddress_1_), .Y(latchW__abc_1281_new_n18_));
AND2X2 AND2X2_137 ( .A(latchW__abc_1281_new_n19_), .B(reset_bF_buf3), .Y(latchW__0LWAddres_2_0__1_));
AND2X2 AND2X2_138 ( .A(AWvalid), .B(\WAddress[2] ), .Y(latchW__abc_1281_new_n21_));
AND2X2 AND2X2_139 ( .A(latchW__abc_1281_new_n13_), .B(LWAddress_2_), .Y(latchW__abc_1281_new_n22_));
AND2X2 AND2X2_14 ( .A(_abc_1210_new_n47_), .B(_abc_1210_new_n36_), .Y(_0Rdata_0_0_));
AND2X2 AND2X2_140 ( .A(latchW__abc_1281_new_n23_), .B(reset_bF_buf2), .Y(latchW__0LWAddres_2_0__2_));
AND2X2 AND2X2_141 ( .A(reset_bF_buf1), .B(maquina_state_0_), .Y(maquina__abc_1295_new_n35_));
AND2X2 AND2X2_142 ( .A(maquina__abc_1295_new_n36_), .B(maquina__abc_1295_new_n37_), .Y(maquina__abc_1295_new_n38_));
AND2X2 AND2X2_143 ( .A(maquina__abc_1295_new_n38_), .B(maquina__abc_1295_new_n35_), .Y(maquina__abc_1295_new_n39_));
AND2X2 AND2X2_144 ( .A(Rready), .B(maquina_state_9_), .Y(maquina__abc_1295_new_n41_));
AND2X2 AND2X2_145 ( .A(maquina_state_10_), .B(Bready), .Y(maquina__abc_1295_new_n43_));
AND2X2 AND2X2_146 ( .A(reset_bF_buf6), .B(maquina_state_2_), .Y(maquina__abc_1295_new_n47_));
AND2X2 AND2X2_147 ( .A(maquina__abc_1295_new_n47_), .B(maquina__abc_1295_new_n46_), .Y(maquina__abc_1295_new_n48_));
AND2X2 AND2X2_148 ( .A(maquina__abc_1295_new_n36_), .B(AWvalid), .Y(maquina__abc_1295_new_n49_));
AND2X2 AND2X2_149 ( .A(maquina__abc_1295_new_n49_), .B(maquina__abc_1295_new_n35_), .Y(maquina__abc_1295_new_n50_));
AND2X2 AND2X2_15 ( .A(decor__abc_1242_new_n13_), .B(decor__abc_1242_new_n14_), .Y(decor__abc_1242_new_n15_));
AND2X2 AND2X2_150 ( .A(reset_bF_buf5), .B(maquina_vel), .Y(maquina__abc_1295_new_n52_));
AND2X2 AND2X2_151 ( .A(maquina__abc_1295_new_n52_), .B(maquina_state_5_), .Y(maquina__abc_1295_new_n53_));
AND2X2 AND2X2_152 ( .A(maquina__abc_1295_new_n56_), .B(reset_bF_buf4), .Y(maquina__abc_1295_new_n57_));
AND2X2 AND2X2_153 ( .A(maquina__abc_1295_new_n57_), .B(maquina__abc_1295_new_n55_), .Y(maquina__abc_1295_new_n58_));
AND2X2 AND2X2_154 ( .A(maquina__abc_1295_new_n52_), .B(maquina_state_8_), .Y(maquina__abc_1295_new_n60_));
AND2X2 AND2X2_155 ( .A(maquina__abc_1295_new_n63_), .B(reset_bF_buf3), .Y(maquina__abc_1295_new_n64_));
AND2X2 AND2X2_156 ( .A(maquina__abc_1295_new_n64_), .B(maquina__abc_1295_new_n62_), .Y(maquina__abc_1295_new_n65_));
AND2X2 AND2X2_157 ( .A(maquina__abc_1295_new_n68_), .B(maquina__abc_1295_new_n69_), .Y(maquina__abc_1295_new_n70_));
AND2X2 AND2X2_158 ( .A(maquina__abc_1295_new_n70_), .B(maquina__abc_1295_new_n67_), .Y(maquina__abc_1295_new_n71_));
AND2X2 AND2X2_159 ( .A(maquina__abc_1295_new_n72_), .B(maquina_state_10_), .Y(maquina__abc_1295_new_n73_));
AND2X2 AND2X2_16 ( .A(decor__abc_1242_new_n16_), .B(_auto_iopadmap_cc_368_execute_1371), .Y(decor__abc_1242_new_n17_));
AND2X2 AND2X2_160 ( .A(maquina__abc_1295_new_n74_), .B(maquina__abc_1295_new_n75_), .Y(maquina__abc_1295_new_n76_));
AND2X2 AND2X2_161 ( .A(maquina__abc_1295_new_n76_), .B(maquina__abc_1295_new_n73_), .Y(maquina__abc_1295_new_n77_));
AND2X2 AND2X2_162 ( .A(maquina__abc_1295_new_n71_), .B(maquina__abc_1295_new_n77_), .Y(_auto_iopadmap_cc_368_execute_1375));
AND2X2 AND2X2_163 ( .A(maquina__abc_1295_new_n79_), .B(maquina__abc_1295_new_n67_), .Y(maquina__abc_1295_new_n80_));
AND2X2 AND2X2_164 ( .A(maquina__abc_1295_new_n81_), .B(maquina__abc_1295_new_n76_), .Y(_auto_iopadmap_cc_368_execute_1439));
AND2X2 AND2X2_165 ( .A(maquina__abc_1295_new_n71_), .B(maquina__abc_1295_new_n83_), .Y(maquina__abc_1295_new_n84_));
AND2X2 AND2X2_166 ( .A(maquina__abc_1295_new_n85_), .B(maquina__abc_1295_new_n76_), .Y(_auto_iopadmap_cc_368_execute_1373));
AND2X2 AND2X2_167 ( .A(maquina__abc_1295_new_n67_), .B(maquina_state_9_), .Y(maquina__abc_1295_new_n88_));
AND2X2 AND2X2_168 ( .A(maquina__abc_1295_new_n89_), .B(maquina__abc_1295_new_n68_), .Y(maquina__abc_1295_new_n90_));
AND2X2 AND2X2_169 ( .A(maquina__abc_1295_new_n90_), .B(maquina__abc_1295_new_n88_), .Y(maquina__abc_1295_new_n91_));
AND2X2 AND2X2_17 ( .A(decor__abc_1242_new_n15_), .B(decor__abc_1242_new_n17_), .Y(flip1_R1));
AND2X2 AND2X2_170 ( .A(maquina__abc_1295_new_n93_), .B(maquina__abc_1295_new_n76_), .Y(maquina__abc_1295_new_n94_));
AND2X2 AND2X2_171 ( .A(maquina__abc_1295_new_n94_), .B(maquina__abc_1295_new_n91_), .Y(maquina__abc_1295_new_n95_));
AND2X2 AND2X2_172 ( .A(maquina__abc_1295_new_n95_), .B(maquina__abc_1295_new_n87_), .Y(_auto_iopadmap_cc_368_execute_1419));
AND2X2 AND2X2_173 ( .A(maquina__abc_1295_new_n84_), .B(maquina__abc_1295_new_n97_), .Y(maquina__abc_1295_new_n98_));
AND2X2 AND2X2_174 ( .A(maquina__abc_1295_new_n99_), .B(maquina__abc_1295_new_n74_), .Y(_auto_iopadmap_cc_368_execute_1371));
AND2X2 AND2X2_175 ( .A(maquina__abc_1295_new_n101_), .B(reset_bF_buf2), .Y(maquina__abc_1295_new_n102_));
AND2X2 AND2X2_176 ( .A(maquina__abc_1295_new_n102_), .B(maquina_state_5_), .Y(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_477));
AND2X2 AND2X2_177 ( .A(maquina__abc_1295_new_n35_), .B(ARvalid), .Y(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_498));
AND2X2 AND2X2_178 ( .A(reset_bF_buf1), .B(maquina_state_7_), .Y(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_494));
AND2X2 AND2X2_179 ( .A(reset_bF_buf0), .B(maquina_state_6_), .Y(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_490));
AND2X2 AND2X2_18 ( .A(decor__abc_1242_new_n13_), .B(LRAddress_0_), .Y(decor__abc_1242_new_n19_));
AND2X2 AND2X2_180 ( .A(reset_bF_buf6), .B(maquina_state_1_), .Y(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_502));
AND2X2 AND2X2_181 ( .A(maquina__abc_1295_new_n102_), .B(maquina_state_8_), .Y(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_506));
AND2X2 AND2X2_182 ( .A(maquina__abc_1295_new_n47_), .B(Wvalid), .Y(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_510));
AND2X2 AND2X2_19 ( .A(decor__abc_1242_new_n17_), .B(decor__abc_1242_new_n19_), .Y(flip2_R1));
AND2X2 AND2X2_2 ( .A(\Wdata[2] ), .B(Wvalid), .Y(_abc_1210_new_n21_));
AND2X2 AND2X2_20 ( .A(decor__abc_1242_new_n14_), .B(LRAddress_1_), .Y(decor__abc_1242_new_n21_));
AND2X2 AND2X2_21 ( .A(decor__abc_1242_new_n17_), .B(decor__abc_1242_new_n21_), .Y(flip3_R1));
AND2X2 AND2X2_22 ( .A(LRAddress_1_), .B(LRAddress_0_), .Y(decor__abc_1242_new_n23_));
AND2X2 AND2X2_23 ( .A(decor__abc_1242_new_n17_), .B(decor__abc_1242_new_n23_), .Y(flip4_R1));
AND2X2 AND2X2_24 ( .A(LRAddress_2_), .B(_auto_iopadmap_cc_368_execute_1371), .Y(decor__abc_1242_new_n25_));
AND2X2 AND2X2_25 ( .A(decor__abc_1242_new_n15_), .B(decor__abc_1242_new_n25_), .Y(flip5_R1));
AND2X2 AND2X2_26 ( .A(decor__abc_1242_new_n19_), .B(decor__abc_1242_new_n25_), .Y(flip6_R1));
AND2X2 AND2X2_27 ( .A(decor__abc_1242_new_n21_), .B(decor__abc_1242_new_n25_), .Y(flip7_R1));
AND2X2 AND2X2_28 ( .A(decor__abc_1242_new_n23_), .B(decor__abc_1242_new_n25_), .Y(flip8_R1));
AND2X2 AND2X2_29 ( .A(decow__abc_1242_new_n13_), .B(decow__abc_1242_new_n14_), .Y(decow__abc_1242_new_n15_));
AND2X2 AND2X2_3 ( .A(LRAddress_0_), .B(\pindata[7] ), .Y(_abc_1210_new_n25_));
AND2X2 AND2X2_30 ( .A(decow__abc_1242_new_n16_), .B(_auto_iopadmap_cc_368_execute_1373), .Y(decow__abc_1242_new_n17_));
AND2X2 AND2X2_31 ( .A(decow__abc_1242_new_n15_), .B(decow__abc_1242_new_n17_), .Y(flip1_W1));
AND2X2 AND2X2_32 ( .A(decow__abc_1242_new_n13_), .B(LWAddress_0_), .Y(decow__abc_1242_new_n19_));
AND2X2 AND2X2_33 ( .A(decow__abc_1242_new_n17_), .B(decow__abc_1242_new_n19_), .Y(flip2_W1));
AND2X2 AND2X2_34 ( .A(decow__abc_1242_new_n14_), .B(LWAddress_1_), .Y(decow__abc_1242_new_n21_));
AND2X2 AND2X2_35 ( .A(decow__abc_1242_new_n17_), .B(decow__abc_1242_new_n21_), .Y(flip3_W1));
AND2X2 AND2X2_36 ( .A(LWAddress_1_), .B(LWAddress_0_), .Y(decow__abc_1242_new_n23_));
AND2X2 AND2X2_37 ( .A(decow__abc_1242_new_n17_), .B(decow__abc_1242_new_n23_), .Y(flip4_W1));
AND2X2 AND2X2_38 ( .A(LWAddress_2_), .B(_auto_iopadmap_cc_368_execute_1373), .Y(decow__abc_1242_new_n25_));
AND2X2 AND2X2_39 ( .A(decow__abc_1242_new_n15_), .B(decow__abc_1242_new_n25_), .Y(flip5_W1));
AND2X2 AND2X2_4 ( .A(_abc_1210_new_n27_), .B(\pindata[6] ), .Y(_abc_1210_new_n28_));
AND2X2 AND2X2_40 ( .A(decow__abc_1242_new_n19_), .B(decow__abc_1242_new_n25_), .Y(flip6_W1));
AND2X2 AND2X2_41 ( .A(decow__abc_1242_new_n21_), .B(decow__abc_1242_new_n25_), .Y(flip7_W1));
AND2X2 AND2X2_42 ( .A(decow__abc_1242_new_n23_), .B(decow__abc_1242_new_n25_), .Y(flip8_W1));
AND2X2 AND2X2_43 ( .A(flip1__abc_1260_new_n9_), .B(flip1_Tx), .Y(flip1__abc_1260_new_n10_));
AND2X2 AND2X2_44 ( .A(flip1__abc_1260_new_n8_), .B(flip1_R1), .Y(flip1__abc_1260_new_n12_));
AND2X2 AND2X2_45 ( .A(flip1__abc_1260_new_n9_), .B(reset_bF_buf3), .Y(flip1__abc_1260_new_n16_));
AND2X2 AND2X2_46 ( .A(flip1__abc_1260_new_n15_), .B(flip1__abc_1260_new_n16_), .Y(flip1__0Rx_0_0_));
AND2X2 AND2X2_47 ( .A(flip2__abc_1260_new_n9_), .B(flip2_Tx), .Y(flip2__abc_1260_new_n10_));
AND2X2 AND2X2_48 ( .A(flip2__abc_1260_new_n8_), .B(flip2_R1), .Y(flip2__abc_1260_new_n12_));
AND2X2 AND2X2_49 ( .A(flip2__abc_1260_new_n9_), .B(reset_bF_buf1), .Y(flip2__abc_1260_new_n16_));
AND2X2 AND2X2_5 ( .A(LRAddress_0_), .B(\pindata[5] ), .Y(_abc_1210_new_n31_));
AND2X2 AND2X2_50 ( .A(flip2__abc_1260_new_n15_), .B(flip2__abc_1260_new_n16_), .Y(flip2__0Rx_0_0_));
AND2X2 AND2X2_51 ( .A(flip3__abc_1260_new_n9_), .B(flip3_Tx), .Y(flip3__abc_1260_new_n10_));
AND2X2 AND2X2_52 ( .A(flip3__abc_1260_new_n8_), .B(flip3_R1), .Y(flip3__abc_1260_new_n12_));
AND2X2 AND2X2_53 ( .A(flip3__abc_1260_new_n9_), .B(reset_bF_buf6), .Y(flip3__abc_1260_new_n16_));
AND2X2 AND2X2_54 ( .A(flip3__abc_1260_new_n15_), .B(flip3__abc_1260_new_n16_), .Y(flip3__0Rx_0_0_));
AND2X2 AND2X2_55 ( .A(flip4__abc_1260_new_n9_), .B(flip4_Tx), .Y(flip4__abc_1260_new_n10_));
AND2X2 AND2X2_56 ( .A(flip4__abc_1260_new_n8_), .B(flip4_R1), .Y(flip4__abc_1260_new_n12_));
AND2X2 AND2X2_57 ( .A(flip4__abc_1260_new_n9_), .B(reset_bF_buf4), .Y(flip4__abc_1260_new_n16_));
AND2X2 AND2X2_58 ( .A(flip4__abc_1260_new_n15_), .B(flip4__abc_1260_new_n16_), .Y(flip4__0Rx_0_0_));
AND2X2 AND2X2_59 ( .A(flip5__abc_1260_new_n9_), .B(flip5_Tx), .Y(flip5__abc_1260_new_n10_));
AND2X2 AND2X2_6 ( .A(_abc_1210_new_n27_), .B(\pindata[4] ), .Y(_abc_1210_new_n32_));
AND2X2 AND2X2_60 ( .A(flip5__abc_1260_new_n8_), .B(flip5_R1), .Y(flip5__abc_1260_new_n12_));
AND2X2 AND2X2_61 ( .A(flip5__abc_1260_new_n9_), .B(reset_bF_buf2), .Y(flip5__abc_1260_new_n16_));
AND2X2 AND2X2_62 ( .A(flip5__abc_1260_new_n15_), .B(flip5__abc_1260_new_n16_), .Y(flip5__0Rx_0_0_));
AND2X2 AND2X2_63 ( .A(flip6__abc_1260_new_n9_), .B(flip6_Tx), .Y(flip6__abc_1260_new_n10_));
AND2X2 AND2X2_64 ( .A(flip6__abc_1260_new_n8_), .B(flip6_R1), .Y(flip6__abc_1260_new_n12_));
AND2X2 AND2X2_65 ( .A(flip6__abc_1260_new_n9_), .B(reset_bF_buf0), .Y(flip6__abc_1260_new_n16_));
AND2X2 AND2X2_66 ( .A(flip6__abc_1260_new_n15_), .B(flip6__abc_1260_new_n16_), .Y(flip6__0Rx_0_0_));
AND2X2 AND2X2_67 ( .A(flip7__abc_1260_new_n9_), .B(flip7_Tx), .Y(flip7__abc_1260_new_n10_));
AND2X2 AND2X2_68 ( .A(flip7__abc_1260_new_n8_), .B(flip7_R1), .Y(flip7__abc_1260_new_n12_));
AND2X2 AND2X2_69 ( .A(flip7__abc_1260_new_n9_), .B(reset_bF_buf5), .Y(flip7__abc_1260_new_n16_));
AND2X2 AND2X2_7 ( .A(_abc_1210_new_n30_), .B(_abc_1210_new_n34_), .Y(_abc_1210_new_n35_));
AND2X2 AND2X2_70 ( .A(flip7__abc_1260_new_n15_), .B(flip7__abc_1260_new_n16_), .Y(flip7__0Rx_0_0_));
AND2X2 AND2X2_71 ( .A(flip8__abc_1260_new_n9_), .B(flip8_Tx), .Y(flip8__abc_1260_new_n10_));
AND2X2 AND2X2_72 ( .A(flip8__abc_1260_new_n8_), .B(flip8_R1), .Y(flip8__abc_1260_new_n12_));
AND2X2 AND2X2_73 ( .A(flip8__abc_1260_new_n9_), .B(reset_bF_buf3), .Y(flip8__abc_1260_new_n16_));
AND2X2 AND2X2_74 ( .A(flip8__abc_1260_new_n15_), .B(flip8__abc_1260_new_n16_), .Y(flip8__0Rx_0_0_));
AND2X2 AND2X2_75 ( .A(\Wdata[0] ), .B(flip1_W1), .Y(flipw1__abc_1271_new_n9_));
AND2X2 AND2X2_76 ( .A(flipw1__abc_1271_new_n10_), .B(flipw1_outdata), .Y(flipw1__abc_1271_new_n11_));
AND2X2 AND2X2_77 ( .A(flipw1__abc_1271_new_n12_), .B(reset_bF_buf2), .Y(flipw1__0outdata_0_0_));
AND2X2 AND2X2_78 ( .A(flip1_W1), .B(\Wdata[1] ), .Y(flipw1__abc_1271_new_n14_));
AND2X2 AND2X2_79 ( .A(flipw1__abc_1271_new_n10_), .B(flipw1_DS), .Y(flipw1__abc_1271_new_n15_));
AND2X2 AND2X2_8 ( .A(LRAddress_0_), .B(\pindata[3] ), .Y(_abc_1210_new_n37_));
AND2X2 AND2X2_80 ( .A(flipw1__abc_1271_new_n16_), .B(reset_bF_buf1), .Y(flipw1__0DS_0_0_));
AND2X2 AND2X2_81 ( .A(\Wdata[0] ), .B(flip2_W1), .Y(flipw2__abc_1271_new_n9_));
AND2X2 AND2X2_82 ( .A(flipw2__abc_1271_new_n10_), .B(flipw2_outdata), .Y(flipw2__abc_1271_new_n11_));
AND2X2 AND2X2_83 ( .A(flipw2__abc_1271_new_n12_), .B(reset_bF_buf0), .Y(flipw2__0outdata_0_0_));
AND2X2 AND2X2_84 ( .A(flip2_W1), .B(\Wdata[1] ), .Y(flipw2__abc_1271_new_n14_));
AND2X2 AND2X2_85 ( .A(flipw2__abc_1271_new_n10_), .B(flipw2_DS), .Y(flipw2__abc_1271_new_n15_));
AND2X2 AND2X2_86 ( .A(flipw2__abc_1271_new_n16_), .B(reset_bF_buf6), .Y(flipw2__0DS_0_0_));
AND2X2 AND2X2_87 ( .A(\Wdata[0] ), .B(flip3_W1), .Y(flipw3__abc_1271_new_n9_));
AND2X2 AND2X2_88 ( .A(flipw3__abc_1271_new_n10_), .B(flipw3_outdata), .Y(flipw3__abc_1271_new_n11_));
AND2X2 AND2X2_89 ( .A(flipw3__abc_1271_new_n12_), .B(reset_bF_buf5), .Y(flipw3__0outdata_0_0_));
AND2X2 AND2X2_9 ( .A(_abc_1210_new_n27_), .B(\pindata[2] ), .Y(_abc_1210_new_n38_));
AND2X2 AND2X2_90 ( .A(flip3_W1), .B(\Wdata[1] ), .Y(flipw3__abc_1271_new_n14_));
AND2X2 AND2X2_91 ( .A(flipw3__abc_1271_new_n10_), .B(flipw3_DS), .Y(flipw3__abc_1271_new_n15_));
AND2X2 AND2X2_92 ( .A(flipw3__abc_1271_new_n16_), .B(reset_bF_buf4), .Y(flipw3__0DS_0_0_));
AND2X2 AND2X2_93 ( .A(\Wdata[0] ), .B(flip4_W1), .Y(flipw4__abc_1271_new_n9_));
AND2X2 AND2X2_94 ( .A(flipw4__abc_1271_new_n10_), .B(flipw4_outdata), .Y(flipw4__abc_1271_new_n11_));
AND2X2 AND2X2_95 ( .A(flipw4__abc_1271_new_n12_), .B(reset_bF_buf3), .Y(flipw4__0outdata_0_0_));
AND2X2 AND2X2_96 ( .A(flip4_W1), .B(\Wdata[1] ), .Y(flipw4__abc_1271_new_n14_));
AND2X2 AND2X2_97 ( .A(flipw4__abc_1271_new_n10_), .B(flipw4_DS), .Y(flipw4__abc_1271_new_n15_));
AND2X2 AND2X2_98 ( .A(flipw4__abc_1271_new_n16_), .B(reset_bF_buf2), .Y(flipw4__0DS_0_0_));
AND2X2 AND2X2_99 ( .A(\Wdata[0] ), .B(flip5_W1), .Y(flipw5__abc_1271_new_n9_));
BUFX2 BUFX2_1 ( .A(_auto_iopadmap_cc_368_execute_1371), .Y(ARready));
BUFX2 BUFX2_10 ( .A(flipw7_DS), .Y(\DSE[6] ));
BUFX2 BUFX2_11 ( .A(flipw8_DS), .Y(\DSE[7] ));
BUFX2 BUFX2_12 ( .A(_auto_iopadmap_cc_368_execute_1386_0_), .Y(\Rdata[0] ));
BUFX2 BUFX2_13 ( .A(1'h0), .Y(\Rdata[1] ));
BUFX2 BUFX2_14 ( .A(1'h0), .Y(\Rdata[2] ));
BUFX2 BUFX2_15 ( .A(1'h0), .Y(\Rdata[3] ));
BUFX2 BUFX2_16 ( .A(1'h0), .Y(\Rdata[4] ));
BUFX2 BUFX2_17 ( .A(1'h0), .Y(\Rdata[5] ));
BUFX2 BUFX2_18 ( .A(1'h0), .Y(\Rdata[6] ));
BUFX2 BUFX2_19 ( .A(1'h0), .Y(\Rdata[7] ));
BUFX2 BUFX2_2 ( .A(_auto_iopadmap_cc_368_execute_1373), .Y(AWready));
BUFX2 BUFX2_20 ( .A(1'h0), .Y(\Rdata[8] ));
BUFX2 BUFX2_21 ( .A(1'h0), .Y(\Rdata[9] ));
BUFX2 BUFX2_22 ( .A(1'h0), .Y(\Rdata[10] ));
BUFX2 BUFX2_23 ( .A(1'h0), .Y(\Rdata[11] ));
BUFX2 BUFX2_24 ( .A(1'h0), .Y(\Rdata[12] ));
BUFX2 BUFX2_25 ( .A(1'h0), .Y(\Rdata[13] ));
BUFX2 BUFX2_26 ( .A(1'h0), .Y(\Rdata[14] ));
BUFX2 BUFX2_27 ( .A(1'h0), .Y(\Rdata[15] ));
BUFX2 BUFX2_28 ( .A(1'h0), .Y(\Rdata[16] ));
BUFX2 BUFX2_29 ( .A(1'h0), .Y(\Rdata[17] ));
BUFX2 BUFX2_3 ( .A(_auto_iopadmap_cc_368_execute_1375), .Y(Bvalid));
BUFX2 BUFX2_30 ( .A(1'h0), .Y(\Rdata[18] ));
BUFX2 BUFX2_31 ( .A(1'h0), .Y(\Rdata[19] ));
BUFX2 BUFX2_32 ( .A(1'h0), .Y(\Rdata[20] ));
BUFX2 BUFX2_33 ( .A(1'h0), .Y(\Rdata[21] ));
BUFX2 BUFX2_34 ( .A(1'h0), .Y(\Rdata[22] ));
BUFX2 BUFX2_35 ( .A(1'h0), .Y(\Rdata[23] ));
BUFX2 BUFX2_36 ( .A(1'h0), .Y(\Rdata[24] ));
BUFX2 BUFX2_37 ( .A(1'h0), .Y(\Rdata[25] ));
BUFX2 BUFX2_38 ( .A(1'h0), .Y(\Rdata[26] ));
BUFX2 BUFX2_39 ( .A(1'h0), .Y(\Rdata[27] ));
BUFX2 BUFX2_4 ( .A(flipw1_DS), .Y(\DSE[0] ));
BUFX2 BUFX2_40 ( .A(1'h0), .Y(\Rdata[28] ));
BUFX2 BUFX2_41 ( .A(1'h0), .Y(\Rdata[29] ));
BUFX2 BUFX2_42 ( .A(1'h0), .Y(\Rdata[30] ));
BUFX2 BUFX2_43 ( .A(1'h0), .Y(\Rdata[31] ));
BUFX2 BUFX2_44 ( .A(_auto_iopadmap_cc_368_execute_1419), .Y(Rvalid));
BUFX2 BUFX2_45 ( .A(flip1_Rx), .Y(\Rx[0] ));
BUFX2 BUFX2_46 ( .A(flip2_Rx), .Y(\Rx[1] ));
BUFX2 BUFX2_47 ( .A(flip3_Rx), .Y(\Rx[2] ));
BUFX2 BUFX2_48 ( .A(flip4_Rx), .Y(\Rx[3] ));
BUFX2 BUFX2_49 ( .A(flip5_Rx), .Y(\Rx[4] ));
BUFX2 BUFX2_5 ( .A(flipw2_DS), .Y(\DSE[1] ));
BUFX2 BUFX2_50 ( .A(flip6_Rx), .Y(\Rx[5] ));
BUFX2 BUFX2_51 ( .A(flip7_Rx), .Y(\Rx[6] ));
BUFX2 BUFX2_52 ( .A(flip8_Rx), .Y(\Rx[7] ));
BUFX2 BUFX2_53 ( .A(flip1_Tx), .Y(\Tx[0] ));
BUFX2 BUFX2_54 ( .A(flip2_Tx), .Y(\Tx[1] ));
BUFX2 BUFX2_55 ( .A(flip3_Tx), .Y(\Tx[2] ));
BUFX2 BUFX2_56 ( .A(flip4_Tx), .Y(\Tx[3] ));
BUFX2 BUFX2_57 ( .A(flip5_Tx), .Y(\Tx[4] ));
BUFX2 BUFX2_58 ( .A(flip6_Tx), .Y(\Tx[5] ));
BUFX2 BUFX2_59 ( .A(flip7_Tx), .Y(\Tx[6] ));
BUFX2 BUFX2_6 ( .A(flipw3_DS), .Y(\DSE[2] ));
BUFX2 BUFX2_60 ( .A(flip8_Tx), .Y(\Tx[7] ));
BUFX2 BUFX2_61 ( .A(_auto_iopadmap_cc_368_execute_1439), .Y(Wready));
BUFX2 BUFX2_62 ( .A(flipw1_outdata), .Y(\datanw[0] ));
BUFX2 BUFX2_63 ( .A(flipw2_outdata), .Y(\datanw[1] ));
BUFX2 BUFX2_64 ( .A(flipw3_outdata), .Y(\datanw[2] ));
BUFX2 BUFX2_65 ( .A(flipw4_outdata), .Y(\datanw[3] ));
BUFX2 BUFX2_66 ( .A(flipw5_outdata), .Y(\datanw[4] ));
BUFX2 BUFX2_67 ( .A(flipw6_outdata), .Y(\datanw[5] ));
BUFX2 BUFX2_68 ( .A(flipw7_outdata), .Y(\datanw[6] ));
BUFX2 BUFX2_69 ( .A(flipw8_outdata), .Y(\datanw[7] ));
BUFX2 BUFX2_7 ( .A(flipw4_DS), .Y(\DSE[3] ));
BUFX2 BUFX2_8 ( .A(flipw5_DS), .Y(\DSE[4] ));
BUFX2 BUFX2_9 ( .A(flipw6_DS), .Y(\DSE[5] ));
BUFX4 BUFX4_1 ( .A(clock), .Y(clock_bF_buf6));
BUFX4 BUFX4_10 ( .A(reset), .Y(reset_bF_buf4));
BUFX4 BUFX4_11 ( .A(reset), .Y(reset_bF_buf3));
BUFX4 BUFX4_12 ( .A(reset), .Y(reset_bF_buf2));
BUFX4 BUFX4_13 ( .A(reset), .Y(reset_bF_buf1));
BUFX4 BUFX4_14 ( .A(reset), .Y(reset_bF_buf0));
BUFX4 BUFX4_2 ( .A(clock), .Y(clock_bF_buf5));
BUFX4 BUFX4_3 ( .A(clock), .Y(clock_bF_buf4));
BUFX4 BUFX4_4 ( .A(clock), .Y(clock_bF_buf3));
BUFX4 BUFX4_5 ( .A(clock), .Y(clock_bF_buf2));
BUFX4 BUFX4_6 ( .A(clock), .Y(clock_bF_buf1));
BUFX4 BUFX4_7 ( .A(clock), .Y(clock_bF_buf0));
BUFX4 BUFX4_8 ( .A(reset), .Y(reset_bF_buf6));
BUFX4 BUFX4_9 ( .A(reset), .Y(reset_bF_buf5));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock_bF_buf6), .D(_0Rdata_0_0_), .Q(_auto_iopadmap_cc_368_execute_1386_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock_bF_buf4), .D(flip4__0Tx_0_0_), .Q(flip4_Tx));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock_bF_buf3), .D(flip5__0Rx_0_0_), .Q(flip5_Rx));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock_bF_buf2), .D(flip5__0Tx_0_0_), .Q(flip5_Tx));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock_bF_buf1), .D(flip6__0Rx_0_0_), .Q(flip6_Rx));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock_bF_buf0), .D(flip6__0Tx_0_0_), .Q(flip6_Tx));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock_bF_buf6), .D(flip7__0Rx_0_0_), .Q(flip7_Rx));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock_bF_buf5), .D(flip7__0Tx_0_0_), .Q(flip7_Tx));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock_bF_buf4), .D(flip8__0Rx_0_0_), .Q(flip8_Rx));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock_bF_buf3), .D(flip8__0Tx_0_0_), .Q(flip8_Tx));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock_bF_buf2), .D(flipw1__0DS_0_0_), .Q(flipw1_DS));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock_bF_buf5), .D(_0vel_0_0_), .Q(maquina_vel));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock_bF_buf1), .D(flipw1__0outdata_0_0_), .Q(flipw1_outdata));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock_bF_buf0), .D(flipw2__0DS_0_0_), .Q(flipw2_DS));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock_bF_buf6), .D(flipw2__0outdata_0_0_), .Q(flipw2_outdata));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock_bF_buf5), .D(flipw3__0DS_0_0_), .Q(flipw3_DS));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock_bF_buf4), .D(flipw3__0outdata_0_0_), .Q(flipw3_outdata));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock_bF_buf3), .D(flipw4__0DS_0_0_), .Q(flipw4_DS));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock_bF_buf2), .D(flipw4__0outdata_0_0_), .Q(flipw4_outdata));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock_bF_buf1), .D(flipw5__0DS_0_0_), .Q(flipw5_DS));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock_bF_buf0), .D(flipw5__0outdata_0_0_), .Q(flipw5_outdata));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock_bF_buf6), .D(flipw6__0DS_0_0_), .Q(flipw6_DS));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock_bF_buf4), .D(flip1__0Rx_0_0_), .Q(flip1_Rx));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock_bF_buf5), .D(flipw6__0outdata_0_0_), .Q(flipw6_outdata));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock_bF_buf4), .D(flipw7__0DS_0_0_), .Q(flipw7_DS));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock_bF_buf3), .D(flipw7__0outdata_0_0_), .Q(flipw7_outdata));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock_bF_buf2), .D(flipw8__0DS_0_0_), .Q(flipw8_DS));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock_bF_buf1), .D(flipw8__0outdata_0_0_), .Q(flipw8_outdata));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock_bF_buf0), .D(latchR__0LWAddres_2_0__0_), .Q(LRAddress_0_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock_bF_buf6), .D(latchR__0LWAddres_2_0__1_), .Q(LRAddress_1_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock_bF_buf5), .D(latchR__0LWAddres_2_0__2_), .Q(LRAddress_2_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock_bF_buf4), .D(latchW__0LWAddres_2_0__0_), .Q(LWAddress_0_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock_bF_buf3), .D(latchW__0LWAddres_2_0__1_), .Q(LWAddress_1_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock_bF_buf3), .D(flip1__0Tx_0_0_), .Q(flip1_Tx));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock_bF_buf2), .D(latchW__0LWAddres_2_0__2_), .Q(LWAddress_2_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock_bF_buf1), .D(maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_0_), .Q(maquina_state_0_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock_bF_buf0), .D(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_477), .Q(maquina_state_1_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock_bF_buf6), .D(maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_2_), .Q(maquina_state_2_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock_bF_buf5), .D(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_490), .Q(maquina_state_3_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock_bF_buf4), .D(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_494), .Q(maquina_state_4_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock_bF_buf3), .D(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_498), .Q(maquina_state_5_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock_bF_buf2), .D(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_502), .Q(maquina_state_6_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock_bF_buf1), .D(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_506), .Q(maquina_state_7_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock_bF_buf0), .D(maquina__abc_1144_auto_fsm_map_cc_118_implement_pattern_cache_510), .Q(maquina_state_8_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock_bF_buf2), .D(flip2__0Rx_0_0_), .Q(flip2_Rx));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock_bF_buf6), .D(maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_9_), .Q(maquina_state_9_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock_bF_buf5), .D(maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_10_), .Q(maquina_state_10_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock_bF_buf1), .D(flip2__0Tx_0_0_), .Q(flip2_Tx));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock_bF_buf0), .D(flip3__0Rx_0_0_), .Q(flip3_Rx));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock_bF_buf6), .D(flip3__0Tx_0_0_), .Q(flip3_Tx));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock_bF_buf5), .D(flip4__0Rx_0_0_), .Q(flip4_Rx));
INVX1 INVX1_1 ( .A(Wvalid), .Y(_abc_1210_new_n18_));
INVX1 INVX1_10 ( .A(LWAddress_0_), .Y(decow__abc_1242_new_n14_));
INVX1 INVX1_11 ( .A(LWAddress_2_), .Y(decow__abc_1242_new_n16_));
INVX1 INVX1_12 ( .A(flip1_W1), .Y(flip1__abc_1260_new_n8_));
INVX1 INVX1_13 ( .A(reset_bF_buf4), .Y(flip1__abc_1260_new_n11_));
INVX1 INVX1_14 ( .A(flip2_W1), .Y(flip2__abc_1260_new_n8_));
INVX1 INVX1_15 ( .A(reset_bF_buf2), .Y(flip2__abc_1260_new_n11_));
INVX1 INVX1_16 ( .A(flip3_W1), .Y(flip3__abc_1260_new_n8_));
INVX1 INVX1_17 ( .A(reset_bF_buf0), .Y(flip3__abc_1260_new_n11_));
INVX1 INVX1_18 ( .A(flip4_W1), .Y(flip4__abc_1260_new_n8_));
INVX1 INVX1_19 ( .A(reset_bF_buf5), .Y(flip4__abc_1260_new_n11_));
INVX1 INVX1_2 ( .A(reset_bF_buf6), .Y(_abc_1210_new_n20_));
INVX1 INVX1_20 ( .A(flip5_W1), .Y(flip5__abc_1260_new_n8_));
INVX1 INVX1_21 ( .A(reset_bF_buf3), .Y(flip5__abc_1260_new_n11_));
INVX1 INVX1_22 ( .A(flip6_W1), .Y(flip6__abc_1260_new_n8_));
INVX1 INVX1_23 ( .A(reset_bF_buf1), .Y(flip6__abc_1260_new_n11_));
INVX1 INVX1_24 ( .A(flip7_W1), .Y(flip7__abc_1260_new_n8_));
INVX1 INVX1_25 ( .A(reset_bF_buf6), .Y(flip7__abc_1260_new_n11_));
INVX1 INVX1_26 ( .A(flip8_W1), .Y(flip8__abc_1260_new_n8_));
INVX1 INVX1_27 ( .A(reset_bF_buf4), .Y(flip8__abc_1260_new_n11_));
INVX1 INVX1_28 ( .A(flip1_W1), .Y(flipw1__abc_1271_new_n10_));
INVX1 INVX1_29 ( .A(flip2_W1), .Y(flipw2__abc_1271_new_n10_));
INVX1 INVX1_3 ( .A(LRAddress_2_), .Y(_abc_1210_new_n24_));
INVX1 INVX1_30 ( .A(flip3_W1), .Y(flipw3__abc_1271_new_n10_));
INVX1 INVX1_31 ( .A(flip4_W1), .Y(flipw4__abc_1271_new_n10_));
INVX1 INVX1_32 ( .A(flip5_W1), .Y(flipw5__abc_1271_new_n10_));
INVX1 INVX1_33 ( .A(flip6_W1), .Y(flipw6__abc_1271_new_n10_));
INVX1 INVX1_34 ( .A(flip7_W1), .Y(flipw7__abc_1271_new_n10_));
INVX1 INVX1_35 ( .A(flip8_W1), .Y(flipw8__abc_1271_new_n10_));
INVX1 INVX1_36 ( .A(ARvalid), .Y(latchR__abc_1281_new_n13_));
INVX1 INVX1_37 ( .A(AWvalid), .Y(latchW__abc_1281_new_n13_));
INVX1 INVX1_38 ( .A(ARvalid), .Y(maquina__abc_1295_new_n36_));
INVX1 INVX1_39 ( .A(AWvalid), .Y(maquina__abc_1295_new_n37_));
INVX1 INVX1_4 ( .A(LRAddress_1_), .Y(_abc_1210_new_n26_));
INVX1 INVX1_40 ( .A(reset_bF_buf0), .Y(maquina__abc_1295_new_n40_));
INVX1 INVX1_41 ( .A(Wvalid), .Y(maquina__abc_1295_new_n46_));
INVX1 INVX1_42 ( .A(Rready), .Y(maquina__abc_1295_new_n54_));
INVX1 INVX1_43 ( .A(Bready), .Y(maquina__abc_1295_new_n61_));
INVX1 INVX1_44 ( .A(maquina_state_2_), .Y(maquina__abc_1295_new_n67_));
INVX1 INVX1_45 ( .A(maquina_state_8_), .Y(maquina__abc_1295_new_n68_));
INVX1 INVX1_46 ( .A(maquina_state_7_), .Y(maquina__abc_1295_new_n69_));
INVX1 INVX1_47 ( .A(maquina_state_4_), .Y(maquina__abc_1295_new_n72_));
INVX1 INVX1_48 ( .A(maquina_state_0_), .Y(maquina__abc_1295_new_n74_));
INVX1 INVX1_49 ( .A(maquina_state_5_), .Y(maquina__abc_1295_new_n75_));
INVX1 INVX1_5 ( .A(LRAddress_0_), .Y(_abc_1210_new_n27_));
INVX1 INVX1_50 ( .A(maquina__abc_1295_new_n63_), .Y(maquina__abc_1295_new_n83_));
INVX1 INVX1_51 ( .A(maquina__abc_1295_new_n84_), .Y(maquina__abc_1295_new_n85_));
INVX1 INVX1_52 ( .A(maquina__abc_1295_new_n79_), .Y(maquina__abc_1295_new_n87_));
INVX1 INVX1_53 ( .A(maquina_state_3_), .Y(maquina__abc_1295_new_n89_));
INVX1 INVX1_54 ( .A(maquina__abc_1295_new_n92_), .Y(maquina__abc_1295_new_n93_));
INVX1 INVX1_55 ( .A(maquina_vel), .Y(maquina__abc_1295_new_n101_));
INVX1 INVX1_6 ( .A(LRAddress_1_), .Y(decor__abc_1242_new_n13_));
INVX1 INVX1_7 ( .A(LRAddress_0_), .Y(decor__abc_1242_new_n14_));
INVX1 INVX1_8 ( .A(LRAddress_2_), .Y(decor__abc_1242_new_n16_));
INVX1 INVX1_9 ( .A(LWAddress_1_), .Y(decow__abc_1242_new_n13_));
OR2X2 OR2X2_1 ( .A(_abc_1210_new_n21_), .B(_abc_1210_new_n20_), .Y(_abc_1210_new_n22_));
OR2X2 OR2X2_10 ( .A(_abc_1210_new_n42_), .B(_abc_1210_new_n41_), .Y(_abc_1210_new_n43_));
OR2X2 OR2X2_11 ( .A(_abc_1210_new_n43_), .B(LRAddress_1_), .Y(_abc_1210_new_n44_));
OR2X2 OR2X2_12 ( .A(_abc_1210_new_n45_), .B(LRAddress_2_), .Y(_abc_1210_new_n46_));
OR2X2 OR2X2_13 ( .A(flip1__abc_1260_new_n8_), .B(flip1_R1), .Y(flip1__abc_1260_new_n9_));
OR2X2 OR2X2_14 ( .A(flip1__abc_1260_new_n12_), .B(flip1__abc_1260_new_n11_), .Y(flip1__abc_1260_new_n13_));
OR2X2 OR2X2_15 ( .A(flip1__abc_1260_new_n10_), .B(flip1__abc_1260_new_n13_), .Y(flip1__0Tx_0_0_));
OR2X2 OR2X2_16 ( .A(flip1__abc_1260_new_n12_), .B(flip1_Rx), .Y(flip1__abc_1260_new_n15_));
OR2X2 OR2X2_17 ( .A(flip2__abc_1260_new_n8_), .B(flip2_R1), .Y(flip2__abc_1260_new_n9_));
OR2X2 OR2X2_18 ( .A(flip2__abc_1260_new_n12_), .B(flip2__abc_1260_new_n11_), .Y(flip2__abc_1260_new_n13_));
OR2X2 OR2X2_19 ( .A(flip2__abc_1260_new_n10_), .B(flip2__abc_1260_new_n13_), .Y(flip2__0Tx_0_0_));
OR2X2 OR2X2_2 ( .A(_abc_1210_new_n22_), .B(_abc_1210_new_n19_), .Y(_0vel_0_0_));
OR2X2 OR2X2_20 ( .A(flip2__abc_1260_new_n12_), .B(flip2_Rx), .Y(flip2__abc_1260_new_n15_));
OR2X2 OR2X2_21 ( .A(flip3__abc_1260_new_n8_), .B(flip3_R1), .Y(flip3__abc_1260_new_n9_));
OR2X2 OR2X2_22 ( .A(flip3__abc_1260_new_n12_), .B(flip3__abc_1260_new_n11_), .Y(flip3__abc_1260_new_n13_));
OR2X2 OR2X2_23 ( .A(flip3__abc_1260_new_n10_), .B(flip3__abc_1260_new_n13_), .Y(flip3__0Tx_0_0_));
OR2X2 OR2X2_24 ( .A(flip3__abc_1260_new_n12_), .B(flip3_Rx), .Y(flip3__abc_1260_new_n15_));
OR2X2 OR2X2_25 ( .A(flip4__abc_1260_new_n8_), .B(flip4_R1), .Y(flip4__abc_1260_new_n9_));
OR2X2 OR2X2_26 ( .A(flip4__abc_1260_new_n12_), .B(flip4__abc_1260_new_n11_), .Y(flip4__abc_1260_new_n13_));
OR2X2 OR2X2_27 ( .A(flip4__abc_1260_new_n10_), .B(flip4__abc_1260_new_n13_), .Y(flip4__0Tx_0_0_));
OR2X2 OR2X2_28 ( .A(flip4__abc_1260_new_n12_), .B(flip4_Rx), .Y(flip4__abc_1260_new_n15_));
OR2X2 OR2X2_29 ( .A(flip5__abc_1260_new_n8_), .B(flip5_R1), .Y(flip5__abc_1260_new_n9_));
OR2X2 OR2X2_3 ( .A(_abc_1210_new_n28_), .B(_abc_1210_new_n26_), .Y(_abc_1210_new_n29_));
OR2X2 OR2X2_30 ( .A(flip5__abc_1260_new_n12_), .B(flip5__abc_1260_new_n11_), .Y(flip5__abc_1260_new_n13_));
OR2X2 OR2X2_31 ( .A(flip5__abc_1260_new_n10_), .B(flip5__abc_1260_new_n13_), .Y(flip5__0Tx_0_0_));
OR2X2 OR2X2_32 ( .A(flip5__abc_1260_new_n12_), .B(flip5_Rx), .Y(flip5__abc_1260_new_n15_));
OR2X2 OR2X2_33 ( .A(flip6__abc_1260_new_n8_), .B(flip6_R1), .Y(flip6__abc_1260_new_n9_));
OR2X2 OR2X2_34 ( .A(flip6__abc_1260_new_n12_), .B(flip6__abc_1260_new_n11_), .Y(flip6__abc_1260_new_n13_));
OR2X2 OR2X2_35 ( .A(flip6__abc_1260_new_n10_), .B(flip6__abc_1260_new_n13_), .Y(flip6__0Tx_0_0_));
OR2X2 OR2X2_36 ( .A(flip6__abc_1260_new_n12_), .B(flip6_Rx), .Y(flip6__abc_1260_new_n15_));
OR2X2 OR2X2_37 ( .A(flip7__abc_1260_new_n8_), .B(flip7_R1), .Y(flip7__abc_1260_new_n9_));
OR2X2 OR2X2_38 ( .A(flip7__abc_1260_new_n12_), .B(flip7__abc_1260_new_n11_), .Y(flip7__abc_1260_new_n13_));
OR2X2 OR2X2_39 ( .A(flip7__abc_1260_new_n10_), .B(flip7__abc_1260_new_n13_), .Y(flip7__0Tx_0_0_));
OR2X2 OR2X2_4 ( .A(_abc_1210_new_n29_), .B(_abc_1210_new_n25_), .Y(_abc_1210_new_n30_));
OR2X2 OR2X2_40 ( .A(flip7__abc_1260_new_n12_), .B(flip7_Rx), .Y(flip7__abc_1260_new_n15_));
OR2X2 OR2X2_41 ( .A(flip8__abc_1260_new_n8_), .B(flip8_R1), .Y(flip8__abc_1260_new_n9_));
OR2X2 OR2X2_42 ( .A(flip8__abc_1260_new_n12_), .B(flip8__abc_1260_new_n11_), .Y(flip8__abc_1260_new_n13_));
OR2X2 OR2X2_43 ( .A(flip8__abc_1260_new_n10_), .B(flip8__abc_1260_new_n13_), .Y(flip8__0Tx_0_0_));
OR2X2 OR2X2_44 ( .A(flip8__abc_1260_new_n12_), .B(flip8_Rx), .Y(flip8__abc_1260_new_n15_));
OR2X2 OR2X2_45 ( .A(flipw1__abc_1271_new_n11_), .B(flipw1__abc_1271_new_n9_), .Y(flipw1__abc_1271_new_n12_));
OR2X2 OR2X2_46 ( .A(flipw1__abc_1271_new_n15_), .B(flipw1__abc_1271_new_n14_), .Y(flipw1__abc_1271_new_n16_));
OR2X2 OR2X2_47 ( .A(flipw2__abc_1271_new_n11_), .B(flipw2__abc_1271_new_n9_), .Y(flipw2__abc_1271_new_n12_));
OR2X2 OR2X2_48 ( .A(flipw2__abc_1271_new_n15_), .B(flipw2__abc_1271_new_n14_), .Y(flipw2__abc_1271_new_n16_));
OR2X2 OR2X2_49 ( .A(flipw3__abc_1271_new_n11_), .B(flipw3__abc_1271_new_n9_), .Y(flipw3__abc_1271_new_n12_));
OR2X2 OR2X2_5 ( .A(_abc_1210_new_n32_), .B(_abc_1210_new_n31_), .Y(_abc_1210_new_n33_));
OR2X2 OR2X2_50 ( .A(flipw3__abc_1271_new_n15_), .B(flipw3__abc_1271_new_n14_), .Y(flipw3__abc_1271_new_n16_));
OR2X2 OR2X2_51 ( .A(flipw4__abc_1271_new_n11_), .B(flipw4__abc_1271_new_n9_), .Y(flipw4__abc_1271_new_n12_));
OR2X2 OR2X2_52 ( .A(flipw4__abc_1271_new_n15_), .B(flipw4__abc_1271_new_n14_), .Y(flipw4__abc_1271_new_n16_));
OR2X2 OR2X2_53 ( .A(flipw5__abc_1271_new_n11_), .B(flipw5__abc_1271_new_n9_), .Y(flipw5__abc_1271_new_n12_));
OR2X2 OR2X2_54 ( .A(flipw5__abc_1271_new_n15_), .B(flipw5__abc_1271_new_n14_), .Y(flipw5__abc_1271_new_n16_));
OR2X2 OR2X2_55 ( .A(flipw6__abc_1271_new_n11_), .B(flipw6__abc_1271_new_n9_), .Y(flipw6__abc_1271_new_n12_));
OR2X2 OR2X2_56 ( .A(flipw6__abc_1271_new_n15_), .B(flipw6__abc_1271_new_n14_), .Y(flipw6__abc_1271_new_n16_));
OR2X2 OR2X2_57 ( .A(flipw7__abc_1271_new_n11_), .B(flipw7__abc_1271_new_n9_), .Y(flipw7__abc_1271_new_n12_));
OR2X2 OR2X2_58 ( .A(flipw7__abc_1271_new_n15_), .B(flipw7__abc_1271_new_n14_), .Y(flipw7__abc_1271_new_n16_));
OR2X2 OR2X2_59 ( .A(flipw8__abc_1271_new_n11_), .B(flipw8__abc_1271_new_n9_), .Y(flipw8__abc_1271_new_n12_));
OR2X2 OR2X2_6 ( .A(_abc_1210_new_n33_), .B(LRAddress_1_), .Y(_abc_1210_new_n34_));
OR2X2 OR2X2_60 ( .A(flipw8__abc_1271_new_n15_), .B(flipw8__abc_1271_new_n14_), .Y(flipw8__abc_1271_new_n16_));
OR2X2 OR2X2_61 ( .A(latchR__abc_1281_new_n14_), .B(latchR__abc_1281_new_n12_), .Y(latchR__abc_1281_new_n15_));
OR2X2 OR2X2_62 ( .A(latchR__abc_1281_new_n18_), .B(latchR__abc_1281_new_n17_), .Y(latchR__abc_1281_new_n19_));
OR2X2 OR2X2_63 ( .A(latchR__abc_1281_new_n22_), .B(latchR__abc_1281_new_n21_), .Y(latchR__abc_1281_new_n23_));
OR2X2 OR2X2_64 ( .A(latchW__abc_1281_new_n14_), .B(latchW__abc_1281_new_n12_), .Y(latchW__abc_1281_new_n15_));
OR2X2 OR2X2_65 ( .A(latchW__abc_1281_new_n18_), .B(latchW__abc_1281_new_n17_), .Y(latchW__abc_1281_new_n19_));
OR2X2 OR2X2_66 ( .A(latchW__abc_1281_new_n22_), .B(latchW__abc_1281_new_n21_), .Y(latchW__abc_1281_new_n23_));
OR2X2 OR2X2_67 ( .A(maquina__abc_1295_new_n41_), .B(maquina__abc_1295_new_n40_), .Y(maquina__abc_1295_new_n42_));
OR2X2 OR2X2_68 ( .A(maquina__abc_1295_new_n42_), .B(maquina__abc_1295_new_n43_), .Y(maquina__abc_1295_new_n44_));
OR2X2 OR2X2_69 ( .A(maquina__abc_1295_new_n44_), .B(maquina__abc_1295_new_n39_), .Y(maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_0_));
OR2X2 OR2X2_7 ( .A(_abc_1210_new_n35_), .B(_abc_1210_new_n24_), .Y(_abc_1210_new_n36_));
OR2X2 OR2X2_70 ( .A(maquina__abc_1295_new_n50_), .B(maquina__abc_1295_new_n48_), .Y(maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_2_));
OR2X2 OR2X2_71 ( .A(maquina__abc_1295_new_n54_), .B(maquina_state_3_), .Y(maquina__abc_1295_new_n55_));
OR2X2 OR2X2_72 ( .A(maquina_state_9_), .B(maquina_state_3_), .Y(maquina__abc_1295_new_n56_));
OR2X2 OR2X2_73 ( .A(maquina__abc_1295_new_n58_), .B(maquina__abc_1295_new_n53_), .Y(maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_9_));
OR2X2 OR2X2_74 ( .A(maquina__abc_1295_new_n61_), .B(maquina_state_4_), .Y(maquina__abc_1295_new_n62_));
OR2X2 OR2X2_75 ( .A(maquina_state_10_), .B(maquina_state_4_), .Y(maquina__abc_1295_new_n63_));
OR2X2 OR2X2_76 ( .A(maquina__abc_1295_new_n65_), .B(maquina__abc_1295_new_n60_), .Y(maquina__abc_1144_auto_fsm_map_cc_170_map_fsm_456_10_));
OR2X2 OR2X2_77 ( .A(maquina__abc_1295_new_n63_), .B(maquina_state_7_), .Y(maquina__abc_1295_new_n79_));
OR2X2 OR2X2_78 ( .A(maquina__abc_1295_new_n80_), .B(maquina_state_8_), .Y(maquina__abc_1295_new_n81_));
OR2X2 OR2X2_79 ( .A(maquina_state_6_), .B(maquina_state_1_), .Y(maquina__abc_1295_new_n92_));
OR2X2 OR2X2_8 ( .A(_abc_1210_new_n38_), .B(_abc_1210_new_n26_), .Y(_abc_1210_new_n39_));
OR2X2 OR2X2_80 ( .A(maquina__abc_1295_new_n56_), .B(maquina__abc_1295_new_n92_), .Y(maquina__abc_1295_new_n97_));
OR2X2 OR2X2_81 ( .A(maquina__abc_1295_new_n98_), .B(maquina_state_5_), .Y(maquina__abc_1295_new_n99_));
OR2X2 OR2X2_9 ( .A(_abc_1210_new_n39_), .B(_abc_1210_new_n37_), .Y(_abc_1210_new_n40_));


endmodule