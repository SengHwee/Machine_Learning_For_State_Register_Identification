module uart(clk, rst, rx, transmit, \tx_byte[0] , \tx_byte[1] , \tx_byte[2] , \tx_byte[3] , \tx_byte[4] , \tx_byte[5] , \tx_byte[6] , \tx_byte[7] , tx, received, \rx_byte[0] , \rx_byte[1] , \rx_byte[2] , \rx_byte[3] , \rx_byte[4] , \rx_byte[5] , \rx_byte[6] , \rx_byte[7] , is_receiving, is_transmitting, recv_error);

wire _0recv_state_2_0__0_; 
wire _0recv_state_2_0__1_; 
wire _0recv_state_2_0__2_; 
wire _0rx_bits_remaining_3_0__0_; 
wire _0rx_bits_remaining_3_0__1_; 
wire _0rx_bits_remaining_3_0__2_; 
wire _0rx_bits_remaining_3_0__3_; 
wire _0rx_clk_divider_10_0__0_; 
wire _0rx_clk_divider_10_0__10_; 
wire _0rx_clk_divider_10_0__1_; 
wire _0rx_clk_divider_10_0__2_; 
wire _0rx_clk_divider_10_0__3_; 
wire _0rx_clk_divider_10_0__4_; 
wire _0rx_clk_divider_10_0__5_; 
wire _0rx_clk_divider_10_0__6_; 
wire _0rx_clk_divider_10_0__7_; 
wire _0rx_clk_divider_10_0__8_; 
wire _0rx_clk_divider_10_0__9_; 
wire _0rx_countdown_5_0__0_; 
wire _0rx_countdown_5_0__1_; 
wire _0rx_countdown_5_0__2_; 
wire _0rx_countdown_5_0__3_; 
wire _0rx_countdown_5_0__4_; 
wire _0rx_countdown_5_0__5_; 
wire _0rx_data_7_0__0_; 
wire _0rx_data_7_0__1_; 
wire _0rx_data_7_0__2_; 
wire _0rx_data_7_0__3_; 
wire _0rx_data_7_0__4_; 
wire _0rx_data_7_0__5_; 
wire _0rx_data_7_0__6_; 
wire _0rx_data_7_0__7_; 
wire _0tx_bits_remaining_3_0__0_; 
wire _0tx_bits_remaining_3_0__1_; 
wire _0tx_bits_remaining_3_0__2_; 
wire _0tx_bits_remaining_3_0__3_; 
wire _0tx_clk_divider_10_0__0_; 
wire _0tx_clk_divider_10_0__10_; 
wire _0tx_clk_divider_10_0__1_; 
wire _0tx_clk_divider_10_0__2_; 
wire _0tx_clk_divider_10_0__3_; 
wire _0tx_clk_divider_10_0__4_; 
wire _0tx_clk_divider_10_0__5_; 
wire _0tx_clk_divider_10_0__6_; 
wire _0tx_clk_divider_10_0__7_; 
wire _0tx_clk_divider_10_0__8_; 
wire _0tx_clk_divider_10_0__9_; 
wire _0tx_countdown_5_0__0_; 
wire _0tx_countdown_5_0__1_; 
wire _0tx_countdown_5_0__2_; 
wire _0tx_countdown_5_0__3_; 
wire _0tx_countdown_5_0__4_; 
wire _0tx_countdown_5_0__5_; 
wire _0tx_data_7_0__0_; 
wire _0tx_data_7_0__1_; 
wire _0tx_data_7_0__2_; 
wire _0tx_data_7_0__3_; 
wire _0tx_data_7_0__4_; 
wire _0tx_data_7_0__5_; 
wire _0tx_data_7_0__6_; 
wire _0tx_data_7_0__7_; 
wire _0tx_out_0_0_; 
wire _0tx_state_1_0__0_; 
wire _0tx_state_1_0__1_; 
wire _abc_2284_new_n144_; 
wire _abc_2284_new_n145_; 
wire _abc_2284_new_n147_; 
wire _abc_2284_new_n148_; 
wire _abc_2284_new_n150_; 
wire _abc_2284_new_n152_; 
wire _abc_2284_new_n154_; 
wire _abc_2284_new_n155_; 
wire _abc_2284_new_n156_; 
wire _abc_2284_new_n157_; 
wire _abc_2284_new_n158_; 
wire _abc_2284_new_n159_; 
wire _abc_2284_new_n160_; 
wire _abc_2284_new_n161_; 
wire _abc_2284_new_n162_; 
wire _abc_2284_new_n163_; 
wire _abc_2284_new_n164_; 
wire _abc_2284_new_n165_; 
wire _abc_2284_new_n166_; 
wire _abc_2284_new_n167_; 
wire _abc_2284_new_n168_; 
wire _abc_2284_new_n169_; 
wire _abc_2284_new_n170_; 
wire _abc_2284_new_n171_; 
wire _abc_2284_new_n172_; 
wire _abc_2284_new_n173_; 
wire _abc_2284_new_n174_; 
wire _abc_2284_new_n175_; 
wire _abc_2284_new_n176_; 
wire _abc_2284_new_n177_; 
wire _abc_2284_new_n178_; 
wire _abc_2284_new_n179_; 
wire _abc_2284_new_n180_; 
wire _abc_2284_new_n181_; 
wire _abc_2284_new_n182_; 
wire _abc_2284_new_n183_; 
wire _abc_2284_new_n184_; 
wire _abc_2284_new_n185_; 
wire _abc_2284_new_n186_; 
wire _abc_2284_new_n187_; 
wire _abc_2284_new_n188_; 
wire _abc_2284_new_n189_; 
wire _abc_2284_new_n190_; 
wire _abc_2284_new_n191_; 
wire _abc_2284_new_n192_; 
wire _abc_2284_new_n193_; 
wire _abc_2284_new_n194_; 
wire _abc_2284_new_n195_; 
wire _abc_2284_new_n196_; 
wire _abc_2284_new_n197_; 
wire _abc_2284_new_n198_; 
wire _abc_2284_new_n199_; 
wire _abc_2284_new_n200_; 
wire _abc_2284_new_n201_; 
wire _abc_2284_new_n202_; 
wire _abc_2284_new_n203_; 
wire _abc_2284_new_n204_; 
wire _abc_2284_new_n205_; 
wire _abc_2284_new_n206_; 
wire _abc_2284_new_n207_; 
wire _abc_2284_new_n208_; 
wire _abc_2284_new_n209_; 
wire _abc_2284_new_n210_; 
wire _abc_2284_new_n211_; 
wire _abc_2284_new_n212_; 
wire _abc_2284_new_n213_; 
wire _abc_2284_new_n214_; 
wire _abc_2284_new_n215_; 
wire _abc_2284_new_n216_; 
wire _abc_2284_new_n217_; 
wire _abc_2284_new_n218_; 
wire _abc_2284_new_n219_; 
wire _abc_2284_new_n220_; 
wire _abc_2284_new_n221_; 
wire _abc_2284_new_n222_; 
wire _abc_2284_new_n223_; 
wire _abc_2284_new_n224_; 
wire _abc_2284_new_n225_; 
wire _abc_2284_new_n226_; 
wire _abc_2284_new_n227_; 
wire _abc_2284_new_n228_; 
wire _abc_2284_new_n229_; 
wire _abc_2284_new_n230_; 
wire _abc_2284_new_n231_; 
wire _abc_2284_new_n232_; 
wire _abc_2284_new_n233_; 
wire _abc_2284_new_n234_; 
wire _abc_2284_new_n235_; 
wire _abc_2284_new_n236_; 
wire _abc_2284_new_n237_; 
wire _abc_2284_new_n238_; 
wire _abc_2284_new_n239_; 
wire _abc_2284_new_n240_; 
wire _abc_2284_new_n241_; 
wire _abc_2284_new_n242_; 
wire _abc_2284_new_n243_; 
wire _abc_2284_new_n244_; 
wire _abc_2284_new_n245_; 
wire _abc_2284_new_n246_; 
wire _abc_2284_new_n247_; 
wire _abc_2284_new_n248_; 
wire _abc_2284_new_n249_; 
wire _abc_2284_new_n250_; 
wire _abc_2284_new_n251_; 
wire _abc_2284_new_n252_; 
wire _abc_2284_new_n253_; 
wire _abc_2284_new_n254_; 
wire _abc_2284_new_n255_; 
wire _abc_2284_new_n256_; 
wire _abc_2284_new_n257_; 
wire _abc_2284_new_n258_; 
wire _abc_2284_new_n259_; 
wire _abc_2284_new_n260_; 
wire _abc_2284_new_n261_; 
wire _abc_2284_new_n262_; 
wire _abc_2284_new_n264_; 
wire _abc_2284_new_n265_; 
wire _abc_2284_new_n266_; 
wire _abc_2284_new_n267_; 
wire _abc_2284_new_n268_; 
wire _abc_2284_new_n269_; 
wire _abc_2284_new_n270_; 
wire _abc_2284_new_n272_; 
wire _abc_2284_new_n273_; 
wire _abc_2284_new_n274_; 
wire _abc_2284_new_n275_; 
wire _abc_2284_new_n276_; 
wire _abc_2284_new_n277_; 
wire _abc_2284_new_n278_; 
wire _abc_2284_new_n280_; 
wire _abc_2284_new_n281_; 
wire _abc_2284_new_n282_; 
wire _abc_2284_new_n283_; 
wire _abc_2284_new_n284_; 
wire _abc_2284_new_n285_; 
wire _abc_2284_new_n286_; 
wire _abc_2284_new_n288_; 
wire _abc_2284_new_n289_; 
wire _abc_2284_new_n290_; 
wire _abc_2284_new_n291_; 
wire _abc_2284_new_n292_; 
wire _abc_2284_new_n293_; 
wire _abc_2284_new_n294_; 
wire _abc_2284_new_n296_; 
wire _abc_2284_new_n297_; 
wire _abc_2284_new_n298_; 
wire _abc_2284_new_n299_; 
wire _abc_2284_new_n300_; 
wire _abc_2284_new_n301_; 
wire _abc_2284_new_n302_; 
wire _abc_2284_new_n304_; 
wire _abc_2284_new_n305_; 
wire _abc_2284_new_n306_; 
wire _abc_2284_new_n307_; 
wire _abc_2284_new_n308_; 
wire _abc_2284_new_n309_; 
wire _abc_2284_new_n310_; 
wire _abc_2284_new_n312_; 
wire _abc_2284_new_n313_; 
wire _abc_2284_new_n314_; 
wire _abc_2284_new_n315_; 
wire _abc_2284_new_n316_; 
wire _abc_2284_new_n317_; 
wire _abc_2284_new_n319_; 
wire _abc_2284_new_n320_; 
wire _abc_2284_new_n321_; 
wire _abc_2284_new_n322_; 
wire _abc_2284_new_n323_; 
wire _abc_2284_new_n324_; 
wire _abc_2284_new_n325_; 
wire _abc_2284_new_n326_; 
wire _abc_2284_new_n327_; 
wire _abc_2284_new_n328_; 
wire _abc_2284_new_n330_; 
wire _abc_2284_new_n331_; 
wire _abc_2284_new_n332_; 
wire _abc_2284_new_n333_; 
wire _abc_2284_new_n334_; 
wire _abc_2284_new_n335_; 
wire _abc_2284_new_n336_; 
wire _abc_2284_new_n337_; 
wire _abc_2284_new_n339_; 
wire _abc_2284_new_n340_; 
wire _abc_2284_new_n341_; 
wire _abc_2284_new_n342_; 
wire _abc_2284_new_n343_; 
wire _abc_2284_new_n344_; 
wire _abc_2284_new_n345_; 
wire _abc_2284_new_n346_; 
wire _abc_2284_new_n347_; 
wire _abc_2284_new_n349_; 
wire _abc_2284_new_n350_; 
wire _abc_2284_new_n351_; 
wire _abc_2284_new_n352_; 
wire _abc_2284_new_n353_; 
wire _abc_2284_new_n354_; 
wire _abc_2284_new_n355_; 
wire _abc_2284_new_n356_; 
wire _abc_2284_new_n360_; 
wire _abc_2284_new_n362_; 
wire _abc_2284_new_n363_; 
wire _abc_2284_new_n367_; 
wire _abc_2284_new_n369_; 
wire _abc_2284_new_n371_; 
wire _abc_2284_new_n372_; 
wire _abc_2284_new_n373_; 
wire _abc_2284_new_n374_; 
wire _abc_2284_new_n376_; 
wire _abc_2284_new_n377_; 
wire _abc_2284_new_n378_; 
wire _abc_2284_new_n379_; 
wire _abc_2284_new_n380_; 
wire _abc_2284_new_n381_; 
wire _abc_2284_new_n382_; 
wire _abc_2284_new_n383_; 
wire _abc_2284_new_n384_; 
wire _abc_2284_new_n385_; 
wire _abc_2284_new_n386_; 
wire _abc_2284_new_n387_; 
wire _abc_2284_new_n388_; 
wire _abc_2284_new_n389_; 
wire _abc_2284_new_n390_; 
wire _abc_2284_new_n391_; 
wire _abc_2284_new_n392_; 
wire _abc_2284_new_n393_; 
wire _abc_2284_new_n394_; 
wire _abc_2284_new_n395_; 
wire _abc_2284_new_n396_; 
wire _abc_2284_new_n397_; 
wire _abc_2284_new_n398_; 
wire _abc_2284_new_n399_; 
wire _abc_2284_new_n400_; 
wire _abc_2284_new_n401_; 
wire _abc_2284_new_n402_; 
wire _abc_2284_new_n403_; 
wire _abc_2284_new_n404_; 
wire _abc_2284_new_n405_; 
wire _abc_2284_new_n406_; 
wire _abc_2284_new_n407_; 
wire _abc_2284_new_n408_; 
wire _abc_2284_new_n409_; 
wire _abc_2284_new_n410_; 
wire _abc_2284_new_n411_; 
wire _abc_2284_new_n412_; 
wire _abc_2284_new_n413_; 
wire _abc_2284_new_n414_; 
wire _abc_2284_new_n415_; 
wire _abc_2284_new_n416_; 
wire _abc_2284_new_n417_; 
wire _abc_2284_new_n418_; 
wire _abc_2284_new_n419_; 
wire _abc_2284_new_n420_; 
wire _abc_2284_new_n421_; 
wire _abc_2284_new_n422_; 
wire _abc_2284_new_n423_; 
wire _abc_2284_new_n424_; 
wire _abc_2284_new_n425_; 
wire _abc_2284_new_n426_; 
wire _abc_2284_new_n428_; 
wire _abc_2284_new_n429_; 
wire _abc_2284_new_n430_; 
wire _abc_2284_new_n431_; 
wire _abc_2284_new_n432_; 
wire _abc_2284_new_n433_; 
wire _abc_2284_new_n434_; 
wire _abc_2284_new_n435_; 
wire _abc_2284_new_n436_; 
wire _abc_2284_new_n437_; 
wire _abc_2284_new_n438_; 
wire _abc_2284_new_n439_; 
wire _abc_2284_new_n440_; 
wire _abc_2284_new_n441_; 
wire _abc_2284_new_n442_; 
wire _abc_2284_new_n443_; 
wire _abc_2284_new_n444_; 
wire _abc_2284_new_n445_; 
wire _abc_2284_new_n447_; 
wire _abc_2284_new_n448_; 
wire _abc_2284_new_n449_; 
wire _abc_2284_new_n450_; 
wire _abc_2284_new_n451_; 
wire _abc_2284_new_n452_; 
wire _abc_2284_new_n453_; 
wire _abc_2284_new_n454_; 
wire _abc_2284_new_n455_; 
wire _abc_2284_new_n456_; 
wire _abc_2284_new_n457_; 
wire _abc_2284_new_n458_; 
wire _abc_2284_new_n459_; 
wire _abc_2284_new_n460_; 
wire _abc_2284_new_n461_; 
wire _abc_2284_new_n462_; 
wire _abc_2284_new_n463_; 
wire _abc_2284_new_n464_; 
wire _abc_2284_new_n465_; 
wire _abc_2284_new_n466_; 
wire _abc_2284_new_n467_; 
wire _abc_2284_new_n468_; 
wire _abc_2284_new_n469_; 
wire _abc_2284_new_n470_; 
wire _abc_2284_new_n471_; 
wire _abc_2284_new_n472_; 
wire _abc_2284_new_n473_; 
wire _abc_2284_new_n474_; 
wire _abc_2284_new_n475_; 
wire _abc_2284_new_n476_; 
wire _abc_2284_new_n477_; 
wire _abc_2284_new_n478_; 
wire _abc_2284_new_n479_; 
wire _abc_2284_new_n481_; 
wire _abc_2284_new_n483_; 
wire _abc_2284_new_n484_; 
wire _abc_2284_new_n487_; 
wire _abc_2284_new_n488_; 
wire _abc_2284_new_n489_; 
wire _abc_2284_new_n490_; 
wire _abc_2284_new_n491_; 
wire _abc_2284_new_n492_; 
wire _abc_2284_new_n493_; 
wire _abc_2284_new_n494_; 
wire _abc_2284_new_n495_; 
wire _abc_2284_new_n496_; 
wire _abc_2284_new_n497_; 
wire _abc_2284_new_n498_; 
wire _abc_2284_new_n499_; 
wire _abc_2284_new_n500_; 
wire _abc_2284_new_n501_; 
wire _abc_2284_new_n502_; 
wire _abc_2284_new_n503_; 
wire _abc_2284_new_n504_; 
wire _abc_2284_new_n505_; 
wire _abc_2284_new_n506_; 
wire _abc_2284_new_n507_; 
wire _abc_2284_new_n508_; 
wire _abc_2284_new_n509_; 
wire _abc_2284_new_n510_; 
wire _abc_2284_new_n511_; 
wire _abc_2284_new_n512_; 
wire _abc_2284_new_n514_; 
wire _abc_2284_new_n515_; 
wire _abc_2284_new_n516_; 
wire _abc_2284_new_n517_; 
wire _abc_2284_new_n518_; 
wire _abc_2284_new_n520_; 
wire _abc_2284_new_n521_; 
wire _abc_2284_new_n522_; 
wire _abc_2284_new_n523_; 
wire _abc_2284_new_n525_; 
wire _abc_2284_new_n526_; 
wire _abc_2284_new_n527_; 
wire _abc_2284_new_n528_; 
wire _abc_2284_new_n529_; 
wire _abc_2284_new_n531_; 
wire _abc_2284_new_n532_; 
wire _abc_2284_new_n533_; 
wire _abc_2284_new_n535_; 
wire _abc_2284_new_n536_; 
wire _abc_2284_new_n537_; 
wire _abc_2284_new_n538_; 
wire _abc_2284_new_n539_; 
wire _abc_2284_new_n541_; 
wire _abc_2284_new_n542_; 
wire _abc_2284_new_n543_; 
wire _abc_2284_new_n544_; 
wire _abc_2284_new_n545_; 
wire _abc_2284_new_n546_; 
wire _abc_2284_new_n547_; 
wire _abc_2284_new_n550_; 
wire _abc_2284_new_n551_; 
wire _abc_2284_new_n553_; 
wire _abc_2284_new_n555_; 
wire _abc_2284_new_n556_; 
wire _abc_2284_new_n558_; 
wire _abc_2284_new_n559_; 
wire _abc_2284_new_n560_; 
wire _abc_2284_new_n562_; 
wire _abc_2284_new_n565_; 
wire _abc_2284_new_n566_; 
wire _abc_2284_new_n568_; 
wire _abc_2284_new_n570_; 
wire _abc_2284_new_n574_; 
wire _abc_2284_new_n575_; 
wire _abc_2284_new_n577_; 
wire _abc_2284_new_n579_; 
wire _abc_2284_new_n581_; 
wire _abc_2284_new_n583_; 
wire _abc_2284_new_n587_; 
wire _abc_2284_new_n590_; 
wire _abc_2284_new_n592_; 
wire _abc_2284_new_n593_; 
wire _abc_2284_new_n595_; 
wire _abc_2284_new_n597_; 
wire _abc_2284_new_n599_; 
wire _abc_2284_new_n601_; 
wire _abc_2284_new_n603_; 
wire _abc_2284_new_n605_; 
wire _abc_2284_new_n607_; 
input clk;
output is_receiving;
output is_transmitting;
output received;
output recv_error;
wire recv_state_0_; 
wire recv_state_1_; 
wire recv_state_2_; 
input rst;
input rx;
wire rx_bits_remaining_0_; 
wire rx_bits_remaining_1_; 
wire rx_bits_remaining_2_; 
wire rx_bits_remaining_3_; 
output \rx_byte[0] ;
output \rx_byte[1] ;
output \rx_byte[2] ;
output \rx_byte[3] ;
output \rx_byte[4] ;
output \rx_byte[5] ;
output \rx_byte[6] ;
output \rx_byte[7] ;
wire rx_clk_divider_0_; 
wire rx_clk_divider_10_; 
wire rx_clk_divider_1_; 
wire rx_clk_divider_2_; 
wire rx_clk_divider_3_; 
wire rx_clk_divider_4_; 
wire rx_clk_divider_5_; 
wire rx_clk_divider_6_; 
wire rx_clk_divider_7_; 
wire rx_clk_divider_8_; 
wire rx_clk_divider_9_; 
wire rx_countdown_0_; 
wire rx_countdown_1_; 
wire rx_countdown_2_; 
wire rx_countdown_3_; 
wire rx_countdown_4_; 
wire rx_countdown_5_; 
input transmit;
output tx;
wire tx_bits_remaining_0_; 
wire tx_bits_remaining_1_; 
wire tx_bits_remaining_2_; 
wire tx_bits_remaining_3_; 
input \tx_byte[0] ;
input \tx_byte[1] ;
input \tx_byte[2] ;
input \tx_byte[3] ;
input \tx_byte[4] ;
input \tx_byte[5] ;
input \tx_byte[6] ;
input \tx_byte[7] ;
wire tx_clk_divider_0_; 
wire tx_clk_divider_10_; 
wire tx_clk_divider_1_; 
wire tx_clk_divider_2_; 
wire tx_clk_divider_3_; 
wire tx_clk_divider_4_; 
wire tx_clk_divider_5_; 
wire tx_clk_divider_6_; 
wire tx_clk_divider_7_; 
wire tx_clk_divider_8_; 
wire tx_clk_divider_9_; 
wire tx_countdown_0_; 
wire tx_countdown_1_; 
wire tx_countdown_2_; 
wire tx_countdown_3_; 
wire tx_countdown_4_; 
wire tx_countdown_5_; 
wire tx_data_0_; 
wire tx_data_1_; 
wire tx_data_2_; 
wire tx_data_3_; 
wire tx_data_4_; 
wire tx_data_5_; 
wire tx_data_6_; 
wire tx_data_7_; 
wire tx_state_0_; 
wire tx_state_1_; 
AND2X2 AND2X2_1 ( .A(_abc_2284_new_n158_), .B(_abc_2284_new_n159_), .Y(_abc_2284_new_n160_));
AND2X2 AND2X2_10 ( .A(tx_clk_divider_1_), .B(tx_clk_divider_0_), .Y(_abc_2284_new_n550_));
AND2X2 AND2X2_11 ( .A(_abc_2284_new_n173_), .B(_abc_2284_new_n174_), .Y(_abc_2284_new_n568_));
AND2X2 AND2X2_12 ( .A(_abc_2284_new_n396_), .B(_abc_2284_new_n397_), .Y(_abc_2284_new_n587_));
AND2X2 AND2X2_2 ( .A(_abc_2284_new_n161_), .B(_abc_2284_new_n162_), .Y(_abc_2284_new_n163_));
AND2X2 AND2X2_3 ( .A(_abc_2284_new_n191_), .B(_abc_2284_new_n176_), .Y(_abc_2284_new_n192_));
AND2X2 AND2X2_4 ( .A(_abc_2284_new_n183_), .B(tx_clk_divider_6_), .Y(_abc_2284_new_n203_));
AND2X2 AND2X2_5 ( .A(_abc_2284_new_n227_), .B(_abc_2284_new_n349_), .Y(_0tx_countdown_5_0__5_));
AND2X2 AND2X2_6 ( .A(_abc_2284_new_n377_), .B(_abc_2284_new_n378_), .Y(_abc_2284_new_n379_));
AND2X2 AND2X2_7 ( .A(_abc_2284_new_n430_), .B(_abc_2284_new_n433_), .Y(_abc_2284_new_n434_));
AND2X2 AND2X2_8 ( .A(_abc_2284_new_n399_), .B(_abc_2284_new_n410_), .Y(_abc_2284_new_n449_));
AND2X2 AND2X2_9 ( .A(_abc_2284_new_n465_), .B(_abc_2284_new_n469_), .Y(_abc_2284_new_n497_));
AOI21X1 AOI21X1_1 ( .A(_abc_2284_new_n166_), .B(_abc_2284_new_n170_), .C(_abc_2284_new_n175_), .Y(_abc_2284_new_n176_));
AOI21X1 AOI21X1_10 ( .A(_abc_2284_new_n399_), .B(_abc_2284_new_n410_), .C(_abc_2284_new_n452_), .Y(_abc_2284_new_n453_));
AOI21X1 AOI21X1_11 ( .A(_abc_2284_new_n449_), .B(_abc_2284_new_n451_), .C(_abc_2284_new_n453_), .Y(_abc_2284_new_n454_));
AOI21X1 AOI21X1_12 ( .A(_abc_2284_new_n399_), .B(_abc_2284_new_n410_), .C(_abc_2284_new_n463_), .Y(_abc_2284_new_n464_));
AOI21X1 AOI21X1_13 ( .A(_abc_2284_new_n449_), .B(_abc_2284_new_n462_), .C(_abc_2284_new_n464_), .Y(_abc_2284_new_n465_));
AOI21X1 AOI21X1_14 ( .A(_abc_2284_new_n399_), .B(_abc_2284_new_n410_), .C(_abc_2284_new_n458_), .Y(_abc_2284_new_n468_));
AOI21X1 AOI21X1_15 ( .A(_abc_2284_new_n449_), .B(_abc_2284_new_n467_), .C(_abc_2284_new_n468_), .Y(_abc_2284_new_n469_));
AOI21X1 AOI21X1_16 ( .A(_abc_2284_new_n478_), .B(_abc_2284_new_n474_), .C(_abc_2284_new_n477_), .Y(_abc_2284_new_n479_));
AOI21X1 AOI21X1_17 ( .A(_abc_2284_new_n496_), .B(_abc_2284_new_n497_), .C(_abc_2284_new_n422_), .Y(_abc_2284_new_n501_));
AOI21X1 AOI21X1_18 ( .A(_abc_2284_new_n508_), .B(_abc_2284_new_n474_), .C(_abc_2284_new_n511_), .Y(_abc_2284_new_n512_));
AOI21X1 AOI21X1_19 ( .A(_abc_2284_new_n471_), .B(_abc_2284_new_n487_), .C(_abc_2284_new_n509_), .Y(_abc_2284_new_n523_));
AOI21X1 AOI21X1_2 ( .A(_abc_2284_new_n191_), .B(_abc_2284_new_n176_), .C(_abc_2284_new_n194_), .Y(_abc_2284_new_n195_));
AOI21X1 AOI21X1_20 ( .A(_abc_2284_new_n167_), .B(_abc_2284_new_n556_), .C(_abc_2284_new_n258_), .Y(_0tx_clk_divider_10_0__3_));
AOI21X1 AOI21X1_21 ( .A(_abc_2284_new_n562_), .B(_abc_2284_new_n183_), .C(_abc_2284_new_n258_), .Y(_0tx_clk_divider_10_0__5_));
AOI21X1 AOI21X1_22 ( .A(_abc_2284_new_n182_), .B(_abc_2284_new_n184_), .C(_abc_2284_new_n258_), .Y(_0tx_clk_divider_10_0__6_));
AOI21X1 AOI21X1_23 ( .A(_abc_2284_new_n565_), .B(_abc_2284_new_n566_), .C(_abc_2284_new_n258_), .Y(_0tx_clk_divider_10_0__7_));
AOI21X1 AOI21X1_24 ( .A(_abc_2284_new_n570_), .B(_abc_2284_new_n165_), .C(_abc_2284_new_n258_), .Y(_0tx_clk_divider_10_0__9_));
AOI21X1 AOI21X1_25 ( .A(rx_clk_divider_1_), .B(rx_clk_divider_0_), .C(_abc_2284_new_n428_), .Y(_abc_2284_new_n575_));
AOI21X1 AOI21X1_26 ( .A(_abc_2284_new_n403_), .B(_abc_2284_new_n579_), .C(_abc_2284_new_n428_), .Y(_0rx_clk_divider_10_0__3_));
AOI21X1 AOI21X1_27 ( .A(_abc_2284_new_n391_), .B(_abc_2284_new_n583_), .C(_abc_2284_new_n428_), .Y(_0rx_clk_divider_10_0__5_));
AOI21X1 AOI21X1_28 ( .A(_abc_2284_new_n402_), .B(_abc_2284_new_n404_), .C(_abc_2284_new_n428_), .Y(_0rx_clk_divider_10_0__6_));
AOI21X1 AOI21X1_3 ( .A(_abc_2284_new_n192_), .B(_abc_2284_new_n193_), .C(_abc_2284_new_n195_), .Y(_abc_2284_new_n196_));
AOI21X1 AOI21X1_4 ( .A(_abc_2284_new_n191_), .B(_abc_2284_new_n176_), .C(_abc_2284_new_n214_), .Y(_abc_2284_new_n215_));
AOI21X1 AOI21X1_5 ( .A(_abc_2284_new_n192_), .B(_abc_2284_new_n213_), .C(_abc_2284_new_n215_), .Y(_abc_2284_new_n216_));
AOI21X1 AOI21X1_6 ( .A(_abc_2284_new_n197_), .B(_abc_2284_new_n207_), .C(_abc_2284_new_n244_), .Y(_abc_2284_new_n245_));
AOI21X1 AOI21X1_7 ( .A(_abc_2284_new_n389_), .B(_abc_2284_new_n393_), .C(_abc_2284_new_n398_), .Y(_abc_2284_new_n399_));
AOI21X1 AOI21X1_8 ( .A(_abc_2284_new_n377_), .B(_abc_2284_new_n378_), .C(_abc_2284_new_n380_), .Y(_abc_2284_new_n407_));
AOI21X1 AOI21X1_9 ( .A(rx), .B(_abc_2284_new_n419_), .C(_abc_2284_new_n425_), .Y(_abc_2284_new_n426_));
AOI22X1 AOI22X1_1 ( .A(_abc_2284_new_n258_), .B(\tx_byte[0] ), .C(tx_data_0_), .D(_abc_2284_new_n261_), .Y(_abc_2284_new_n262_));
AOI22X1 AOI22X1_10 ( .A(_abc_2284_new_n327_), .B(_abc_2284_new_n155_), .C(_abc_2284_new_n260_), .D(_abc_2284_new_n369_), .Y(_0tx_state_1_0__1_));
AOI22X1 AOI22X1_11 ( .A(rx_bits_remaining_3_), .B(_abc_2284_new_n447_), .C(_abc_2284_new_n474_), .D(_abc_2284_new_n478_), .Y(_abc_2284_new_n547_));
AOI22X1 AOI22X1_2 ( .A(_abc_2284_new_n258_), .B(\tx_byte[1] ), .C(tx_data_1_), .D(_abc_2284_new_n261_), .Y(_abc_2284_new_n270_));
AOI22X1 AOI22X1_3 ( .A(_abc_2284_new_n258_), .B(\tx_byte[2] ), .C(tx_data_2_), .D(_abc_2284_new_n261_), .Y(_abc_2284_new_n278_));
AOI22X1 AOI22X1_4 ( .A(_abc_2284_new_n258_), .B(\tx_byte[3] ), .C(tx_data_3_), .D(_abc_2284_new_n261_), .Y(_abc_2284_new_n286_));
AOI22X1 AOI22X1_5 ( .A(_abc_2284_new_n258_), .B(\tx_byte[4] ), .C(tx_data_4_), .D(_abc_2284_new_n261_), .Y(_abc_2284_new_n294_));
AOI22X1 AOI22X1_6 ( .A(_abc_2284_new_n258_), .B(\tx_byte[5] ), .C(tx_data_5_), .D(_abc_2284_new_n261_), .Y(_abc_2284_new_n302_));
AOI22X1 AOI22X1_7 ( .A(_abc_2284_new_n258_), .B(\tx_byte[6] ), .C(tx_data_6_), .D(_abc_2284_new_n261_), .Y(_abc_2284_new_n310_));
AOI22X1 AOI22X1_8 ( .A(_abc_2284_new_n323_), .B(_abc_2284_new_n324_), .C(_abc_2284_new_n319_), .D(_abc_2284_new_n328_), .Y(_0tx_bits_remaining_3_0__0_));
AOI22X1 AOI22X1_9 ( .A(_abc_2284_new_n331_), .B(_abc_2284_new_n362_), .C(_abc_2284_new_n216_), .D(_abc_2284_new_n363_), .Y(_0tx_countdown_5_0__3_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_0rx_clk_divider_10_0__6_), .Q(rx_clk_divider_6_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(_0tx_clk_divider_10_0__4_), .Q(tx_clk_divider_4_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(_0tx_clk_divider_10_0__5_), .Q(tx_clk_divider_5_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(_0tx_clk_divider_10_0__6_), .Q(tx_clk_divider_6_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(_0tx_clk_divider_10_0__7_), .Q(tx_clk_divider_7_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(_0tx_clk_divider_10_0__8_), .Q(tx_clk_divider_8_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(_0tx_clk_divider_10_0__9_), .Q(tx_clk_divider_9_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(_0tx_clk_divider_10_0__10_), .Q(tx_clk_divider_10_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(_0recv_state_2_0__0_), .Q(recv_state_0_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(_0recv_state_2_0__1_), .Q(recv_state_1_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(_0recv_state_2_0__2_), .Q(recv_state_2_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_0rx_clk_divider_10_0__7_), .Q(rx_clk_divider_7_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(_0rx_countdown_5_0__0_), .Q(rx_countdown_0_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(_0rx_countdown_5_0__1_), .Q(rx_countdown_1_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(_0rx_countdown_5_0__2_), .Q(rx_countdown_2_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(_0rx_countdown_5_0__3_), .Q(rx_countdown_3_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(_0rx_countdown_5_0__4_), .Q(rx_countdown_4_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(_0rx_countdown_5_0__5_), .Q(rx_countdown_5_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(_0rx_bits_remaining_3_0__0_), .Q(rx_bits_remaining_0_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(_0rx_bits_remaining_3_0__1_), .Q(rx_bits_remaining_1_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(_0rx_bits_remaining_3_0__2_), .Q(rx_bits_remaining_2_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(_0rx_bits_remaining_3_0__3_), .Q(rx_bits_remaining_3_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_0rx_clk_divider_10_0__8_), .Q(rx_clk_divider_8_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(_0rx_data_7_0__0_), .Q(\rx_byte[0] ));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(_0rx_data_7_0__1_), .Q(\rx_byte[1] ));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(_0rx_data_7_0__2_), .Q(\rx_byte[2] ));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(_0rx_data_7_0__3_), .Q(\rx_byte[3] ));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(_0rx_data_7_0__4_), .Q(\rx_byte[4] ));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(_0rx_data_7_0__5_), .Q(\rx_byte[5] ));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(_0rx_data_7_0__6_), .Q(\rx_byte[6] ));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(_0rx_data_7_0__7_), .Q(\rx_byte[7] ));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(_0tx_out_0_0_), .Q(tx));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(_0tx_state_1_0__0_), .Q(tx_state_0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_0rx_clk_divider_10_0__9_), .Q(rx_clk_divider_9_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(_0tx_state_1_0__1_), .Q(tx_state_1_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(_0tx_countdown_5_0__0_), .Q(tx_countdown_0_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(_0tx_countdown_5_0__1_), .Q(tx_countdown_1_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(_0tx_countdown_5_0__2_), .Q(tx_countdown_2_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(_0tx_countdown_5_0__3_), .Q(tx_countdown_3_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(_0tx_countdown_5_0__4_), .Q(tx_countdown_4_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(_0tx_countdown_5_0__5_), .Q(tx_countdown_5_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(_0tx_bits_remaining_3_0__0_), .Q(tx_bits_remaining_0_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(_0tx_bits_remaining_3_0__1_), .Q(tx_bits_remaining_1_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(_0tx_bits_remaining_3_0__2_), .Q(tx_bits_remaining_2_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_0rx_clk_divider_10_0__10_), .Q(rx_clk_divider_10_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(_0tx_bits_remaining_3_0__3_), .Q(tx_bits_remaining_3_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(_0tx_data_7_0__0_), .Q(tx_data_0_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(_0tx_data_7_0__1_), .Q(tx_data_1_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(_0tx_data_7_0__2_), .Q(tx_data_2_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(_0tx_data_7_0__3_), .Q(tx_data_3_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(_0tx_data_7_0__4_), .Q(tx_data_4_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(_0tx_data_7_0__5_), .Q(tx_data_5_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(_0tx_data_7_0__6_), .Q(tx_data_6_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(_0tx_data_7_0__7_), .Q(tx_data_7_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(_0rx_clk_divider_10_0__0_), .Q(rx_clk_divider_0_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(_0tx_clk_divider_10_0__0_), .Q(tx_clk_divider_0_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(_0rx_clk_divider_10_0__1_), .Q(rx_clk_divider_1_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(_0rx_clk_divider_10_0__2_), .Q(rx_clk_divider_2_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(_0rx_clk_divider_10_0__3_), .Q(rx_clk_divider_3_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(_0rx_clk_divider_10_0__4_), .Q(rx_clk_divider_4_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(_0rx_clk_divider_10_0__5_), .Q(rx_clk_divider_5_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(_0tx_clk_divider_10_0__1_), .Q(tx_clk_divider_1_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(_0tx_clk_divider_10_0__2_), .Q(tx_clk_divider_2_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(_0tx_clk_divider_10_0__3_), .Q(tx_clk_divider_3_));
INVX1 INVX1_1 ( .A(recv_state_1_), .Y(_abc_2284_new_n144_));
INVX1 INVX1_10 ( .A(tx_clk_divider_6_), .Y(_abc_2284_new_n181_));
INVX1 INVX1_11 ( .A(tx_clk_divider_5_), .Y(_abc_2284_new_n186_));
INVX1 INVX1_12 ( .A(tx_clk_divider_4_), .Y(_abc_2284_new_n187_));
INVX1 INVX1_13 ( .A(tx_countdown_1_), .Y(_abc_2284_new_n194_));
INVX1 INVX1_14 ( .A(tx_countdown_0_), .Y(_abc_2284_new_n198_));
INVX1 INVX1_15 ( .A(_abc_2284_new_n175_), .Y(_abc_2284_new_n200_));
INVX1 INVX1_16 ( .A(_abc_2284_new_n190_), .Y(_abc_2284_new_n205_));
INVX1 INVX1_17 ( .A(tx_countdown_2_), .Y(_abc_2284_new_n210_));
INVX1 INVX1_18 ( .A(tx_countdown_3_), .Y(_abc_2284_new_n214_));
INVX1 INVX1_19 ( .A(tx_countdown_4_), .Y(_abc_2284_new_n228_));
INVX1 INVX1_2 ( .A(tx_state_1_), .Y(_abc_2284_new_n147_));
INVX1 INVX1_20 ( .A(tx_data_1_), .Y(_abc_2284_new_n237_));
INVX1 INVX1_21 ( .A(tx_data_0_), .Y(_abc_2284_new_n241_));
INVX1 INVX1_22 ( .A(transmit), .Y(_abc_2284_new_n254_));
INVX1 INVX1_23 ( .A(rst), .Y(_abc_2284_new_n255_));
INVX1 INVX1_24 ( .A(_abc_2284_new_n256_), .Y(_abc_2284_new_n257_));
INVX1 INVX1_25 ( .A(_abc_2284_new_n259_), .Y(_abc_2284_new_n260_));
INVX1 INVX1_26 ( .A(tx_data_2_), .Y(_abc_2284_new_n264_));
INVX1 INVX1_27 ( .A(tx_data_3_), .Y(_abc_2284_new_n272_));
INVX1 INVX1_28 ( .A(tx_data_4_), .Y(_abc_2284_new_n280_));
INVX1 INVX1_29 ( .A(tx_data_5_), .Y(_abc_2284_new_n288_));
INVX1 INVX1_3 ( .A(tx_state_0_), .Y(_abc_2284_new_n148_));
INVX1 INVX1_30 ( .A(tx_data_6_), .Y(_abc_2284_new_n296_));
INVX1 INVX1_31 ( .A(tx_data_7_), .Y(_abc_2284_new_n304_));
INVX1 INVX1_32 ( .A(tx_bits_remaining_0_), .Y(_abc_2284_new_n319_));
INVX1 INVX1_33 ( .A(_abc_2284_new_n236_), .Y(_abc_2284_new_n320_));
INVX1 INVX1_34 ( .A(_abc_2284_new_n156_), .Y(_abc_2284_new_n321_));
INVX1 INVX1_35 ( .A(tx_bits_remaining_1_), .Y(_abc_2284_new_n330_));
INVX1 INVX1_36 ( .A(_abc_2284_new_n261_), .Y(_abc_2284_new_n331_));
INVX1 INVX1_37 ( .A(tx_bits_remaining_2_), .Y(_abc_2284_new_n340_));
INVX1 INVX1_38 ( .A(_abc_2284_new_n258_), .Y(_abc_2284_new_n349_));
INVX1 INVX1_39 ( .A(_abc_2284_new_n234_), .Y(_abc_2284_new_n350_));
INVX1 INVX1_4 ( .A(_abc_2284_new_n154_), .Y(_abc_2284_new_n155_));
INVX1 INVX1_40 ( .A(tx_bits_remaining_3_), .Y(_abc_2284_new_n353_));
INVX1 INVX1_41 ( .A(rx_clk_divider_10_), .Y(_abc_2284_new_n376_));
INVX1 INVX1_42 ( .A(rx_clk_divider_4_), .Y(_abc_2284_new_n380_));
INVX1 INVX1_43 ( .A(rx_clk_divider_5_), .Y(_abc_2284_new_n381_));
INVX1 INVX1_44 ( .A(rx_clk_divider_6_), .Y(_abc_2284_new_n383_));
INVX1 INVX1_45 ( .A(rx_clk_divider_7_), .Y(_abc_2284_new_n384_));
INVX1 INVX1_46 ( .A(rx_clk_divider_9_), .Y(_abc_2284_new_n394_));
INVX1 INVX1_47 ( .A(rx_clk_divider_8_), .Y(_abc_2284_new_n395_));
INVX1 INVX1_48 ( .A(rx_clk_divider_1_), .Y(_abc_2284_new_n400_));
INVX1 INVX1_49 ( .A(_abc_2284_new_n407_), .Y(_abc_2284_new_n408_));
INVX1 INVX1_5 ( .A(tx_clk_divider_10_), .Y(_abc_2284_new_n157_));
INVX1 INVX1_50 ( .A(rx_countdown_0_), .Y(_abc_2284_new_n412_));
INVX1 INVX1_51 ( .A(recv_state_2_), .Y(_abc_2284_new_n416_));
INVX1 INVX1_52 ( .A(_abc_2284_new_n418_), .Y(_abc_2284_new_n419_));
INVX1 INVX1_53 ( .A(_abc_2284_new_n428_), .Y(_abc_2284_new_n429_));
INVX1 INVX1_54 ( .A(_abc_2284_new_n406_), .Y(_abc_2284_new_n435_));
INVX1 INVX1_55 ( .A(rx_clk_divider_0_), .Y(_abc_2284_new_n436_));
INVX1 INVX1_56 ( .A(_abc_2284_new_n447_), .Y(_abc_2284_new_n448_));
INVX1 INVX1_57 ( .A(rx_countdown_2_), .Y(_abc_2284_new_n452_));
INVX1 INVX1_58 ( .A(rx_countdown_4_), .Y(_abc_2284_new_n457_));
INVX1 INVX1_59 ( .A(rx_countdown_3_), .Y(_abc_2284_new_n458_));
INVX1 INVX1_6 ( .A(tx_clk_divider_9_), .Y(_abc_2284_new_n171_));
INVX1 INVX1_60 ( .A(rx_countdown_5_), .Y(_abc_2284_new_n463_));
INVX1 INVX1_61 ( .A(_abc_2284_new_n423_), .Y(_abc_2284_new_n473_));
INVX1 INVX1_62 ( .A(_abc_2284_new_n451_), .Y(_abc_2284_new_n475_));
INVX1 INVX1_63 ( .A(_abc_2284_new_n445_), .Y(_abc_2284_new_n481_));
INVX1 INVX1_64 ( .A(_abc_2284_new_n439_), .Y(_abc_2284_new_n490_));
INVX1 INVX1_65 ( .A(rx_bits_remaining_1_), .Y(_abc_2284_new_n502_));
INVX1 INVX1_66 ( .A(rx), .Y(_abc_2284_new_n507_));
INVX1 INVX1_67 ( .A(_abc_2284_new_n474_), .Y(_abc_2284_new_n516_));
INVX1 INVX1_68 ( .A(rx_bits_remaining_0_), .Y(_abc_2284_new_n525_));
INVX1 INVX1_69 ( .A(rx_bits_remaining_2_), .Y(_abc_2284_new_n535_));
INVX1 INVX1_7 ( .A(tx_clk_divider_8_), .Y(_abc_2284_new_n172_));
INVX1 INVX1_70 ( .A(rx_bits_remaining_3_), .Y(_abc_2284_new_n541_));
INVX1 INVX1_71 ( .A(_abc_2284_new_n159_), .Y(_abc_2284_new_n555_));
INVX1 INVX1_72 ( .A(_abc_2284_new_n188_), .Y(_abc_2284_new_n558_));
INVX1 INVX1_73 ( .A(_abc_2284_new_n169_), .Y(_abc_2284_new_n565_));
INVX1 INVX1_74 ( .A(_abc_2284_new_n378_), .Y(_abc_2284_new_n574_));
INVX1 INVX1_75 ( .A(\rx_byte[0] ), .Y(_abc_2284_new_n592_));
INVX1 INVX1_76 ( .A(\rx_byte[1] ), .Y(_abc_2284_new_n593_));
INVX1 INVX1_77 ( .A(\rx_byte[2] ), .Y(_abc_2284_new_n595_));
INVX1 INVX1_78 ( .A(\rx_byte[3] ), .Y(_abc_2284_new_n597_));
INVX1 INVX1_79 ( .A(\rx_byte[4] ), .Y(_abc_2284_new_n599_));
INVX1 INVX1_8 ( .A(_abc_2284_new_n178_), .Y(_abc_2284_new_n179_));
INVX1 INVX1_80 ( .A(\rx_byte[5] ), .Y(_abc_2284_new_n601_));
INVX1 INVX1_81 ( .A(\rx_byte[6] ), .Y(_abc_2284_new_n603_));
INVX1 INVX1_82 ( .A(\rx_byte[7] ), .Y(_abc_2284_new_n605_));
INVX1 INVX1_9 ( .A(tx_clk_divider_7_), .Y(_abc_2284_new_n180_));
MUX2X1 MUX2X1_1 ( .A(tx_countdown_4_), .B(_abc_2284_new_n230_), .S(_abc_2284_new_n222_), .Y(_abc_2284_new_n325_));
MUX2X1 MUX2X1_2 ( .A(rx_countdown_4_), .B(_abc_2284_new_n483_), .S(_abc_2284_new_n413_), .Y(_abc_2284_new_n484_));
MUX2X1 MUX2X1_3 ( .A(_abc_2284_new_n592_), .B(_abc_2284_new_n593_), .S(_abc_2284_new_n472_), .Y(_0rx_data_7_0__0_));
MUX2X1 MUX2X1_4 ( .A(_abc_2284_new_n593_), .B(_abc_2284_new_n595_), .S(_abc_2284_new_n472_), .Y(_0rx_data_7_0__1_));
MUX2X1 MUX2X1_5 ( .A(_abc_2284_new_n595_), .B(_abc_2284_new_n597_), .S(_abc_2284_new_n472_), .Y(_0rx_data_7_0__2_));
MUX2X1 MUX2X1_6 ( .A(_abc_2284_new_n597_), .B(_abc_2284_new_n599_), .S(_abc_2284_new_n472_), .Y(_0rx_data_7_0__3_));
MUX2X1 MUX2X1_7 ( .A(_abc_2284_new_n599_), .B(_abc_2284_new_n601_), .S(_abc_2284_new_n472_), .Y(_0rx_data_7_0__4_));
MUX2X1 MUX2X1_8 ( .A(_abc_2284_new_n601_), .B(_abc_2284_new_n603_), .S(_abc_2284_new_n472_), .Y(_0rx_data_7_0__5_));
MUX2X1 MUX2X1_9 ( .A(_abc_2284_new_n603_), .B(_abc_2284_new_n605_), .S(_abc_2284_new_n472_), .Y(_0rx_data_7_0__6_));
NAND2X1 NAND2X1_1 ( .A(_abc_2284_new_n144_), .B(_abc_2284_new_n145_), .Y(is_receiving));
NAND2X1 NAND2X1_10 ( .A(tx_clk_divider_4_), .B(_abc_2284_new_n167_), .Y(_abc_2284_new_n189_));
NAND2X1 NAND2X1_11 ( .A(_abc_2284_new_n170_), .B(_abc_2284_new_n166_), .Y(_abc_2284_new_n199_));
NAND2X1 NAND2X1_12 ( .A(_abc_2284_new_n199_), .B(_abc_2284_new_n200_), .Y(_abc_2284_new_n201_));
NAND2X1 NAND2X1_13 ( .A(_abc_2284_new_n197_), .B(_abc_2284_new_n207_), .Y(_abc_2284_new_n208_));
NAND2X1 NAND2X1_14 ( .A(_abc_2284_new_n208_), .B(_abc_2284_new_n196_), .Y(_abc_2284_new_n209_));
NAND2X1 NAND2X1_15 ( .A(_abc_2284_new_n210_), .B(_abc_2284_new_n211_), .Y(_abc_2284_new_n212_));
NAND2X1 NAND2X1_16 ( .A(_abc_2284_new_n176_), .B(_abc_2284_new_n191_), .Y(_abc_2284_new_n222_));
NAND2X1 NAND2X1_17 ( .A(tx_countdown_4_), .B(_abc_2284_new_n223_), .Y(_abc_2284_new_n229_));
NAND2X1 NAND2X1_18 ( .A(_abc_2284_new_n229_), .B(_abc_2284_new_n224_), .Y(_abc_2284_new_n230_));
NAND2X1 NAND2X1_19 ( .A(_abc_2284_new_n234_), .B(_abc_2284_new_n235_), .Y(_abc_2284_new_n236_));
NAND2X1 NAND2X1_2 ( .A(_abc_2284_new_n147_), .B(_abc_2284_new_n148_), .Y(is_transmitting));
NAND2X1 NAND2X1_20 ( .A(_abc_2284_new_n237_), .B(_abc_2284_new_n236_), .Y(_abc_2284_new_n238_));
NAND2X1 NAND2X1_21 ( .A(_abc_2284_new_n242_), .B(_abc_2284_new_n243_), .Y(_abc_2284_new_n244_));
NAND2X1 NAND2X1_22 ( .A(_abc_2284_new_n246_), .B(_abc_2284_new_n247_), .Y(_abc_2284_new_n248_));
NAND2X1 NAND2X1_23 ( .A(_abc_2284_new_n241_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n252_));
NAND2X1 NAND2X1_24 ( .A(_abc_2284_new_n262_), .B(_abc_2284_new_n253_), .Y(_0tx_data_7_0__0_));
NAND2X1 NAND2X1_25 ( .A(_abc_2284_new_n264_), .B(_abc_2284_new_n236_), .Y(_abc_2284_new_n265_));
NAND2X1 NAND2X1_26 ( .A(_abc_2284_new_n237_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n268_));
NAND2X1 NAND2X1_27 ( .A(_abc_2284_new_n270_), .B(_abc_2284_new_n269_), .Y(_0tx_data_7_0__1_));
NAND2X1 NAND2X1_28 ( .A(_abc_2284_new_n272_), .B(_abc_2284_new_n236_), .Y(_abc_2284_new_n273_));
NAND2X1 NAND2X1_29 ( .A(_abc_2284_new_n264_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n276_));
NAND2X1 NAND2X1_3 ( .A(recv_state_1_), .B(recv_state_2_), .Y(_abc_2284_new_n150_));
NAND2X1 NAND2X1_30 ( .A(_abc_2284_new_n278_), .B(_abc_2284_new_n277_), .Y(_0tx_data_7_0__2_));
NAND2X1 NAND2X1_31 ( .A(_abc_2284_new_n280_), .B(_abc_2284_new_n236_), .Y(_abc_2284_new_n281_));
NAND2X1 NAND2X1_32 ( .A(_abc_2284_new_n272_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n284_));
NAND2X1 NAND2X1_33 ( .A(_abc_2284_new_n286_), .B(_abc_2284_new_n285_), .Y(_0tx_data_7_0__3_));
NAND2X1 NAND2X1_34 ( .A(_abc_2284_new_n288_), .B(_abc_2284_new_n236_), .Y(_abc_2284_new_n289_));
NAND2X1 NAND2X1_35 ( .A(_abc_2284_new_n280_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n292_));
NAND2X1 NAND2X1_36 ( .A(_abc_2284_new_n294_), .B(_abc_2284_new_n293_), .Y(_0tx_data_7_0__4_));
NAND2X1 NAND2X1_37 ( .A(_abc_2284_new_n296_), .B(_abc_2284_new_n236_), .Y(_abc_2284_new_n297_));
NAND2X1 NAND2X1_38 ( .A(_abc_2284_new_n288_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n300_));
NAND2X1 NAND2X1_39 ( .A(_abc_2284_new_n302_), .B(_abc_2284_new_n301_), .Y(_0tx_data_7_0__5_));
NAND2X1 NAND2X1_4 ( .A(recv_state_0_), .B(recv_state_2_), .Y(_abc_2284_new_n152_));
NAND2X1 NAND2X1_40 ( .A(_abc_2284_new_n304_), .B(_abc_2284_new_n236_), .Y(_abc_2284_new_n305_));
NAND2X1 NAND2X1_41 ( .A(_abc_2284_new_n296_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n308_));
NAND2X1 NAND2X1_42 ( .A(_abc_2284_new_n310_), .B(_abc_2284_new_n309_), .Y(_0tx_data_7_0__6_));
NAND2X1 NAND2X1_43 ( .A(_abc_2284_new_n254_), .B(_abc_2284_new_n304_), .Y(_abc_2284_new_n312_));
NAND2X1 NAND2X1_44 ( .A(tx_data_7_), .B(_abc_2284_new_n259_), .Y(_abc_2284_new_n317_));
NAND2X1 NAND2X1_45 ( .A(_abc_2284_new_n322_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n323_));
NAND2X1 NAND2X1_46 ( .A(_abc_2284_new_n322_), .B(_abc_2284_new_n327_), .Y(_abc_2284_new_n328_));
NAND2X1 NAND2X1_47 ( .A(tx_bits_remaining_0_), .B(_abc_2284_new_n330_), .Y(_abc_2284_new_n332_));
NAND2X1 NAND2X1_48 ( .A(tx_bits_remaining_1_), .B(_abc_2284_new_n319_), .Y(_abc_2284_new_n333_));
NAND2X1 NAND2X1_49 ( .A(_abc_2284_new_n330_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n336_));
NAND2X1 NAND2X1_5 ( .A(_abc_2284_new_n157_), .B(_abc_2284_new_n165_), .Y(_abc_2284_new_n166_));
NAND2X1 NAND2X1_50 ( .A(tx_bits_remaining_2_), .B(_abc_2284_new_n234_), .Y(_abc_2284_new_n342_));
NAND2X1 NAND2X1_51 ( .A(_abc_2284_new_n340_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n345_));
NAND2X1 NAND2X1_52 ( .A(tx_bits_remaining_2_), .B(_abc_2284_new_n259_), .Y(_abc_2284_new_n347_));
NAND2X1 NAND2X1_53 ( .A(_abc_2284_new_n353_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n354_));
NAND2X1 NAND2X1_54 ( .A(_abc_2284_new_n320_), .B(_abc_2284_new_n327_), .Y(_abc_2284_new_n369_));
NAND2X1 NAND2X1_55 ( .A(_abc_2284_new_n241_), .B(_abc_2284_new_n236_), .Y(_abc_2284_new_n371_));
NAND2X1 NAND2X1_56 ( .A(tx), .B(_abc_2284_new_n261_), .Y(_abc_2284_new_n374_));
NAND2X1 NAND2X1_57 ( .A(_abc_2284_new_n380_), .B(_abc_2284_new_n381_), .Y(_abc_2284_new_n382_));
NAND2X1 NAND2X1_58 ( .A(_abc_2284_new_n383_), .B(_abc_2284_new_n384_), .Y(_abc_2284_new_n385_));
NAND2X1 NAND2X1_59 ( .A(_abc_2284_new_n376_), .B(_abc_2284_new_n388_), .Y(_abc_2284_new_n389_));
NAND2X1 NAND2X1_6 ( .A(_abc_2284_new_n158_), .B(_abc_2284_new_n159_), .Y(_abc_2284_new_n167_));
NAND2X1 NAND2X1_60 ( .A(_abc_2284_new_n377_), .B(_abc_2284_new_n378_), .Y(_abc_2284_new_n403_));
NAND2X1 NAND2X1_61 ( .A(_abc_2284_new_n410_), .B(_abc_2284_new_n399_), .Y(_abc_2284_new_n413_));
NAND2X1 NAND2X1_62 ( .A(_abc_2284_new_n412_), .B(_abc_2284_new_n413_), .Y(_abc_2284_new_n414_));
NAND2X1 NAND2X1_63 ( .A(_abc_2284_new_n411_), .B(_abc_2284_new_n414_), .Y(_abc_2284_new_n415_));
NAND2X1 NAND2X1_64 ( .A(recv_state_2_), .B(_abc_2284_new_n255_), .Y(_abc_2284_new_n420_));
NAND2X1 NAND2X1_65 ( .A(recv_state_0_), .B(_abc_2284_new_n255_), .Y(_abc_2284_new_n422_));
NAND2X1 NAND2X1_66 ( .A(_abc_2284_new_n379_), .B(_abc_2284_new_n386_), .Y(_abc_2284_new_n430_));
NAND2X1 NAND2X1_67 ( .A(_abc_2284_new_n388_), .B(_abc_2284_new_n431_), .Y(_abc_2284_new_n432_));
NAND2X1 NAND2X1_68 ( .A(_abc_2284_new_n440_), .B(_abc_2284_new_n434_), .Y(_abc_2284_new_n441_));
NAND2X1 NAND2X1_69 ( .A(_abc_2284_new_n145_), .B(_abc_2284_new_n421_), .Y(_abc_2284_new_n447_));
NAND2X1 NAND2X1_7 ( .A(_abc_2284_new_n161_), .B(_abc_2284_new_n162_), .Y(_abc_2284_new_n168_));
NAND2X1 NAND2X1_70 ( .A(_abc_2284_new_n452_), .B(_abc_2284_new_n458_), .Y(_abc_2284_new_n459_));
NAND2X1 NAND2X1_71 ( .A(_abc_2284_new_n457_), .B(_abc_2284_new_n460_), .Y(_abc_2284_new_n461_));
NAND2X1 NAND2X1_72 ( .A(_abc_2284_new_n465_), .B(_abc_2284_new_n469_), .Y(_abc_2284_new_n470_));
NAND2X1 NAND2X1_73 ( .A(_abc_2284_new_n448_), .B(_abc_2284_new_n471_), .Y(_abc_2284_new_n472_));
NAND2X1 NAND2X1_74 ( .A(rx_countdown_2_), .B(_abc_2284_new_n413_), .Y(_abc_2284_new_n476_));
NAND2X1 NAND2X1_75 ( .A(rx_countdown_0_), .B(_abc_2284_new_n493_), .Y(_abc_2284_new_n494_));
NAND2X1 NAND2X1_76 ( .A(recv_state_1_), .B(_abc_2284_new_n509_), .Y(_abc_2284_new_n510_));
NAND2X1 NAND2X1_77 ( .A(_abc_2284_new_n497_), .B(_abc_2284_new_n496_), .Y(_abc_2284_new_n514_));
NAND2X1 NAND2X1_78 ( .A(rx_bits_remaining_0_), .B(_abc_2284_new_n471_), .Y(_abc_2284_new_n527_));
NAND2X1 NAND2X1_79 ( .A(_abc_2284_new_n535_), .B(_abc_2284_new_n536_), .Y(_abc_2284_new_n542_));
NAND2X1 NAND2X1_8 ( .A(tx_clk_divider_0_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n177_));
NAND2X1 NAND2X1_80 ( .A(_abc_2284_new_n543_), .B(_abc_2284_new_n471_), .Y(_abc_2284_new_n544_));
NAND2X1 NAND2X1_81 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n546_), .Y(_0rx_bits_remaining_3_0__3_));
NAND2X1 NAND2X1_82 ( .A(_abc_2284_new_n393_), .B(_abc_2284_new_n389_), .Y(_abc_2284_new_n590_));
NAND2X1 NAND2X1_9 ( .A(tx_clk_divider_6_), .B(_abc_2284_new_n183_), .Y(_abc_2284_new_n184_));
NAND3X1 NAND3X1_1 ( .A(_abc_2284_new_n164_), .B(_abc_2284_new_n160_), .C(_abc_2284_new_n163_), .Y(_abc_2284_new_n165_));
NAND3X1 NAND3X1_10 ( .A(tx_countdown_0_), .B(_abc_2284_new_n176_), .C(_abc_2284_new_n191_), .Y(_abc_2284_new_n197_));
NAND3X1 NAND3X1_11 ( .A(_abc_2284_new_n178_), .B(_abc_2284_new_n205_), .C(_abc_2284_new_n204_), .Y(_abc_2284_new_n206_));
NAND3X1 NAND3X1_12 ( .A(_abc_2284_new_n176_), .B(_abc_2284_new_n217_), .C(_abc_2284_new_n191_), .Y(_abc_2284_new_n218_));
NAND3X1 NAND3X1_13 ( .A(_abc_2284_new_n218_), .B(_abc_2284_new_n219_), .C(_abc_2284_new_n216_), .Y(_abc_2284_new_n220_));
NAND3X1 NAND3X1_14 ( .A(_abc_2284_new_n210_), .B(_abc_2284_new_n214_), .C(_abc_2284_new_n211_), .Y(_abc_2284_new_n223_));
NAND3X1 NAND3X1_15 ( .A(_abc_2284_new_n176_), .B(_abc_2284_new_n230_), .C(_abc_2284_new_n191_), .Y(_abc_2284_new_n231_));
NAND3X1 NAND3X1_16 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n239_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n240_));
NAND3X1 NAND3X1_17 ( .A(_abc_2284_new_n176_), .B(_abc_2284_new_n193_), .C(_abc_2284_new_n191_), .Y(_abc_2284_new_n242_));
NAND3X1 NAND3X1_18 ( .A(_abc_2284_new_n176_), .B(_abc_2284_new_n213_), .C(_abc_2284_new_n191_), .Y(_abc_2284_new_n246_));
NAND3X1 NAND3X1_19 ( .A(_abc_2284_new_n245_), .B(_abc_2284_new_n250_), .C(_abc_2284_new_n233_), .Y(_abc_2284_new_n251_));
NAND3X1 NAND3X1_2 ( .A(tx_clk_divider_10_), .B(_abc_2284_new_n164_), .C(_abc_2284_new_n169_), .Y(_abc_2284_new_n170_));
NAND3X1 NAND3X1_20 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n252_), .C(_abc_2284_new_n240_), .Y(_abc_2284_new_n253_));
NAND3X1 NAND3X1_21 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n266_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n267_));
NAND3X1 NAND3X1_22 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n268_), .C(_abc_2284_new_n267_), .Y(_abc_2284_new_n269_));
NAND3X1 NAND3X1_23 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n274_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n275_));
NAND3X1 NAND3X1_24 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n276_), .C(_abc_2284_new_n275_), .Y(_abc_2284_new_n277_));
NAND3X1 NAND3X1_25 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n282_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n283_));
NAND3X1 NAND3X1_26 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n284_), .C(_abc_2284_new_n283_), .Y(_abc_2284_new_n285_));
NAND3X1 NAND3X1_27 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n290_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n291_));
NAND3X1 NAND3X1_28 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n292_), .C(_abc_2284_new_n291_), .Y(_abc_2284_new_n293_));
NAND3X1 NAND3X1_29 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n298_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n299_));
NAND3X1 NAND3X1_3 ( .A(_abc_2284_new_n172_), .B(_abc_2284_new_n160_), .C(_abc_2284_new_n163_), .Y(_abc_2284_new_n173_));
NAND3X1 NAND3X1_30 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n300_), .C(_abc_2284_new_n299_), .Y(_abc_2284_new_n301_));
NAND3X1 NAND3X1_31 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n306_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n307_));
NAND3X1 NAND3X1_32 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n308_), .C(_abc_2284_new_n307_), .Y(_abc_2284_new_n309_));
NAND3X1 NAND3X1_33 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n315_));
NAND3X1 NAND3X1_34 ( .A(tx_data_7_), .B(_abc_2284_new_n156_), .C(_abc_2284_new_n315_), .Y(_abc_2284_new_n316_));
NAND3X1 NAND3X1_35 ( .A(_abc_2284_new_n314_), .B(_abc_2284_new_n317_), .C(_abc_2284_new_n316_), .Y(_0tx_data_7_0__7_));
NAND3X1 NAND3X1_36 ( .A(_abc_2284_new_n196_), .B(_abc_2284_new_n208_), .C(_abc_2284_new_n325_), .Y(_abc_2284_new_n326_));
NAND3X1 NAND3X1_37 ( .A(_abc_2284_new_n332_), .B(_abc_2284_new_n333_), .C(_abc_2284_new_n236_), .Y(_abc_2284_new_n334_));
NAND3X1 NAND3X1_38 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n334_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n335_));
NAND3X1 NAND3X1_39 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n336_), .C(_abc_2284_new_n335_), .Y(_abc_2284_new_n337_));
NAND3X1 NAND3X1_4 ( .A(_abc_2284_new_n171_), .B(_abc_2284_new_n174_), .C(_abc_2284_new_n173_), .Y(_abc_2284_new_n175_));
NAND3X1 NAND3X1_40 ( .A(tx_bits_remaining_2_), .B(_abc_2284_new_n254_), .C(_abc_2284_new_n256_), .Y(_abc_2284_new_n339_));
NAND3X1 NAND3X1_41 ( .A(_abc_2284_new_n341_), .B(_abc_2284_new_n342_), .C(_abc_2284_new_n236_), .Y(_abc_2284_new_n343_));
NAND3X1 NAND3X1_42 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n343_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n344_));
NAND3X1 NAND3X1_43 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n345_), .C(_abc_2284_new_n344_), .Y(_abc_2284_new_n346_));
NAND3X1 NAND3X1_44 ( .A(_abc_2284_new_n339_), .B(_abc_2284_new_n347_), .C(_abc_2284_new_n346_), .Y(_0tx_bits_remaining_3_0__2_));
NAND3X1 NAND3X1_45 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n351_), .C(_abc_2284_new_n221_), .Y(_abc_2284_new_n352_));
NAND3X1 NAND3X1_46 ( .A(_abc_2284_new_n156_), .B(_abc_2284_new_n354_), .C(_abc_2284_new_n352_), .Y(_abc_2284_new_n355_));
NAND3X1 NAND3X1_47 ( .A(_abc_2284_new_n349_), .B(_abc_2284_new_n356_), .C(_abc_2284_new_n355_), .Y(_0tx_bits_remaining_3_0__3_));
NAND3X1 NAND3X1_48 ( .A(_abc_2284_new_n320_), .B(_abc_2284_new_n156_), .C(_abc_2284_new_n327_), .Y(_abc_2284_new_n363_));
NAND3X1 NAND3X1_49 ( .A(_abc_2284_new_n379_), .B(_abc_2284_new_n387_), .C(_abc_2284_new_n386_), .Y(_abc_2284_new_n388_));
NAND3X1 NAND3X1_5 ( .A(_abc_2284_new_n181_), .B(_abc_2284_new_n161_), .C(_abc_2284_new_n160_), .Y(_abc_2284_new_n182_));
NAND3X1 NAND3X1_50 ( .A(_abc_2284_new_n377_), .B(_abc_2284_new_n378_), .C(_abc_2284_new_n390_), .Y(_abc_2284_new_n391_));
NAND3X1 NAND3X1_51 ( .A(rx_clk_divider_10_), .B(_abc_2284_new_n387_), .C(_abc_2284_new_n392_), .Y(_abc_2284_new_n393_));
NAND3X1 NAND3X1_52 ( .A(_abc_2284_new_n395_), .B(_abc_2284_new_n379_), .C(_abc_2284_new_n386_), .Y(_abc_2284_new_n396_));
NAND3X1 NAND3X1_53 ( .A(_abc_2284_new_n394_), .B(_abc_2284_new_n397_), .C(_abc_2284_new_n396_), .Y(_abc_2284_new_n398_));
NAND3X1 NAND3X1_54 ( .A(_abc_2284_new_n400_), .B(rx_clk_divider_0_), .C(_abc_2284_new_n377_), .Y(_abc_2284_new_n401_));
NAND3X1 NAND3X1_55 ( .A(_abc_2284_new_n383_), .B(_abc_2284_new_n390_), .C(_abc_2284_new_n379_), .Y(_abc_2284_new_n402_));
NAND3X1 NAND3X1_56 ( .A(_abc_2284_new_n384_), .B(_abc_2284_new_n404_), .C(_abc_2284_new_n402_), .Y(_abc_2284_new_n405_));
NAND3X1 NAND3X1_57 ( .A(_abc_2284_new_n380_), .B(_abc_2284_new_n377_), .C(_abc_2284_new_n378_), .Y(_abc_2284_new_n406_));
NAND3X1 NAND3X1_58 ( .A(_abc_2284_new_n381_), .B(_abc_2284_new_n406_), .C(_abc_2284_new_n408_), .Y(_abc_2284_new_n409_));
NAND3X1 NAND3X1_59 ( .A(rx_countdown_0_), .B(_abc_2284_new_n410_), .C(_abc_2284_new_n399_), .Y(_abc_2284_new_n411_));
NAND3X1 NAND3X1_6 ( .A(_abc_2284_new_n158_), .B(_abc_2284_new_n159_), .C(_abc_2284_new_n161_), .Y(_abc_2284_new_n183_));
NAND3X1 NAND3X1_60 ( .A(_abc_2284_new_n377_), .B(_abc_2284_new_n438_), .C(_abc_2284_new_n437_), .Y(_abc_2284_new_n439_));
NAND3X1 NAND3X1_61 ( .A(_abc_2284_new_n376_), .B(_abc_2284_new_n412_), .C(_abc_2284_new_n442_), .Y(_abc_2284_new_n443_));
NAND3X1 NAND3X1_62 ( .A(_abc_2284_new_n455_), .B(_abc_2284_new_n454_), .C(_abc_2284_new_n415_), .Y(_abc_2284_new_n456_));
NAND3X1 NAND3X1_63 ( .A(_abc_2284_new_n406_), .B(_abc_2284_new_n408_), .C(_abc_2284_new_n490_), .Y(_abc_2284_new_n491_));
NAND3X1 NAND3X1_64 ( .A(_abc_2284_new_n376_), .B(_abc_2284_new_n492_), .C(_abc_2284_new_n488_), .Y(_abc_2284_new_n493_));
NAND3X1 NAND3X1_65 ( .A(_abc_2284_new_n455_), .B(_abc_2284_new_n494_), .C(_abc_2284_new_n443_), .Y(_abc_2284_new_n495_));
NAND3X1 NAND3X1_66 ( .A(rx), .B(_abc_2284_new_n497_), .C(_abc_2284_new_n496_), .Y(_abc_2284_new_n498_));
NAND3X1 NAND3X1_67 ( .A(_abc_2284_new_n487_), .B(_abc_2284_new_n499_), .C(_abc_2284_new_n498_), .Y(_abc_2284_new_n500_));
NAND3X1 NAND3X1_68 ( .A(rx_bits_remaining_0_), .B(_abc_2284_new_n502_), .C(_abc_2284_new_n503_), .Y(_abc_2284_new_n504_));
NAND3X1 NAND3X1_69 ( .A(_abc_2284_new_n507_), .B(_abc_2284_new_n497_), .C(_abc_2284_new_n496_), .Y(_abc_2284_new_n508_));
NAND3X1 NAND3X1_7 ( .A(_abc_2284_new_n180_), .B(_abc_2284_new_n184_), .C(_abc_2284_new_n182_), .Y(_abc_2284_new_n185_));
NAND3X1 NAND3X1_70 ( .A(_abc_2284_new_n500_), .B(_abc_2284_new_n512_), .C(_abc_2284_new_n506_), .Y(_0recv_state_2_0__0_));
NAND3X1 NAND3X1_71 ( .A(_abc_2284_new_n510_), .B(_abc_2284_new_n515_), .C(_abc_2284_new_n518_), .Y(_0recv_state_2_0__1_));
NAND3X1 NAND3X1_72 ( .A(_abc_2284_new_n521_), .B(_abc_2284_new_n417_), .C(_abc_2284_new_n514_), .Y(_abc_2284_new_n522_));
NAND3X1 NAND3X1_73 ( .A(_abc_2284_new_n522_), .B(_abc_2284_new_n523_), .C(_abc_2284_new_n520_), .Y(_0recv_state_2_0__2_));
NAND3X1 NAND3X1_74 ( .A(_abc_2284_new_n448_), .B(_abc_2284_new_n528_), .C(_abc_2284_new_n527_), .Y(_abc_2284_new_n529_));
NAND3X1 NAND3X1_75 ( .A(_abc_2284_new_n448_), .B(_abc_2284_new_n545_), .C(_abc_2284_new_n544_), .Y(_abc_2284_new_n546_));
NAND3X1 NAND3X1_76 ( .A(_abc_2284_new_n349_), .B(_abc_2284_new_n551_), .C(_abc_2284_new_n222_), .Y(_0tx_clk_divider_10_0__1_));
NAND3X1 NAND3X1_77 ( .A(_abc_2284_new_n553_), .B(_abc_2284_new_n349_), .C(_abc_2284_new_n222_), .Y(_0tx_clk_divider_10_0__2_));
NAND3X1 NAND3X1_78 ( .A(_abc_2284_new_n560_), .B(_abc_2284_new_n349_), .C(_abc_2284_new_n222_), .Y(_0tx_clk_divider_10_0__4_));
NAND3X1 NAND3X1_79 ( .A(_abc_2284_new_n568_), .B(_abc_2284_new_n349_), .C(_abc_2284_new_n222_), .Y(_0tx_clk_divider_10_0__8_));
NAND3X1 NAND3X1_8 ( .A(_abc_2284_new_n187_), .B(_abc_2284_new_n158_), .C(_abc_2284_new_n159_), .Y(_abc_2284_new_n188_));
NAND3X1 NAND3X1_80 ( .A(_abc_2284_new_n199_), .B(_abc_2284_new_n349_), .C(_abc_2284_new_n222_), .Y(_0tx_clk_divider_10_0__10_));
NAND3X1 NAND3X1_81 ( .A(_abc_2284_new_n574_), .B(_abc_2284_new_n575_), .C(_abc_2284_new_n493_), .Y(_0rx_clk_divider_10_0__1_));
NAND3X1 NAND3X1_82 ( .A(_abc_2284_new_n577_), .B(_abc_2284_new_n429_), .C(_abc_2284_new_n493_), .Y(_0rx_clk_divider_10_0__2_));
NAND3X1 NAND3X1_83 ( .A(_abc_2284_new_n581_), .B(_abc_2284_new_n429_), .C(_abc_2284_new_n493_), .Y(_0rx_clk_divider_10_0__4_));
NAND3X1 NAND3X1_84 ( .A(_abc_2284_new_n587_), .B(_abc_2284_new_n429_), .C(_abc_2284_new_n493_), .Y(_0rx_clk_divider_10_0__8_));
NAND3X1 NAND3X1_85 ( .A(_abc_2284_new_n590_), .B(_abc_2284_new_n429_), .C(_abc_2284_new_n413_), .Y(_0rx_clk_divider_10_0__10_));
NAND3X1 NAND3X1_9 ( .A(_abc_2284_new_n186_), .B(_abc_2284_new_n188_), .C(_abc_2284_new_n189_), .Y(_abc_2284_new_n190_));
NOR2X1 NOR2X1_1 ( .A(recv_state_0_), .B(recv_state_2_), .Y(_abc_2284_new_n145_));
NOR2X1 NOR2X1_10 ( .A(tx_clk_divider_8_), .B(tx_clk_divider_9_), .Y(_abc_2284_new_n164_));
NOR2X1 NOR2X1_11 ( .A(_abc_2284_new_n167_), .B(_abc_2284_new_n168_), .Y(_abc_2284_new_n169_));
NOR2X1 NOR2X1_12 ( .A(tx_clk_divider_1_), .B(_abc_2284_new_n177_), .Y(_abc_2284_new_n178_));
NOR2X1 NOR2X1_13 ( .A(tx_clk_divider_6_), .B(_abc_2284_new_n183_), .Y(_abc_2284_new_n202_));
NOR2X1 NOR2X1_14 ( .A(tx_countdown_0_), .B(tx_countdown_1_), .Y(_abc_2284_new_n211_));
NOR2X1 NOR2X1_15 ( .A(_abc_2284_new_n209_), .B(_abc_2284_new_n220_), .Y(_abc_2284_new_n221_));
NOR2X1 NOR2X1_16 ( .A(_abc_2284_new_n232_), .B(_abc_2284_new_n227_), .Y(_abc_2284_new_n233_));
NOR2X1 NOR2X1_17 ( .A(tx_bits_remaining_1_), .B(tx_bits_remaining_0_), .Y(_abc_2284_new_n234_));
NOR2X1 NOR2X1_18 ( .A(tx_bits_remaining_3_), .B(tx_bits_remaining_2_), .Y(_abc_2284_new_n235_));
NOR2X1 NOR2X1_19 ( .A(_abc_2284_new_n248_), .B(_abc_2284_new_n249_), .Y(_abc_2284_new_n250_));
NOR2X1 NOR2X1_2 ( .A(recv_state_0_), .B(_abc_2284_new_n150_), .Y(received));
NOR2X1 NOR2X1_20 ( .A(_abc_2284_new_n254_), .B(_abc_2284_new_n257_), .Y(_abc_2284_new_n258_));
NOR2X1 NOR2X1_21 ( .A(rst), .B(_abc_2284_new_n147_), .Y(_abc_2284_new_n259_));
NOR2X1 NOR2X1_22 ( .A(_abc_2284_new_n320_), .B(_abc_2284_new_n321_), .Y(_abc_2284_new_n322_));
NOR2X1 NOR2X1_23 ( .A(_abc_2284_new_n319_), .B(_abc_2284_new_n261_), .Y(_abc_2284_new_n324_));
NOR2X1 NOR2X1_24 ( .A(_abc_2284_new_n258_), .B(_abc_2284_new_n208_), .Y(_0tx_countdown_5_0__0_));
NOR2X1 NOR2X1_25 ( .A(_abc_2284_new_n258_), .B(_abc_2284_new_n196_), .Y(_0tx_countdown_5_0__1_));
NOR2X1 NOR2X1_26 ( .A(_abc_2284_new_n258_), .B(_abc_2284_new_n249_), .Y(_abc_2284_new_n360_));
NOR2X1 NOR2X1_27 ( .A(_abc_2284_new_n258_), .B(_abc_2284_new_n325_), .Y(_0tx_countdown_5_0__4_));
NOR2X1 NOR2X1_28 ( .A(_abc_2284_new_n371_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n372_));
NOR2X1 NOR2X1_29 ( .A(rx_clk_divider_2_), .B(rx_clk_divider_3_), .Y(_abc_2284_new_n377_));
NOR2X1 NOR2X1_3 ( .A(recv_state_1_), .B(_abc_2284_new_n152_), .Y(recv_error));
NOR2X1 NOR2X1_30 ( .A(rx_clk_divider_1_), .B(rx_clk_divider_0_), .Y(_abc_2284_new_n378_));
NOR2X1 NOR2X1_31 ( .A(_abc_2284_new_n382_), .B(_abc_2284_new_n385_), .Y(_abc_2284_new_n386_));
NOR2X1 NOR2X1_32 ( .A(rx_clk_divider_8_), .B(rx_clk_divider_9_), .Y(_abc_2284_new_n387_));
NOR2X1 NOR2X1_33 ( .A(rx_clk_divider_4_), .B(rx_clk_divider_5_), .Y(_abc_2284_new_n390_));
NOR2X1 NOR2X1_34 ( .A(rst), .B(_abc_2284_new_n144_), .Y(_abc_2284_new_n421_));
NOR2X1 NOR2X1_35 ( .A(recv_state_2_), .B(_abc_2284_new_n422_), .Y(_abc_2284_new_n423_));
NOR2X1 NOR2X1_36 ( .A(_abc_2284_new_n421_), .B(_abc_2284_new_n423_), .Y(_abc_2284_new_n424_));
NOR2X1 NOR2X1_37 ( .A(_abc_2284_new_n426_), .B(_abc_2284_new_n415_), .Y(_0rx_countdown_5_0__0_));
NOR2X1 NOR2X1_38 ( .A(rx), .B(_abc_2284_new_n418_), .Y(_abc_2284_new_n428_));
NOR2X1 NOR2X1_39 ( .A(rx_clk_divider_1_), .B(_abc_2284_new_n436_), .Y(_abc_2284_new_n437_));
NOR2X1 NOR2X1_4 ( .A(rst), .B(_abc_2284_new_n148_), .Y(_abc_2284_new_n154_));
NOR2X1 NOR2X1_40 ( .A(_abc_2284_new_n441_), .B(_abc_2284_new_n432_), .Y(_abc_2284_new_n442_));
NOR2X1 NOR2X1_41 ( .A(_abc_2284_new_n419_), .B(_abc_2284_new_n425_), .Y(_abc_2284_new_n445_));
NOR2X1 NOR2X1_42 ( .A(rx_countdown_1_), .B(rx_countdown_4_), .Y(_abc_2284_new_n455_));
NOR2X1 NOR2X1_43 ( .A(_abc_2284_new_n450_), .B(_abc_2284_new_n459_), .Y(_abc_2284_new_n460_));
NOR2X1 NOR2X1_44 ( .A(_abc_2284_new_n470_), .B(_abc_2284_new_n456_), .Y(_abc_2284_new_n471_));
NOR2X1 NOR2X1_45 ( .A(recv_state_1_), .B(_abc_2284_new_n473_), .Y(_abc_2284_new_n474_));
NOR2X1 NOR2X1_46 ( .A(_abc_2284_new_n426_), .B(_abc_2284_new_n484_), .Y(_0rx_countdown_5_0__4_));
NOR2X1 NOR2X1_47 ( .A(_abc_2284_new_n426_), .B(_abc_2284_new_n465_), .Y(_0rx_countdown_5_0__5_));
NOR2X1 NOR2X1_48 ( .A(_abc_2284_new_n144_), .B(_abc_2284_new_n473_), .Y(_abc_2284_new_n487_));
NOR2X1 NOR2X1_49 ( .A(_abc_2284_new_n489_), .B(_abc_2284_new_n491_), .Y(_abc_2284_new_n492_));
NOR2X1 NOR2X1_5 ( .A(tx_state_1_), .B(_abc_2284_new_n155_), .Y(_abc_2284_new_n156_));
NOR2X1 NOR2X1_50 ( .A(_abc_2284_new_n477_), .B(_abc_2284_new_n495_), .Y(_abc_2284_new_n496_));
NOR2X1 NOR2X1_51 ( .A(rx_bits_remaining_2_), .B(rx_bits_remaining_3_), .Y(_abc_2284_new_n503_));
NOR2X1 NOR2X1_52 ( .A(rst), .B(_abc_2284_new_n152_), .Y(_abc_2284_new_n509_));
NOR2X1 NOR2X1_53 ( .A(rst), .B(_abc_2284_new_n416_), .Y(_abc_2284_new_n521_));
NOR2X1 NOR2X1_54 ( .A(rx_bits_remaining_0_), .B(rx_bits_remaining_1_), .Y(_abc_2284_new_n536_));
NOR2X1 NOR2X1_55 ( .A(tx_clk_divider_0_), .B(_abc_2284_new_n258_), .Y(_0tx_clk_divider_10_0__0_));
NOR2X1 NOR2X1_56 ( .A(_abc_2284_new_n159_), .B(_abc_2284_new_n550_), .Y(_abc_2284_new_n551_));
NOR2X1 NOR2X1_57 ( .A(_abc_2284_new_n187_), .B(_abc_2284_new_n160_), .Y(_abc_2284_new_n559_));
NOR2X1 NOR2X1_58 ( .A(_abc_2284_new_n558_), .B(_abc_2284_new_n559_), .Y(_abc_2284_new_n560_));
NOR2X1 NOR2X1_59 ( .A(rx_clk_divider_0_), .B(_abc_2284_new_n428_), .Y(_0rx_clk_divider_10_0__0_));
NOR2X1 NOR2X1_6 ( .A(tx_clk_divider_2_), .B(tx_clk_divider_3_), .Y(_abc_2284_new_n158_));
NOR2X1 NOR2X1_60 ( .A(_abc_2284_new_n407_), .B(_abc_2284_new_n435_), .Y(_abc_2284_new_n581_));
NOR2X1 NOR2X1_61 ( .A(_abc_2284_new_n428_), .B(_abc_2284_new_n434_), .Y(_0rx_clk_divider_10_0__7_));
NOR2X1 NOR2X1_62 ( .A(_abc_2284_new_n428_), .B(_abc_2284_new_n488_), .Y(_0rx_clk_divider_10_0__9_));
NOR2X1 NOR2X1_7 ( .A(tx_clk_divider_1_), .B(tx_clk_divider_0_), .Y(_abc_2284_new_n159_));
NOR2X1 NOR2X1_8 ( .A(tx_clk_divider_4_), .B(tx_clk_divider_5_), .Y(_abc_2284_new_n161_));
NOR2X1 NOR2X1_9 ( .A(tx_clk_divider_6_), .B(tx_clk_divider_7_), .Y(_abc_2284_new_n162_));
NOR3X1 NOR3X1_1 ( .A(_abc_2284_new_n179_), .B(_abc_2284_new_n190_), .C(_abc_2284_new_n185_), .Y(_abc_2284_new_n191_));
NOR3X1 NOR3X1_2 ( .A(tx_clk_divider_7_), .B(_abc_2284_new_n202_), .C(_abc_2284_new_n203_), .Y(_abc_2284_new_n204_));
NOR3X1 NOR3X1_3 ( .A(_abc_2284_new_n227_), .B(_abc_2284_new_n220_), .C(_abc_2284_new_n326_), .Y(_abc_2284_new_n327_));
NOR3X1 NOR3X1_4 ( .A(tx_state_1_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n251_), .Y(_abc_2284_new_n367_));
NOR3X1 NOR3X1_5 ( .A(_abc_2284_new_n401_), .B(_abc_2284_new_n409_), .C(_abc_2284_new_n405_), .Y(_abc_2284_new_n410_));
NOR3X1 NOR3X1_6 ( .A(rx_clk_divider_5_), .B(rx_clk_divider_6_), .C(rx_clk_divider_8_), .Y(_abc_2284_new_n438_));
NOR3X1 NOR3X1_7 ( .A(_abc_2284_new_n407_), .B(_abc_2284_new_n439_), .C(_abc_2284_new_n435_), .Y(_abc_2284_new_n440_));
NOR3X1 NOR3X1_8 ( .A(rx), .B(_abc_2284_new_n470_), .C(_abc_2284_new_n456_), .Y(_abc_2284_new_n478_));
NOR3X1 NOR3X1_9 ( .A(_abc_2284_new_n504_), .B(_abc_2284_new_n470_), .C(_abc_2284_new_n456_), .Y(_abc_2284_new_n505_));
OAI21X1 OAI21X1_1 ( .A(_abc_2284_new_n167_), .B(_abc_2284_new_n168_), .C(tx_clk_divider_8_), .Y(_abc_2284_new_n174_));
OAI21X1 OAI21X1_10 ( .A(_abc_2284_new_n210_), .B(_abc_2284_new_n192_), .C(_abc_2284_new_n218_), .Y(_abc_2284_new_n249_));
OAI21X1 OAI21X1_11 ( .A(tx_state_1_), .B(tx_state_0_), .C(_abc_2284_new_n255_), .Y(_abc_2284_new_n256_));
OAI21X1 OAI21X1_12 ( .A(transmit), .B(_abc_2284_new_n154_), .C(_abc_2284_new_n260_), .Y(_abc_2284_new_n261_));
OAI21X1 OAI21X1_13 ( .A(tx_data_1_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n265_), .Y(_abc_2284_new_n266_));
OAI21X1 OAI21X1_14 ( .A(tx_data_2_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n273_), .Y(_abc_2284_new_n274_));
OAI21X1 OAI21X1_15 ( .A(tx_data_3_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n281_), .Y(_abc_2284_new_n282_));
OAI21X1 OAI21X1_16 ( .A(tx_data_4_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n289_), .Y(_abc_2284_new_n290_));
OAI21X1 OAI21X1_17 ( .A(tx_data_5_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n297_), .Y(_abc_2284_new_n298_));
OAI21X1 OAI21X1_18 ( .A(tx_data_6_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n305_), .Y(_abc_2284_new_n306_));
OAI21X1 OAI21X1_19 ( .A(_abc_2284_new_n254_), .B(\tx_byte[7] ), .C(_abc_2284_new_n312_), .Y(_abc_2284_new_n313_));
OAI21X1 OAI21X1_2 ( .A(_abc_2284_new_n206_), .B(_abc_2284_new_n201_), .C(_abc_2284_new_n198_), .Y(_abc_2284_new_n207_));
OAI21X1 OAI21X1_20 ( .A(_abc_2284_new_n330_), .B(_abc_2284_new_n331_), .C(_abc_2284_new_n337_), .Y(_0tx_bits_remaining_3_0__1_));
OAI21X1 OAI21X1_21 ( .A(tx_bits_remaining_1_), .B(tx_bits_remaining_0_), .C(_abc_2284_new_n340_), .Y(_abc_2284_new_n341_));
OAI21X1 OAI21X1_22 ( .A(tx_bits_remaining_2_), .B(_abc_2284_new_n350_), .C(tx_bits_remaining_3_), .Y(_abc_2284_new_n351_));
OAI21X1 OAI21X1_23 ( .A(_abc_2284_new_n259_), .B(_abc_2284_new_n155_), .C(tx_bits_remaining_3_), .Y(_abc_2284_new_n356_));
OAI21X1 OAI21X1_24 ( .A(_abc_2284_new_n321_), .B(_abc_2284_new_n315_), .C(_abc_2284_new_n360_), .Y(_0tx_countdown_5_0__2_));
OAI21X1 OAI21X1_25 ( .A(_abc_2284_new_n320_), .B(_abc_2284_new_n251_), .C(_abc_2284_new_n156_), .Y(_abc_2284_new_n362_));
OAI21X1 OAI21X1_26 ( .A(_abc_2284_new_n155_), .B(_abc_2284_new_n367_), .C(_abc_2284_new_n349_), .Y(_0tx_state_1_0__0_));
OAI21X1 OAI21X1_27 ( .A(tx), .B(_abc_2284_new_n327_), .C(_abc_2284_new_n156_), .Y(_abc_2284_new_n373_));
OAI21X1 OAI21X1_28 ( .A(_abc_2284_new_n372_), .B(_abc_2284_new_n373_), .C(_abc_2284_new_n374_), .Y(_0tx_out_0_0_));
OAI21X1 OAI21X1_29 ( .A(_abc_2284_new_n385_), .B(_abc_2284_new_n391_), .C(_abc_2284_new_n387_), .Y(_abc_2284_new_n392_));
OAI21X1 OAI21X1_3 ( .A(_abc_2284_new_n206_), .B(_abc_2284_new_n201_), .C(tx_countdown_2_), .Y(_abc_2284_new_n219_));
OAI21X1 OAI21X1_30 ( .A(_abc_2284_new_n385_), .B(_abc_2284_new_n391_), .C(rx_clk_divider_8_), .Y(_abc_2284_new_n397_));
OAI21X1 OAI21X1_31 ( .A(_abc_2284_new_n382_), .B(_abc_2284_new_n403_), .C(rx_clk_divider_6_), .Y(_abc_2284_new_n404_));
OAI21X1 OAI21X1_32 ( .A(recv_state_1_), .B(recv_state_0_), .C(_abc_2284_new_n255_), .Y(_abc_2284_new_n417_));
OAI21X1 OAI21X1_33 ( .A(_abc_2284_new_n416_), .B(rst), .C(_abc_2284_new_n417_), .Y(_abc_2284_new_n418_));
OAI21X1 OAI21X1_34 ( .A(recv_state_0_), .B(_abc_2284_new_n420_), .C(_abc_2284_new_n424_), .Y(_abc_2284_new_n425_));
OAI21X1 OAI21X1_35 ( .A(rx_clk_divider_8_), .B(_abc_2284_new_n430_), .C(rx_clk_divider_9_), .Y(_abc_2284_new_n431_));
OAI21X1 OAI21X1_36 ( .A(rx_clk_divider_6_), .B(_abc_2284_new_n391_), .C(rx_clk_divider_7_), .Y(_abc_2284_new_n433_));
OAI21X1 OAI21X1_37 ( .A(_abc_2284_new_n445_), .B(_abc_2284_new_n444_), .C(_abc_2284_new_n429_), .Y(_0rx_countdown_5_0__1_));
OAI21X1 OAI21X1_38 ( .A(rx_countdown_2_), .B(_abc_2284_new_n450_), .C(rx_countdown_3_), .Y(_abc_2284_new_n466_));
OAI21X1 OAI21X1_39 ( .A(_abc_2284_new_n450_), .B(_abc_2284_new_n459_), .C(_abc_2284_new_n466_), .Y(_abc_2284_new_n467_));
OAI21X1 OAI21X1_4 ( .A(_abc_2284_new_n206_), .B(_abc_2284_new_n201_), .C(tx_countdown_5_), .Y(_abc_2284_new_n226_));
OAI21X1 OAI21X1_40 ( .A(_abc_2284_new_n413_), .B(_abc_2284_new_n475_), .C(_abc_2284_new_n476_), .Y(_abc_2284_new_n477_));
OAI21X1 OAI21X1_41 ( .A(_abc_2284_new_n426_), .B(_abc_2284_new_n479_), .C(_abc_2284_new_n472_), .Y(_0rx_countdown_5_0__2_));
OAI21X1 OAI21X1_42 ( .A(_abc_2284_new_n426_), .B(_abc_2284_new_n469_), .C(_abc_2284_new_n481_), .Y(_0rx_countdown_5_0__3_));
OAI21X1 OAI21X1_43 ( .A(_abc_2284_new_n391_), .B(_abc_2284_new_n385_), .C(_abc_2284_new_n433_), .Y(_abc_2284_new_n489_));
OAI21X1 OAI21X1_44 ( .A(_abc_2284_new_n470_), .B(_abc_2284_new_n456_), .C(_abc_2284_new_n422_), .Y(_abc_2284_new_n499_));
OAI21X1 OAI21X1_45 ( .A(_abc_2284_new_n505_), .B(_abc_2284_new_n501_), .C(_abc_2284_new_n448_), .Y(_abc_2284_new_n506_));
OAI21X1 OAI21X1_46 ( .A(rx), .B(_abc_2284_new_n418_), .C(_abc_2284_new_n510_), .Y(_abc_2284_new_n511_));
OAI21X1 OAI21X1_47 ( .A(rx), .B(_abc_2284_new_n514_), .C(_abc_2284_new_n487_), .Y(_abc_2284_new_n515_));
OAI21X1 OAI21X1_48 ( .A(recv_state_1_), .B(_abc_2284_new_n473_), .C(_abc_2284_new_n447_), .Y(_abc_2284_new_n517_));
OAI21X1 OAI21X1_49 ( .A(_abc_2284_new_n516_), .B(_abc_2284_new_n478_), .C(_abc_2284_new_n517_), .Y(_abc_2284_new_n518_));
OAI21X1 OAI21X1_5 ( .A(_abc_2284_new_n222_), .B(_abc_2284_new_n225_), .C(_abc_2284_new_n226_), .Y(_abc_2284_new_n227_));
OAI21X1 OAI21X1_50 ( .A(_abc_2284_new_n516_), .B(_abc_2284_new_n508_), .C(_abc_2284_new_n447_), .Y(_abc_2284_new_n526_));
OAI21X1 OAI21X1_51 ( .A(_abc_2284_new_n470_), .B(_abc_2284_new_n456_), .C(_abc_2284_new_n525_), .Y(_abc_2284_new_n528_));
OAI21X1 OAI21X1_52 ( .A(_abc_2284_new_n525_), .B(_abc_2284_new_n526_), .C(_abc_2284_new_n529_), .Y(_0rx_bits_remaining_3_0__0_));
OAI21X1 OAI21X1_53 ( .A(_abc_2284_new_n470_), .B(_abc_2284_new_n456_), .C(_abc_2284_new_n502_), .Y(_abc_2284_new_n532_));
OAI21X1 OAI21X1_54 ( .A(_abc_2284_new_n531_), .B(_abc_2284_new_n514_), .C(_abc_2284_new_n532_), .Y(_abc_2284_new_n533_));
OAI21X1 OAI21X1_55 ( .A(_abc_2284_new_n470_), .B(_abc_2284_new_n456_), .C(_abc_2284_new_n535_), .Y(_abc_2284_new_n538_));
OAI21X1 OAI21X1_56 ( .A(_abc_2284_new_n537_), .B(_abc_2284_new_n514_), .C(_abc_2284_new_n538_), .Y(_abc_2284_new_n539_));
OAI21X1 OAI21X1_57 ( .A(_abc_2284_new_n470_), .B(_abc_2284_new_n456_), .C(_abc_2284_new_n541_), .Y(_abc_2284_new_n545_));
OAI21X1 OAI21X1_58 ( .A(tx_clk_divider_2_), .B(_abc_2284_new_n555_), .C(tx_clk_divider_3_), .Y(_abc_2284_new_n556_));
OAI21X1 OAI21X1_59 ( .A(tx_clk_divider_4_), .B(_abc_2284_new_n167_), .C(tx_clk_divider_5_), .Y(_abc_2284_new_n562_));
OAI21X1 OAI21X1_6 ( .A(_abc_2284_new_n228_), .B(_abc_2284_new_n192_), .C(_abc_2284_new_n231_), .Y(_abc_2284_new_n232_));
OAI21X1 OAI21X1_60 ( .A(tx_clk_divider_6_), .B(_abc_2284_new_n183_), .C(tx_clk_divider_7_), .Y(_abc_2284_new_n566_));
OAI21X1 OAI21X1_61 ( .A(tx_clk_divider_8_), .B(_abc_2284_new_n565_), .C(tx_clk_divider_9_), .Y(_abc_2284_new_n570_));
OAI21X1 OAI21X1_62 ( .A(rx_clk_divider_2_), .B(_abc_2284_new_n574_), .C(rx_clk_divider_3_), .Y(_abc_2284_new_n579_));
OAI21X1 OAI21X1_63 ( .A(rx_clk_divider_4_), .B(_abc_2284_new_n403_), .C(rx_clk_divider_5_), .Y(_abc_2284_new_n583_));
OAI21X1 OAI21X1_64 ( .A(_abc_2284_new_n447_), .B(_abc_2284_new_n514_), .C(\rx_byte[7] ), .Y(_abc_2284_new_n607_));
OAI21X1 OAI21X1_65 ( .A(_abc_2284_new_n507_), .B(_abc_2284_new_n472_), .C(_abc_2284_new_n607_), .Y(_0rx_data_7_0__7_));
OAI21X1 OAI21X1_7 ( .A(tx_data_0_), .B(_abc_2284_new_n236_), .C(_abc_2284_new_n238_), .Y(_abc_2284_new_n239_));
OAI21X1 OAI21X1_8 ( .A(_abc_2284_new_n206_), .B(_abc_2284_new_n201_), .C(tx_countdown_1_), .Y(_abc_2284_new_n243_));
OAI21X1 OAI21X1_9 ( .A(_abc_2284_new_n206_), .B(_abc_2284_new_n201_), .C(tx_countdown_3_), .Y(_abc_2284_new_n247_));
OAI22X1 OAI22X1_1 ( .A(_abc_2284_new_n447_), .B(_abc_2284_new_n533_), .C(_abc_2284_new_n502_), .D(_abc_2284_new_n526_), .Y(_0rx_bits_remaining_3_0__1_));
OAI22X1 OAI22X1_2 ( .A(_abc_2284_new_n447_), .B(_abc_2284_new_n539_), .C(_abc_2284_new_n535_), .D(_abc_2284_new_n526_), .Y(_0rx_bits_remaining_3_0__2_));
OR2X2 OR2X2_1 ( .A(_abc_2284_new_n223_), .B(tx_countdown_4_), .Y(_abc_2284_new_n224_));
OR2X2 OR2X2_2 ( .A(_abc_2284_new_n313_), .B(_abc_2284_new_n257_), .Y(_abc_2284_new_n314_));
OR2X2 OR2X2_3 ( .A(rx_countdown_0_), .B(rx_countdown_1_), .Y(_abc_2284_new_n450_));
OR2X2 OR2X2_4 ( .A(_abc_2284_new_n498_), .B(_abc_2284_new_n516_), .Y(_abc_2284_new_n520_));
XNOR2X1 XNOR2X1_1 ( .A(tx_countdown_0_), .B(tx_countdown_1_), .Y(_abc_2284_new_n193_));
XNOR2X1 XNOR2X1_10 ( .A(_abc_2284_new_n542_), .B(_abc_2284_new_n541_), .Y(_abc_2284_new_n543_));
XNOR2X1 XNOR2X1_11 ( .A(_abc_2284_new_n159_), .B(tx_clk_divider_2_), .Y(_abc_2284_new_n553_));
XNOR2X1 XNOR2X1_12 ( .A(_abc_2284_new_n378_), .B(rx_clk_divider_2_), .Y(_abc_2284_new_n577_));
XNOR2X1 XNOR2X1_2 ( .A(_abc_2284_new_n212_), .B(tx_countdown_3_), .Y(_abc_2284_new_n213_));
XNOR2X1 XNOR2X1_3 ( .A(_abc_2284_new_n211_), .B(_abc_2284_new_n210_), .Y(_abc_2284_new_n217_));
XNOR2X1 XNOR2X1_4 ( .A(_abc_2284_new_n450_), .B(rx_countdown_2_), .Y(_abc_2284_new_n451_));
XNOR2X1 XNOR2X1_5 ( .A(_abc_2284_new_n461_), .B(rx_countdown_5_), .Y(_abc_2284_new_n462_));
XNOR2X1 XNOR2X1_6 ( .A(_abc_2284_new_n460_), .B(_abc_2284_new_n457_), .Y(_abc_2284_new_n483_));
XNOR2X1 XNOR2X1_7 ( .A(_abc_2284_new_n396_), .B(_abc_2284_new_n394_), .Y(_abc_2284_new_n488_));
XNOR2X1 XNOR2X1_8 ( .A(rx_bits_remaining_0_), .B(rx_bits_remaining_1_), .Y(_abc_2284_new_n531_));
XNOR2X1 XNOR2X1_9 ( .A(_abc_2284_new_n536_), .B(_abc_2284_new_n535_), .Y(_abc_2284_new_n537_));
XOR2X1 XOR2X1_1 ( .A(_abc_2284_new_n224_), .B(tx_countdown_5_), .Y(_abc_2284_new_n225_));
XOR2X1 XOR2X1_2 ( .A(_abc_2284_new_n443_), .B(rx_countdown_1_), .Y(_abc_2284_new_n444_));


endmodule