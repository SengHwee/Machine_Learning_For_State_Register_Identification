module mc_top(clk_i, rst_i, \wb_data_i[0] , \wb_data_i[1] , \wb_data_i[2] , \wb_data_i[3] , \wb_data_i[4] , \wb_data_i[5] , \wb_data_i[6] , \wb_data_i[7] , \wb_data_i[8] , \wb_data_i[9] , \wb_data_i[10] , \wb_data_i[11] , \wb_data_i[12] , \wb_data_i[13] , \wb_data_i[14] , \wb_data_i[15] , \wb_data_i[16] , \wb_data_i[17] , \wb_data_i[18] , \wb_data_i[19] , \wb_data_i[20] , \wb_data_i[21] , \wb_data_i[22] , \wb_data_i[23] , \wb_data_i[24] , \wb_data_i[25] , \wb_data_i[26] , \wb_data_i[27] , \wb_data_i[28] , \wb_data_i[29] , \wb_data_i[30] , \wb_data_i[31] , \wb_addr_i[0] , \wb_addr_i[1] , \wb_addr_i[2] , \wb_addr_i[3] , \wb_addr_i[4] , \wb_addr_i[5] , \wb_addr_i[6] , \wb_addr_i[7] , \wb_addr_i[8] , \wb_addr_i[9] , \wb_addr_i[10] , \wb_addr_i[11] , \wb_addr_i[12] , \wb_addr_i[13] , \wb_addr_i[14] , \wb_addr_i[15] , \wb_addr_i[16] , \wb_addr_i[17] , \wb_addr_i[18] , \wb_addr_i[19] , \wb_addr_i[20] , \wb_addr_i[21] , \wb_addr_i[22] , \wb_addr_i[23] , \wb_addr_i[24] , \wb_addr_i[25] , \wb_addr_i[26] , \wb_addr_i[27] , \wb_addr_i[28] , \wb_addr_i[29] , \wb_addr_i[30] , \wb_addr_i[31] , \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] , \wb_sel_i[3] , wb_we_i, wb_cyc_i, wb_stb_i, susp_req_i, resume_req_i, mc_clk_i, mc_br_pad_i, mc_ack_pad_i, \mc_data_pad_i[0] , \mc_data_pad_i[1] , \mc_data_pad_i[2] , \mc_data_pad_i[3] , \mc_data_pad_i[4] , \mc_data_pad_i[5] , \mc_data_pad_i[6] , \mc_data_pad_i[7] , \mc_data_pad_i[8] , \mc_data_pad_i[9] , \mc_data_pad_i[10] , \mc_data_pad_i[11] , \mc_data_pad_i[12] , \mc_data_pad_i[13] , \mc_data_pad_i[14] , \mc_data_pad_i[15] , \mc_data_pad_i[16] , \mc_data_pad_i[17] , \mc_data_pad_i[18] , \mc_data_pad_i[19] , \mc_data_pad_i[20] , \mc_data_pad_i[21] , \mc_data_pad_i[22] , \mc_data_pad_i[23] , \mc_data_pad_i[24] , \mc_data_pad_i[25] , \mc_data_pad_i[26] , \mc_data_pad_i[27] , \mc_data_pad_i[28] , \mc_data_pad_i[29] , \mc_data_pad_i[30] , \mc_data_pad_i[31] , \mc_dp_pad_i[0] , \mc_dp_pad_i[1] , \mc_dp_pad_i[2] , \mc_dp_pad_i[3] , mc_sts_pad_i, \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] , \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] , \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] , \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] , \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] , \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] , \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] , \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] , wb_ack_o, wb_err_o, suspended_o, \poc_o[0] , \poc_o[1] , \poc_o[2] , \poc_o[3] , \poc_o[4] , \poc_o[5] , \poc_o[6] , \poc_o[7] , \poc_o[8] , \poc_o[9] , \poc_o[10] , \poc_o[11] , \poc_o[12] , \poc_o[13] , \poc_o[14] , \poc_o[15] , \poc_o[16] , \poc_o[17] , \poc_o[18] , \poc_o[19] , \poc_o[20] , \poc_o[21] , \poc_o[22] , \poc_o[23] , \poc_o[24] , \poc_o[25] , \poc_o[26] , \poc_o[27] , \poc_o[28] , \poc_o[29] , \poc_o[30] , \poc_o[31] , mc_bg_pad_o, \mc_addr_pad_o[0] , \mc_addr_pad_o[1] , \mc_addr_pad_o[2] , \mc_addr_pad_o[3] , \mc_addr_pad_o[4] , \mc_addr_pad_o[5] , \mc_addr_pad_o[6] , \mc_addr_pad_o[7] , \mc_addr_pad_o[8] , \mc_addr_pad_o[9] , \mc_addr_pad_o[10] , \mc_addr_pad_o[11] , \mc_addr_pad_o[12] , \mc_addr_pad_o[13] , \mc_addr_pad_o[14] , \mc_addr_pad_o[15] , \mc_addr_pad_o[16] , \mc_addr_pad_o[17] , \mc_addr_pad_o[18] , \mc_addr_pad_o[19] , \mc_addr_pad_o[20] , \mc_addr_pad_o[21] , \mc_addr_pad_o[22] , \mc_addr_pad_o[23] , \mc_data_pad_o[0] , \mc_data_pad_o[1] , \mc_data_pad_o[2] , \mc_data_pad_o[3] , \mc_data_pad_o[4] , \mc_data_pad_o[5] , \mc_data_pad_o[6] , \mc_data_pad_o[7] , \mc_data_pad_o[8] , \mc_data_pad_o[9] , \mc_data_pad_o[10] , \mc_data_pad_o[11] , \mc_data_pad_o[12] , \mc_data_pad_o[13] , \mc_data_pad_o[14] , \mc_data_pad_o[15] , \mc_data_pad_o[16] , \mc_data_pad_o[17] , \mc_data_pad_o[18] , \mc_data_pad_o[19] , \mc_data_pad_o[20] , \mc_data_pad_o[21] , \mc_data_pad_o[22] , \mc_data_pad_o[23] , \mc_data_pad_o[24] , \mc_data_pad_o[25] , \mc_data_pad_o[26] , \mc_data_pad_o[27] , \mc_data_pad_o[28] , \mc_data_pad_o[29] , \mc_data_pad_o[30] , \mc_data_pad_o[31] , \mc_dp_pad_o[0] , \mc_dp_pad_o[1] , \mc_dp_pad_o[2] , \mc_dp_pad_o[3] , mc_doe_pad_doe_o, \mc_dqm_pad_o[0] , \mc_dqm_pad_o[1] , \mc_dqm_pad_o[2] , \mc_dqm_pad_o[3] , mc_oe_pad_o_, mc_we_pad_o_, mc_cas_pad_o_, mc_ras_pad_o_, mc_cke_pad_o_, \mc_cs_pad_o_[0] , \mc_cs_pad_o_[1] , \mc_cs_pad_o_[2] , \mc_cs_pad_o_[3] , \mc_cs_pad_o_[4] , \mc_cs_pad_o_[5] , \mc_cs_pad_o_[6] , \mc_cs_pad_o_[7] , mc_rp_pad_o_, mc_vpen_pad_o, mc_adsc_pad_o_, mc_adv_pad_o_, mc_zz_pad_o, mc_coe_pad_coe_o);

wire _abc_81086_new_n236_; 
wire _abc_81086_new_n238_; 
wire _abc_81086_new_n239_; 
wire _abc_81086_new_n240_; 
wire _abc_81086_new_n241_; 
wire _abc_81086_new_n243_; 
wire _abc_81086_new_n244_; 
wire _abc_81086_new_n245_; 
wire _abc_81086_new_n247_; 
wire _abc_81086_new_n248_; 
wire _abc_81086_new_n249_; 
wire _abc_81086_new_n251_; 
wire _abc_81086_new_n252_; 
wire _abc_81086_new_n253_; 
wire _abc_81086_new_n255_; 
wire _abc_81086_new_n256_; 
wire _abc_81086_new_n257_; 
wire _abc_81086_new_n259_; 
wire _abc_81086_new_n260_; 
wire _abc_81086_new_n261_; 
wire _abc_81086_new_n263_; 
wire _abc_81086_new_n264_; 
wire _abc_81086_new_n265_; 
wire _abc_81086_new_n267_; 
wire _abc_81086_new_n268_; 
wire _abc_81086_new_n269_; 
wire _abc_81086_new_n271_; 
wire _abc_81086_new_n272_; 
wire _abc_81086_new_n274_; 
wire _abc_81086_new_n275_; 
wire _abc_81086_new_n277_; 
wire _abc_81086_new_n278_; 
wire _abc_81086_new_n280_; 
wire _abc_81086_new_n281_; 
wire _abc_81086_new_n283_; 
wire _abc_81086_new_n284_; 
wire _abc_81086_new_n286_; 
wire _abc_81086_new_n287_; 
wire _abc_81086_new_n289_; 
wire _abc_81086_new_n290_; 
wire _abc_81086_new_n292_; 
wire _abc_81086_new_n293_; 
wire _abc_81086_new_n295_; 
wire _abc_81086_new_n296_; 
wire _abc_81086_new_n298_; 
wire _abc_81086_new_n299_; 
wire _abc_81086_new_n301_; 
wire _abc_81086_new_n302_; 
wire _abc_81086_new_n304_; 
wire _abc_81086_new_n305_; 
wire _abc_81086_new_n307_; 
wire _abc_81086_new_n308_; 
wire _abc_81086_new_n310_; 
wire _abc_81086_new_n311_; 
wire _abc_81086_new_n313_; 
wire _abc_81086_new_n314_; 
wire _abc_81086_new_n316_; 
wire _abc_81086_new_n317_; 
wire _abc_81086_new_n319_; 
wire _abc_81086_new_n320_; 
wire _abc_81086_new_n322_; 
wire _abc_81086_new_n323_; 
wire _abc_81086_new_n325_; 
wire _abc_81086_new_n326_; 
wire _abc_81086_new_n328_; 
wire _abc_81086_new_n329_; 
wire _abc_81086_new_n331_; 
wire _abc_81086_new_n332_; 
wire _abc_81086_new_n334_; 
wire _abc_81086_new_n335_; 
wire _abc_81086_new_n337_; 
wire _abc_81086_new_n338_; 
wire _abc_81086_new_n340_; 
wire _abc_81086_new_n341_; 
wire _abc_81086_new_n343_; 
wire _abc_81086_new_n344_; 
wire _abc_81086_new_n346_; 
wire _abc_81086_new_n347_; 
wire _abc_81086_new_n349_; 
wire _abc_81086_new_n350_; 
wire _abc_81086_new_n352_; 
wire _abc_81086_new_n353_; 
wire _abc_81086_new_n370_; 
wire _abc_81086_new_n371_; 
wire _abc_81086_new_n373_; 
wire _abc_81086_new_n374_; 
wire _abc_81086_new_n376_; 
wire _abc_81086_new_n377_; 
wire _abc_81086_new_n379_; 
wire _abc_81086_new_n380_; 
wire _abc_81086_new_n382_; 
wire _abc_81086_new_n383_; 
wire _abc_81086_new_n385_; 
wire _abc_81086_new_n386_; 
wire _abc_81086_new_n388_; 
wire _abc_81086_new_n389_; 
wire _abc_81086_new_n394_; 
wire _abc_81086_new_n395_; 
wire _abc_81086_new_n397_; 
wire _abc_81086_new_n398_; 
wire _abc_81086_new_n463_; 
wire _abc_81086_new_n464_; 
wire _abc_81086_new_n465_; 
wire bank_adr_0_; 
wire bank_adr_1_; 
wire bank_clr; 
wire bank_clr_all; 
wire bank_open; 
wire bank_set; 
wire cas_; 
input clk_i;
wire cmd_a10; 
wire cs_0_; 
wire cs_1_; 
wire cs_2_; 
wire cs_3_; 
wire cs_4_; 
wire cs_5_; 
wire cs_6_; 
wire cs_7_; 
wire cs_en; 
wire cs_le; 
wire cs_le_d; 
wire cs_need_rfr_0_; 
wire cs_need_rfr_1_; 
wire cs_need_rfr_2_; 
wire cs_need_rfr_3_; 
wire cs_need_rfr_4_; 
wire cs_need_rfr_5_; 
wire cs_need_rfr_6_; 
wire cs_need_rfr_7_; 
wire csc_10_; 
wire csc_1_; 
wire csc_2_; 
wire csc_3_; 
wire csc_4_; 
wire csc_5_; 
wire csc_6_; 
wire csc_7_; 
wire csc_9_; 
wire csc_s_1_; 
wire csc_s_2_; 
wire csc_s_3_; 
wire csc_s_4_; 
wire csc_s_5_; 
wire csc_s_6_; 
wire csc_s_7_; 
wire data_oe; 
wire dv; 
wire err; 
wire fs; 
wire init_ack; 
wire init_req; 
wire lmr_ack; 
wire lmr_req; 
wire lmr_sel; 
input mc_ack_pad_i;
wire mc_ack_r; 
wire mc_addr_d_0_; 
wire mc_addr_d_10_; 
wire mc_addr_d_11_; 
wire mc_addr_d_12_; 
wire mc_addr_d_13_; 
wire mc_addr_d_14_; 
wire mc_addr_d_15_; 
wire mc_addr_d_16_; 
wire mc_addr_d_17_; 
wire mc_addr_d_18_; 
wire mc_addr_d_19_; 
wire mc_addr_d_1_; 
wire mc_addr_d_20_; 
wire mc_addr_d_21_; 
wire mc_addr_d_22_; 
wire mc_addr_d_23_; 
wire mc_addr_d_2_; 
wire mc_addr_d_3_; 
wire mc_addr_d_4_; 
wire mc_addr_d_5_; 
wire mc_addr_d_6_; 
wire mc_addr_d_7_; 
wire mc_addr_d_8_; 
wire mc_addr_d_9_; 
output \mc_addr_pad_o[0] ;
output \mc_addr_pad_o[10] ;
output \mc_addr_pad_o[11] ;
output \mc_addr_pad_o[12] ;
output \mc_addr_pad_o[13] ;
output \mc_addr_pad_o[14] ;
output \mc_addr_pad_o[15] ;
output \mc_addr_pad_o[16] ;
output \mc_addr_pad_o[17] ;
output \mc_addr_pad_o[18] ;
output \mc_addr_pad_o[19] ;
output \mc_addr_pad_o[1] ;
output \mc_addr_pad_o[20] ;
output \mc_addr_pad_o[21] ;
output \mc_addr_pad_o[22] ;
output \mc_addr_pad_o[23] ;
output \mc_addr_pad_o[2] ;
output \mc_addr_pad_o[3] ;
output \mc_addr_pad_o[4] ;
output \mc_addr_pad_o[5] ;
output \mc_addr_pad_o[6] ;
output \mc_addr_pad_o[7] ;
output \mc_addr_pad_o[8] ;
output \mc_addr_pad_o[9] ;
wire mc_adsc_d; 
output mc_adsc_pad_o_;
wire mc_adv_d; 
output mc_adv_pad_o_;
wire mc_bg_d; 
output mc_bg_pad_o;
input mc_br_pad_i;
wire mc_br_r; 
wire mc_c_oe_d; 
output mc_cas_pad_o_;
output mc_cke_pad_o_;
input mc_clk_i;
output mc_coe_pad_coe_o;
output \mc_cs_pad_o_[0] ;
output \mc_cs_pad_o_[1] ;
output \mc_cs_pad_o_[2] ;
output \mc_cs_pad_o_[3] ;
output \mc_cs_pad_o_[4] ;
output \mc_cs_pad_o_[5] ;
output \mc_cs_pad_o_[6] ;
output \mc_cs_pad_o_[7] ;
wire mc_data_ir_0_; 
wire mc_data_ir_10_; 
wire mc_data_ir_11_; 
wire mc_data_ir_12_; 
wire mc_data_ir_13_; 
wire mc_data_ir_14_; 
wire mc_data_ir_15_; 
wire mc_data_ir_16_; 
wire mc_data_ir_17_; 
wire mc_data_ir_18_; 
wire mc_data_ir_19_; 
wire mc_data_ir_1_; 
wire mc_data_ir_20_; 
wire mc_data_ir_21_; 
wire mc_data_ir_22_; 
wire mc_data_ir_23_; 
wire mc_data_ir_24_; 
wire mc_data_ir_25_; 
wire mc_data_ir_26_; 
wire mc_data_ir_27_; 
wire mc_data_ir_28_; 
wire mc_data_ir_29_; 
wire mc_data_ir_2_; 
wire mc_data_ir_30_; 
wire mc_data_ir_31_; 
wire mc_data_ir_32_; 
wire mc_data_ir_33_; 
wire mc_data_ir_34_; 
wire mc_data_ir_35_; 
wire mc_data_ir_3_; 
wire mc_data_ir_4_; 
wire mc_data_ir_5_; 
wire mc_data_ir_6_; 
wire mc_data_ir_7_; 
wire mc_data_ir_8_; 
wire mc_data_ir_9_; 
wire mc_data_od_0_; 
wire mc_data_od_10_; 
wire mc_data_od_11_; 
wire mc_data_od_12_; 
wire mc_data_od_13_; 
wire mc_data_od_14_; 
wire mc_data_od_15_; 
wire mc_data_od_16_; 
wire mc_data_od_17_; 
wire mc_data_od_18_; 
wire mc_data_od_19_; 
wire mc_data_od_1_; 
wire mc_data_od_20_; 
wire mc_data_od_21_; 
wire mc_data_od_22_; 
wire mc_data_od_23_; 
wire mc_data_od_24_; 
wire mc_data_od_25_; 
wire mc_data_od_26_; 
wire mc_data_od_27_; 
wire mc_data_od_28_; 
wire mc_data_od_29_; 
wire mc_data_od_2_; 
wire mc_data_od_30_; 
wire mc_data_od_31_; 
wire mc_data_od_3_; 
wire mc_data_od_4_; 
wire mc_data_od_5_; 
wire mc_data_od_6_; 
wire mc_data_od_7_; 
wire mc_data_od_8_; 
wire mc_data_od_9_; 
input \mc_data_pad_i[0] ;
input \mc_data_pad_i[10] ;
input \mc_data_pad_i[11] ;
input \mc_data_pad_i[12] ;
input \mc_data_pad_i[13] ;
input \mc_data_pad_i[14] ;
input \mc_data_pad_i[15] ;
input \mc_data_pad_i[16] ;
input \mc_data_pad_i[17] ;
input \mc_data_pad_i[18] ;
input \mc_data_pad_i[19] ;
input \mc_data_pad_i[1] ;
input \mc_data_pad_i[20] ;
input \mc_data_pad_i[21] ;
input \mc_data_pad_i[22] ;
input \mc_data_pad_i[23] ;
input \mc_data_pad_i[24] ;
input \mc_data_pad_i[25] ;
input \mc_data_pad_i[26] ;
input \mc_data_pad_i[27] ;
input \mc_data_pad_i[28] ;
input \mc_data_pad_i[29] ;
input \mc_data_pad_i[2] ;
input \mc_data_pad_i[30] ;
input \mc_data_pad_i[31] ;
input \mc_data_pad_i[3] ;
input \mc_data_pad_i[4] ;
input \mc_data_pad_i[5] ;
input \mc_data_pad_i[6] ;
input \mc_data_pad_i[7] ;
input \mc_data_pad_i[8] ;
input \mc_data_pad_i[9] ;
output \mc_data_pad_o[0] ;
output \mc_data_pad_o[10] ;
output \mc_data_pad_o[11] ;
output \mc_data_pad_o[12] ;
output \mc_data_pad_o[13] ;
output \mc_data_pad_o[14] ;
output \mc_data_pad_o[15] ;
output \mc_data_pad_o[16] ;
output \mc_data_pad_o[17] ;
output \mc_data_pad_o[18] ;
output \mc_data_pad_o[19] ;
output \mc_data_pad_o[1] ;
output \mc_data_pad_o[20] ;
output \mc_data_pad_o[21] ;
output \mc_data_pad_o[22] ;
output \mc_data_pad_o[23] ;
output \mc_data_pad_o[24] ;
output \mc_data_pad_o[25] ;
output \mc_data_pad_o[26] ;
output \mc_data_pad_o[27] ;
output \mc_data_pad_o[28] ;
output \mc_data_pad_o[29] ;
output \mc_data_pad_o[2] ;
output \mc_data_pad_o[30] ;
output \mc_data_pad_o[31] ;
output \mc_data_pad_o[3] ;
output \mc_data_pad_o[4] ;
output \mc_data_pad_o[5] ;
output \mc_data_pad_o[6] ;
output \mc_data_pad_o[7] ;
output \mc_data_pad_o[8] ;
output \mc_data_pad_o[9] ;
output mc_doe_pad_doe_o;
wire mc_dp_od_0_; 
wire mc_dp_od_1_; 
wire mc_dp_od_2_; 
wire mc_dp_od_3_; 
input \mc_dp_pad_i[0] ;
input \mc_dp_pad_i[1] ;
input \mc_dp_pad_i[2] ;
input \mc_dp_pad_i[3] ;
output \mc_dp_pad_o[0] ;
output \mc_dp_pad_o[1] ;
output \mc_dp_pad_o[2] ;
output \mc_dp_pad_o[3] ;
output \mc_dqm_pad_o[0] ;
output \mc_dqm_pad_o[1] ;
output \mc_dqm_pad_o[2] ;
output \mc_dqm_pad_o[3] ;
output mc_oe_pad_o_;
output mc_ras_pad_o_;
output mc_rp_pad_o_;
wire mc_sts_ir; 
input mc_sts_pad_i;
output mc_vpen_pad_o;
output mc_we_pad_o_;
output mc_zz_pad_o;
wire mem_ack; 
wire mem_ack_r; 
wire mem_dout_0_; 
wire mem_dout_10_; 
wire mem_dout_11_; 
wire mem_dout_12_; 
wire mem_dout_13_; 
wire mem_dout_14_; 
wire mem_dout_15_; 
wire mem_dout_16_; 
wire mem_dout_17_; 
wire mem_dout_18_; 
wire mem_dout_19_; 
wire mem_dout_1_; 
wire mem_dout_20_; 
wire mem_dout_21_; 
wire mem_dout_22_; 
wire mem_dout_23_; 
wire mem_dout_24_; 
wire mem_dout_25_; 
wire mem_dout_26_; 
wire mem_dout_27_; 
wire mem_dout_28_; 
wire mem_dout_29_; 
wire mem_dout_2_; 
wire mem_dout_30_; 
wire mem_dout_31_; 
wire mem_dout_3_; 
wire mem_dout_4_; 
wire mem_dout_5_; 
wire mem_dout_6_; 
wire mem_dout_7_; 
wire mem_dout_8_; 
wire mem_dout_9_; 
wire next_adr; 
wire not_mem_cyc; 
wire obct_cs_0_; 
wire obct_cs_1_; 
wire obct_cs_2_; 
wire obct_cs_3_; 
wire obct_cs_4_; 
wire obct_cs_5_; 
wire obct_cs_6_; 
wire obct_cs_7_; 
wire oe_; 
wire pack_le0; 
wire pack_le1; 
wire pack_le2; 
wire page_size_10_; 
wire page_size_8_; 
wire page_size_9_; 
wire par_err; 
output \poc_o[0] ;
output \poc_o[10] ;
output \poc_o[11] ;
output \poc_o[12] ;
output \poc_o[13] ;
output \poc_o[14] ;
output \poc_o[15] ;
output \poc_o[16] ;
output \poc_o[17] ;
output \poc_o[18] ;
output \poc_o[19] ;
output \poc_o[1] ;
output \poc_o[20] ;
output \poc_o[21] ;
output \poc_o[22] ;
output \poc_o[23] ;
output \poc_o[24] ;
output \poc_o[25] ;
output \poc_o[26] ;
output \poc_o[27] ;
output \poc_o[28] ;
output \poc_o[29] ;
output \poc_o[2] ;
output \poc_o[30] ;
output \poc_o[31] ;
output \poc_o[3] ;
output \poc_o[4] ;
output \poc_o[5] ;
output \poc_o[6] ;
output \poc_o[7] ;
output \poc_o[8] ;
output \poc_o[9] ;
wire ras_; 
wire ref_int_0_; 
wire ref_int_1_; 
wire ref_int_2_; 
input resume_req_i;
wire rf_dout_0_; 
wire rf_dout_10_; 
wire rf_dout_11_; 
wire rf_dout_12_; 
wire rf_dout_13_; 
wire rf_dout_14_; 
wire rf_dout_15_; 
wire rf_dout_16_; 
wire rf_dout_17_; 
wire rf_dout_18_; 
wire rf_dout_19_; 
wire rf_dout_1_; 
wire rf_dout_20_; 
wire rf_dout_21_; 
wire rf_dout_22_; 
wire rf_dout_23_; 
wire rf_dout_24_; 
wire rf_dout_25_; 
wire rf_dout_26_; 
wire rf_dout_27_; 
wire rf_dout_28_; 
wire rf_dout_29_; 
wire rf_dout_2_; 
wire rf_dout_30_; 
wire rf_dout_31_; 
wire rf_dout_3_; 
wire rf_dout_4_; 
wire rf_dout_5_; 
wire rf_dout_6_; 
wire rf_dout_7_; 
wire rf_dout_8_; 
wire rf_dout_9_; 
wire rfr_ack; 
wire rfr_ps_val_0_; 
wire rfr_ps_val_1_; 
wire rfr_ps_val_2_; 
wire rfr_ps_val_3_; 
wire rfr_ps_val_4_; 
wire rfr_ps_val_5_; 
wire rfr_ps_val_6_; 
wire rfr_ps_val_7_; 
wire rfr_req; 
wire row_adr_0_; 
wire row_adr_10_; 
wire row_adr_11_; 
wire row_adr_12_; 
wire row_adr_1_; 
wire row_adr_2_; 
wire row_adr_3_; 
wire row_adr_4_; 
wire row_adr_5_; 
wire row_adr_6_; 
wire row_adr_7_; 
wire row_adr_8_; 
wire row_adr_9_; 
wire row_same; 
wire row_sel; 
input rst_i;
wire sp_csc_10_; 
wire sp_csc_1_; 
wire sp_csc_2_; 
wire sp_csc_3_; 
wire sp_csc_4_; 
wire sp_csc_5_; 
wire sp_csc_6_; 
wire sp_csc_7_; 
wire sp_csc_9_; 
wire sp_tms_0_; 
wire sp_tms_10_; 
wire sp_tms_11_; 
wire sp_tms_12_; 
wire sp_tms_13_; 
wire sp_tms_14_; 
wire sp_tms_15_; 
wire sp_tms_16_; 
wire sp_tms_17_; 
wire sp_tms_18_; 
wire sp_tms_19_; 
wire sp_tms_1_; 
wire sp_tms_20_; 
wire sp_tms_21_; 
wire sp_tms_22_; 
wire sp_tms_23_; 
wire sp_tms_24_; 
wire sp_tms_25_; 
wire sp_tms_26_; 
wire sp_tms_27_; 
wire sp_tms_2_; 
wire sp_tms_3_; 
wire sp_tms_4_; 
wire sp_tms_5_; 
wire sp_tms_6_; 
wire sp_tms_7_; 
wire sp_tms_8_; 
wire sp_tms_9_; 
wire spec_req_cs_0_; 
wire spec_req_cs_1_; 
wire spec_req_cs_2_; 
wire spec_req_cs_3_; 
wire spec_req_cs_4_; 
wire spec_req_cs_5_; 
wire spec_req_cs_6_; 
wire spec_req_cs_7_; 
input susp_req_i;
wire susp_sel; 
output suspended_o;
wire tms_0_; 
wire tms_10_; 
wire tms_11_; 
wire tms_12_; 
wire tms_13_; 
wire tms_14_; 
wire tms_15_; 
wire tms_16_; 
wire tms_17_; 
wire tms_18_; 
wire tms_19_; 
wire tms_1_; 
wire tms_20_; 
wire tms_21_; 
wire tms_22_; 
wire tms_23_; 
wire tms_24_; 
wire tms_25_; 
wire tms_26_; 
wire tms_27_; 
wire tms_2_; 
wire tms_3_; 
wire tms_4_; 
wire tms_5_; 
wire tms_6_; 
wire tms_7_; 
wire tms_8_; 
wire tms_9_; 
wire tms_s_0_; 
wire tms_s_10_; 
wire tms_s_11_; 
wire tms_s_12_; 
wire tms_s_13_; 
wire tms_s_14_; 
wire tms_s_15_; 
wire tms_s_16_; 
wire tms_s_17_; 
wire tms_s_18_; 
wire tms_s_19_; 
wire tms_s_1_; 
wire tms_s_20_; 
wire tms_s_21_; 
wire tms_s_22_; 
wire tms_s_23_; 
wire tms_s_24_; 
wire tms_s_25_; 
wire tms_s_26_; 
wire tms_s_27_; 
wire tms_s_2_; 
wire tms_s_3_; 
wire tms_s_4_; 
wire tms_s_5_; 
wire tms_s_6_; 
wire tms_s_7_; 
wire tms_s_8_; 
wire tms_s_9_; 
wire u0__0cs_7_0__0_; 
wire u0__0cs_7_0__1_; 
wire u0__0cs_7_0__2_; 
wire u0__0cs_7_0__3_; 
wire u0__0cs_7_0__4_; 
wire u0__0cs_7_0__5_; 
wire u0__0cs_7_0__6_; 
wire u0__0cs_7_0__7_; 
wire u0__0csc_31_0__10_; 
wire u0__0csc_31_0__11_; 
wire u0__0csc_31_0__1_; 
wire u0__0csc_31_0__2_; 
wire u0__0csc_31_0__3_; 
wire u0__0csc_31_0__4_; 
wire u0__0csc_31_0__5_; 
wire u0__0csc_31_0__6_; 
wire u0__0csc_31_0__7_; 
wire u0__0csc_31_0__9_; 
wire u0__0csc_mask_r_10_0__0_; 
wire u0__0csc_mask_r_10_0__10_; 
wire u0__0csc_mask_r_10_0__1_; 
wire u0__0csc_mask_r_10_0__2_; 
wire u0__0csc_mask_r_10_0__3_; 
wire u0__0csc_mask_r_10_0__4_; 
wire u0__0csc_mask_r_10_0__5_; 
wire u0__0csc_mask_r_10_0__6_; 
wire u0__0csc_mask_r_10_0__7_; 
wire u0__0csc_mask_r_10_0__8_; 
wire u0__0csc_mask_r_10_0__9_; 
wire u0__0csr_r2_7_0__0_; 
wire u0__0csr_r2_7_0__1_; 
wire u0__0csr_r2_7_0__2_; 
wire u0__0csr_r2_7_0__3_; 
wire u0__0csr_r2_7_0__4_; 
wire u0__0csr_r2_7_0__5_; 
wire u0__0csr_r2_7_0__6_; 
wire u0__0csr_r2_7_0__7_; 
wire u0__0csr_r_10_1__0_; 
wire u0__0csr_r_10_1__1_; 
wire u0__0csr_r_10_1__2_; 
wire u0__0csr_r_10_1__3_; 
wire u0__0csr_r_10_1__4_; 
wire u0__0csr_r_10_1__5_; 
wire u0__0csr_r_10_1__6_; 
wire u0__0csr_r_10_1__7_; 
wire u0__0csr_r_10_1__8_; 
wire u0__0csr_r_10_1__9_; 
wire u0__0init_req_0_0_; 
wire u0__0lmr_req_0_0_; 
wire u0__0poc_31_0__0_; 
wire u0__0poc_31_0__10_; 
wire u0__0poc_31_0__11_; 
wire u0__0poc_31_0__12_; 
wire u0__0poc_31_0__13_; 
wire u0__0poc_31_0__14_; 
wire u0__0poc_31_0__15_; 
wire u0__0poc_31_0__16_; 
wire u0__0poc_31_0__17_; 
wire u0__0poc_31_0__18_; 
wire u0__0poc_31_0__19_; 
wire u0__0poc_31_0__1_; 
wire u0__0poc_31_0__20_; 
wire u0__0poc_31_0__21_; 
wire u0__0poc_31_0__22_; 
wire u0__0poc_31_0__23_; 
wire u0__0poc_31_0__24_; 
wire u0__0poc_31_0__25_; 
wire u0__0poc_31_0__26_; 
wire u0__0poc_31_0__27_; 
wire u0__0poc_31_0__28_; 
wire u0__0poc_31_0__29_; 
wire u0__0poc_31_0__2_; 
wire u0__0poc_31_0__30_; 
wire u0__0poc_31_0__31_; 
wire u0__0poc_31_0__3_; 
wire u0__0poc_31_0__4_; 
wire u0__0poc_31_0__5_; 
wire u0__0poc_31_0__6_; 
wire u0__0poc_31_0__7_; 
wire u0__0poc_31_0__8_; 
wire u0__0poc_31_0__9_; 
wire u0__0rf_we_0_0_; 
wire u0__0sp_csc_31_0__10_; 
wire u0__0sp_csc_31_0__1_; 
wire u0__0sp_csc_31_0__2_; 
wire u0__0sp_csc_31_0__3_; 
wire u0__0sp_csc_31_0__4_; 
wire u0__0sp_csc_31_0__5_; 
wire u0__0sp_csc_31_0__6_; 
wire u0__0sp_csc_31_0__7_; 
wire u0__0sp_csc_31_0__9_; 
wire u0__0sp_tms_31_0__0_; 
wire u0__0sp_tms_31_0__10_; 
wire u0__0sp_tms_31_0__11_; 
wire u0__0sp_tms_31_0__12_; 
wire u0__0sp_tms_31_0__13_; 
wire u0__0sp_tms_31_0__14_; 
wire u0__0sp_tms_31_0__15_; 
wire u0__0sp_tms_31_0__16_; 
wire u0__0sp_tms_31_0__17_; 
wire u0__0sp_tms_31_0__18_; 
wire u0__0sp_tms_31_0__19_; 
wire u0__0sp_tms_31_0__1_; 
wire u0__0sp_tms_31_0__20_; 
wire u0__0sp_tms_31_0__21_; 
wire u0__0sp_tms_31_0__22_; 
wire u0__0sp_tms_31_0__23_; 
wire u0__0sp_tms_31_0__24_; 
wire u0__0sp_tms_31_0__25_; 
wire u0__0sp_tms_31_0__26_; 
wire u0__0sp_tms_31_0__27_; 
wire u0__0sp_tms_31_0__2_; 
wire u0__0sp_tms_31_0__3_; 
wire u0__0sp_tms_31_0__4_; 
wire u0__0sp_tms_31_0__5_; 
wire u0__0sp_tms_31_0__6_; 
wire u0__0sp_tms_31_0__7_; 
wire u0__0sp_tms_31_0__8_; 
wire u0__0sp_tms_31_0__9_; 
wire u0__0spec_req_cs_7_0__0_; 
wire u0__0spec_req_cs_7_0__1_; 
wire u0__0spec_req_cs_7_0__2_; 
wire u0__0spec_req_cs_7_0__3_; 
wire u0__0spec_req_cs_7_0__4_; 
wire u0__0spec_req_cs_7_0__5_; 
wire u0__0spec_req_cs_7_0__6_; 
wire u0__0spec_req_cs_7_0__7_; 
wire u0__0sreq_cs_le_0_0_; 
wire u0__0tms_31_0__0_; 
wire u0__0tms_31_0__10_; 
wire u0__0tms_31_0__11_; 
wire u0__0tms_31_0__12_; 
wire u0__0tms_31_0__13_; 
wire u0__0tms_31_0__14_; 
wire u0__0tms_31_0__15_; 
wire u0__0tms_31_0__16_; 
wire u0__0tms_31_0__17_; 
wire u0__0tms_31_0__18_; 
wire u0__0tms_31_0__19_; 
wire u0__0tms_31_0__1_; 
wire u0__0tms_31_0__20_; 
wire u0__0tms_31_0__21_; 
wire u0__0tms_31_0__22_; 
wire u0__0tms_31_0__23_; 
wire u0__0tms_31_0__24_; 
wire u0__0tms_31_0__25_; 
wire u0__0tms_31_0__26_; 
wire u0__0tms_31_0__27_; 
wire u0__0tms_31_0__2_; 
wire u0__0tms_31_0__3_; 
wire u0__0tms_31_0__4_; 
wire u0__0tms_31_0__5_; 
wire u0__0tms_31_0__6_; 
wire u0__0tms_31_0__7_; 
wire u0__0tms_31_0__8_; 
wire u0__0tms_31_0__9_; 
wire u0__0wp_err_0_0_; 
wire u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602; 
wire u0__abc_74894_new_n1100_; 
wire u0__abc_74894_new_n1101_; 
wire u0__abc_74894_new_n1102_; 
wire u0__abc_74894_new_n1103_; 
wire u0__abc_74894_new_n1104_; 
wire u0__abc_74894_new_n1106_; 
wire u0__abc_74894_new_n1107_; 
wire u0__abc_74894_new_n1108_; 
wire u0__abc_74894_new_n1109_; 
wire u0__abc_74894_new_n1110_; 
wire u0__abc_74894_new_n1112_; 
wire u0__abc_74894_new_n1113_; 
wire u0__abc_74894_new_n1114_; 
wire u0__abc_74894_new_n1115_; 
wire u0__abc_74894_new_n1116_; 
wire u0__abc_74894_new_n1117_; 
wire u0__abc_74894_new_n1119_; 
wire u0__abc_74894_new_n1120_; 
wire u0__abc_74894_new_n1121_; 
wire u0__abc_74894_new_n1122_; 
wire u0__abc_74894_new_n1123_; 
wire u0__abc_74894_new_n1125_; 
wire u0__abc_74894_new_n1126_; 
wire u0__abc_74894_new_n1127_; 
wire u0__abc_74894_new_n1128_; 
wire u0__abc_74894_new_n1129_; 
wire u0__abc_74894_new_n1130_; 
wire u0__abc_74894_new_n1131_; 
wire u0__abc_74894_new_n1132_; 
wire u0__abc_74894_new_n1134_; 
wire u0__abc_74894_new_n1135_; 
wire u0__abc_74894_new_n1136_; 
wire u0__abc_74894_new_n1137_; 
wire u0__abc_74894_new_n1138_; 
wire u0__abc_74894_new_n1140_; 
wire u0__abc_74894_new_n1141_; 
wire u0__abc_74894_new_n1142_; 
wire u0__abc_74894_new_n1143_; 
wire u0__abc_74894_new_n1144_; 
wire u0__abc_74894_new_n1145_; 
wire u0__abc_74894_new_n1147_; 
wire u0__abc_74894_new_n1148_; 
wire u0__abc_74894_new_n1149_; 
wire u0__abc_74894_new_n1150_; 
wire u0__abc_74894_new_n1151_; 
wire u0__abc_74894_new_n1152_; 
wire u0__abc_74894_new_n1154_; 
wire u0__abc_74894_new_n1155_; 
wire u0__abc_74894_new_n1156_; 
wire u0__abc_74894_new_n1157_; 
wire u0__abc_74894_new_n1158_; 
wire u0__abc_74894_new_n1159_; 
wire u0__abc_74894_new_n1160_; 
wire u0__abc_74894_new_n1161_; 
wire u0__abc_74894_new_n1162_; 
wire u0__abc_74894_new_n1163_; 
wire u0__abc_74894_new_n1164_; 
wire u0__abc_74894_new_n1165_; 
wire u0__abc_74894_new_n1166_; 
wire u0__abc_74894_new_n1167_; 
wire u0__abc_74894_new_n1168_; 
wire u0__abc_74894_new_n1169_; 
wire u0__abc_74894_new_n1170_; 
wire u0__abc_74894_new_n1171_; 
wire u0__abc_74894_new_n1172_; 
wire u0__abc_74894_new_n1173_; 
wire u0__abc_74894_new_n1174_; 
wire u0__abc_74894_new_n1176_; 
wire u0__abc_74894_new_n1177_; 
wire u0__abc_74894_new_n1178_; 
wire u0__abc_74894_new_n1179_; 
wire u0__abc_74894_new_n1180_; 
wire u0__abc_74894_new_n1181_; 
wire u0__abc_74894_new_n1182_; 
wire u0__abc_74894_new_n1183_; 
wire u0__abc_74894_new_n1184_; 
wire u0__abc_74894_new_n1185_; 
wire u0__abc_74894_new_n1186_; 
wire u0__abc_74894_new_n1187_; 
wire u0__abc_74894_new_n1188_; 
wire u0__abc_74894_new_n1189_; 
wire u0__abc_74894_new_n1190_; 
wire u0__abc_74894_new_n1191_; 
wire u0__abc_74894_new_n1192_; 
wire u0__abc_74894_new_n1193_; 
wire u0__abc_74894_new_n1194_; 
wire u0__abc_74894_new_n1196_; 
wire u0__abc_74894_new_n1197_; 
wire u0__abc_74894_new_n1198_; 
wire u0__abc_74894_new_n1199_; 
wire u0__abc_74894_new_n1200_; 
wire u0__abc_74894_new_n1201_; 
wire u0__abc_74894_new_n1202_; 
wire u0__abc_74894_new_n1203_; 
wire u0__abc_74894_new_n1204_; 
wire u0__abc_74894_new_n1205_; 
wire u0__abc_74894_new_n1206_; 
wire u0__abc_74894_new_n1207_; 
wire u0__abc_74894_new_n1208_; 
wire u0__abc_74894_new_n1209_; 
wire u0__abc_74894_new_n1210_; 
wire u0__abc_74894_new_n1211_; 
wire u0__abc_74894_new_n1212_; 
wire u0__abc_74894_new_n1213_; 
wire u0__abc_74894_new_n1214_; 
wire u0__abc_74894_new_n1216_; 
wire u0__abc_74894_new_n1217_; 
wire u0__abc_74894_new_n1218_; 
wire u0__abc_74894_new_n1219_; 
wire u0__abc_74894_new_n1220_; 
wire u0__abc_74894_new_n1221_; 
wire u0__abc_74894_new_n1222_; 
wire u0__abc_74894_new_n1223_; 
wire u0__abc_74894_new_n1224_; 
wire u0__abc_74894_new_n1225_; 
wire u0__abc_74894_new_n1226_; 
wire u0__abc_74894_new_n1227_; 
wire u0__abc_74894_new_n1228_; 
wire u0__abc_74894_new_n1229_; 
wire u0__abc_74894_new_n1230_; 
wire u0__abc_74894_new_n1231_; 
wire u0__abc_74894_new_n1232_; 
wire u0__abc_74894_new_n1233_; 
wire u0__abc_74894_new_n1234_; 
wire u0__abc_74894_new_n1236_; 
wire u0__abc_74894_new_n1237_; 
wire u0__abc_74894_new_n1238_; 
wire u0__abc_74894_new_n1239_; 
wire u0__abc_74894_new_n1240_; 
wire u0__abc_74894_new_n1241_; 
wire u0__abc_74894_new_n1242_; 
wire u0__abc_74894_new_n1243_; 
wire u0__abc_74894_new_n1244_; 
wire u0__abc_74894_new_n1245_; 
wire u0__abc_74894_new_n1246_; 
wire u0__abc_74894_new_n1247_; 
wire u0__abc_74894_new_n1248_; 
wire u0__abc_74894_new_n1249_; 
wire u0__abc_74894_new_n1250_; 
wire u0__abc_74894_new_n1251_; 
wire u0__abc_74894_new_n1252_; 
wire u0__abc_74894_new_n1253_; 
wire u0__abc_74894_new_n1254_; 
wire u0__abc_74894_new_n1256_; 
wire u0__abc_74894_new_n1257_; 
wire u0__abc_74894_new_n1258_; 
wire u0__abc_74894_new_n1259_; 
wire u0__abc_74894_new_n1260_; 
wire u0__abc_74894_new_n1261_; 
wire u0__abc_74894_new_n1262_; 
wire u0__abc_74894_new_n1263_; 
wire u0__abc_74894_new_n1264_; 
wire u0__abc_74894_new_n1265_; 
wire u0__abc_74894_new_n1266_; 
wire u0__abc_74894_new_n1267_; 
wire u0__abc_74894_new_n1268_; 
wire u0__abc_74894_new_n1269_; 
wire u0__abc_74894_new_n1270_; 
wire u0__abc_74894_new_n1271_; 
wire u0__abc_74894_new_n1272_; 
wire u0__abc_74894_new_n1273_; 
wire u0__abc_74894_new_n1274_; 
wire u0__abc_74894_new_n1276_; 
wire u0__abc_74894_new_n1277_; 
wire u0__abc_74894_new_n1278_; 
wire u0__abc_74894_new_n1279_; 
wire u0__abc_74894_new_n1280_; 
wire u0__abc_74894_new_n1281_; 
wire u0__abc_74894_new_n1282_; 
wire u0__abc_74894_new_n1283_; 
wire u0__abc_74894_new_n1284_; 
wire u0__abc_74894_new_n1285_; 
wire u0__abc_74894_new_n1286_; 
wire u0__abc_74894_new_n1287_; 
wire u0__abc_74894_new_n1288_; 
wire u0__abc_74894_new_n1289_; 
wire u0__abc_74894_new_n1290_; 
wire u0__abc_74894_new_n1291_; 
wire u0__abc_74894_new_n1292_; 
wire u0__abc_74894_new_n1293_; 
wire u0__abc_74894_new_n1294_; 
wire u0__abc_74894_new_n1296_; 
wire u0__abc_74894_new_n1297_; 
wire u0__abc_74894_new_n1298_; 
wire u0__abc_74894_new_n1299_; 
wire u0__abc_74894_new_n1300_; 
wire u0__abc_74894_new_n1301_; 
wire u0__abc_74894_new_n1302_; 
wire u0__abc_74894_new_n1303_; 
wire u0__abc_74894_new_n1304_; 
wire u0__abc_74894_new_n1305_; 
wire u0__abc_74894_new_n1306_; 
wire u0__abc_74894_new_n1307_; 
wire u0__abc_74894_new_n1308_; 
wire u0__abc_74894_new_n1309_; 
wire u0__abc_74894_new_n1310_; 
wire u0__abc_74894_new_n1311_; 
wire u0__abc_74894_new_n1312_; 
wire u0__abc_74894_new_n1313_; 
wire u0__abc_74894_new_n1314_; 
wire u0__abc_74894_new_n1316_; 
wire u0__abc_74894_new_n1317_; 
wire u0__abc_74894_new_n1318_; 
wire u0__abc_74894_new_n1319_; 
wire u0__abc_74894_new_n1320_; 
wire u0__abc_74894_new_n1321_; 
wire u0__abc_74894_new_n1322_; 
wire u0__abc_74894_new_n1323_; 
wire u0__abc_74894_new_n1324_; 
wire u0__abc_74894_new_n1325_; 
wire u0__abc_74894_new_n1326_; 
wire u0__abc_74894_new_n1327_; 
wire u0__abc_74894_new_n1328_; 
wire u0__abc_74894_new_n1329_; 
wire u0__abc_74894_new_n1330_; 
wire u0__abc_74894_new_n1331_; 
wire u0__abc_74894_new_n1332_; 
wire u0__abc_74894_new_n1333_; 
wire u0__abc_74894_new_n1334_; 
wire u0__abc_74894_new_n1336_; 
wire u0__abc_74894_new_n1337_; 
wire u0__abc_74894_new_n1338_; 
wire u0__abc_74894_new_n1339_; 
wire u0__abc_74894_new_n1340_; 
wire u0__abc_74894_new_n1341_; 
wire u0__abc_74894_new_n1342_; 
wire u0__abc_74894_new_n1343_; 
wire u0__abc_74894_new_n1344_; 
wire u0__abc_74894_new_n1345_; 
wire u0__abc_74894_new_n1346_; 
wire u0__abc_74894_new_n1347_; 
wire u0__abc_74894_new_n1348_; 
wire u0__abc_74894_new_n1349_; 
wire u0__abc_74894_new_n1350_; 
wire u0__abc_74894_new_n1351_; 
wire u0__abc_74894_new_n1352_; 
wire u0__abc_74894_new_n1353_; 
wire u0__abc_74894_new_n1354_; 
wire u0__abc_74894_new_n1356_; 
wire u0__abc_74894_new_n1357_; 
wire u0__abc_74894_new_n1358_; 
wire u0__abc_74894_new_n1359_; 
wire u0__abc_74894_new_n1360_; 
wire u0__abc_74894_new_n1361_; 
wire u0__abc_74894_new_n1362_; 
wire u0__abc_74894_new_n1363_; 
wire u0__abc_74894_new_n1364_; 
wire u0__abc_74894_new_n1365_; 
wire u0__abc_74894_new_n1366_; 
wire u0__abc_74894_new_n1367_; 
wire u0__abc_74894_new_n1368_; 
wire u0__abc_74894_new_n1369_; 
wire u0__abc_74894_new_n1370_; 
wire u0__abc_74894_new_n1371_; 
wire u0__abc_74894_new_n1372_; 
wire u0__abc_74894_new_n1373_; 
wire u0__abc_74894_new_n1374_; 
wire u0__abc_74894_new_n1376_; 
wire u0__abc_74894_new_n1377_; 
wire u0__abc_74894_new_n1378_; 
wire u0__abc_74894_new_n1379_; 
wire u0__abc_74894_new_n1380_; 
wire u0__abc_74894_new_n1381_; 
wire u0__abc_74894_new_n1382_; 
wire u0__abc_74894_new_n1383_; 
wire u0__abc_74894_new_n1384_; 
wire u0__abc_74894_new_n1385_; 
wire u0__abc_74894_new_n1386_; 
wire u0__abc_74894_new_n1387_; 
wire u0__abc_74894_new_n1388_; 
wire u0__abc_74894_new_n1389_; 
wire u0__abc_74894_new_n1390_; 
wire u0__abc_74894_new_n1391_; 
wire u0__abc_74894_new_n1392_; 
wire u0__abc_74894_new_n1393_; 
wire u0__abc_74894_new_n1394_; 
wire u0__abc_74894_new_n1396_; 
wire u0__abc_74894_new_n1397_; 
wire u0__abc_74894_new_n1398_; 
wire u0__abc_74894_new_n1399_; 
wire u0__abc_74894_new_n1400_; 
wire u0__abc_74894_new_n1401_; 
wire u0__abc_74894_new_n1402_; 
wire u0__abc_74894_new_n1403_; 
wire u0__abc_74894_new_n1404_; 
wire u0__abc_74894_new_n1405_; 
wire u0__abc_74894_new_n1406_; 
wire u0__abc_74894_new_n1407_; 
wire u0__abc_74894_new_n1408_; 
wire u0__abc_74894_new_n1409_; 
wire u0__abc_74894_new_n1410_; 
wire u0__abc_74894_new_n1411_; 
wire u0__abc_74894_new_n1412_; 
wire u0__abc_74894_new_n1413_; 
wire u0__abc_74894_new_n1414_; 
wire u0__abc_74894_new_n1416_; 
wire u0__abc_74894_new_n1417_; 
wire u0__abc_74894_new_n1418_; 
wire u0__abc_74894_new_n1419_; 
wire u0__abc_74894_new_n1420_; 
wire u0__abc_74894_new_n1421_; 
wire u0__abc_74894_new_n1422_; 
wire u0__abc_74894_new_n1423_; 
wire u0__abc_74894_new_n1424_; 
wire u0__abc_74894_new_n1425_; 
wire u0__abc_74894_new_n1426_; 
wire u0__abc_74894_new_n1427_; 
wire u0__abc_74894_new_n1428_; 
wire u0__abc_74894_new_n1429_; 
wire u0__abc_74894_new_n1430_; 
wire u0__abc_74894_new_n1431_; 
wire u0__abc_74894_new_n1432_; 
wire u0__abc_74894_new_n1433_; 
wire u0__abc_74894_new_n1434_; 
wire u0__abc_74894_new_n1436_; 
wire u0__abc_74894_new_n1437_; 
wire u0__abc_74894_new_n1438_; 
wire u0__abc_74894_new_n1439_; 
wire u0__abc_74894_new_n1440_; 
wire u0__abc_74894_new_n1441_; 
wire u0__abc_74894_new_n1442_; 
wire u0__abc_74894_new_n1443_; 
wire u0__abc_74894_new_n1444_; 
wire u0__abc_74894_new_n1445_; 
wire u0__abc_74894_new_n1446_; 
wire u0__abc_74894_new_n1447_; 
wire u0__abc_74894_new_n1448_; 
wire u0__abc_74894_new_n1449_; 
wire u0__abc_74894_new_n1450_; 
wire u0__abc_74894_new_n1451_; 
wire u0__abc_74894_new_n1452_; 
wire u0__abc_74894_new_n1453_; 
wire u0__abc_74894_new_n1454_; 
wire u0__abc_74894_new_n1456_; 
wire u0__abc_74894_new_n1457_; 
wire u0__abc_74894_new_n1458_; 
wire u0__abc_74894_new_n1459_; 
wire u0__abc_74894_new_n1460_; 
wire u0__abc_74894_new_n1461_; 
wire u0__abc_74894_new_n1462_; 
wire u0__abc_74894_new_n1463_; 
wire u0__abc_74894_new_n1464_; 
wire u0__abc_74894_new_n1465_; 
wire u0__abc_74894_new_n1466_; 
wire u0__abc_74894_new_n1467_; 
wire u0__abc_74894_new_n1468_; 
wire u0__abc_74894_new_n1469_; 
wire u0__abc_74894_new_n1470_; 
wire u0__abc_74894_new_n1471_; 
wire u0__abc_74894_new_n1472_; 
wire u0__abc_74894_new_n1473_; 
wire u0__abc_74894_new_n1474_; 
wire u0__abc_74894_new_n1476_; 
wire u0__abc_74894_new_n1477_; 
wire u0__abc_74894_new_n1478_; 
wire u0__abc_74894_new_n1479_; 
wire u0__abc_74894_new_n1480_; 
wire u0__abc_74894_new_n1481_; 
wire u0__abc_74894_new_n1482_; 
wire u0__abc_74894_new_n1483_; 
wire u0__abc_74894_new_n1484_; 
wire u0__abc_74894_new_n1485_; 
wire u0__abc_74894_new_n1486_; 
wire u0__abc_74894_new_n1487_; 
wire u0__abc_74894_new_n1488_; 
wire u0__abc_74894_new_n1489_; 
wire u0__abc_74894_new_n1490_; 
wire u0__abc_74894_new_n1491_; 
wire u0__abc_74894_new_n1492_; 
wire u0__abc_74894_new_n1493_; 
wire u0__abc_74894_new_n1494_; 
wire u0__abc_74894_new_n1496_; 
wire u0__abc_74894_new_n1497_; 
wire u0__abc_74894_new_n1498_; 
wire u0__abc_74894_new_n1499_; 
wire u0__abc_74894_new_n1500_; 
wire u0__abc_74894_new_n1501_; 
wire u0__abc_74894_new_n1502_; 
wire u0__abc_74894_new_n1503_; 
wire u0__abc_74894_new_n1504_; 
wire u0__abc_74894_new_n1505_; 
wire u0__abc_74894_new_n1506_; 
wire u0__abc_74894_new_n1507_; 
wire u0__abc_74894_new_n1508_; 
wire u0__abc_74894_new_n1509_; 
wire u0__abc_74894_new_n1510_; 
wire u0__abc_74894_new_n1511_; 
wire u0__abc_74894_new_n1512_; 
wire u0__abc_74894_new_n1513_; 
wire u0__abc_74894_new_n1514_; 
wire u0__abc_74894_new_n1516_; 
wire u0__abc_74894_new_n1517_; 
wire u0__abc_74894_new_n1518_; 
wire u0__abc_74894_new_n1519_; 
wire u0__abc_74894_new_n1520_; 
wire u0__abc_74894_new_n1521_; 
wire u0__abc_74894_new_n1522_; 
wire u0__abc_74894_new_n1523_; 
wire u0__abc_74894_new_n1524_; 
wire u0__abc_74894_new_n1525_; 
wire u0__abc_74894_new_n1526_; 
wire u0__abc_74894_new_n1527_; 
wire u0__abc_74894_new_n1528_; 
wire u0__abc_74894_new_n1529_; 
wire u0__abc_74894_new_n1530_; 
wire u0__abc_74894_new_n1531_; 
wire u0__abc_74894_new_n1532_; 
wire u0__abc_74894_new_n1533_; 
wire u0__abc_74894_new_n1534_; 
wire u0__abc_74894_new_n1536_; 
wire u0__abc_74894_new_n1537_; 
wire u0__abc_74894_new_n1538_; 
wire u0__abc_74894_new_n1539_; 
wire u0__abc_74894_new_n1540_; 
wire u0__abc_74894_new_n1541_; 
wire u0__abc_74894_new_n1542_; 
wire u0__abc_74894_new_n1543_; 
wire u0__abc_74894_new_n1544_; 
wire u0__abc_74894_new_n1545_; 
wire u0__abc_74894_new_n1546_; 
wire u0__abc_74894_new_n1547_; 
wire u0__abc_74894_new_n1548_; 
wire u0__abc_74894_new_n1549_; 
wire u0__abc_74894_new_n1550_; 
wire u0__abc_74894_new_n1551_; 
wire u0__abc_74894_new_n1552_; 
wire u0__abc_74894_new_n1553_; 
wire u0__abc_74894_new_n1554_; 
wire u0__abc_74894_new_n1556_; 
wire u0__abc_74894_new_n1557_; 
wire u0__abc_74894_new_n1558_; 
wire u0__abc_74894_new_n1559_; 
wire u0__abc_74894_new_n1560_; 
wire u0__abc_74894_new_n1561_; 
wire u0__abc_74894_new_n1562_; 
wire u0__abc_74894_new_n1563_; 
wire u0__abc_74894_new_n1564_; 
wire u0__abc_74894_new_n1565_; 
wire u0__abc_74894_new_n1566_; 
wire u0__abc_74894_new_n1567_; 
wire u0__abc_74894_new_n1568_; 
wire u0__abc_74894_new_n1569_; 
wire u0__abc_74894_new_n1570_; 
wire u0__abc_74894_new_n1571_; 
wire u0__abc_74894_new_n1572_; 
wire u0__abc_74894_new_n1573_; 
wire u0__abc_74894_new_n1574_; 
wire u0__abc_74894_new_n1576_; 
wire u0__abc_74894_new_n1577_; 
wire u0__abc_74894_new_n1578_; 
wire u0__abc_74894_new_n1579_; 
wire u0__abc_74894_new_n1580_; 
wire u0__abc_74894_new_n1581_; 
wire u0__abc_74894_new_n1582_; 
wire u0__abc_74894_new_n1583_; 
wire u0__abc_74894_new_n1584_; 
wire u0__abc_74894_new_n1585_; 
wire u0__abc_74894_new_n1586_; 
wire u0__abc_74894_new_n1587_; 
wire u0__abc_74894_new_n1588_; 
wire u0__abc_74894_new_n1589_; 
wire u0__abc_74894_new_n1590_; 
wire u0__abc_74894_new_n1591_; 
wire u0__abc_74894_new_n1592_; 
wire u0__abc_74894_new_n1593_; 
wire u0__abc_74894_new_n1594_; 
wire u0__abc_74894_new_n1596_; 
wire u0__abc_74894_new_n1597_; 
wire u0__abc_74894_new_n1598_; 
wire u0__abc_74894_new_n1599_; 
wire u0__abc_74894_new_n1600_; 
wire u0__abc_74894_new_n1601_; 
wire u0__abc_74894_new_n1602_; 
wire u0__abc_74894_new_n1603_; 
wire u0__abc_74894_new_n1604_; 
wire u0__abc_74894_new_n1605_; 
wire u0__abc_74894_new_n1606_; 
wire u0__abc_74894_new_n1607_; 
wire u0__abc_74894_new_n1608_; 
wire u0__abc_74894_new_n1609_; 
wire u0__abc_74894_new_n1610_; 
wire u0__abc_74894_new_n1611_; 
wire u0__abc_74894_new_n1612_; 
wire u0__abc_74894_new_n1613_; 
wire u0__abc_74894_new_n1614_; 
wire u0__abc_74894_new_n1616_; 
wire u0__abc_74894_new_n1617_; 
wire u0__abc_74894_new_n1618_; 
wire u0__abc_74894_new_n1619_; 
wire u0__abc_74894_new_n1620_; 
wire u0__abc_74894_new_n1621_; 
wire u0__abc_74894_new_n1622_; 
wire u0__abc_74894_new_n1623_; 
wire u0__abc_74894_new_n1624_; 
wire u0__abc_74894_new_n1625_; 
wire u0__abc_74894_new_n1626_; 
wire u0__abc_74894_new_n1627_; 
wire u0__abc_74894_new_n1628_; 
wire u0__abc_74894_new_n1629_; 
wire u0__abc_74894_new_n1630_; 
wire u0__abc_74894_new_n1631_; 
wire u0__abc_74894_new_n1632_; 
wire u0__abc_74894_new_n1633_; 
wire u0__abc_74894_new_n1634_; 
wire u0__abc_74894_new_n1636_; 
wire u0__abc_74894_new_n1637_; 
wire u0__abc_74894_new_n1638_; 
wire u0__abc_74894_new_n1639_; 
wire u0__abc_74894_new_n1640_; 
wire u0__abc_74894_new_n1641_; 
wire u0__abc_74894_new_n1642_; 
wire u0__abc_74894_new_n1643_; 
wire u0__abc_74894_new_n1644_; 
wire u0__abc_74894_new_n1645_; 
wire u0__abc_74894_new_n1646_; 
wire u0__abc_74894_new_n1647_; 
wire u0__abc_74894_new_n1648_; 
wire u0__abc_74894_new_n1649_; 
wire u0__abc_74894_new_n1650_; 
wire u0__abc_74894_new_n1651_; 
wire u0__abc_74894_new_n1652_; 
wire u0__abc_74894_new_n1653_; 
wire u0__abc_74894_new_n1654_; 
wire u0__abc_74894_new_n1656_; 
wire u0__abc_74894_new_n1657_; 
wire u0__abc_74894_new_n1658_; 
wire u0__abc_74894_new_n1659_; 
wire u0__abc_74894_new_n1660_; 
wire u0__abc_74894_new_n1661_; 
wire u0__abc_74894_new_n1662_; 
wire u0__abc_74894_new_n1663_; 
wire u0__abc_74894_new_n1664_; 
wire u0__abc_74894_new_n1665_; 
wire u0__abc_74894_new_n1666_; 
wire u0__abc_74894_new_n1667_; 
wire u0__abc_74894_new_n1668_; 
wire u0__abc_74894_new_n1669_; 
wire u0__abc_74894_new_n1670_; 
wire u0__abc_74894_new_n1671_; 
wire u0__abc_74894_new_n1672_; 
wire u0__abc_74894_new_n1673_; 
wire u0__abc_74894_new_n1674_; 
wire u0__abc_74894_new_n1676_; 
wire u0__abc_74894_new_n1677_; 
wire u0__abc_74894_new_n1678_; 
wire u0__abc_74894_new_n1679_; 
wire u0__abc_74894_new_n1680_; 
wire u0__abc_74894_new_n1681_; 
wire u0__abc_74894_new_n1682_; 
wire u0__abc_74894_new_n1683_; 
wire u0__abc_74894_new_n1684_; 
wire u0__abc_74894_new_n1685_; 
wire u0__abc_74894_new_n1686_; 
wire u0__abc_74894_new_n1687_; 
wire u0__abc_74894_new_n1688_; 
wire u0__abc_74894_new_n1689_; 
wire u0__abc_74894_new_n1690_; 
wire u0__abc_74894_new_n1691_; 
wire u0__abc_74894_new_n1692_; 
wire u0__abc_74894_new_n1693_; 
wire u0__abc_74894_new_n1694_; 
wire u0__abc_74894_new_n1696_; 
wire u0__abc_74894_new_n1697_; 
wire u0__abc_74894_new_n1698_; 
wire u0__abc_74894_new_n1699_; 
wire u0__abc_74894_new_n1700_; 
wire u0__abc_74894_new_n1701_; 
wire u0__abc_74894_new_n1702_; 
wire u0__abc_74894_new_n1703_; 
wire u0__abc_74894_new_n1704_; 
wire u0__abc_74894_new_n1705_; 
wire u0__abc_74894_new_n1706_; 
wire u0__abc_74894_new_n1707_; 
wire u0__abc_74894_new_n1708_; 
wire u0__abc_74894_new_n1709_; 
wire u0__abc_74894_new_n1710_; 
wire u0__abc_74894_new_n1711_; 
wire u0__abc_74894_new_n1712_; 
wire u0__abc_74894_new_n1713_; 
wire u0__abc_74894_new_n1714_; 
wire u0__abc_74894_new_n1717_; 
wire u0__abc_74894_new_n1737_; 
wire u0__abc_74894_new_n1757_; 
wire u0__abc_74894_new_n1796_; 
wire u0__abc_74894_new_n1811_; 
wire u0__abc_74894_new_n1817_; 
wire u0__abc_74894_new_n1818_; 
wire u0__abc_74894_new_n1819_; 
wire u0__abc_74894_new_n1820_; 
wire u0__abc_74894_new_n1821_; 
wire u0__abc_74894_new_n1822_; 
wire u0__abc_74894_new_n1823_; 
wire u0__abc_74894_new_n1824_; 
wire u0__abc_74894_new_n1825_; 
wire u0__abc_74894_new_n1826_; 
wire u0__abc_74894_new_n1827_; 
wire u0__abc_74894_new_n1828_; 
wire u0__abc_74894_new_n1829_; 
wire u0__abc_74894_new_n1830_; 
wire u0__abc_74894_new_n1831_; 
wire u0__abc_74894_new_n1832_; 
wire u0__abc_74894_new_n1833_; 
wire u0__abc_74894_new_n1834_; 
wire u0__abc_74894_new_n1835_; 
wire u0__abc_74894_new_n1837_; 
wire u0__abc_74894_new_n1838_; 
wire u0__abc_74894_new_n1839_; 
wire u0__abc_74894_new_n1840_; 
wire u0__abc_74894_new_n1841_; 
wire u0__abc_74894_new_n1842_; 
wire u0__abc_74894_new_n1843_; 
wire u0__abc_74894_new_n1844_; 
wire u0__abc_74894_new_n1845_; 
wire u0__abc_74894_new_n1846_; 
wire u0__abc_74894_new_n1847_; 
wire u0__abc_74894_new_n1848_; 
wire u0__abc_74894_new_n1849_; 
wire u0__abc_74894_new_n1850_; 
wire u0__abc_74894_new_n1851_; 
wire u0__abc_74894_new_n1852_; 
wire u0__abc_74894_new_n1853_; 
wire u0__abc_74894_new_n1854_; 
wire u0__abc_74894_new_n1855_; 
wire u0__abc_74894_new_n1857_; 
wire u0__abc_74894_new_n1858_; 
wire u0__abc_74894_new_n1859_; 
wire u0__abc_74894_new_n1860_; 
wire u0__abc_74894_new_n1861_; 
wire u0__abc_74894_new_n1862_; 
wire u0__abc_74894_new_n1863_; 
wire u0__abc_74894_new_n1864_; 
wire u0__abc_74894_new_n1865_; 
wire u0__abc_74894_new_n1866_; 
wire u0__abc_74894_new_n1867_; 
wire u0__abc_74894_new_n1868_; 
wire u0__abc_74894_new_n1869_; 
wire u0__abc_74894_new_n1870_; 
wire u0__abc_74894_new_n1871_; 
wire u0__abc_74894_new_n1872_; 
wire u0__abc_74894_new_n1873_; 
wire u0__abc_74894_new_n1874_; 
wire u0__abc_74894_new_n1875_; 
wire u0__abc_74894_new_n1877_; 
wire u0__abc_74894_new_n1878_; 
wire u0__abc_74894_new_n1879_; 
wire u0__abc_74894_new_n1880_; 
wire u0__abc_74894_new_n1881_; 
wire u0__abc_74894_new_n1882_; 
wire u0__abc_74894_new_n1883_; 
wire u0__abc_74894_new_n1884_; 
wire u0__abc_74894_new_n1885_; 
wire u0__abc_74894_new_n1886_; 
wire u0__abc_74894_new_n1887_; 
wire u0__abc_74894_new_n1888_; 
wire u0__abc_74894_new_n1889_; 
wire u0__abc_74894_new_n1890_; 
wire u0__abc_74894_new_n1891_; 
wire u0__abc_74894_new_n1892_; 
wire u0__abc_74894_new_n1893_; 
wire u0__abc_74894_new_n1894_; 
wire u0__abc_74894_new_n1895_; 
wire u0__abc_74894_new_n1897_; 
wire u0__abc_74894_new_n1898_; 
wire u0__abc_74894_new_n1899_; 
wire u0__abc_74894_new_n1900_; 
wire u0__abc_74894_new_n1901_; 
wire u0__abc_74894_new_n1902_; 
wire u0__abc_74894_new_n1903_; 
wire u0__abc_74894_new_n1904_; 
wire u0__abc_74894_new_n1905_; 
wire u0__abc_74894_new_n1906_; 
wire u0__abc_74894_new_n1907_; 
wire u0__abc_74894_new_n1908_; 
wire u0__abc_74894_new_n1909_; 
wire u0__abc_74894_new_n1910_; 
wire u0__abc_74894_new_n1911_; 
wire u0__abc_74894_new_n1912_; 
wire u0__abc_74894_new_n1913_; 
wire u0__abc_74894_new_n1914_; 
wire u0__abc_74894_new_n1915_; 
wire u0__abc_74894_new_n1917_; 
wire u0__abc_74894_new_n1918_; 
wire u0__abc_74894_new_n1919_; 
wire u0__abc_74894_new_n1920_; 
wire u0__abc_74894_new_n1921_; 
wire u0__abc_74894_new_n1922_; 
wire u0__abc_74894_new_n1923_; 
wire u0__abc_74894_new_n1924_; 
wire u0__abc_74894_new_n1925_; 
wire u0__abc_74894_new_n1926_; 
wire u0__abc_74894_new_n1927_; 
wire u0__abc_74894_new_n1928_; 
wire u0__abc_74894_new_n1929_; 
wire u0__abc_74894_new_n1930_; 
wire u0__abc_74894_new_n1931_; 
wire u0__abc_74894_new_n1932_; 
wire u0__abc_74894_new_n1933_; 
wire u0__abc_74894_new_n1934_; 
wire u0__abc_74894_new_n1935_; 
wire u0__abc_74894_new_n1937_; 
wire u0__abc_74894_new_n1938_; 
wire u0__abc_74894_new_n1939_; 
wire u0__abc_74894_new_n1940_; 
wire u0__abc_74894_new_n1941_; 
wire u0__abc_74894_new_n1942_; 
wire u0__abc_74894_new_n1943_; 
wire u0__abc_74894_new_n1944_; 
wire u0__abc_74894_new_n1945_; 
wire u0__abc_74894_new_n1946_; 
wire u0__abc_74894_new_n1947_; 
wire u0__abc_74894_new_n1948_; 
wire u0__abc_74894_new_n1949_; 
wire u0__abc_74894_new_n1950_; 
wire u0__abc_74894_new_n1951_; 
wire u0__abc_74894_new_n1952_; 
wire u0__abc_74894_new_n1953_; 
wire u0__abc_74894_new_n1954_; 
wire u0__abc_74894_new_n1955_; 
wire u0__abc_74894_new_n1958_; 
wire u0__abc_74894_new_n1973_; 
wire u0__abc_74894_new_n1977_; 
wire u0__abc_74894_new_n1978_; 
wire u0__abc_74894_new_n1979_; 
wire u0__abc_74894_new_n1980_; 
wire u0__abc_74894_new_n1981_; 
wire u0__abc_74894_new_n1982_; 
wire u0__abc_74894_new_n1983_; 
wire u0__abc_74894_new_n1984_; 
wire u0__abc_74894_new_n1985_; 
wire u0__abc_74894_new_n1986_; 
wire u0__abc_74894_new_n1987_; 
wire u0__abc_74894_new_n1988_; 
wire u0__abc_74894_new_n1989_; 
wire u0__abc_74894_new_n1990_; 
wire u0__abc_74894_new_n1991_; 
wire u0__abc_74894_new_n1992_; 
wire u0__abc_74894_new_n1993_; 
wire u0__abc_74894_new_n1994_; 
wire u0__abc_74894_new_n1995_; 
wire u0__abc_74894_new_n1997_; 
wire u0__abc_74894_new_n1998_; 
wire u0__abc_74894_new_n1999_; 
wire u0__abc_74894_new_n2000_; 
wire u0__abc_74894_new_n2001_; 
wire u0__abc_74894_new_n2002_; 
wire u0__abc_74894_new_n2003_; 
wire u0__abc_74894_new_n2004_; 
wire u0__abc_74894_new_n2005_; 
wire u0__abc_74894_new_n2006_; 
wire u0__abc_74894_new_n2007_; 
wire u0__abc_74894_new_n2008_; 
wire u0__abc_74894_new_n2009_; 
wire u0__abc_74894_new_n2010_; 
wire u0__abc_74894_new_n2011_; 
wire u0__abc_74894_new_n2012_; 
wire u0__abc_74894_new_n2013_; 
wire u0__abc_74894_new_n2014_; 
wire u0__abc_74894_new_n2015_; 
wire u0__abc_74894_new_n2018_; 
wire u0__abc_74894_new_n2020_; 
wire u0__abc_74894_new_n2031_; 
wire u0__abc_74894_new_n2058_; 
wire u0__abc_74894_new_n2073_; 
wire u0__abc_74894_new_n2078_; 
wire u0__abc_74894_new_n2111_; 
wire u0__abc_74894_new_n2133_; 
wire u0__abc_74894_new_n2151_; 
wire u0__abc_74894_new_n2171_; 
wire u0__abc_74894_new_n2178_; 
wire u0__abc_74894_new_n2193_; 
wire u0__abc_74894_new_n2218_; 
wire u0__abc_74894_new_n2273_; 
wire u0__abc_74894_new_n2437_; 
wire u0__abc_74894_new_n2438_; 
wire u0__abc_74894_new_n2439_; 
wire u0__abc_74894_new_n2440_; 
wire u0__abc_74894_new_n2441_; 
wire u0__abc_74894_new_n2442_; 
wire u0__abc_74894_new_n2443_; 
wire u0__abc_74894_new_n2444_; 
wire u0__abc_74894_new_n2445_; 
wire u0__abc_74894_new_n2446_; 
wire u0__abc_74894_new_n2447_; 
wire u0__abc_74894_new_n2448_; 
wire u0__abc_74894_new_n2449_; 
wire u0__abc_74894_new_n2450_; 
wire u0__abc_74894_new_n2451_; 
wire u0__abc_74894_new_n2452_; 
wire u0__abc_74894_new_n2453_; 
wire u0__abc_74894_new_n2454_; 
wire u0__abc_74894_new_n2455_; 
wire u0__abc_74894_new_n2456_; 
wire u0__abc_74894_new_n2457_; 
wire u0__abc_74894_new_n2458_; 
wire u0__abc_74894_new_n2460_; 
wire u0__abc_74894_new_n2461_; 
wire u0__abc_74894_new_n2462_; 
wire u0__abc_74894_new_n2463_; 
wire u0__abc_74894_new_n2464_; 
wire u0__abc_74894_new_n2465_; 
wire u0__abc_74894_new_n2466_; 
wire u0__abc_74894_new_n2467_; 
wire u0__abc_74894_new_n2468_; 
wire u0__abc_74894_new_n2469_; 
wire u0__abc_74894_new_n2470_; 
wire u0__abc_74894_new_n2471_; 
wire u0__abc_74894_new_n2472_; 
wire u0__abc_74894_new_n2473_; 
wire u0__abc_74894_new_n2474_; 
wire u0__abc_74894_new_n2476_; 
wire u0__abc_74894_new_n2477_; 
wire u0__abc_74894_new_n2478_; 
wire u0__abc_74894_new_n2479_; 
wire u0__abc_74894_new_n2480_; 
wire u0__abc_74894_new_n2481_; 
wire u0__abc_74894_new_n2482_; 
wire u0__abc_74894_new_n2483_; 
wire u0__abc_74894_new_n2484_; 
wire u0__abc_74894_new_n2485_; 
wire u0__abc_74894_new_n2486_; 
wire u0__abc_74894_new_n2487_; 
wire u0__abc_74894_new_n2488_; 
wire u0__abc_74894_new_n2489_; 
wire u0__abc_74894_new_n2490_; 
wire u0__abc_74894_new_n2492_; 
wire u0__abc_74894_new_n2493_; 
wire u0__abc_74894_new_n2494_; 
wire u0__abc_74894_new_n2495_; 
wire u0__abc_74894_new_n2496_; 
wire u0__abc_74894_new_n2497_; 
wire u0__abc_74894_new_n2498_; 
wire u0__abc_74894_new_n2499_; 
wire u0__abc_74894_new_n2500_; 
wire u0__abc_74894_new_n2501_; 
wire u0__abc_74894_new_n2502_; 
wire u0__abc_74894_new_n2503_; 
wire u0__abc_74894_new_n2504_; 
wire u0__abc_74894_new_n2505_; 
wire u0__abc_74894_new_n2506_; 
wire u0__abc_74894_new_n2508_; 
wire u0__abc_74894_new_n2509_; 
wire u0__abc_74894_new_n2510_; 
wire u0__abc_74894_new_n2511_; 
wire u0__abc_74894_new_n2512_; 
wire u0__abc_74894_new_n2513_; 
wire u0__abc_74894_new_n2514_; 
wire u0__abc_74894_new_n2515_; 
wire u0__abc_74894_new_n2516_; 
wire u0__abc_74894_new_n2517_; 
wire u0__abc_74894_new_n2518_; 
wire u0__abc_74894_new_n2519_; 
wire u0__abc_74894_new_n2520_; 
wire u0__abc_74894_new_n2521_; 
wire u0__abc_74894_new_n2522_; 
wire u0__abc_74894_new_n2524_; 
wire u0__abc_74894_new_n2525_; 
wire u0__abc_74894_new_n2526_; 
wire u0__abc_74894_new_n2527_; 
wire u0__abc_74894_new_n2528_; 
wire u0__abc_74894_new_n2529_; 
wire u0__abc_74894_new_n2530_; 
wire u0__abc_74894_new_n2531_; 
wire u0__abc_74894_new_n2532_; 
wire u0__abc_74894_new_n2533_; 
wire u0__abc_74894_new_n2534_; 
wire u0__abc_74894_new_n2535_; 
wire u0__abc_74894_new_n2536_; 
wire u0__abc_74894_new_n2537_; 
wire u0__abc_74894_new_n2538_; 
wire u0__abc_74894_new_n2540_; 
wire u0__abc_74894_new_n2541_; 
wire u0__abc_74894_new_n2542_; 
wire u0__abc_74894_new_n2543_; 
wire u0__abc_74894_new_n2544_; 
wire u0__abc_74894_new_n2545_; 
wire u0__abc_74894_new_n2546_; 
wire u0__abc_74894_new_n2547_; 
wire u0__abc_74894_new_n2548_; 
wire u0__abc_74894_new_n2549_; 
wire u0__abc_74894_new_n2550_; 
wire u0__abc_74894_new_n2551_; 
wire u0__abc_74894_new_n2552_; 
wire u0__abc_74894_new_n2553_; 
wire u0__abc_74894_new_n2554_; 
wire u0__abc_74894_new_n2556_; 
wire u0__abc_74894_new_n2557_; 
wire u0__abc_74894_new_n2558_; 
wire u0__abc_74894_new_n2559_; 
wire u0__abc_74894_new_n2560_; 
wire u0__abc_74894_new_n2561_; 
wire u0__abc_74894_new_n2562_; 
wire u0__abc_74894_new_n2563_; 
wire u0__abc_74894_new_n2564_; 
wire u0__abc_74894_new_n2565_; 
wire u0__abc_74894_new_n2566_; 
wire u0__abc_74894_new_n2567_; 
wire u0__abc_74894_new_n2568_; 
wire u0__abc_74894_new_n2569_; 
wire u0__abc_74894_new_n2570_; 
wire u0__abc_74894_new_n2572_; 
wire u0__abc_74894_new_n2573_; 
wire u0__abc_74894_new_n2574_; 
wire u0__abc_74894_new_n2575_; 
wire u0__abc_74894_new_n2576_; 
wire u0__abc_74894_new_n2577_; 
wire u0__abc_74894_new_n2578_; 
wire u0__abc_74894_new_n2579_; 
wire u0__abc_74894_new_n2580_; 
wire u0__abc_74894_new_n2581_; 
wire u0__abc_74894_new_n2582_; 
wire u0__abc_74894_new_n2583_; 
wire u0__abc_74894_new_n2584_; 
wire u0__abc_74894_new_n2585_; 
wire u0__abc_74894_new_n2586_; 
wire u0__abc_74894_new_n2588_; 
wire u0__abc_74894_new_n2589_; 
wire u0__abc_74894_new_n2590_; 
wire u0__abc_74894_new_n2591_; 
wire u0__abc_74894_new_n2592_; 
wire u0__abc_74894_new_n2593_; 
wire u0__abc_74894_new_n2594_; 
wire u0__abc_74894_new_n2595_; 
wire u0__abc_74894_new_n2596_; 
wire u0__abc_74894_new_n2597_; 
wire u0__abc_74894_new_n2598_; 
wire u0__abc_74894_new_n2599_; 
wire u0__abc_74894_new_n2600_; 
wire u0__abc_74894_new_n2601_; 
wire u0__abc_74894_new_n2602_; 
wire u0__abc_74894_new_n2604_; 
wire u0__abc_74894_new_n2605_; 
wire u0__abc_74894_new_n2606_; 
wire u0__abc_74894_new_n2607_; 
wire u0__abc_74894_new_n2608_; 
wire u0__abc_74894_new_n2609_; 
wire u0__abc_74894_new_n2610_; 
wire u0__abc_74894_new_n2611_; 
wire u0__abc_74894_new_n2612_; 
wire u0__abc_74894_new_n2613_; 
wire u0__abc_74894_new_n2614_; 
wire u0__abc_74894_new_n2615_; 
wire u0__abc_74894_new_n2616_; 
wire u0__abc_74894_new_n2617_; 
wire u0__abc_74894_new_n2618_; 
wire u0__abc_74894_new_n2620_; 
wire u0__abc_74894_new_n2621_; 
wire u0__abc_74894_new_n2622_; 
wire u0__abc_74894_new_n2623_; 
wire u0__abc_74894_new_n2624_; 
wire u0__abc_74894_new_n2625_; 
wire u0__abc_74894_new_n2626_; 
wire u0__abc_74894_new_n2627_; 
wire u0__abc_74894_new_n2628_; 
wire u0__abc_74894_new_n2629_; 
wire u0__abc_74894_new_n2630_; 
wire u0__abc_74894_new_n2631_; 
wire u0__abc_74894_new_n2632_; 
wire u0__abc_74894_new_n2633_; 
wire u0__abc_74894_new_n2634_; 
wire u0__abc_74894_new_n2636_; 
wire u0__abc_74894_new_n2637_; 
wire u0__abc_74894_new_n2638_; 
wire u0__abc_74894_new_n2639_; 
wire u0__abc_74894_new_n2640_; 
wire u0__abc_74894_new_n2641_; 
wire u0__abc_74894_new_n2642_; 
wire u0__abc_74894_new_n2643_; 
wire u0__abc_74894_new_n2644_; 
wire u0__abc_74894_new_n2645_; 
wire u0__abc_74894_new_n2646_; 
wire u0__abc_74894_new_n2647_; 
wire u0__abc_74894_new_n2648_; 
wire u0__abc_74894_new_n2649_; 
wire u0__abc_74894_new_n2650_; 
wire u0__abc_74894_new_n2652_; 
wire u0__abc_74894_new_n2653_; 
wire u0__abc_74894_new_n2654_; 
wire u0__abc_74894_new_n2655_; 
wire u0__abc_74894_new_n2656_; 
wire u0__abc_74894_new_n2657_; 
wire u0__abc_74894_new_n2658_; 
wire u0__abc_74894_new_n2659_; 
wire u0__abc_74894_new_n2660_; 
wire u0__abc_74894_new_n2661_; 
wire u0__abc_74894_new_n2662_; 
wire u0__abc_74894_new_n2663_; 
wire u0__abc_74894_new_n2664_; 
wire u0__abc_74894_new_n2665_; 
wire u0__abc_74894_new_n2666_; 
wire u0__abc_74894_new_n2668_; 
wire u0__abc_74894_new_n2669_; 
wire u0__abc_74894_new_n2670_; 
wire u0__abc_74894_new_n2671_; 
wire u0__abc_74894_new_n2672_; 
wire u0__abc_74894_new_n2673_; 
wire u0__abc_74894_new_n2674_; 
wire u0__abc_74894_new_n2675_; 
wire u0__abc_74894_new_n2676_; 
wire u0__abc_74894_new_n2677_; 
wire u0__abc_74894_new_n2678_; 
wire u0__abc_74894_new_n2679_; 
wire u0__abc_74894_new_n2680_; 
wire u0__abc_74894_new_n2681_; 
wire u0__abc_74894_new_n2682_; 
wire u0__abc_74894_new_n2684_; 
wire u0__abc_74894_new_n2685_; 
wire u0__abc_74894_new_n2686_; 
wire u0__abc_74894_new_n2687_; 
wire u0__abc_74894_new_n2688_; 
wire u0__abc_74894_new_n2689_; 
wire u0__abc_74894_new_n2690_; 
wire u0__abc_74894_new_n2691_; 
wire u0__abc_74894_new_n2692_; 
wire u0__abc_74894_new_n2693_; 
wire u0__abc_74894_new_n2694_; 
wire u0__abc_74894_new_n2695_; 
wire u0__abc_74894_new_n2696_; 
wire u0__abc_74894_new_n2697_; 
wire u0__abc_74894_new_n2698_; 
wire u0__abc_74894_new_n2700_; 
wire u0__abc_74894_new_n2701_; 
wire u0__abc_74894_new_n2702_; 
wire u0__abc_74894_new_n2703_; 
wire u0__abc_74894_new_n2704_; 
wire u0__abc_74894_new_n2705_; 
wire u0__abc_74894_new_n2706_; 
wire u0__abc_74894_new_n2707_; 
wire u0__abc_74894_new_n2708_; 
wire u0__abc_74894_new_n2709_; 
wire u0__abc_74894_new_n2710_; 
wire u0__abc_74894_new_n2711_; 
wire u0__abc_74894_new_n2712_; 
wire u0__abc_74894_new_n2713_; 
wire u0__abc_74894_new_n2714_; 
wire u0__abc_74894_new_n2716_; 
wire u0__abc_74894_new_n2717_; 
wire u0__abc_74894_new_n2718_; 
wire u0__abc_74894_new_n2719_; 
wire u0__abc_74894_new_n2720_; 
wire u0__abc_74894_new_n2721_; 
wire u0__abc_74894_new_n2722_; 
wire u0__abc_74894_new_n2723_; 
wire u0__abc_74894_new_n2724_; 
wire u0__abc_74894_new_n2725_; 
wire u0__abc_74894_new_n2726_; 
wire u0__abc_74894_new_n2727_; 
wire u0__abc_74894_new_n2728_; 
wire u0__abc_74894_new_n2729_; 
wire u0__abc_74894_new_n2730_; 
wire u0__abc_74894_new_n2732_; 
wire u0__abc_74894_new_n2733_; 
wire u0__abc_74894_new_n2734_; 
wire u0__abc_74894_new_n2735_; 
wire u0__abc_74894_new_n2736_; 
wire u0__abc_74894_new_n2737_; 
wire u0__abc_74894_new_n2738_; 
wire u0__abc_74894_new_n2739_; 
wire u0__abc_74894_new_n2740_; 
wire u0__abc_74894_new_n2741_; 
wire u0__abc_74894_new_n2742_; 
wire u0__abc_74894_new_n2743_; 
wire u0__abc_74894_new_n2744_; 
wire u0__abc_74894_new_n2745_; 
wire u0__abc_74894_new_n2746_; 
wire u0__abc_74894_new_n2748_; 
wire u0__abc_74894_new_n2749_; 
wire u0__abc_74894_new_n2750_; 
wire u0__abc_74894_new_n2751_; 
wire u0__abc_74894_new_n2752_; 
wire u0__abc_74894_new_n2753_; 
wire u0__abc_74894_new_n2754_; 
wire u0__abc_74894_new_n2755_; 
wire u0__abc_74894_new_n2756_; 
wire u0__abc_74894_new_n2757_; 
wire u0__abc_74894_new_n2758_; 
wire u0__abc_74894_new_n2759_; 
wire u0__abc_74894_new_n2760_; 
wire u0__abc_74894_new_n2761_; 
wire u0__abc_74894_new_n2762_; 
wire u0__abc_74894_new_n2764_; 
wire u0__abc_74894_new_n2765_; 
wire u0__abc_74894_new_n2766_; 
wire u0__abc_74894_new_n2767_; 
wire u0__abc_74894_new_n2768_; 
wire u0__abc_74894_new_n2769_; 
wire u0__abc_74894_new_n2770_; 
wire u0__abc_74894_new_n2771_; 
wire u0__abc_74894_new_n2772_; 
wire u0__abc_74894_new_n2773_; 
wire u0__abc_74894_new_n2774_; 
wire u0__abc_74894_new_n2775_; 
wire u0__abc_74894_new_n2776_; 
wire u0__abc_74894_new_n2777_; 
wire u0__abc_74894_new_n2778_; 
wire u0__abc_74894_new_n2780_; 
wire u0__abc_74894_new_n2781_; 
wire u0__abc_74894_new_n2782_; 
wire u0__abc_74894_new_n2783_; 
wire u0__abc_74894_new_n2784_; 
wire u0__abc_74894_new_n2785_; 
wire u0__abc_74894_new_n2786_; 
wire u0__abc_74894_new_n2787_; 
wire u0__abc_74894_new_n2788_; 
wire u0__abc_74894_new_n2789_; 
wire u0__abc_74894_new_n2790_; 
wire u0__abc_74894_new_n2791_; 
wire u0__abc_74894_new_n2792_; 
wire u0__abc_74894_new_n2793_; 
wire u0__abc_74894_new_n2794_; 
wire u0__abc_74894_new_n2796_; 
wire u0__abc_74894_new_n2797_; 
wire u0__abc_74894_new_n2798_; 
wire u0__abc_74894_new_n2799_; 
wire u0__abc_74894_new_n2800_; 
wire u0__abc_74894_new_n2801_; 
wire u0__abc_74894_new_n2802_; 
wire u0__abc_74894_new_n2803_; 
wire u0__abc_74894_new_n2804_; 
wire u0__abc_74894_new_n2805_; 
wire u0__abc_74894_new_n2806_; 
wire u0__abc_74894_new_n2807_; 
wire u0__abc_74894_new_n2808_; 
wire u0__abc_74894_new_n2809_; 
wire u0__abc_74894_new_n2810_; 
wire u0__abc_74894_new_n2812_; 
wire u0__abc_74894_new_n2813_; 
wire u0__abc_74894_new_n2814_; 
wire u0__abc_74894_new_n2815_; 
wire u0__abc_74894_new_n2816_; 
wire u0__abc_74894_new_n2817_; 
wire u0__abc_74894_new_n2818_; 
wire u0__abc_74894_new_n2819_; 
wire u0__abc_74894_new_n2820_; 
wire u0__abc_74894_new_n2821_; 
wire u0__abc_74894_new_n2822_; 
wire u0__abc_74894_new_n2823_; 
wire u0__abc_74894_new_n2824_; 
wire u0__abc_74894_new_n2825_; 
wire u0__abc_74894_new_n2826_; 
wire u0__abc_74894_new_n2828_; 
wire u0__abc_74894_new_n2829_; 
wire u0__abc_74894_new_n2830_; 
wire u0__abc_74894_new_n2831_; 
wire u0__abc_74894_new_n2832_; 
wire u0__abc_74894_new_n2833_; 
wire u0__abc_74894_new_n2834_; 
wire u0__abc_74894_new_n2835_; 
wire u0__abc_74894_new_n2836_; 
wire u0__abc_74894_new_n2837_; 
wire u0__abc_74894_new_n2838_; 
wire u0__abc_74894_new_n2839_; 
wire u0__abc_74894_new_n2840_; 
wire u0__abc_74894_new_n2841_; 
wire u0__abc_74894_new_n2842_; 
wire u0__abc_74894_new_n2844_; 
wire u0__abc_74894_new_n2845_; 
wire u0__abc_74894_new_n2846_; 
wire u0__abc_74894_new_n2847_; 
wire u0__abc_74894_new_n2848_; 
wire u0__abc_74894_new_n2849_; 
wire u0__abc_74894_new_n2850_; 
wire u0__abc_74894_new_n2851_; 
wire u0__abc_74894_new_n2852_; 
wire u0__abc_74894_new_n2853_; 
wire u0__abc_74894_new_n2854_; 
wire u0__abc_74894_new_n2855_; 
wire u0__abc_74894_new_n2856_; 
wire u0__abc_74894_new_n2857_; 
wire u0__abc_74894_new_n2858_; 
wire u0__abc_74894_new_n2860_; 
wire u0__abc_74894_new_n2861_; 
wire u0__abc_74894_new_n2862_; 
wire u0__abc_74894_new_n2863_; 
wire u0__abc_74894_new_n2864_; 
wire u0__abc_74894_new_n2865_; 
wire u0__abc_74894_new_n2866_; 
wire u0__abc_74894_new_n2867_; 
wire u0__abc_74894_new_n2868_; 
wire u0__abc_74894_new_n2869_; 
wire u0__abc_74894_new_n2870_; 
wire u0__abc_74894_new_n2871_; 
wire u0__abc_74894_new_n2872_; 
wire u0__abc_74894_new_n2873_; 
wire u0__abc_74894_new_n2874_; 
wire u0__abc_74894_new_n2876_; 
wire u0__abc_74894_new_n2877_; 
wire u0__abc_74894_new_n2878_; 
wire u0__abc_74894_new_n2879_; 
wire u0__abc_74894_new_n2880_; 
wire u0__abc_74894_new_n2881_; 
wire u0__abc_74894_new_n2882_; 
wire u0__abc_74894_new_n2883_; 
wire u0__abc_74894_new_n2884_; 
wire u0__abc_74894_new_n2885_; 
wire u0__abc_74894_new_n2886_; 
wire u0__abc_74894_new_n2887_; 
wire u0__abc_74894_new_n2888_; 
wire u0__abc_74894_new_n2889_; 
wire u0__abc_74894_new_n2890_; 
wire u0__abc_74894_new_n2970_; 
wire u0__abc_74894_new_n2973_; 
wire u0__abc_74894_new_n2974_; 
wire u0__abc_74894_new_n2975_; 
wire u0__abc_74894_new_n2976_; 
wire u0__abc_74894_new_n2977_; 
wire u0__abc_74894_new_n2978_; 
wire u0__abc_74894_new_n2979_; 
wire u0__abc_74894_new_n2980_; 
wire u0__abc_74894_new_n2981_; 
wire u0__abc_74894_new_n2982_; 
wire u0__abc_74894_new_n2983_; 
wire u0__abc_74894_new_n2984_; 
wire u0__abc_74894_new_n2985_; 
wire u0__abc_74894_new_n2986_; 
wire u0__abc_74894_new_n2987_; 
wire u0__abc_74894_new_n2989_; 
wire u0__abc_74894_new_n2990_; 
wire u0__abc_74894_new_n2991_; 
wire u0__abc_74894_new_n2992_; 
wire u0__abc_74894_new_n2993_; 
wire u0__abc_74894_new_n2994_; 
wire u0__abc_74894_new_n2995_; 
wire u0__abc_74894_new_n2996_; 
wire u0__abc_74894_new_n2997_; 
wire u0__abc_74894_new_n2998_; 
wire u0__abc_74894_new_n2999_; 
wire u0__abc_74894_new_n3000_; 
wire u0__abc_74894_new_n3001_; 
wire u0__abc_74894_new_n3002_; 
wire u0__abc_74894_new_n3003_; 
wire u0__abc_74894_new_n3005_; 
wire u0__abc_74894_new_n3006_; 
wire u0__abc_74894_new_n3007_; 
wire u0__abc_74894_new_n3008_; 
wire u0__abc_74894_new_n3009_; 
wire u0__abc_74894_new_n3010_; 
wire u0__abc_74894_new_n3011_; 
wire u0__abc_74894_new_n3012_; 
wire u0__abc_74894_new_n3013_; 
wire u0__abc_74894_new_n3014_; 
wire u0__abc_74894_new_n3015_; 
wire u0__abc_74894_new_n3016_; 
wire u0__abc_74894_new_n3017_; 
wire u0__abc_74894_new_n3018_; 
wire u0__abc_74894_new_n3019_; 
wire u0__abc_74894_new_n3021_; 
wire u0__abc_74894_new_n3022_; 
wire u0__abc_74894_new_n3023_; 
wire u0__abc_74894_new_n3024_; 
wire u0__abc_74894_new_n3025_; 
wire u0__abc_74894_new_n3026_; 
wire u0__abc_74894_new_n3027_; 
wire u0__abc_74894_new_n3028_; 
wire u0__abc_74894_new_n3029_; 
wire u0__abc_74894_new_n3030_; 
wire u0__abc_74894_new_n3031_; 
wire u0__abc_74894_new_n3032_; 
wire u0__abc_74894_new_n3033_; 
wire u0__abc_74894_new_n3034_; 
wire u0__abc_74894_new_n3035_; 
wire u0__abc_74894_new_n3037_; 
wire u0__abc_74894_new_n3038_; 
wire u0__abc_74894_new_n3039_; 
wire u0__abc_74894_new_n3040_; 
wire u0__abc_74894_new_n3041_; 
wire u0__abc_74894_new_n3042_; 
wire u0__abc_74894_new_n3043_; 
wire u0__abc_74894_new_n3044_; 
wire u0__abc_74894_new_n3045_; 
wire u0__abc_74894_new_n3046_; 
wire u0__abc_74894_new_n3047_; 
wire u0__abc_74894_new_n3048_; 
wire u0__abc_74894_new_n3049_; 
wire u0__abc_74894_new_n3050_; 
wire u0__abc_74894_new_n3051_; 
wire u0__abc_74894_new_n3053_; 
wire u0__abc_74894_new_n3054_; 
wire u0__abc_74894_new_n3055_; 
wire u0__abc_74894_new_n3056_; 
wire u0__abc_74894_new_n3057_; 
wire u0__abc_74894_new_n3058_; 
wire u0__abc_74894_new_n3059_; 
wire u0__abc_74894_new_n3060_; 
wire u0__abc_74894_new_n3061_; 
wire u0__abc_74894_new_n3062_; 
wire u0__abc_74894_new_n3063_; 
wire u0__abc_74894_new_n3064_; 
wire u0__abc_74894_new_n3065_; 
wire u0__abc_74894_new_n3066_; 
wire u0__abc_74894_new_n3067_; 
wire u0__abc_74894_new_n3069_; 
wire u0__abc_74894_new_n3070_; 
wire u0__abc_74894_new_n3071_; 
wire u0__abc_74894_new_n3072_; 
wire u0__abc_74894_new_n3073_; 
wire u0__abc_74894_new_n3074_; 
wire u0__abc_74894_new_n3075_; 
wire u0__abc_74894_new_n3076_; 
wire u0__abc_74894_new_n3077_; 
wire u0__abc_74894_new_n3078_; 
wire u0__abc_74894_new_n3079_; 
wire u0__abc_74894_new_n3080_; 
wire u0__abc_74894_new_n3081_; 
wire u0__abc_74894_new_n3082_; 
wire u0__abc_74894_new_n3083_; 
wire u0__abc_74894_new_n3101_; 
wire u0__abc_74894_new_n3102_; 
wire u0__abc_74894_new_n3103_; 
wire u0__abc_74894_new_n3104_; 
wire u0__abc_74894_new_n3105_; 
wire u0__abc_74894_new_n3106_; 
wire u0__abc_74894_new_n3107_; 
wire u0__abc_74894_new_n3108_; 
wire u0__abc_74894_new_n3109_; 
wire u0__abc_74894_new_n3110_; 
wire u0__abc_74894_new_n3111_; 
wire u0__abc_74894_new_n3112_; 
wire u0__abc_74894_new_n3113_; 
wire u0__abc_74894_new_n3114_; 
wire u0__abc_74894_new_n3115_; 
wire u0__abc_74894_new_n3117_; 
wire u0__abc_74894_new_n3118_; 
wire u0__abc_74894_new_n3119_; 
wire u0__abc_74894_new_n3120_; 
wire u0__abc_74894_new_n3121_; 
wire u0__abc_74894_new_n3122_; 
wire u0__abc_74894_new_n3123_; 
wire u0__abc_74894_new_n3124_; 
wire u0__abc_74894_new_n3125_; 
wire u0__abc_74894_new_n3126_; 
wire u0__abc_74894_new_n3127_; 
wire u0__abc_74894_new_n3128_; 
wire u0__abc_74894_new_n3129_; 
wire u0__abc_74894_new_n3130_; 
wire u0__abc_74894_new_n3131_; 
wire u0__abc_74894_new_n3133_; 
wire u0__abc_74894_new_n3134_; 
wire u0__abc_74894_new_n3135_; 
wire u0__abc_74894_new_n3136_; 
wire u0__abc_74894_new_n3137_; 
wire u0__abc_74894_new_n3138_; 
wire u0__abc_74894_new_n3139_; 
wire u0__abc_74894_new_n3140_; 
wire u0__abc_74894_new_n3141_; 
wire u0__abc_74894_new_n3142_; 
wire u0__abc_74894_new_n3143_; 
wire u0__abc_74894_new_n3144_; 
wire u0__abc_74894_new_n3145_; 
wire u0__abc_74894_new_n3146_; 
wire u0__abc_74894_new_n3147_; 
wire u0__abc_74894_new_n3469_; 
wire u0__abc_74894_new_n3470_; 
wire u0__abc_74894_new_n3471_; 
wire u0__abc_74894_new_n3472_; 
wire u0__abc_74894_new_n3473_; 
wire u0__abc_74894_new_n3474_; 
wire u0__abc_74894_new_n3475_; 
wire u0__abc_74894_new_n3476_; 
wire u0__abc_74894_new_n3477_; 
wire u0__abc_74894_new_n3479_; 
wire u0__abc_74894_new_n3481_; 
wire u0__abc_74894_new_n3483_; 
wire u0__abc_74894_new_n3485_; 
wire u0__abc_74894_new_n3487_; 
wire u0__abc_74894_new_n3489_; 
wire u0__abc_74894_new_n3491_; 
wire u0__abc_74894_new_n3493_; 
wire u0__abc_74894_new_n3494_; 
wire u0__abc_74894_new_n3496_; 
wire u0__abc_74894_new_n3497_; 
wire u0__abc_74894_new_n3499_; 
wire u0__abc_74894_new_n3500_; 
wire u0__abc_74894_new_n3502_; 
wire u0__abc_74894_new_n3503_; 
wire u0__abc_74894_new_n3505_; 
wire u0__abc_74894_new_n3506_; 
wire u0__abc_74894_new_n3508_; 
wire u0__abc_74894_new_n3509_; 
wire u0__abc_74894_new_n3511_; 
wire u0__abc_74894_new_n3512_; 
wire u0__abc_74894_new_n3514_; 
wire u0__abc_74894_new_n3515_; 
wire u0__abc_74894_new_n3517_; 
wire u0__abc_74894_new_n3518_; 
wire u0__abc_74894_new_n3520_; 
wire u0__abc_74894_new_n3521_; 
wire u0__abc_74894_new_n3523_; 
wire u0__abc_74894_new_n3524_; 
wire u0__abc_74894_new_n3526_; 
wire u0__abc_74894_new_n3527_; 
wire u0__abc_74894_new_n3529_; 
wire u0__abc_74894_new_n3530_; 
wire u0__abc_74894_new_n3532_; 
wire u0__abc_74894_new_n3533_; 
wire u0__abc_74894_new_n3535_; 
wire u0__abc_74894_new_n3536_; 
wire u0__abc_74894_new_n3538_; 
wire u0__abc_74894_new_n3539_; 
wire u0__abc_74894_new_n3541_; 
wire u0__abc_74894_new_n3542_; 
wire u0__abc_74894_new_n3544_; 
wire u0__abc_74894_new_n3545_; 
wire u0__abc_74894_new_n3547_; 
wire u0__abc_74894_new_n3548_; 
wire u0__abc_74894_new_n3550_; 
wire u0__abc_74894_new_n3551_; 
wire u0__abc_74894_new_n3553_; 
wire u0__abc_74894_new_n3554_; 
wire u0__abc_74894_new_n3556_; 
wire u0__abc_74894_new_n3557_; 
wire u0__abc_74894_new_n3559_; 
wire u0__abc_74894_new_n3560_; 
wire u0__abc_74894_new_n3562_; 
wire u0__abc_74894_new_n3563_; 
wire u0__abc_74894_new_n3565_; 
wire u0__abc_74894_new_n3566_; 
wire u0__abc_74894_new_n3568_; 
wire u0__abc_74894_new_n3569_; 
wire u0__abc_74894_new_n3571_; 
wire u0__abc_74894_new_n3572_; 
wire u0__abc_74894_new_n3574_; 
wire u0__abc_74894_new_n3575_; 
wire u0__abc_74894_new_n3577_; 
wire u0__abc_74894_new_n3578_; 
wire u0__abc_74894_new_n3580_; 
wire u0__abc_74894_new_n3581_; 
wire u0__abc_74894_new_n3583_; 
wire u0__abc_74894_new_n3584_; 
wire u0__abc_74894_new_n3586_; 
wire u0__abc_74894_new_n3587_; 
wire u0__abc_74894_new_n3589_; 
wire u0__abc_74894_new_n3590_; 
wire u0__abc_74894_new_n3592_; 
wire u0__abc_74894_new_n3593_; 
wire u0__abc_74894_new_n3594_; 
wire u0__abc_74894_new_n3595_; 
wire u0__abc_74894_new_n3596_; 
wire u0__abc_74894_new_n3597_; 
wire u0__abc_74894_new_n3598_; 
wire u0__abc_74894_new_n3599_; 
wire u0__abc_74894_new_n3601_; 
wire u0__abc_74894_new_n3602_; 
wire u0__abc_74894_new_n3604_; 
wire u0__abc_74894_new_n3605_; 
wire u0__abc_74894_new_n3607_; 
wire u0__abc_74894_new_n3608_; 
wire u0__abc_74894_new_n3610_; 
wire u0__abc_74894_new_n3611_; 
wire u0__abc_74894_new_n3613_; 
wire u0__abc_74894_new_n3614_; 
wire u0__abc_74894_new_n3616_; 
wire u0__abc_74894_new_n3617_; 
wire u0__abc_74894_new_n3619_; 
wire u0__abc_74894_new_n3620_; 
wire u0__abc_74894_new_n3622_; 
wire u0__abc_74894_new_n3623_; 
wire u0__abc_74894_new_n3625_; 
wire u0__abc_74894_new_n3626_; 
wire u0__abc_74894_new_n3628_; 
wire u0__abc_74894_new_n3629_; 
wire u0__abc_74894_new_n3631_; 
wire u0__abc_74894_new_n3632_; 
wire u0__abc_74894_new_n3633_; 
wire u0__abc_74894_new_n3634_; 
wire u0__abc_74894_new_n3635_; 
wire u0__abc_74894_new_n3637_; 
wire u0__abc_74894_new_n3638_; 
wire u0__abc_74894_new_n3640_; 
wire u0__abc_74894_new_n3641_; 
wire u0__abc_74894_new_n3643_; 
wire u0__abc_74894_new_n3644_; 
wire u0__abc_74894_new_n3646_; 
wire u0__abc_74894_new_n3647_; 
wire u0__abc_74894_new_n3649_; 
wire u0__abc_74894_new_n3650_; 
wire u0__abc_74894_new_n3652_; 
wire u0__abc_74894_new_n3653_; 
wire u0__abc_74894_new_n3655_; 
wire u0__abc_74894_new_n3656_; 
wire u0__abc_74894_new_n3658_; 
wire u0__abc_74894_new_n3659_; 
wire u0__abc_74894_new_n3661_; 
wire u0__abc_74894_new_n3662_; 
wire u0__abc_74894_new_n3664_; 
wire u0__abc_74894_new_n3665_; 
wire u0__abc_74894_new_n3667_; 
wire u0__abc_74894_new_n3668_; 
wire u0__abc_74894_new_n3670_; 
wire u0__abc_74894_new_n3671_; 
wire u0__abc_74894_new_n3673_; 
wire u0__abc_74894_new_n3674_; 
wire u0__abc_74894_new_n3676_; 
wire u0__abc_74894_new_n3677_; 
wire u0__abc_74894_new_n3679_; 
wire u0__abc_74894_new_n3680_; 
wire u0__abc_74894_new_n3682_; 
wire u0__abc_74894_new_n3683_; 
wire u0__abc_74894_new_n3685_; 
wire u0__abc_74894_new_n3686_; 
wire u0__abc_74894_new_n3688_; 
wire u0__abc_74894_new_n3689_; 
wire u0__abc_74894_new_n3690_; 
wire u0__abc_74894_new_n3691_; 
wire u0__abc_74894_new_n3692_; 
wire u0__abc_74894_new_n3693_; 
wire u0__abc_74894_new_n3694_; 
wire u0__abc_74894_new_n3695_; 
wire u0__abc_74894_new_n3696_; 
wire u0__abc_74894_new_n3697_; 
wire u0__abc_74894_new_n3698_; 
wire u0__abc_74894_new_n3699_; 
wire u0__abc_74894_new_n3700_; 
wire u0__abc_74894_new_n3701_; 
wire u0__abc_74894_new_n3702_; 
wire u0__abc_74894_new_n3703_; 
wire u0__abc_74894_new_n3704_; 
wire u0__abc_74894_new_n3705_; 
wire u0__abc_74894_new_n3706_; 
wire u0__abc_74894_new_n3707_; 
wire u0__abc_74894_new_n3708_; 
wire u0__abc_74894_new_n3709_; 
wire u0__abc_74894_new_n3710_; 
wire u0__abc_74894_new_n3711_; 
wire u0__abc_74894_new_n3712_; 
wire u0__abc_74894_new_n3713_; 
wire u0__abc_74894_new_n3714_; 
wire u0__abc_74894_new_n3715_; 
wire u0__abc_74894_new_n3716_; 
wire u0__abc_74894_new_n3717_; 
wire u0__abc_74894_new_n3718_; 
wire u0__abc_74894_new_n3719_; 
wire u0__abc_74894_new_n3720_; 
wire u0__abc_74894_new_n3721_; 
wire u0__abc_74894_new_n3722_; 
wire u0__abc_74894_new_n3723_; 
wire u0__abc_74894_new_n3724_; 
wire u0__abc_74894_new_n3725_; 
wire u0__abc_74894_new_n3726_; 
wire u0__abc_74894_new_n3727_; 
wire u0__abc_74894_new_n3728_; 
wire u0__abc_74894_new_n3729_; 
wire u0__abc_74894_new_n3730_; 
wire u0__abc_74894_new_n3731_; 
wire u0__abc_74894_new_n3732_; 
wire u0__abc_74894_new_n3733_; 
wire u0__abc_74894_new_n3734_; 
wire u0__abc_74894_new_n3735_; 
wire u0__abc_74894_new_n3736_; 
wire u0__abc_74894_new_n3737_; 
wire u0__abc_74894_new_n3738_; 
wire u0__abc_74894_new_n3739_; 
wire u0__abc_74894_new_n3740_; 
wire u0__abc_74894_new_n3741_; 
wire u0__abc_74894_new_n3742_; 
wire u0__abc_74894_new_n3743_; 
wire u0__abc_74894_new_n3744_; 
wire u0__abc_74894_new_n3745_; 
wire u0__abc_74894_new_n3746_; 
wire u0__abc_74894_new_n3747_; 
wire u0__abc_74894_new_n3748_; 
wire u0__abc_74894_new_n3749_; 
wire u0__abc_74894_new_n3750_; 
wire u0__abc_74894_new_n3751_; 
wire u0__abc_74894_new_n3752_; 
wire u0__abc_74894_new_n3753_; 
wire u0__abc_74894_new_n3754_; 
wire u0__abc_74894_new_n3756_; 
wire u0__abc_74894_new_n3757_; 
wire u0__abc_74894_new_n3758_; 
wire u0__abc_74894_new_n3759_; 
wire u0__abc_74894_new_n3760_; 
wire u0__abc_74894_new_n3761_; 
wire u0__abc_74894_new_n3762_; 
wire u0__abc_74894_new_n3763_; 
wire u0__abc_74894_new_n3764_; 
wire u0__abc_74894_new_n3765_; 
wire u0__abc_74894_new_n3766_; 
wire u0__abc_74894_new_n3767_; 
wire u0__abc_74894_new_n3768_; 
wire u0__abc_74894_new_n3769_; 
wire u0__abc_74894_new_n3770_; 
wire u0__abc_74894_new_n3771_; 
wire u0__abc_74894_new_n3772_; 
wire u0__abc_74894_new_n3773_; 
wire u0__abc_74894_new_n3774_; 
wire u0__abc_74894_new_n3775_; 
wire u0__abc_74894_new_n3776_; 
wire u0__abc_74894_new_n3778_; 
wire u0__abc_74894_new_n3779_; 
wire u0__abc_74894_new_n3780_; 
wire u0__abc_74894_new_n3781_; 
wire u0__abc_74894_new_n3782_; 
wire u0__abc_74894_new_n3783_; 
wire u0__abc_74894_new_n3784_; 
wire u0__abc_74894_new_n3785_; 
wire u0__abc_74894_new_n3786_; 
wire u0__abc_74894_new_n3787_; 
wire u0__abc_74894_new_n3788_; 
wire u0__abc_74894_new_n3789_; 
wire u0__abc_74894_new_n3790_; 
wire u0__abc_74894_new_n3791_; 
wire u0__abc_74894_new_n3792_; 
wire u0__abc_74894_new_n3793_; 
wire u0__abc_74894_new_n3794_; 
wire u0__abc_74894_new_n3795_; 
wire u0__abc_74894_new_n3797_; 
wire u0__abc_74894_new_n3798_; 
wire u0__abc_74894_new_n3799_; 
wire u0__abc_74894_new_n3800_; 
wire u0__abc_74894_new_n3801_; 
wire u0__abc_74894_new_n3802_; 
wire u0__abc_74894_new_n3803_; 
wire u0__abc_74894_new_n3804_; 
wire u0__abc_74894_new_n3805_; 
wire u0__abc_74894_new_n3806_; 
wire u0__abc_74894_new_n3807_; 
wire u0__abc_74894_new_n3808_; 
wire u0__abc_74894_new_n3809_; 
wire u0__abc_74894_new_n3810_; 
wire u0__abc_74894_new_n3811_; 
wire u0__abc_74894_new_n3812_; 
wire u0__abc_74894_new_n3813_; 
wire u0__abc_74894_new_n3814_; 
wire u0__abc_74894_new_n3815_; 
wire u0__abc_74894_new_n3816_; 
wire u0__abc_74894_new_n3817_; 
wire u0__abc_74894_new_n3818_; 
wire u0__abc_74894_new_n3819_; 
wire u0__abc_74894_new_n3820_; 
wire u0__abc_74894_new_n3822_; 
wire u0__abc_74894_new_n3823_; 
wire u0__abc_74894_new_n3824_; 
wire u0__abc_74894_new_n3825_; 
wire u0__abc_74894_new_n3826_; 
wire u0__abc_74894_new_n3827_; 
wire u0__abc_74894_new_n3828_; 
wire u0__abc_74894_new_n3829_; 
wire u0__abc_74894_new_n3830_; 
wire u0__abc_74894_new_n3831_; 
wire u0__abc_74894_new_n3832_; 
wire u0__abc_74894_new_n3833_; 
wire u0__abc_74894_new_n3834_; 
wire u0__abc_74894_new_n3835_; 
wire u0__abc_74894_new_n3836_; 
wire u0__abc_74894_new_n3837_; 
wire u0__abc_74894_new_n3838_; 
wire u0__abc_74894_new_n3840_; 
wire u0__abc_74894_new_n3841_; 
wire u0__abc_74894_new_n3842_; 
wire u0__abc_74894_new_n3843_; 
wire u0__abc_74894_new_n3844_; 
wire u0__abc_74894_new_n3845_; 
wire u0__abc_74894_new_n3846_; 
wire u0__abc_74894_new_n3847_; 
wire u0__abc_74894_new_n3848_; 
wire u0__abc_74894_new_n3849_; 
wire u0__abc_74894_new_n3850_; 
wire u0__abc_74894_new_n3851_; 
wire u0__abc_74894_new_n3852_; 
wire u0__abc_74894_new_n3853_; 
wire u0__abc_74894_new_n3854_; 
wire u0__abc_74894_new_n3855_; 
wire u0__abc_74894_new_n3856_; 
wire u0__abc_74894_new_n3857_; 
wire u0__abc_74894_new_n3858_; 
wire u0__abc_74894_new_n3859_; 
wire u0__abc_74894_new_n3860_; 
wire u0__abc_74894_new_n3861_; 
wire u0__abc_74894_new_n3863_; 
wire u0__abc_74894_new_n3864_; 
wire u0__abc_74894_new_n3865_; 
wire u0__abc_74894_new_n3866_; 
wire u0__abc_74894_new_n3867_; 
wire u0__abc_74894_new_n3868_; 
wire u0__abc_74894_new_n3869_; 
wire u0__abc_74894_new_n3870_; 
wire u0__abc_74894_new_n3871_; 
wire u0__abc_74894_new_n3872_; 
wire u0__abc_74894_new_n3873_; 
wire u0__abc_74894_new_n3874_; 
wire u0__abc_74894_new_n3875_; 
wire u0__abc_74894_new_n3876_; 
wire u0__abc_74894_new_n3877_; 
wire u0__abc_74894_new_n3878_; 
wire u0__abc_74894_new_n3879_; 
wire u0__abc_74894_new_n3881_; 
wire u0__abc_74894_new_n3882_; 
wire u0__abc_74894_new_n3883_; 
wire u0__abc_74894_new_n3884_; 
wire u0__abc_74894_new_n3885_; 
wire u0__abc_74894_new_n3886_; 
wire u0__abc_74894_new_n3887_; 
wire u0__abc_74894_new_n3888_; 
wire u0__abc_74894_new_n3889_; 
wire u0__abc_74894_new_n3890_; 
wire u0__abc_74894_new_n3891_; 
wire u0__abc_74894_new_n3892_; 
wire u0__abc_74894_new_n3893_; 
wire u0__abc_74894_new_n3894_; 
wire u0__abc_74894_new_n3895_; 
wire u0__abc_74894_new_n3896_; 
wire u0__abc_74894_new_n3897_; 
wire u0__abc_74894_new_n3898_; 
wire u0__abc_74894_new_n3900_; 
wire u0__abc_74894_new_n3901_; 
wire u0__abc_74894_new_n3902_; 
wire u0__abc_74894_new_n3903_; 
wire u0__abc_74894_new_n3904_; 
wire u0__abc_74894_new_n3905_; 
wire u0__abc_74894_new_n3906_; 
wire u0__abc_74894_new_n3907_; 
wire u0__abc_74894_new_n3908_; 
wire u0__abc_74894_new_n3909_; 
wire u0__abc_74894_new_n3910_; 
wire u0__abc_74894_new_n3911_; 
wire u0__abc_74894_new_n3912_; 
wire u0__abc_74894_new_n3913_; 
wire u0__abc_74894_new_n3914_; 
wire u0__abc_74894_new_n3915_; 
wire u0__abc_74894_new_n3916_; 
wire u0__abc_74894_new_n3918_; 
wire u0__abc_74894_new_n3919_; 
wire u0__abc_74894_new_n3920_; 
wire u0__abc_74894_new_n3921_; 
wire u0__abc_74894_new_n3922_; 
wire u0__abc_74894_new_n3923_; 
wire u0__abc_74894_new_n3924_; 
wire u0__abc_74894_new_n3925_; 
wire u0__abc_74894_new_n3926_; 
wire u0__abc_74894_new_n3927_; 
wire u0__abc_74894_new_n3928_; 
wire u0__abc_74894_new_n3929_; 
wire u0__abc_74894_new_n3930_; 
wire u0__abc_74894_new_n3931_; 
wire u0__abc_74894_new_n3932_; 
wire u0__abc_74894_new_n3933_; 
wire u0__abc_74894_new_n3934_; 
wire u0__abc_74894_new_n3935_; 
wire u0__abc_74894_new_n3936_; 
wire u0__abc_74894_new_n3937_; 
wire u0__abc_74894_new_n3939_; 
wire u0__abc_74894_new_n3940_; 
wire u0__abc_74894_new_n3941_; 
wire u0__abc_74894_new_n3942_; 
wire u0__abc_74894_new_n3943_; 
wire u0__abc_74894_new_n3944_; 
wire u0__abc_74894_new_n3945_; 
wire u0__abc_74894_new_n3946_; 
wire u0__abc_74894_new_n3947_; 
wire u0__abc_74894_new_n3948_; 
wire u0__abc_74894_new_n3949_; 
wire u0__abc_74894_new_n3950_; 
wire u0__abc_74894_new_n3951_; 
wire u0__abc_74894_new_n3952_; 
wire u0__abc_74894_new_n3953_; 
wire u0__abc_74894_new_n3954_; 
wire u0__abc_74894_new_n3955_; 
wire u0__abc_74894_new_n3957_; 
wire u0__abc_74894_new_n3958_; 
wire u0__abc_74894_new_n3959_; 
wire u0__abc_74894_new_n3960_; 
wire u0__abc_74894_new_n3961_; 
wire u0__abc_74894_new_n3962_; 
wire u0__abc_74894_new_n3963_; 
wire u0__abc_74894_new_n3964_; 
wire u0__abc_74894_new_n3965_; 
wire u0__abc_74894_new_n3966_; 
wire u0__abc_74894_new_n3967_; 
wire u0__abc_74894_new_n3968_; 
wire u0__abc_74894_new_n3969_; 
wire u0__abc_74894_new_n3970_; 
wire u0__abc_74894_new_n3971_; 
wire u0__abc_74894_new_n3972_; 
wire u0__abc_74894_new_n3973_; 
wire u0__abc_74894_new_n3974_; 
wire u0__abc_74894_new_n3976_; 
wire u0__abc_74894_new_n3977_; 
wire u0__abc_74894_new_n3978_; 
wire u0__abc_74894_new_n3979_; 
wire u0__abc_74894_new_n3980_; 
wire u0__abc_74894_new_n3981_; 
wire u0__abc_74894_new_n3982_; 
wire u0__abc_74894_new_n3983_; 
wire u0__abc_74894_new_n3984_; 
wire u0__abc_74894_new_n3985_; 
wire u0__abc_74894_new_n3986_; 
wire u0__abc_74894_new_n3987_; 
wire u0__abc_74894_new_n3988_; 
wire u0__abc_74894_new_n3989_; 
wire u0__abc_74894_new_n3990_; 
wire u0__abc_74894_new_n3991_; 
wire u0__abc_74894_new_n3992_; 
wire u0__abc_74894_new_n3993_; 
wire u0__abc_74894_new_n3995_; 
wire u0__abc_74894_new_n3996_; 
wire u0__abc_74894_new_n3997_; 
wire u0__abc_74894_new_n3998_; 
wire u0__abc_74894_new_n3999_; 
wire u0__abc_74894_new_n4000_; 
wire u0__abc_74894_new_n4001_; 
wire u0__abc_74894_new_n4002_; 
wire u0__abc_74894_new_n4003_; 
wire u0__abc_74894_new_n4004_; 
wire u0__abc_74894_new_n4005_; 
wire u0__abc_74894_new_n4006_; 
wire u0__abc_74894_new_n4007_; 
wire u0__abc_74894_new_n4008_; 
wire u0__abc_74894_new_n4009_; 
wire u0__abc_74894_new_n4010_; 
wire u0__abc_74894_new_n4011_; 
wire u0__abc_74894_new_n4012_; 
wire u0__abc_74894_new_n4013_; 
wire u0__abc_74894_new_n4014_; 
wire u0__abc_74894_new_n4015_; 
wire u0__abc_74894_new_n4017_; 
wire u0__abc_74894_new_n4018_; 
wire u0__abc_74894_new_n4019_; 
wire u0__abc_74894_new_n4020_; 
wire u0__abc_74894_new_n4021_; 
wire u0__abc_74894_new_n4022_; 
wire u0__abc_74894_new_n4023_; 
wire u0__abc_74894_new_n4024_; 
wire u0__abc_74894_new_n4025_; 
wire u0__abc_74894_new_n4026_; 
wire u0__abc_74894_new_n4027_; 
wire u0__abc_74894_new_n4028_; 
wire u0__abc_74894_new_n4029_; 
wire u0__abc_74894_new_n4030_; 
wire u0__abc_74894_new_n4031_; 
wire u0__abc_74894_new_n4032_; 
wire u0__abc_74894_new_n4033_; 
wire u0__abc_74894_new_n4034_; 
wire u0__abc_74894_new_n4035_; 
wire u0__abc_74894_new_n4036_; 
wire u0__abc_74894_new_n4037_; 
wire u0__abc_74894_new_n4039_; 
wire u0__abc_74894_new_n4040_; 
wire u0__abc_74894_new_n4041_; 
wire u0__abc_74894_new_n4042_; 
wire u0__abc_74894_new_n4043_; 
wire u0__abc_74894_new_n4044_; 
wire u0__abc_74894_new_n4045_; 
wire u0__abc_74894_new_n4046_; 
wire u0__abc_74894_new_n4047_; 
wire u0__abc_74894_new_n4048_; 
wire u0__abc_74894_new_n4049_; 
wire u0__abc_74894_new_n4050_; 
wire u0__abc_74894_new_n4051_; 
wire u0__abc_74894_new_n4052_; 
wire u0__abc_74894_new_n4053_; 
wire u0__abc_74894_new_n4054_; 
wire u0__abc_74894_new_n4055_; 
wire u0__abc_74894_new_n4056_; 
wire u0__abc_74894_new_n4057_; 
wire u0__abc_74894_new_n4058_; 
wire u0__abc_74894_new_n4059_; 
wire u0__abc_74894_new_n4061_; 
wire u0__abc_74894_new_n4062_; 
wire u0__abc_74894_new_n4063_; 
wire u0__abc_74894_new_n4064_; 
wire u0__abc_74894_new_n4065_; 
wire u0__abc_74894_new_n4066_; 
wire u0__abc_74894_new_n4067_; 
wire u0__abc_74894_new_n4068_; 
wire u0__abc_74894_new_n4069_; 
wire u0__abc_74894_new_n4070_; 
wire u0__abc_74894_new_n4071_; 
wire u0__abc_74894_new_n4072_; 
wire u0__abc_74894_new_n4073_; 
wire u0__abc_74894_new_n4074_; 
wire u0__abc_74894_new_n4075_; 
wire u0__abc_74894_new_n4076_; 
wire u0__abc_74894_new_n4077_; 
wire u0__abc_74894_new_n4078_; 
wire u0__abc_74894_new_n4079_; 
wire u0__abc_74894_new_n4081_; 
wire u0__abc_74894_new_n4082_; 
wire u0__abc_74894_new_n4083_; 
wire u0__abc_74894_new_n4084_; 
wire u0__abc_74894_new_n4085_; 
wire u0__abc_74894_new_n4086_; 
wire u0__abc_74894_new_n4087_; 
wire u0__abc_74894_new_n4088_; 
wire u0__abc_74894_new_n4089_; 
wire u0__abc_74894_new_n4090_; 
wire u0__abc_74894_new_n4091_; 
wire u0__abc_74894_new_n4092_; 
wire u0__abc_74894_new_n4093_; 
wire u0__abc_74894_new_n4094_; 
wire u0__abc_74894_new_n4095_; 
wire u0__abc_74894_new_n4096_; 
wire u0__abc_74894_new_n4097_; 
wire u0__abc_74894_new_n4098_; 
wire u0__abc_74894_new_n4099_; 
wire u0__abc_74894_new_n4100_; 
wire u0__abc_74894_new_n4101_; 
wire u0__abc_74894_new_n4103_; 
wire u0__abc_74894_new_n4104_; 
wire u0__abc_74894_new_n4105_; 
wire u0__abc_74894_new_n4106_; 
wire u0__abc_74894_new_n4107_; 
wire u0__abc_74894_new_n4108_; 
wire u0__abc_74894_new_n4109_; 
wire u0__abc_74894_new_n4110_; 
wire u0__abc_74894_new_n4111_; 
wire u0__abc_74894_new_n4112_; 
wire u0__abc_74894_new_n4113_; 
wire u0__abc_74894_new_n4114_; 
wire u0__abc_74894_new_n4115_; 
wire u0__abc_74894_new_n4116_; 
wire u0__abc_74894_new_n4117_; 
wire u0__abc_74894_new_n4118_; 
wire u0__abc_74894_new_n4119_; 
wire u0__abc_74894_new_n4120_; 
wire u0__abc_74894_new_n4121_; 
wire u0__abc_74894_new_n4122_; 
wire u0__abc_74894_new_n4123_; 
wire u0__abc_74894_new_n4125_; 
wire u0__abc_74894_new_n4126_; 
wire u0__abc_74894_new_n4127_; 
wire u0__abc_74894_new_n4128_; 
wire u0__abc_74894_new_n4129_; 
wire u0__abc_74894_new_n4130_; 
wire u0__abc_74894_new_n4131_; 
wire u0__abc_74894_new_n4132_; 
wire u0__abc_74894_new_n4133_; 
wire u0__abc_74894_new_n4134_; 
wire u0__abc_74894_new_n4135_; 
wire u0__abc_74894_new_n4136_; 
wire u0__abc_74894_new_n4137_; 
wire u0__abc_74894_new_n4138_; 
wire u0__abc_74894_new_n4139_; 
wire u0__abc_74894_new_n4140_; 
wire u0__abc_74894_new_n4141_; 
wire u0__abc_74894_new_n4142_; 
wire u0__abc_74894_new_n4143_; 
wire u0__abc_74894_new_n4144_; 
wire u0__abc_74894_new_n4145_; 
wire u0__abc_74894_new_n4147_; 
wire u0__abc_74894_new_n4148_; 
wire u0__abc_74894_new_n4149_; 
wire u0__abc_74894_new_n4150_; 
wire u0__abc_74894_new_n4151_; 
wire u0__abc_74894_new_n4152_; 
wire u0__abc_74894_new_n4153_; 
wire u0__abc_74894_new_n4154_; 
wire u0__abc_74894_new_n4155_; 
wire u0__abc_74894_new_n4156_; 
wire u0__abc_74894_new_n4157_; 
wire u0__abc_74894_new_n4158_; 
wire u0__abc_74894_new_n4159_; 
wire u0__abc_74894_new_n4160_; 
wire u0__abc_74894_new_n4161_; 
wire u0__abc_74894_new_n4162_; 
wire u0__abc_74894_new_n4163_; 
wire u0__abc_74894_new_n4164_; 
wire u0__abc_74894_new_n4166_; 
wire u0__abc_74894_new_n4167_; 
wire u0__abc_74894_new_n4168_; 
wire u0__abc_74894_new_n4169_; 
wire u0__abc_74894_new_n4170_; 
wire u0__abc_74894_new_n4171_; 
wire u0__abc_74894_new_n4172_; 
wire u0__abc_74894_new_n4173_; 
wire u0__abc_74894_new_n4174_; 
wire u0__abc_74894_new_n4175_; 
wire u0__abc_74894_new_n4176_; 
wire u0__abc_74894_new_n4177_; 
wire u0__abc_74894_new_n4178_; 
wire u0__abc_74894_new_n4179_; 
wire u0__abc_74894_new_n4180_; 
wire u0__abc_74894_new_n4181_; 
wire u0__abc_74894_new_n4182_; 
wire u0__abc_74894_new_n4183_; 
wire u0__abc_74894_new_n4184_; 
wire u0__abc_74894_new_n4185_; 
wire u0__abc_74894_new_n4186_; 
wire u0__abc_74894_new_n4187_; 
wire u0__abc_74894_new_n4189_; 
wire u0__abc_74894_new_n4190_; 
wire u0__abc_74894_new_n4191_; 
wire u0__abc_74894_new_n4192_; 
wire u0__abc_74894_new_n4193_; 
wire u0__abc_74894_new_n4194_; 
wire u0__abc_74894_new_n4195_; 
wire u0__abc_74894_new_n4196_; 
wire u0__abc_74894_new_n4197_; 
wire u0__abc_74894_new_n4198_; 
wire u0__abc_74894_new_n4199_; 
wire u0__abc_74894_new_n4200_; 
wire u0__abc_74894_new_n4201_; 
wire u0__abc_74894_new_n4202_; 
wire u0__abc_74894_new_n4203_; 
wire u0__abc_74894_new_n4204_; 
wire u0__abc_74894_new_n4205_; 
wire u0__abc_74894_new_n4206_; 
wire u0__abc_74894_new_n4208_; 
wire u0__abc_74894_new_n4209_; 
wire u0__abc_74894_new_n4210_; 
wire u0__abc_74894_new_n4211_; 
wire u0__abc_74894_new_n4212_; 
wire u0__abc_74894_new_n4213_; 
wire u0__abc_74894_new_n4214_; 
wire u0__abc_74894_new_n4215_; 
wire u0__abc_74894_new_n4216_; 
wire u0__abc_74894_new_n4217_; 
wire u0__abc_74894_new_n4218_; 
wire u0__abc_74894_new_n4219_; 
wire u0__abc_74894_new_n4220_; 
wire u0__abc_74894_new_n4221_; 
wire u0__abc_74894_new_n4222_; 
wire u0__abc_74894_new_n4223_; 
wire u0__abc_74894_new_n4224_; 
wire u0__abc_74894_new_n4225_; 
wire u0__abc_74894_new_n4226_; 
wire u0__abc_74894_new_n4228_; 
wire u0__abc_74894_new_n4229_; 
wire u0__abc_74894_new_n4230_; 
wire u0__abc_74894_new_n4231_; 
wire u0__abc_74894_new_n4232_; 
wire u0__abc_74894_new_n4233_; 
wire u0__abc_74894_new_n4234_; 
wire u0__abc_74894_new_n4235_; 
wire u0__abc_74894_new_n4236_; 
wire u0__abc_74894_new_n4237_; 
wire u0__abc_74894_new_n4238_; 
wire u0__abc_74894_new_n4239_; 
wire u0__abc_74894_new_n4240_; 
wire u0__abc_74894_new_n4241_; 
wire u0__abc_74894_new_n4242_; 
wire u0__abc_74894_new_n4243_; 
wire u0__abc_74894_new_n4244_; 
wire u0__abc_74894_new_n4245_; 
wire u0__abc_74894_new_n4246_; 
wire u0__abc_74894_new_n4247_; 
wire u0__abc_74894_new_n4248_; 
wire u0__abc_74894_new_n4249_; 
wire u0__abc_74894_new_n4250_; 
wire u0__abc_74894_new_n4251_; 
wire u0__abc_74894_new_n4252_; 
wire u0__abc_74894_new_n4254_; 
wire u0__abc_74894_new_n4255_; 
wire u0__abc_74894_new_n4256_; 
wire u0__abc_74894_new_n4257_; 
wire u0__abc_74894_new_n4258_; 
wire u0__abc_74894_new_n4259_; 
wire u0__abc_74894_new_n4260_; 
wire u0__abc_74894_new_n4261_; 
wire u0__abc_74894_new_n4262_; 
wire u0__abc_74894_new_n4263_; 
wire u0__abc_74894_new_n4264_; 
wire u0__abc_74894_new_n4265_; 
wire u0__abc_74894_new_n4266_; 
wire u0__abc_74894_new_n4267_; 
wire u0__abc_74894_new_n4268_; 
wire u0__abc_74894_new_n4269_; 
wire u0__abc_74894_new_n4270_; 
wire u0__abc_74894_new_n4271_; 
wire u0__abc_74894_new_n4272_; 
wire u0__abc_74894_new_n4273_; 
wire u0__abc_74894_new_n4274_; 
wire u0__abc_74894_new_n4275_; 
wire u0__abc_74894_new_n4276_; 
wire u0__abc_74894_new_n4277_; 
wire u0__abc_74894_new_n4278_; 
wire u0__abc_74894_new_n4280_; 
wire u0__abc_74894_new_n4281_; 
wire u0__abc_74894_new_n4282_; 
wire u0__abc_74894_new_n4283_; 
wire u0__abc_74894_new_n4284_; 
wire u0__abc_74894_new_n4285_; 
wire u0__abc_74894_new_n4286_; 
wire u0__abc_74894_new_n4287_; 
wire u0__abc_74894_new_n4288_; 
wire u0__abc_74894_new_n4289_; 
wire u0__abc_74894_new_n4290_; 
wire u0__abc_74894_new_n4291_; 
wire u0__abc_74894_new_n4292_; 
wire u0__abc_74894_new_n4293_; 
wire u0__abc_74894_new_n4294_; 
wire u0__abc_74894_new_n4295_; 
wire u0__abc_74894_new_n4296_; 
wire u0__abc_74894_new_n4297_; 
wire u0__abc_74894_new_n4298_; 
wire u0__abc_74894_new_n4299_; 
wire u0__abc_74894_new_n4300_; 
wire u0__abc_74894_new_n4301_; 
wire u0__abc_74894_new_n4302_; 
wire u0__abc_74894_new_n4303_; 
wire u0__abc_74894_new_n4304_; 
wire u0__abc_74894_new_n4306_; 
wire u0__abc_74894_new_n4307_; 
wire u0__abc_74894_new_n4308_; 
wire u0__abc_74894_new_n4309_; 
wire u0__abc_74894_new_n4310_; 
wire u0__abc_74894_new_n4311_; 
wire u0__abc_74894_new_n4312_; 
wire u0__abc_74894_new_n4313_; 
wire u0__abc_74894_new_n4314_; 
wire u0__abc_74894_new_n4315_; 
wire u0__abc_74894_new_n4316_; 
wire u0__abc_74894_new_n4317_; 
wire u0__abc_74894_new_n4318_; 
wire u0__abc_74894_new_n4319_; 
wire u0__abc_74894_new_n4320_; 
wire u0__abc_74894_new_n4321_; 
wire u0__abc_74894_new_n4322_; 
wire u0__abc_74894_new_n4323_; 
wire u0__abc_74894_new_n4324_; 
wire u0__abc_74894_new_n4325_; 
wire u0__abc_74894_new_n4326_; 
wire u0__abc_74894_new_n4327_; 
wire u0__abc_74894_new_n4328_; 
wire u0__abc_74894_new_n4329_; 
wire u0__abc_74894_new_n4330_; 
wire u0__abc_74894_new_n4331_; 
wire u0__abc_74894_new_n4333_; 
wire u0__abc_74894_new_n4334_; 
wire u0__abc_74894_new_n4335_; 
wire u0__abc_74894_new_n4336_; 
wire u0__abc_74894_new_n4337_; 
wire u0__abc_74894_new_n4338_; 
wire u0__abc_74894_new_n4339_; 
wire u0__abc_74894_new_n4340_; 
wire u0__abc_74894_new_n4341_; 
wire u0__abc_74894_new_n4342_; 
wire u0__abc_74894_new_n4343_; 
wire u0__abc_74894_new_n4344_; 
wire u0__abc_74894_new_n4345_; 
wire u0__abc_74894_new_n4346_; 
wire u0__abc_74894_new_n4347_; 
wire u0__abc_74894_new_n4348_; 
wire u0__abc_74894_new_n4349_; 
wire u0__abc_74894_new_n4350_; 
wire u0__abc_74894_new_n4351_; 
wire u0__abc_74894_new_n4352_; 
wire u0__abc_74894_new_n4353_; 
wire u0__abc_74894_new_n4354_; 
wire u0__abc_74894_new_n4355_; 
wire u0__abc_74894_new_n4356_; 
wire u0__abc_74894_new_n4357_; 
wire u0__abc_74894_new_n4359_; 
wire u0__abc_74894_new_n4360_; 
wire u0__abc_74894_new_n4361_; 
wire u0__abc_74894_new_n4362_; 
wire u0__abc_74894_new_n4363_; 
wire u0__abc_74894_new_n4364_; 
wire u0__abc_74894_new_n4365_; 
wire u0__abc_74894_new_n4366_; 
wire u0__abc_74894_new_n4367_; 
wire u0__abc_74894_new_n4368_; 
wire u0__abc_74894_new_n4369_; 
wire u0__abc_74894_new_n4370_; 
wire u0__abc_74894_new_n4371_; 
wire u0__abc_74894_new_n4372_; 
wire u0__abc_74894_new_n4373_; 
wire u0__abc_74894_new_n4374_; 
wire u0__abc_74894_new_n4375_; 
wire u0__abc_74894_new_n4376_; 
wire u0__abc_74894_new_n4377_; 
wire u0__abc_74894_new_n4378_; 
wire u0__abc_74894_new_n4379_; 
wire u0__abc_74894_new_n4380_; 
wire u0__abc_74894_new_n4381_; 
wire u0__abc_74894_new_n4383_; 
wire u0__abc_74894_new_n4384_; 
wire u0__abc_74894_new_n4385_; 
wire u0__abc_74894_new_n4386_; 
wire u0__abc_74894_new_n4387_; 
wire u0__abc_74894_new_n4388_; 
wire u0__abc_74894_new_n4389_; 
wire u0__abc_74894_new_n4390_; 
wire u0__abc_74894_new_n4391_; 
wire u0__abc_74894_new_n4392_; 
wire u0__abc_74894_new_n4393_; 
wire u0__abc_74894_new_n4394_; 
wire u0__abc_74894_new_n4395_; 
wire u0__abc_74894_new_n4396_; 
wire u0__abc_74894_new_n4397_; 
wire u0__abc_74894_new_n4398_; 
wire u0__abc_74894_new_n4399_; 
wire u0__abc_74894_new_n4400_; 
wire u0__abc_74894_new_n4401_; 
wire u0__abc_74894_new_n4402_; 
wire u0__abc_74894_new_n4403_; 
wire u0__abc_74894_new_n4404_; 
wire u0__abc_74894_new_n4405_; 
wire u0__abc_74894_new_n4407_; 
wire u0__abc_74894_new_n4408_; 
wire u0__abc_74894_new_n4409_; 
wire u0__abc_74894_new_n4410_; 
wire u0__abc_74894_new_n4411_; 
wire u0__abc_74894_new_n4412_; 
wire u0__abc_74894_new_n4413_; 
wire u0__abc_74894_new_n4414_; 
wire u0__abc_74894_new_n4415_; 
wire u0__abc_74894_new_n4416_; 
wire u0__abc_74894_new_n4417_; 
wire u0__abc_74894_new_n4418_; 
wire u0__abc_74894_new_n4419_; 
wire u0__abc_74894_new_n4420_; 
wire u0__abc_74894_new_n4421_; 
wire u0__abc_74894_new_n4422_; 
wire u0__abc_74894_new_n4423_; 
wire u0__abc_74894_new_n4424_; 
wire u0__abc_74894_new_n4425_; 
wire u0__abc_74894_new_n4426_; 
wire u0__abc_74894_new_n4427_; 
wire u0__abc_74894_new_n4428_; 
wire u0__abc_74894_new_n4429_; 
wire u0__abc_74894_new_n4431_; 
wire u0__abc_74894_new_n4432_; 
wire u0__abc_74894_new_n4433_; 
wire u0__abc_74894_new_n4437_; 
wire u0__abc_74894_new_n4438_; 
wire u0__abc_74894_new_n4440_; 
wire u0__abc_74894_new_n4441_; 
wire u0__abc_74894_new_n4443_; 
wire u0__abc_74894_new_n4444_; 
wire u0__abc_74894_new_n4446_; 
wire u0__abc_74894_new_n4447_; 
wire u0__abc_74894_new_n4449_; 
wire u0__abc_74894_new_n4450_; 
wire u0__abc_74894_new_n4452_; 
wire u0__abc_74894_new_n4453_; 
wire u0__abc_74894_new_n4455_; 
wire u0__abc_74894_new_n4456_; 
wire u0__abc_74894_new_n4458_; 
wire u0__abc_74894_new_n4459_; 
wire u0__abc_74894_new_n4461_; 
wire u0__abc_74894_new_n4462_; 
wire u0__abc_74894_new_n4463_; 
wire u0__abc_74894_new_n4464_; 
wire u0__abc_74894_new_n4465_; 
wire u0__abc_74894_new_n4467_; 
wire u0__abc_74894_new_n4468_; 
wire u0__abc_74894_new_n4469_; 
wire u0__abc_74894_new_n4470_; 
wire u0__abc_74894_new_n4471_; 
wire u0__abc_74894_new_n4473_; 
wire u0__abc_74894_new_n4474_; 
wire u0__abc_74894_new_n4475_; 
wire u0__abc_74894_new_n4476_; 
wire u0_cs0; 
wire u0_cs1; 
wire u0_csc0_0_; 
wire u0_csc0_10_; 
wire u0_csc0_11_; 
wire u0_csc0_12_; 
wire u0_csc0_13_; 
wire u0_csc0_14_; 
wire u0_csc0_15_; 
wire u0_csc0_16_; 
wire u0_csc0_17_; 
wire u0_csc0_18_; 
wire u0_csc0_19_; 
wire u0_csc0_1_; 
wire u0_csc0_20_; 
wire u0_csc0_21_; 
wire u0_csc0_22_; 
wire u0_csc0_23_; 
wire u0_csc0_24_; 
wire u0_csc0_25_; 
wire u0_csc0_26_; 
wire u0_csc0_27_; 
wire u0_csc0_28_; 
wire u0_csc0_29_; 
wire u0_csc0_2_; 
wire u0_csc0_30_; 
wire u0_csc0_31_; 
wire u0_csc0_3_; 
wire u0_csc0_4_; 
wire u0_csc0_5_; 
wire u0_csc0_6_; 
wire u0_csc0_7_; 
wire u0_csc0_8_; 
wire u0_csc0_9_; 
wire u0_csc1_0_; 
wire u0_csc1_10_; 
wire u0_csc1_11_; 
wire u0_csc1_12_; 
wire u0_csc1_13_; 
wire u0_csc1_14_; 
wire u0_csc1_15_; 
wire u0_csc1_16_; 
wire u0_csc1_17_; 
wire u0_csc1_18_; 
wire u0_csc1_19_; 
wire u0_csc1_1_; 
wire u0_csc1_20_; 
wire u0_csc1_21_; 
wire u0_csc1_22_; 
wire u0_csc1_23_; 
wire u0_csc1_24_; 
wire u0_csc1_25_; 
wire u0_csc1_26_; 
wire u0_csc1_27_; 
wire u0_csc1_28_; 
wire u0_csc1_29_; 
wire u0_csc1_2_; 
wire u0_csc1_30_; 
wire u0_csc1_31_; 
wire u0_csc1_3_; 
wire u0_csc1_4_; 
wire u0_csc1_5_; 
wire u0_csc1_6_; 
wire u0_csc1_7_; 
wire u0_csc1_8_; 
wire u0_csc1_9_; 
wire u0_csc_mask_0_; 
wire u0_csc_mask_10_; 
wire u0_csc_mask_1_; 
wire u0_csc_mask_2_; 
wire u0_csc_mask_3_; 
wire u0_csc_mask_4_; 
wire u0_csc_mask_5_; 
wire u0_csc_mask_6_; 
wire u0_csc_mask_7_; 
wire u0_csc_mask_8_; 
wire u0_csc_mask_9_; 
wire u0_csr_0_; 
wire u0_csr_3_; 
wire u0_csr_4_; 
wire u0_csr_5_; 
wire u0_csr_6_; 
wire u0_csr_7_; 
wire u0_init_ack0; 
wire u0_init_ack1; 
wire u0_init_ack_r; 
wire u0_init_req0; 
wire u0_init_req1; 
wire u0_lmr_ack0; 
wire u0_lmr_ack1; 
wire u0_lmr_ack_r; 
wire u0_lmr_req0; 
wire u0_lmr_req1; 
wire u0_rf_we; 
wire u0_rst_r2; 
wire u0_rst_r3; 
wire u0_sreq_cs_le; 
wire u0_tms0_0_; 
wire u0_tms0_10_; 
wire u0_tms0_11_; 
wire u0_tms0_12_; 
wire u0_tms0_13_; 
wire u0_tms0_14_; 
wire u0_tms0_15_; 
wire u0_tms0_16_; 
wire u0_tms0_17_; 
wire u0_tms0_18_; 
wire u0_tms0_19_; 
wire u0_tms0_1_; 
wire u0_tms0_20_; 
wire u0_tms0_21_; 
wire u0_tms0_22_; 
wire u0_tms0_23_; 
wire u0_tms0_24_; 
wire u0_tms0_25_; 
wire u0_tms0_26_; 
wire u0_tms0_27_; 
wire u0_tms0_28_; 
wire u0_tms0_29_; 
wire u0_tms0_2_; 
wire u0_tms0_30_; 
wire u0_tms0_31_; 
wire u0_tms0_3_; 
wire u0_tms0_4_; 
wire u0_tms0_5_; 
wire u0_tms0_6_; 
wire u0_tms0_7_; 
wire u0_tms0_8_; 
wire u0_tms0_9_; 
wire u0_tms1_0_; 
wire u0_tms1_10_; 
wire u0_tms1_11_; 
wire u0_tms1_12_; 
wire u0_tms1_13_; 
wire u0_tms1_14_; 
wire u0_tms1_15_; 
wire u0_tms1_16_; 
wire u0_tms1_17_; 
wire u0_tms1_18_; 
wire u0_tms1_19_; 
wire u0_tms1_1_; 
wire u0_tms1_20_; 
wire u0_tms1_21_; 
wire u0_tms1_22_; 
wire u0_tms1_23_; 
wire u0_tms1_24_; 
wire u0_tms1_25_; 
wire u0_tms1_26_; 
wire u0_tms1_27_; 
wire u0_tms1_28_; 
wire u0_tms1_29_; 
wire u0_tms1_2_; 
wire u0_tms1_30_; 
wire u0_tms1_31_; 
wire u0_tms1_3_; 
wire u0_tms1_4_; 
wire u0_tms1_5_; 
wire u0_tms1_6_; 
wire u0_tms1_7_; 
wire u0_tms1_8_; 
wire u0_tms1_9_; 
wire u0_u0__0csc_31_0__0_; 
wire u0_u0__0csc_31_0__10_; 
wire u0_u0__0csc_31_0__11_; 
wire u0_u0__0csc_31_0__12_; 
wire u0_u0__0csc_31_0__13_; 
wire u0_u0__0csc_31_0__14_; 
wire u0_u0__0csc_31_0__15_; 
wire u0_u0__0csc_31_0__16_; 
wire u0_u0__0csc_31_0__17_; 
wire u0_u0__0csc_31_0__18_; 
wire u0_u0__0csc_31_0__19_; 
wire u0_u0__0csc_31_0__1_; 
wire u0_u0__0csc_31_0__20_; 
wire u0_u0__0csc_31_0__21_; 
wire u0_u0__0csc_31_0__22_; 
wire u0_u0__0csc_31_0__23_; 
wire u0_u0__0csc_31_0__24_; 
wire u0_u0__0csc_31_0__25_; 
wire u0_u0__0csc_31_0__26_; 
wire u0_u0__0csc_31_0__27_; 
wire u0_u0__0csc_31_0__28_; 
wire u0_u0__0csc_31_0__29_; 
wire u0_u0__0csc_31_0__2_; 
wire u0_u0__0csc_31_0__30_; 
wire u0_u0__0csc_31_0__31_; 
wire u0_u0__0csc_31_0__3_; 
wire u0_u0__0csc_31_0__4_; 
wire u0_u0__0csc_31_0__5_; 
wire u0_u0__0csc_31_0__6_; 
wire u0_u0__0csc_31_0__7_; 
wire u0_u0__0csc_31_0__8_; 
wire u0_u0__0csc_31_0__9_; 
wire u0_u0__0init_req_0_0_; 
wire u0_u0__0init_req_we_0_0_; 
wire u0_u0__0inited_0_0_; 
wire u0_u0__0lmr_req_0_0_; 
wire u0_u0__0lmr_req_we_0_0_; 
wire u0_u0__0tms_31_0__0_; 
wire u0_u0__0tms_31_0__10_; 
wire u0_u0__0tms_31_0__11_; 
wire u0_u0__0tms_31_0__12_; 
wire u0_u0__0tms_31_0__13_; 
wire u0_u0__0tms_31_0__14_; 
wire u0_u0__0tms_31_0__15_; 
wire u0_u0__0tms_31_0__16_; 
wire u0_u0__0tms_31_0__17_; 
wire u0_u0__0tms_31_0__18_; 
wire u0_u0__0tms_31_0__19_; 
wire u0_u0__0tms_31_0__1_; 
wire u0_u0__0tms_31_0__20_; 
wire u0_u0__0tms_31_0__21_; 
wire u0_u0__0tms_31_0__22_; 
wire u0_u0__0tms_31_0__23_; 
wire u0_u0__0tms_31_0__24_; 
wire u0_u0__0tms_31_0__25_; 
wire u0_u0__0tms_31_0__26_; 
wire u0_u0__0tms_31_0__27_; 
wire u0_u0__0tms_31_0__28_; 
wire u0_u0__0tms_31_0__29_; 
wire u0_u0__0tms_31_0__2_; 
wire u0_u0__0tms_31_0__30_; 
wire u0_u0__0tms_31_0__31_; 
wire u0_u0__0tms_31_0__3_; 
wire u0_u0__0tms_31_0__4_; 
wire u0_u0__0tms_31_0__5_; 
wire u0_u0__0tms_31_0__6_; 
wire u0_u0__0tms_31_0__7_; 
wire u0_u0__0tms_31_0__8_; 
wire u0_u0__0tms_31_0__9_; 
wire u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494; 
wire u0_u0__abc_72207_new_n205_; 
wire u0_u0__abc_72207_new_n206_; 
wire u0_u0__abc_72207_new_n207_; 
wire u0_u0__abc_72207_new_n208_; 
wire u0_u0__abc_72207_new_n209_; 
wire u0_u0__abc_72207_new_n210_; 
wire u0_u0__abc_72207_new_n211_; 
wire u0_u0__abc_72207_new_n212_; 
wire u0_u0__abc_72207_new_n214_; 
wire u0_u0__abc_72207_new_n215_; 
wire u0_u0__abc_72207_new_n216_; 
wire u0_u0__abc_72207_new_n217_; 
wire u0_u0__abc_72207_new_n218_; 
wire u0_u0__abc_72207_new_n219_; 
wire u0_u0__abc_72207_new_n220_; 
wire u0_u0__abc_72207_new_n222_; 
wire u0_u0__abc_72207_new_n223_; 
wire u0_u0__abc_72207_new_n225_; 
wire u0_u0__abc_72207_new_n226_; 
wire u0_u0__abc_72207_new_n228_; 
wire u0_u0__abc_72207_new_n229_; 
wire u0_u0__abc_72207_new_n231_; 
wire u0_u0__abc_72207_new_n232_; 
wire u0_u0__abc_72207_new_n234_; 
wire u0_u0__abc_72207_new_n235_; 
wire u0_u0__abc_72207_new_n237_; 
wire u0_u0__abc_72207_new_n238_; 
wire u0_u0__abc_72207_new_n240_; 
wire u0_u0__abc_72207_new_n241_; 
wire u0_u0__abc_72207_new_n243_; 
wire u0_u0__abc_72207_new_n244_; 
wire u0_u0__abc_72207_new_n246_; 
wire u0_u0__abc_72207_new_n247_; 
wire u0_u0__abc_72207_new_n249_; 
wire u0_u0__abc_72207_new_n250_; 
wire u0_u0__abc_72207_new_n252_; 
wire u0_u0__abc_72207_new_n253_; 
wire u0_u0__abc_72207_new_n255_; 
wire u0_u0__abc_72207_new_n256_; 
wire u0_u0__abc_72207_new_n258_; 
wire u0_u0__abc_72207_new_n259_; 
wire u0_u0__abc_72207_new_n261_; 
wire u0_u0__abc_72207_new_n262_; 
wire u0_u0__abc_72207_new_n264_; 
wire u0_u0__abc_72207_new_n265_; 
wire u0_u0__abc_72207_new_n267_; 
wire u0_u0__abc_72207_new_n268_; 
wire u0_u0__abc_72207_new_n270_; 
wire u0_u0__abc_72207_new_n271_; 
wire u0_u0__abc_72207_new_n273_; 
wire u0_u0__abc_72207_new_n274_; 
wire u0_u0__abc_72207_new_n276_; 
wire u0_u0__abc_72207_new_n277_; 
wire u0_u0__abc_72207_new_n279_; 
wire u0_u0__abc_72207_new_n280_; 
wire u0_u0__abc_72207_new_n282_; 
wire u0_u0__abc_72207_new_n283_; 
wire u0_u0__abc_72207_new_n285_; 
wire u0_u0__abc_72207_new_n286_; 
wire u0_u0__abc_72207_new_n288_; 
wire u0_u0__abc_72207_new_n289_; 
wire u0_u0__abc_72207_new_n291_; 
wire u0_u0__abc_72207_new_n292_; 
wire u0_u0__abc_72207_new_n294_; 
wire u0_u0__abc_72207_new_n295_; 
wire u0_u0__abc_72207_new_n297_; 
wire u0_u0__abc_72207_new_n298_; 
wire u0_u0__abc_72207_new_n300_; 
wire u0_u0__abc_72207_new_n301_; 
wire u0_u0__abc_72207_new_n303_; 
wire u0_u0__abc_72207_new_n304_; 
wire u0_u0__abc_72207_new_n306_; 
wire u0_u0__abc_72207_new_n307_; 
wire u0_u0__abc_72207_new_n309_; 
wire u0_u0__abc_72207_new_n310_; 
wire u0_u0__abc_72207_new_n312_; 
wire u0_u0__abc_72207_new_n313_; 
wire u0_u0__abc_72207_new_n315_; 
wire u0_u0__abc_72207_new_n316_; 
wire u0_u0__abc_72207_new_n318_; 
wire u0_u0__abc_72207_new_n319_; 
wire u0_u0__abc_72207_new_n320_; 
wire u0_u0__abc_72207_new_n321_; 
wire u0_u0__abc_72207_new_n322_; 
wire u0_u0__abc_72207_new_n324_; 
wire u0_u0__abc_72207_new_n325_; 
wire u0_u0__abc_72207_new_n326_; 
wire u0_u0__abc_72207_new_n327_; 
wire u0_u0__abc_72207_new_n328_; 
wire u0_u0__abc_72207_new_n329_; 
wire u0_u0__abc_72207_new_n330_; 
wire u0_u0__abc_72207_new_n332_; 
wire u0_u0__abc_72207_new_n333_; 
wire u0_u0__abc_72207_new_n334_; 
wire u0_u0__abc_72207_new_n336_; 
wire u0_u0__abc_72207_new_n337_; 
wire u0_u0__abc_72207_new_n338_; 
wire u0_u0__abc_72207_new_n340_; 
wire u0_u0__abc_72207_new_n342_; 
wire u0_u0__abc_72207_new_n343_; 
wire u0_u0__abc_72207_new_n344_; 
wire u0_u0__abc_72207_new_n345_; 
wire u0_u0__abc_72207_new_n346_; 
wire u0_u0__abc_72207_new_n347_; 
wire u0_u0__abc_72207_new_n349_; 
wire u0_u0__abc_72207_new_n350_; 
wire u0_u0__abc_72207_new_n351_; 
wire u0_u0__abc_72207_new_n352_; 
wire u0_u0__abc_72207_new_n353_; 
wire u0_u0__abc_72207_new_n354_; 
wire u0_u0__abc_72207_new_n356_; 
wire u0_u0__abc_72207_new_n357_; 
wire u0_u0__abc_72207_new_n359_; 
wire u0_u0__abc_72207_new_n360_; 
wire u0_u0__abc_72207_new_n362_; 
wire u0_u0__abc_72207_new_n363_; 
wire u0_u0__abc_72207_new_n365_; 
wire u0_u0__abc_72207_new_n366_; 
wire u0_u0__abc_72207_new_n368_; 
wire u0_u0__abc_72207_new_n369_; 
wire u0_u0__abc_72207_new_n371_; 
wire u0_u0__abc_72207_new_n372_; 
wire u0_u0__abc_72207_new_n374_; 
wire u0_u0__abc_72207_new_n375_; 
wire u0_u0__abc_72207_new_n377_; 
wire u0_u0__abc_72207_new_n378_; 
wire u0_u0__abc_72207_new_n380_; 
wire u0_u0__abc_72207_new_n381_; 
wire u0_u0__abc_72207_new_n383_; 
wire u0_u0__abc_72207_new_n384_; 
wire u0_u0__abc_72207_new_n386_; 
wire u0_u0__abc_72207_new_n387_; 
wire u0_u0__abc_72207_new_n389_; 
wire u0_u0__abc_72207_new_n390_; 
wire u0_u0__abc_72207_new_n392_; 
wire u0_u0__abc_72207_new_n393_; 
wire u0_u0__abc_72207_new_n395_; 
wire u0_u0__abc_72207_new_n396_; 
wire u0_u0__abc_72207_new_n398_; 
wire u0_u0__abc_72207_new_n399_; 
wire u0_u0__abc_72207_new_n401_; 
wire u0_u0__abc_72207_new_n402_; 
wire u0_u0__abc_72207_new_n404_; 
wire u0_u0__abc_72207_new_n405_; 
wire u0_u0__abc_72207_new_n407_; 
wire u0_u0__abc_72207_new_n408_; 
wire u0_u0__abc_72207_new_n410_; 
wire u0_u0__abc_72207_new_n411_; 
wire u0_u0__abc_72207_new_n413_; 
wire u0_u0__abc_72207_new_n414_; 
wire u0_u0__abc_72207_new_n416_; 
wire u0_u0__abc_72207_new_n417_; 
wire u0_u0__abc_72207_new_n419_; 
wire u0_u0__abc_72207_new_n420_; 
wire u0_u0__abc_72207_new_n422_; 
wire u0_u0__abc_72207_new_n423_; 
wire u0_u0__abc_72207_new_n425_; 
wire u0_u0__abc_72207_new_n426_; 
wire u0_u0__abc_72207_new_n428_; 
wire u0_u0__abc_72207_new_n429_; 
wire u0_u0__abc_72207_new_n431_; 
wire u0_u0__abc_72207_new_n432_; 
wire u0_u0__abc_72207_new_n434_; 
wire u0_u0__abc_72207_new_n435_; 
wire u0_u0__abc_72207_new_n436_; 
wire u0_u0__abc_72207_new_n437_; 
wire u0_u0__abc_72207_new_n438_; 
wire u0_u0__abc_72207_new_n439_; 
wire u0_u0__abc_72207_new_n440_; 
wire u0_u0__abc_72207_new_n441_; 
wire u0_u0__abc_72207_new_n442_; 
wire u0_u0__abc_72207_new_n443_; 
wire u0_u0__abc_72207_new_n444_; 
wire u0_u0__abc_72207_new_n445_; 
wire u0_u0__abc_72207_new_n446_; 
wire u0_u0__abc_72207_new_n447_; 
wire u0_u0__abc_72207_new_n448_; 
wire u0_u0__abc_72207_new_n449_; 
wire u0_u0__abc_72207_new_n450_; 
wire u0_u0__abc_72207_new_n451_; 
wire u0_u0__abc_72207_new_n452_; 
wire u0_u0__abc_72207_new_n453_; 
wire u0_u0__abc_72207_new_n454_; 
wire u0_u0__abc_72207_new_n455_; 
wire u0_u0__abc_72207_new_n456_; 
wire u0_u0__abc_72207_new_n457_; 
wire u0_u0__abc_72207_new_n458_; 
wire u0_u0__abc_72207_new_n462_; 
wire u0_u0__abc_72207_new_n463_; 
wire u0_u0__abc_72207_new_n464_; 
wire u0_u0_addr_r_2_; 
wire u0_u0_addr_r_3_; 
wire u0_u0_addr_r_4_; 
wire u0_u0_addr_r_5_; 
wire u0_u0_addr_r_6_; 
wire u0_u0_init_req_we; 
wire u0_u0_inited; 
wire u0_u0_lmr_req_we; 
wire u0_u0_rst_r2; 
wire u0_u0_wp_err; 
wire u0_u1__0csc_31_0__0_; 
wire u0_u1__0csc_31_0__10_; 
wire u0_u1__0csc_31_0__11_; 
wire u0_u1__0csc_31_0__12_; 
wire u0_u1__0csc_31_0__13_; 
wire u0_u1__0csc_31_0__14_; 
wire u0_u1__0csc_31_0__15_; 
wire u0_u1__0csc_31_0__16_; 
wire u0_u1__0csc_31_0__17_; 
wire u0_u1__0csc_31_0__18_; 
wire u0_u1__0csc_31_0__19_; 
wire u0_u1__0csc_31_0__1_; 
wire u0_u1__0csc_31_0__20_; 
wire u0_u1__0csc_31_0__21_; 
wire u0_u1__0csc_31_0__22_; 
wire u0_u1__0csc_31_0__23_; 
wire u0_u1__0csc_31_0__24_; 
wire u0_u1__0csc_31_0__25_; 
wire u0_u1__0csc_31_0__26_; 
wire u0_u1__0csc_31_0__27_; 
wire u0_u1__0csc_31_0__28_; 
wire u0_u1__0csc_31_0__29_; 
wire u0_u1__0csc_31_0__2_; 
wire u0_u1__0csc_31_0__30_; 
wire u0_u1__0csc_31_0__31_; 
wire u0_u1__0csc_31_0__3_; 
wire u0_u1__0csc_31_0__4_; 
wire u0_u1__0csc_31_0__5_; 
wire u0_u1__0csc_31_0__6_; 
wire u0_u1__0csc_31_0__7_; 
wire u0_u1__0csc_31_0__8_; 
wire u0_u1__0csc_31_0__9_; 
wire u0_u1__0init_req_0_0_; 
wire u0_u1__0init_req_we_0_0_; 
wire u0_u1__0inited_0_0_; 
wire u0_u1__0lmr_req_0_0_; 
wire u0_u1__0lmr_req_we_0_0_; 
wire u0_u1__0tms_31_0__0_; 
wire u0_u1__0tms_31_0__10_; 
wire u0_u1__0tms_31_0__11_; 
wire u0_u1__0tms_31_0__12_; 
wire u0_u1__0tms_31_0__13_; 
wire u0_u1__0tms_31_0__14_; 
wire u0_u1__0tms_31_0__15_; 
wire u0_u1__0tms_31_0__16_; 
wire u0_u1__0tms_31_0__17_; 
wire u0_u1__0tms_31_0__18_; 
wire u0_u1__0tms_31_0__19_; 
wire u0_u1__0tms_31_0__1_; 
wire u0_u1__0tms_31_0__20_; 
wire u0_u1__0tms_31_0__21_; 
wire u0_u1__0tms_31_0__22_; 
wire u0_u1__0tms_31_0__23_; 
wire u0_u1__0tms_31_0__24_; 
wire u0_u1__0tms_31_0__25_; 
wire u0_u1__0tms_31_0__26_; 
wire u0_u1__0tms_31_0__27_; 
wire u0_u1__0tms_31_0__28_; 
wire u0_u1__0tms_31_0__29_; 
wire u0_u1__0tms_31_0__2_; 
wire u0_u1__0tms_31_0__30_; 
wire u0_u1__0tms_31_0__31_; 
wire u0_u1__0tms_31_0__3_; 
wire u0_u1__0tms_31_0__4_; 
wire u0_u1__0tms_31_0__5_; 
wire u0_u1__0tms_31_0__6_; 
wire u0_u1__0tms_31_0__7_; 
wire u0_u1__0tms_31_0__8_; 
wire u0_u1__0tms_31_0__9_; 
wire u0_u1__abc_72470_auto_rtlil_cc_1942_NotGate_71506; 
wire u0_u1__abc_72470_new_n201_; 
wire u0_u1__abc_72470_new_n202_; 
wire u0_u1__abc_72470_new_n203_; 
wire u0_u1__abc_72470_new_n204_; 
wire u0_u1__abc_72470_new_n205_; 
wire u0_u1__abc_72470_new_n206_; 
wire u0_u1__abc_72470_new_n207_; 
wire u0_u1__abc_72470_new_n208_; 
wire u0_u1__abc_72470_new_n210_; 
wire u0_u1__abc_72470_new_n211_; 
wire u0_u1__abc_72470_new_n212_; 
wire u0_u1__abc_72470_new_n213_; 
wire u0_u1__abc_72470_new_n214_; 
wire u0_u1__abc_72470_new_n215_; 
wire u0_u1__abc_72470_new_n217_; 
wire u0_u1__abc_72470_new_n218_; 
wire u0_u1__abc_72470_new_n219_; 
wire u0_u1__abc_72470_new_n221_; 
wire u0_u1__abc_72470_new_n222_; 
wire u0_u1__abc_72470_new_n224_; 
wire u0_u1__abc_72470_new_n225_; 
wire u0_u1__abc_72470_new_n227_; 
wire u0_u1__abc_72470_new_n228_; 
wire u0_u1__abc_72470_new_n230_; 
wire u0_u1__abc_72470_new_n231_; 
wire u0_u1__abc_72470_new_n233_; 
wire u0_u1__abc_72470_new_n234_; 
wire u0_u1__abc_72470_new_n236_; 
wire u0_u1__abc_72470_new_n237_; 
wire u0_u1__abc_72470_new_n239_; 
wire u0_u1__abc_72470_new_n240_; 
wire u0_u1__abc_72470_new_n242_; 
wire u0_u1__abc_72470_new_n243_; 
wire u0_u1__abc_72470_new_n245_; 
wire u0_u1__abc_72470_new_n246_; 
wire u0_u1__abc_72470_new_n248_; 
wire u0_u1__abc_72470_new_n249_; 
wire u0_u1__abc_72470_new_n251_; 
wire u0_u1__abc_72470_new_n252_; 
wire u0_u1__abc_72470_new_n254_; 
wire u0_u1__abc_72470_new_n255_; 
wire u0_u1__abc_72470_new_n257_; 
wire u0_u1__abc_72470_new_n258_; 
wire u0_u1__abc_72470_new_n260_; 
wire u0_u1__abc_72470_new_n261_; 
wire u0_u1__abc_72470_new_n263_; 
wire u0_u1__abc_72470_new_n264_; 
wire u0_u1__abc_72470_new_n266_; 
wire u0_u1__abc_72470_new_n267_; 
wire u0_u1__abc_72470_new_n269_; 
wire u0_u1__abc_72470_new_n270_; 
wire u0_u1__abc_72470_new_n272_; 
wire u0_u1__abc_72470_new_n273_; 
wire u0_u1__abc_72470_new_n275_; 
wire u0_u1__abc_72470_new_n276_; 
wire u0_u1__abc_72470_new_n278_; 
wire u0_u1__abc_72470_new_n279_; 
wire u0_u1__abc_72470_new_n281_; 
wire u0_u1__abc_72470_new_n282_; 
wire u0_u1__abc_72470_new_n284_; 
wire u0_u1__abc_72470_new_n285_; 
wire u0_u1__abc_72470_new_n287_; 
wire u0_u1__abc_72470_new_n288_; 
wire u0_u1__abc_72470_new_n290_; 
wire u0_u1__abc_72470_new_n291_; 
wire u0_u1__abc_72470_new_n293_; 
wire u0_u1__abc_72470_new_n294_; 
wire u0_u1__abc_72470_new_n296_; 
wire u0_u1__abc_72470_new_n297_; 
wire u0_u1__abc_72470_new_n299_; 
wire u0_u1__abc_72470_new_n300_; 
wire u0_u1__abc_72470_new_n302_; 
wire u0_u1__abc_72470_new_n303_; 
wire u0_u1__abc_72470_new_n305_; 
wire u0_u1__abc_72470_new_n306_; 
wire u0_u1__abc_72470_new_n308_; 
wire u0_u1__abc_72470_new_n309_; 
wire u0_u1__abc_72470_new_n311_; 
wire u0_u1__abc_72470_new_n312_; 
wire u0_u1__abc_72470_new_n315_; 
wire u0_u1__abc_72470_new_n316_; 
wire u0_u1__abc_72470_new_n318_; 
wire u0_u1__abc_72470_new_n319_; 
wire u0_u1__abc_72470_new_n321_; 
wire u0_u1__abc_72470_new_n322_; 
wire u0_u1__abc_72470_new_n324_; 
wire u0_u1__abc_72470_new_n325_; 
wire u0_u1__abc_72470_new_n327_; 
wire u0_u1__abc_72470_new_n328_; 
wire u0_u1__abc_72470_new_n330_; 
wire u0_u1__abc_72470_new_n331_; 
wire u0_u1__abc_72470_new_n333_; 
wire u0_u1__abc_72470_new_n334_; 
wire u0_u1__abc_72470_new_n336_; 
wire u0_u1__abc_72470_new_n337_; 
wire u0_u1__abc_72470_new_n339_; 
wire u0_u1__abc_72470_new_n340_; 
wire u0_u1__abc_72470_new_n342_; 
wire u0_u1__abc_72470_new_n343_; 
wire u0_u1__abc_72470_new_n345_; 
wire u0_u1__abc_72470_new_n346_; 
wire u0_u1__abc_72470_new_n348_; 
wire u0_u1__abc_72470_new_n349_; 
wire u0_u1__abc_72470_new_n351_; 
wire u0_u1__abc_72470_new_n352_; 
wire u0_u1__abc_72470_new_n354_; 
wire u0_u1__abc_72470_new_n355_; 
wire u0_u1__abc_72470_new_n357_; 
wire u0_u1__abc_72470_new_n358_; 
wire u0_u1__abc_72470_new_n360_; 
wire u0_u1__abc_72470_new_n361_; 
wire u0_u1__abc_72470_new_n363_; 
wire u0_u1__abc_72470_new_n364_; 
wire u0_u1__abc_72470_new_n366_; 
wire u0_u1__abc_72470_new_n367_; 
wire u0_u1__abc_72470_new_n369_; 
wire u0_u1__abc_72470_new_n370_; 
wire u0_u1__abc_72470_new_n372_; 
wire u0_u1__abc_72470_new_n373_; 
wire u0_u1__abc_72470_new_n375_; 
wire u0_u1__abc_72470_new_n376_; 
wire u0_u1__abc_72470_new_n378_; 
wire u0_u1__abc_72470_new_n379_; 
wire u0_u1__abc_72470_new_n381_; 
wire u0_u1__abc_72470_new_n382_; 
wire u0_u1__abc_72470_new_n384_; 
wire u0_u1__abc_72470_new_n385_; 
wire u0_u1__abc_72470_new_n387_; 
wire u0_u1__abc_72470_new_n388_; 
wire u0_u1__abc_72470_new_n390_; 
wire u0_u1__abc_72470_new_n391_; 
wire u0_u1__abc_72470_new_n393_; 
wire u0_u1__abc_72470_new_n394_; 
wire u0_u1__abc_72470_new_n396_; 
wire u0_u1__abc_72470_new_n397_; 
wire u0_u1__abc_72470_new_n399_; 
wire u0_u1__abc_72470_new_n400_; 
wire u0_u1__abc_72470_new_n402_; 
wire u0_u1__abc_72470_new_n403_; 
wire u0_u1__abc_72470_new_n405_; 
wire u0_u1__abc_72470_new_n406_; 
wire u0_u1__abc_72470_new_n408_; 
wire u0_u1__abc_72470_new_n409_; 
wire u0_u1__abc_72470_new_n411_; 
wire u0_u1__abc_72470_new_n412_; 
wire u0_u1__abc_72470_new_n413_; 
wire u0_u1__abc_72470_new_n414_; 
wire u0_u1__abc_72470_new_n415_; 
wire u0_u1__abc_72470_new_n416_; 
wire u0_u1__abc_72470_new_n417_; 
wire u0_u1__abc_72470_new_n418_; 
wire u0_u1__abc_72470_new_n419_; 
wire u0_u1__abc_72470_new_n420_; 
wire u0_u1__abc_72470_new_n421_; 
wire u0_u1__abc_72470_new_n422_; 
wire u0_u1__abc_72470_new_n423_; 
wire u0_u1__abc_72470_new_n424_; 
wire u0_u1__abc_72470_new_n425_; 
wire u0_u1__abc_72470_new_n426_; 
wire u0_u1__abc_72470_new_n427_; 
wire u0_u1__abc_72470_new_n428_; 
wire u0_u1__abc_72470_new_n429_; 
wire u0_u1__abc_72470_new_n430_; 
wire u0_u1__abc_72470_new_n431_; 
wire u0_u1__abc_72470_new_n432_; 
wire u0_u1__abc_72470_new_n433_; 
wire u0_u1__abc_72470_new_n434_; 
wire u0_u1__abc_72470_new_n438_; 
wire u0_u1__abc_72470_new_n439_; 
wire u0_u1__abc_72470_new_n440_; 
wire u0_u1_addr_r_2_; 
wire u0_u1_addr_r_3_; 
wire u0_u1_addr_r_4_; 
wire u0_u1_addr_r_5_; 
wire u0_u1_addr_r_6_; 
wire u0_u1_init_req_we; 
wire u0_u1_inited; 
wire u0_u1_lmr_req_we; 
wire u0_u1_rst_r2; 
wire u0_u1_wp_err; 
wire u0_wb_addr_r_2_; 
wire u0_wb_addr_r_3_; 
wire u0_wb_addr_r_4_; 
wire u0_wb_addr_r_5_; 
wire u0_wb_addr_r_6_; 
wire u0_wp_err; 
wire u1__0acs_addr_23_0__0_; 
wire u1__0acs_addr_23_0__10_; 
wire u1__0acs_addr_23_0__11_; 
wire u1__0acs_addr_23_0__12_; 
wire u1__0acs_addr_23_0__13_; 
wire u1__0acs_addr_23_0__14_; 
wire u1__0acs_addr_23_0__15_; 
wire u1__0acs_addr_23_0__16_; 
wire u1__0acs_addr_23_0__17_; 
wire u1__0acs_addr_23_0__18_; 
wire u1__0acs_addr_23_0__19_; 
wire u1__0acs_addr_23_0__1_; 
wire u1__0acs_addr_23_0__20_; 
wire u1__0acs_addr_23_0__21_; 
wire u1__0acs_addr_23_0__22_; 
wire u1__0acs_addr_23_0__23_; 
wire u1__0acs_addr_23_0__2_; 
wire u1__0acs_addr_23_0__3_; 
wire u1__0acs_addr_23_0__4_; 
wire u1__0acs_addr_23_0__5_; 
wire u1__0acs_addr_23_0__6_; 
wire u1__0acs_addr_23_0__7_; 
wire u1__0acs_addr_23_0__8_; 
wire u1__0acs_addr_23_0__9_; 
wire u1__0bank_adr_1_0__0_; 
wire u1__0bank_adr_1_0__1_; 
wire u1__0col_adr_9_0__0_; 
wire u1__0col_adr_9_0__1_; 
wire u1__0col_adr_9_0__2_; 
wire u1__0col_adr_9_0__3_; 
wire u1__0col_adr_9_0__4_; 
wire u1__0col_adr_9_0__5_; 
wire u1__0col_adr_9_0__6_; 
wire u1__0col_adr_9_0__7_; 
wire u1__0col_adr_9_0__8_; 
wire u1__0col_adr_9_0__9_; 
wire u1__0row_adr_12_0__0_; 
wire u1__0row_adr_12_0__10_; 
wire u1__0row_adr_12_0__11_; 
wire u1__0row_adr_12_0__12_; 
wire u1__0row_adr_12_0__1_; 
wire u1__0row_adr_12_0__2_; 
wire u1__0row_adr_12_0__3_; 
wire u1__0row_adr_12_0__4_; 
wire u1__0row_adr_12_0__5_; 
wire u1__0row_adr_12_0__6_; 
wire u1__0row_adr_12_0__7_; 
wire u1__0row_adr_12_0__8_; 
wire u1__0row_adr_12_0__9_; 
wire u1__0sram_addr_23_0__0_; 
wire u1__0sram_addr_23_0__10_; 
wire u1__0sram_addr_23_0__11_; 
wire u1__0sram_addr_23_0__12_; 
wire u1__0sram_addr_23_0__13_; 
wire u1__0sram_addr_23_0__14_; 
wire u1__0sram_addr_23_0__15_; 
wire u1__0sram_addr_23_0__16_; 
wire u1__0sram_addr_23_0__17_; 
wire u1__0sram_addr_23_0__18_; 
wire u1__0sram_addr_23_0__19_; 
wire u1__0sram_addr_23_0__1_; 
wire u1__0sram_addr_23_0__20_; 
wire u1__0sram_addr_23_0__21_; 
wire u1__0sram_addr_23_0__22_; 
wire u1__0sram_addr_23_0__23_; 
wire u1__0sram_addr_23_0__2_; 
wire u1__0sram_addr_23_0__3_; 
wire u1__0sram_addr_23_0__4_; 
wire u1__0sram_addr_23_0__5_; 
wire u1__0sram_addr_23_0__6_; 
wire u1__0sram_addr_23_0__7_; 
wire u1__0sram_addr_23_0__8_; 
wire u1__0sram_addr_23_0__9_; 
wire u1__abc_72801_new_n258_; 
wire u1__abc_72801_new_n259_; 
wire u1__abc_72801_new_n260_; 
wire u1__abc_72801_new_n261_; 
wire u1__abc_72801_new_n262_; 
wire u1__abc_72801_new_n263_; 
wire u1__abc_72801_new_n264_; 
wire u1__abc_72801_new_n265_; 
wire u1__abc_72801_new_n266_; 
wire u1__abc_72801_new_n267_; 
wire u1__abc_72801_new_n268_; 
wire u1__abc_72801_new_n269_; 
wire u1__abc_72801_new_n270_; 
wire u1__abc_72801_new_n271_; 
wire u1__abc_72801_new_n273_; 
wire u1__abc_72801_new_n274_; 
wire u1__abc_72801_new_n276_; 
wire u1__abc_72801_new_n277_; 
wire u1__abc_72801_new_n278_; 
wire u1__abc_72801_new_n279_; 
wire u1__abc_72801_new_n280_; 
wire u1__abc_72801_new_n281_; 
wire u1__abc_72801_new_n282_; 
wire u1__abc_72801_new_n284_; 
wire u1__abc_72801_new_n285_; 
wire u1__abc_72801_new_n286_; 
wire u1__abc_72801_new_n287_; 
wire u1__abc_72801_new_n288_; 
wire u1__abc_72801_new_n289_; 
wire u1__abc_72801_new_n290_; 
wire u1__abc_72801_new_n291_; 
wire u1__abc_72801_new_n292_; 
wire u1__abc_72801_new_n293_; 
wire u1__abc_72801_new_n294_; 
wire u1__abc_72801_new_n295_; 
wire u1__abc_72801_new_n296_; 
wire u1__abc_72801_new_n297_; 
wire u1__abc_72801_new_n298_; 
wire u1__abc_72801_new_n299_; 
wire u1__abc_72801_new_n300_; 
wire u1__abc_72801_new_n301_; 
wire u1__abc_72801_new_n302_; 
wire u1__abc_72801_new_n303_; 
wire u1__abc_72801_new_n304_; 
wire u1__abc_72801_new_n305_; 
wire u1__abc_72801_new_n307_; 
wire u1__abc_72801_new_n308_; 
wire u1__abc_72801_new_n309_; 
wire u1__abc_72801_new_n310_; 
wire u1__abc_72801_new_n311_; 
wire u1__abc_72801_new_n312_; 
wire u1__abc_72801_new_n313_; 
wire u1__abc_72801_new_n314_; 
wire u1__abc_72801_new_n315_; 
wire u1__abc_72801_new_n316_; 
wire u1__abc_72801_new_n317_; 
wire u1__abc_72801_new_n318_; 
wire u1__abc_72801_new_n319_; 
wire u1__abc_72801_new_n320_; 
wire u1__abc_72801_new_n322_; 
wire u1__abc_72801_new_n323_; 
wire u1__abc_72801_new_n324_; 
wire u1__abc_72801_new_n325_; 
wire u1__abc_72801_new_n326_; 
wire u1__abc_72801_new_n327_; 
wire u1__abc_72801_new_n328_; 
wire u1__abc_72801_new_n329_; 
wire u1__abc_72801_new_n331_; 
wire u1__abc_72801_new_n332_; 
wire u1__abc_72801_new_n333_; 
wire u1__abc_72801_new_n334_; 
wire u1__abc_72801_new_n335_; 
wire u1__abc_72801_new_n336_; 
wire u1__abc_72801_new_n337_; 
wire u1__abc_72801_new_n338_; 
wire u1__abc_72801_new_n339_; 
wire u1__abc_72801_new_n340_; 
wire u1__abc_72801_new_n341_; 
wire u1__abc_72801_new_n342_; 
wire u1__abc_72801_new_n343_; 
wire u1__abc_72801_new_n344_; 
wire u1__abc_72801_new_n346_; 
wire u1__abc_72801_new_n347_; 
wire u1__abc_72801_new_n348_; 
wire u1__abc_72801_new_n349_; 
wire u1__abc_72801_new_n350_; 
wire u1__abc_72801_new_n351_; 
wire u1__abc_72801_new_n352_; 
wire u1__abc_72801_new_n353_; 
wire u1__abc_72801_new_n354_; 
wire u1__abc_72801_new_n355_; 
wire u1__abc_72801_new_n356_; 
wire u1__abc_72801_new_n357_; 
wire u1__abc_72801_new_n359_; 
wire u1__abc_72801_new_n360_; 
wire u1__abc_72801_new_n361_; 
wire u1__abc_72801_new_n362_; 
wire u1__abc_72801_new_n363_; 
wire u1__abc_72801_new_n364_; 
wire u1__abc_72801_new_n365_; 
wire u1__abc_72801_new_n366_; 
wire u1__abc_72801_new_n367_; 
wire u1__abc_72801_new_n368_; 
wire u1__abc_72801_new_n369_; 
wire u1__abc_72801_new_n371_; 
wire u1__abc_72801_new_n372_; 
wire u1__abc_72801_new_n373_; 
wire u1__abc_72801_new_n374_; 
wire u1__abc_72801_new_n375_; 
wire u1__abc_72801_new_n376_; 
wire u1__abc_72801_new_n377_; 
wire u1__abc_72801_new_n378_; 
wire u1__abc_72801_new_n380_; 
wire u1__abc_72801_new_n381_; 
wire u1__abc_72801_new_n382_; 
wire u1__abc_72801_new_n383_; 
wire u1__abc_72801_new_n384_; 
wire u1__abc_72801_new_n385_; 
wire u1__abc_72801_new_n386_; 
wire u1__abc_72801_new_n387_; 
wire u1__abc_72801_new_n389_; 
wire u1__abc_72801_new_n390_; 
wire u1__abc_72801_new_n391_; 
wire u1__abc_72801_new_n392_; 
wire u1__abc_72801_new_n393_; 
wire u1__abc_72801_new_n394_; 
wire u1__abc_72801_new_n395_; 
wire u1__abc_72801_new_n396_; 
wire u1__abc_72801_new_n398_; 
wire u1__abc_72801_new_n399_; 
wire u1__abc_72801_new_n400_; 
wire u1__abc_72801_new_n401_; 
wire u1__abc_72801_new_n402_; 
wire u1__abc_72801_new_n403_; 
wire u1__abc_72801_new_n404_; 
wire u1__abc_72801_new_n405_; 
wire u1__abc_72801_new_n407_; 
wire u1__abc_72801_new_n408_; 
wire u1__abc_72801_new_n409_; 
wire u1__abc_72801_new_n410_; 
wire u1__abc_72801_new_n411_; 
wire u1__abc_72801_new_n412_; 
wire u1__abc_72801_new_n413_; 
wire u1__abc_72801_new_n414_; 
wire u1__abc_72801_new_n415_; 
wire u1__abc_72801_new_n417_; 
wire u1__abc_72801_new_n418_; 
wire u1__abc_72801_new_n419_; 
wire u1__abc_72801_new_n420_; 
wire u1__abc_72801_new_n421_; 
wire u1__abc_72801_new_n422_; 
wire u1__abc_72801_new_n423_; 
wire u1__abc_72801_new_n424_; 
wire u1__abc_72801_new_n425_; 
wire u1__abc_72801_new_n426_; 
wire u1__abc_72801_new_n427_; 
wire u1__abc_72801_new_n428_; 
wire u1__abc_72801_new_n430_; 
wire u1__abc_72801_new_n431_; 
wire u1__abc_72801_new_n432_; 
wire u1__abc_72801_new_n433_; 
wire u1__abc_72801_new_n434_; 
wire u1__abc_72801_new_n435_; 
wire u1__abc_72801_new_n436_; 
wire u1__abc_72801_new_n437_; 
wire u1__abc_72801_new_n438_; 
wire u1__abc_72801_new_n439_; 
wire u1__abc_72801_new_n441_; 
wire u1__abc_72801_new_n442_; 
wire u1__abc_72801_new_n443_; 
wire u1__abc_72801_new_n444_; 
wire u1__abc_72801_new_n445_; 
wire u1__abc_72801_new_n446_; 
wire u1__abc_72801_new_n447_; 
wire u1__abc_72801_new_n448_; 
wire u1__abc_72801_new_n449_; 
wire u1__abc_72801_new_n450_; 
wire u1__abc_72801_new_n451_; 
wire u1__abc_72801_new_n453_; 
wire u1__abc_72801_new_n454_; 
wire u1__abc_72801_new_n455_; 
wire u1__abc_72801_new_n456_; 
wire u1__abc_72801_new_n457_; 
wire u1__abc_72801_new_n458_; 
wire u1__abc_72801_new_n460_; 
wire u1__abc_72801_new_n461_; 
wire u1__abc_72801_new_n462_; 
wire u1__abc_72801_new_n464_; 
wire u1__abc_72801_new_n465_; 
wire u1__abc_72801_new_n467_; 
wire u1__abc_72801_new_n468_; 
wire u1__abc_72801_new_n470_; 
wire u1__abc_72801_new_n471_; 
wire u1__abc_72801_new_n473_; 
wire u1__abc_72801_new_n474_; 
wire u1__abc_72801_new_n476_; 
wire u1__abc_72801_new_n477_; 
wire u1__abc_72801_new_n479_; 
wire u1__abc_72801_new_n480_; 
wire u1__abc_72801_new_n482_; 
wire u1__abc_72801_new_n483_; 
wire u1__abc_72801_new_n485_; 
wire u1__abc_72801_new_n486_; 
wire u1__abc_72801_new_n488_; 
wire u1__abc_72801_new_n489_; 
wire u1__abc_72801_new_n491_; 
wire u1__abc_72801_new_n492_; 
wire u1__abc_72801_new_n493_; 
wire u1__abc_72801_new_n494_; 
wire u1__abc_72801_new_n495_; 
wire u1__abc_72801_new_n496_; 
wire u1__abc_72801_new_n498_; 
wire u1__abc_72801_new_n499_; 
wire u1__abc_72801_new_n500_; 
wire u1__abc_72801_new_n501_; 
wire u1__abc_72801_new_n502_; 
wire u1__abc_72801_new_n503_; 
wire u1__abc_72801_new_n505_; 
wire u1__abc_72801_new_n506_; 
wire u1__abc_72801_new_n507_; 
wire u1__abc_72801_new_n508_; 
wire u1__abc_72801_new_n510_; 
wire u1__abc_72801_new_n511_; 
wire u1__abc_72801_new_n512_; 
wire u1__abc_72801_new_n513_; 
wire u1__abc_72801_new_n515_; 
wire u1__abc_72801_new_n516_; 
wire u1__abc_72801_new_n517_; 
wire u1__abc_72801_new_n518_; 
wire u1__abc_72801_new_n520_; 
wire u1__abc_72801_new_n521_; 
wire u1__abc_72801_new_n522_; 
wire u1__abc_72801_new_n523_; 
wire u1__abc_72801_new_n525_; 
wire u1__abc_72801_new_n526_; 
wire u1__abc_72801_new_n527_; 
wire u1__abc_72801_new_n528_; 
wire u1__abc_72801_new_n530_; 
wire u1__abc_72801_new_n531_; 
wire u1__abc_72801_new_n532_; 
wire u1__abc_72801_new_n533_; 
wire u1__abc_72801_new_n535_; 
wire u1__abc_72801_new_n536_; 
wire u1__abc_72801_new_n537_; 
wire u1__abc_72801_new_n538_; 
wire u1__abc_72801_new_n539_; 
wire u1__abc_72801_new_n541_; 
wire u1__abc_72801_new_n542_; 
wire u1__abc_72801_new_n543_; 
wire u1__abc_72801_new_n544_; 
wire u1__abc_72801_new_n545_; 
wire u1__abc_72801_new_n546_; 
wire u1__abc_72801_new_n548_; 
wire u1__abc_72801_new_n549_; 
wire u1__abc_72801_new_n550_; 
wire u1__abc_72801_new_n551_; 
wire u1__abc_72801_new_n553_; 
wire u1__abc_72801_new_n554_; 
wire u1__abc_72801_new_n555_; 
wire u1__abc_72801_new_n556_; 
wire u1__abc_72801_new_n558_; 
wire u1__abc_72801_new_n559_; 
wire u1__abc_72801_new_n560_; 
wire u1__abc_72801_new_n561_; 
wire u1__abc_72801_new_n563_; 
wire u1__abc_72801_new_n564_; 
wire u1__abc_72801_new_n565_; 
wire u1__abc_72801_new_n566_; 
wire u1__abc_72801_new_n568_; 
wire u1__abc_72801_new_n569_; 
wire u1__abc_72801_new_n570_; 
wire u1__abc_72801_new_n571_; 
wire u1__abc_72801_new_n573_; 
wire u1__abc_72801_new_n574_; 
wire u1__abc_72801_new_n575_; 
wire u1__abc_72801_new_n576_; 
wire u1__abc_72801_new_n577_; 
wire u1__abc_72801_new_n579_; 
wire u1__abc_72801_new_n580_; 
wire u1__abc_72801_new_n581_; 
wire u1__abc_72801_new_n582_; 
wire u1__abc_72801_new_n583_; 
wire u1__abc_72801_new_n585_; 
wire u1__abc_72801_new_n586_; 
wire u1__abc_72801_new_n587_; 
wire u1__abc_72801_new_n588_; 
wire u1__abc_72801_new_n589_; 
wire u1__abc_72801_new_n591_; 
wire u1__abc_72801_new_n592_; 
wire u1__abc_72801_new_n593_; 
wire u1__abc_72801_new_n594_; 
wire u1__abc_72801_new_n596_; 
wire u1__abc_72801_new_n597_; 
wire u1__abc_72801_new_n598_; 
wire u1__abc_72801_new_n599_; 
wire u1__abc_72801_new_n601_; 
wire u1__abc_72801_new_n602_; 
wire u1__abc_72801_new_n603_; 
wire u1__abc_72801_new_n605_; 
wire u1__abc_72801_new_n606_; 
wire u1__abc_72801_new_n607_; 
wire u1__abc_72801_new_n608_; 
wire u1__abc_72801_new_n610_; 
wire u1__abc_72801_new_n611_; 
wire u1__abc_72801_new_n612_; 
wire u1__abc_72801_new_n613_; 
wire u1__abc_72801_new_n615_; 
wire u1__abc_72801_new_n616_; 
wire u1__abc_72801_new_n617_; 
wire u1__abc_72801_new_n618_; 
wire u1__abc_72801_new_n620_; 
wire u1__abc_72801_new_n622_; 
wire u1__abc_72801_new_n624_; 
wire u1__abc_72801_new_n626_; 
wire u1__abc_72801_new_n628_; 
wire u1__abc_72801_new_n630_; 
wire u1__abc_72801_new_n632_; 
wire u1__abc_72801_new_n634_; 
wire u1__abc_72801_new_n636_; 
wire u1__abc_72801_new_n638_; 
wire u1__abc_72801_new_n640_; 
wire u1__abc_72801_new_n642_; 
wire u1__abc_72801_new_n644_; 
wire u1__abc_72801_new_n646_; 
wire u1__abc_72801_new_n648_; 
wire u1__abc_72801_new_n649_; 
wire u1__abc_72801_new_n651_; 
wire u1__abc_72801_new_n652_; 
wire u1__abc_72801_new_n654_; 
wire u1__abc_72801_new_n655_; 
wire u1__abc_72801_new_n657_; 
wire u1__abc_72801_new_n659_; 
wire u1__abc_72801_new_n661_; 
wire u1__abc_72801_new_n663_; 
wire u1__abc_72801_new_n665_; 
wire u1__abc_72801_new_n667_; 
wire u1__abc_72801_new_n669_; 
wire u1__abc_72801_new_n671_; 
wire u1__abc_72801_new_n672_; 
wire u1__abc_72801_new_n673_; 
wire u1__abc_72801_new_n674_; 
wire u1__abc_72801_new_n675_; 
wire u1__abc_72801_new_n676_; 
wire u1__abc_72801_new_n677_; 
wire u1__abc_72801_new_n678_; 
wire u1__abc_72801_new_n679_; 
wire u1__abc_72801_new_n680_; 
wire u1__abc_72801_new_n681_; 
wire u1__abc_72801_new_n682_; 
wire u1__abc_72801_new_n683_; 
wire u1__abc_72801_new_n684_; 
wire u1__abc_72801_new_n685_; 
wire u1__abc_72801_new_n686_; 
wire u1__abc_72801_new_n687_; 
wire u1__abc_72801_new_n688_; 
wire u1__abc_72801_new_n690_; 
wire u1__abc_72801_new_n691_; 
wire u1__abc_72801_new_n692_; 
wire u1__abc_72801_new_n693_; 
wire u1__abc_72801_new_n694_; 
wire u1__abc_72801_new_n695_; 
wire u1__abc_72801_new_n696_; 
wire u1__abc_72801_new_n698_; 
wire u1__abc_72801_new_n699_; 
wire u1__abc_72801_new_n700_; 
wire u1__abc_72801_new_n701_; 
wire u1__abc_72801_new_n702_; 
wire u1__abc_72801_new_n703_; 
wire u1__abc_72801_new_n704_; 
wire u1__abc_72801_new_n705_; 
wire u1__abc_72801_new_n707_; 
wire u1__abc_72801_new_n708_; 
wire u1__abc_72801_new_n709_; 
wire u1__abc_72801_new_n710_; 
wire u1__abc_72801_new_n711_; 
wire u1__abc_72801_new_n712_; 
wire u1__abc_72801_new_n713_; 
wire u1__abc_72801_new_n715_; 
wire u1__abc_72801_new_n716_; 
wire u1__abc_72801_new_n717_; 
wire u1__abc_72801_new_n718_; 
wire u1__abc_72801_new_n719_; 
wire u1__abc_72801_new_n720_; 
wire u1__abc_72801_new_n721_; 
wire u1__abc_72801_new_n723_; 
wire u1__abc_72801_new_n724_; 
wire u1__abc_72801_new_n725_; 
wire u1__abc_72801_new_n726_; 
wire u1__abc_72801_new_n727_; 
wire u1__abc_72801_new_n728_; 
wire u1__abc_72801_new_n729_; 
wire u1__abc_72801_new_n731_; 
wire u1__abc_72801_new_n732_; 
wire u1__abc_72801_new_n733_; 
wire u1__abc_72801_new_n734_; 
wire u1__abc_72801_new_n735_; 
wire u1__abc_72801_new_n736_; 
wire u1__abc_72801_new_n737_; 
wire u1__abc_72801_new_n739_; 
wire u1__abc_72801_new_n740_; 
wire u1__abc_72801_new_n741_; 
wire u1__abc_72801_new_n742_; 
wire u1__abc_72801_new_n743_; 
wire u1__abc_72801_new_n744_; 
wire u1__abc_72801_new_n745_; 
wire u1__abc_72801_new_n747_; 
wire u1__abc_72801_new_n748_; 
wire u1__abc_72801_new_n749_; 
wire u1__abc_72801_new_n750_; 
wire u1__abc_72801_new_n751_; 
wire u1__abc_72801_new_n752_; 
wire u1__abc_72801_new_n753_; 
wire u1__abc_72801_new_n755_; 
wire u1__abc_72801_new_n756_; 
wire u1__abc_72801_new_n757_; 
wire u1__abc_72801_new_n758_; 
wire u1__abc_72801_new_n759_; 
wire u1__abc_72801_new_n760_; 
wire u1__abc_72801_new_n761_; 
wire u1__abc_72801_new_n762_; 
wire u1__abc_72801_new_n764_; 
wire u1__abc_72801_new_n765_; 
wire u1__abc_72801_new_n766_; 
wire u1__abc_72801_new_n767_; 
wire u1__abc_72801_new_n768_; 
wire u1__abc_72801_new_n769_; 
wire u1__abc_72801_new_n770_; 
wire u1__abc_72801_new_n772_; 
wire u1__abc_72801_new_n773_; 
wire u1__abc_72801_new_n774_; 
wire u1__abc_72801_new_n775_; 
wire u1__abc_72801_new_n776_; 
wire u1__abc_72801_new_n777_; 
wire u1__abc_72801_new_n778_; 
wire u1__abc_72801_new_n780_; 
wire u1__abc_72801_new_n781_; 
wire u1__abc_72801_new_n782_; 
wire u1__abc_72801_new_n783_; 
wire u1__abc_72801_new_n785_; 
wire u1__abc_72801_new_n786_; 
wire u1__abc_72801_new_n787_; 
wire u1__abc_72801_new_n788_; 
wire u1__abc_72801_new_n790_; 
wire u1__abc_72801_new_n791_; 
wire u1__abc_72801_new_n792_; 
wire u1__abc_72801_new_n794_; 
wire u1__abc_72801_new_n795_; 
wire u1__abc_72801_new_n796_; 
wire u1__abc_72801_new_n798_; 
wire u1__abc_72801_new_n799_; 
wire u1__abc_72801_new_n801_; 
wire u1__abc_72801_new_n802_; 
wire u1__abc_72801_new_n804_; 
wire u1__abc_72801_new_n805_; 
wire u1__abc_72801_new_n807_; 
wire u1__abc_72801_new_n808_; 
wire u1__abc_72801_new_n810_; 
wire u1__abc_72801_new_n811_; 
wire u1__abc_72801_new_n813_; 
wire u1__abc_72801_new_n814_; 
wire u1__abc_72801_new_n816_; 
wire u1__abc_72801_new_n817_; 
wire u1__abc_72801_new_n819_; 
wire u1__abc_72801_new_n820_; 
wire u1__abc_72801_new_n821_; 
wire u1__abc_72801_new_n822_; 
wire u1__abc_72801_new_n823_; 
wire u1__abc_72801_new_n824_; 
wire u1__abc_72801_new_n825_; 
wire u1__abc_72801_new_n826_; 
wire u1_acs_addr_0_; 
wire u1_acs_addr_10_; 
wire u1_acs_addr_11_; 
wire u1_acs_addr_12_; 
wire u1_acs_addr_13_; 
wire u1_acs_addr_14_; 
wire u1_acs_addr_15_; 
wire u1_acs_addr_16_; 
wire u1_acs_addr_17_; 
wire u1_acs_addr_18_; 
wire u1_acs_addr_19_; 
wire u1_acs_addr_1_; 
wire u1_acs_addr_20_; 
wire u1_acs_addr_21_; 
wire u1_acs_addr_22_; 
wire u1_acs_addr_23_; 
wire u1_acs_addr_2_; 
wire u1_acs_addr_3_; 
wire u1_acs_addr_4_; 
wire u1_acs_addr_5_; 
wire u1_acs_addr_6_; 
wire u1_acs_addr_7_; 
wire u1_acs_addr_8_; 
wire u1_acs_addr_9_; 
wire u1_acs_addr_pl1_0_; 
wire u1_acs_addr_pl1_10_; 
wire u1_acs_addr_pl1_11_; 
wire u1_acs_addr_pl1_12_; 
wire u1_acs_addr_pl1_13_; 
wire u1_acs_addr_pl1_14_; 
wire u1_acs_addr_pl1_15_; 
wire u1_acs_addr_pl1_16_; 
wire u1_acs_addr_pl1_17_; 
wire u1_acs_addr_pl1_18_; 
wire u1_acs_addr_pl1_19_; 
wire u1_acs_addr_pl1_1_; 
wire u1_acs_addr_pl1_20_; 
wire u1_acs_addr_pl1_21_; 
wire u1_acs_addr_pl1_22_; 
wire u1_acs_addr_pl1_23_; 
wire u1_acs_addr_pl1_2_; 
wire u1_acs_addr_pl1_3_; 
wire u1_acs_addr_pl1_4_; 
wire u1_acs_addr_pl1_5_; 
wire u1_acs_addr_pl1_6_; 
wire u1_acs_addr_pl1_7_; 
wire u1_acs_addr_pl1_8_; 
wire u1_acs_addr_pl1_9_; 
wire u1_bas; 
wire u1_col_adr_0_; 
wire u1_col_adr_1_; 
wire u1_col_adr_2_; 
wire u1_col_adr_3_; 
wire u1_col_adr_4_; 
wire u1_col_adr_5_; 
wire u1_col_adr_6_; 
wire u1_col_adr_7_; 
wire u1_col_adr_8_; 
wire u1_col_adr_9_; 
wire u1_sram_addr_0_; 
wire u1_sram_addr_10_; 
wire u1_sram_addr_11_; 
wire u1_sram_addr_12_; 
wire u1_sram_addr_13_; 
wire u1_sram_addr_14_; 
wire u1_sram_addr_15_; 
wire u1_sram_addr_16_; 
wire u1_sram_addr_17_; 
wire u1_sram_addr_18_; 
wire u1_sram_addr_19_; 
wire u1_sram_addr_1_; 
wire u1_sram_addr_20_; 
wire u1_sram_addr_21_; 
wire u1_sram_addr_22_; 
wire u1_sram_addr_23_; 
wire u1_sram_addr_2_; 
wire u1_sram_addr_3_; 
wire u1_sram_addr_4_; 
wire u1_sram_addr_5_; 
wire u1_sram_addr_6_; 
wire u1_sram_addr_7_; 
wire u1_sram_addr_8_; 
wire u1_sram_addr_9_; 
wire u1_u0__0out_r_12_0__0_; 
wire u1_u0__0out_r_12_0__10_; 
wire u1_u0__0out_r_12_0__11_; 
wire u1_u0__0out_r_12_0__12_; 
wire u1_u0__0out_r_12_0__1_; 
wire u1_u0__0out_r_12_0__2_; 
wire u1_u0__0out_r_12_0__3_; 
wire u1_u0__0out_r_12_0__4_; 
wire u1_u0__0out_r_12_0__5_; 
wire u1_u0__0out_r_12_0__6_; 
wire u1_u0__0out_r_12_0__7_; 
wire u1_u0__0out_r_12_0__8_; 
wire u1_u0__0out_r_12_0__9_; 
wire u1_u0__abc_72719_new_n100_; 
wire u1_u0__abc_72719_new_n102_; 
wire u1_u0__abc_72719_new_n103_; 
wire u1_u0__abc_72719_new_n104_; 
wire u1_u0__abc_72719_new_n107_; 
wire u1_u0__abc_72719_new_n108_; 
wire u1_u0__abc_72719_new_n109_; 
wire u1_u0__abc_72719_new_n111_; 
wire u1_u0__abc_72719_new_n112_; 
wire u1_u0__abc_72719_new_n113_; 
wire u1_u0__abc_72719_new_n114_; 
wire u1_u0__abc_72719_new_n115_; 
wire u1_u0__abc_72719_new_n116_; 
wire u1_u0__abc_72719_new_n119_; 
wire u1_u0__abc_72719_new_n120_; 
wire u1_u0__abc_72719_new_n121_; 
wire u1_u0__abc_72719_new_n123_; 
wire u1_u0__abc_72719_new_n124_; 
wire u1_u0__abc_72719_new_n125_; 
wire u1_u0__abc_72719_new_n126_; 
wire u1_u0__abc_72719_new_n127_; 
wire u1_u0__abc_72719_new_n129_; 
wire u1_u0__abc_72719_new_n52_; 
wire u1_u0__abc_72719_new_n54_; 
wire u1_u0__abc_72719_new_n56_; 
wire u1_u0__abc_72719_new_n57_; 
wire u1_u0__abc_72719_new_n58_; 
wire u1_u0__abc_72719_new_n60_; 
wire u1_u0__abc_72719_new_n61_; 
wire u1_u0__abc_72719_new_n62_; 
wire u1_u0__abc_72719_new_n65_; 
wire u1_u0__abc_72719_new_n66_; 
wire u1_u0__abc_72719_new_n67_; 
wire u1_u0__abc_72719_new_n68_; 
wire u1_u0__abc_72719_new_n69_; 
wire u1_u0__abc_72719_new_n70_; 
wire u1_u0__abc_72719_new_n71_; 
wire u1_u0__abc_72719_new_n74_; 
wire u1_u0__abc_72719_new_n75_; 
wire u1_u0__abc_72719_new_n76_; 
wire u1_u0__abc_72719_new_n77_; 
wire u1_u0__abc_72719_new_n78_; 
wire u1_u0__abc_72719_new_n81_; 
wire u1_u0__abc_72719_new_n82_; 
wire u1_u0__abc_72719_new_n83_; 
wire u1_u0__abc_72719_new_n84_; 
wire u1_u0__abc_72719_new_n85_; 
wire u1_u0__abc_72719_new_n86_; 
wire u1_u0__abc_72719_new_n89_; 
wire u1_u0__abc_72719_new_n91_; 
wire u1_u0__abc_72719_new_n93_; 
wire u1_u0__abc_72719_new_n94_; 
wire u1_u0__abc_72719_new_n95_; 
wire u1_u0__abc_72719_new_n96_; 
wire u1_u0__abc_72719_new_n97_; 
wire u1_u0__abc_72719_new_n99_; 
wire u1_u0_inc_next; 
wire u1_wb_write_go; 
wire u1_wr_cycle; 
wire u1_wr_hold; 
wire u2__0bank_open_0_0_; 
wire u2__0row_same_0_0_; 
wire u2__abc_74202_new_n100_; 
wire u2__abc_74202_new_n101_; 
wire u2__abc_74202_new_n102_; 
wire u2__abc_74202_new_n103_; 
wire u2__abc_74202_new_n104_; 
wire u2__abc_74202_new_n105_; 
wire u2__abc_74202_new_n107_; 
wire u2__abc_74202_new_n108_; 
wire u2__abc_74202_new_n109_; 
wire u2__abc_74202_new_n110_; 
wire u2__abc_74202_new_n111_; 
wire u2__abc_74202_new_n112_; 
wire u2__abc_74202_new_n64_; 
wire u2__abc_74202_new_n65_; 
wire u2__abc_74202_new_n67_; 
wire u2__abc_74202_new_n81_; 
wire u2__abc_74202_new_n90_; 
wire u2__abc_74202_new_n91_; 
wire u2_bank_clr_0; 
wire u2_bank_clr_1; 
wire u2_bank_clr_all_0; 
wire u2_bank_clr_all_1; 
wire u2_bank_open_0; 
wire u2_bank_open_1; 
wire u2_bank_set_0; 
wire u2_bank_set_1; 
wire u2_row_same_0; 
wire u2_row_same_1; 
wire u2_u0__0b0_last_row_12_0__0_; 
wire u2_u0__0b0_last_row_12_0__10_; 
wire u2_u0__0b0_last_row_12_0__11_; 
wire u2_u0__0b0_last_row_12_0__12_; 
wire u2_u0__0b0_last_row_12_0__1_; 
wire u2_u0__0b0_last_row_12_0__2_; 
wire u2_u0__0b0_last_row_12_0__3_; 
wire u2_u0__0b0_last_row_12_0__4_; 
wire u2_u0__0b0_last_row_12_0__5_; 
wire u2_u0__0b0_last_row_12_0__6_; 
wire u2_u0__0b0_last_row_12_0__7_; 
wire u2_u0__0b0_last_row_12_0__8_; 
wire u2_u0__0b0_last_row_12_0__9_; 
wire u2_u0__0b1_last_row_12_0__0_; 
wire u2_u0__0b1_last_row_12_0__10_; 
wire u2_u0__0b1_last_row_12_0__11_; 
wire u2_u0__0b1_last_row_12_0__12_; 
wire u2_u0__0b1_last_row_12_0__1_; 
wire u2_u0__0b1_last_row_12_0__2_; 
wire u2_u0__0b1_last_row_12_0__3_; 
wire u2_u0__0b1_last_row_12_0__4_; 
wire u2_u0__0b1_last_row_12_0__5_; 
wire u2_u0__0b1_last_row_12_0__6_; 
wire u2_u0__0b1_last_row_12_0__7_; 
wire u2_u0__0b1_last_row_12_0__8_; 
wire u2_u0__0b1_last_row_12_0__9_; 
wire u2_u0__0b2_last_row_12_0__0_; 
wire u2_u0__0b2_last_row_12_0__10_; 
wire u2_u0__0b2_last_row_12_0__11_; 
wire u2_u0__0b2_last_row_12_0__12_; 
wire u2_u0__0b2_last_row_12_0__1_; 
wire u2_u0__0b2_last_row_12_0__2_; 
wire u2_u0__0b2_last_row_12_0__3_; 
wire u2_u0__0b2_last_row_12_0__4_; 
wire u2_u0__0b2_last_row_12_0__5_; 
wire u2_u0__0b2_last_row_12_0__6_; 
wire u2_u0__0b2_last_row_12_0__7_; 
wire u2_u0__0b2_last_row_12_0__8_; 
wire u2_u0__0b2_last_row_12_0__9_; 
wire u2_u0__0b3_last_row_12_0__0_; 
wire u2_u0__0b3_last_row_12_0__10_; 
wire u2_u0__0b3_last_row_12_0__11_; 
wire u2_u0__0b3_last_row_12_0__12_; 
wire u2_u0__0b3_last_row_12_0__1_; 
wire u2_u0__0b3_last_row_12_0__2_; 
wire u2_u0__0b3_last_row_12_0__3_; 
wire u2_u0__0b3_last_row_12_0__4_; 
wire u2_u0__0b3_last_row_12_0__5_; 
wire u2_u0__0b3_last_row_12_0__6_; 
wire u2_u0__0b3_last_row_12_0__7_; 
wire u2_u0__0b3_last_row_12_0__8_; 
wire u2_u0__0b3_last_row_12_0__9_; 
wire u2_u0__0bank0_open_0_0_; 
wire u2_u0__0bank1_open_0_0_; 
wire u2_u0__0bank2_open_0_0_; 
wire u2_u0__0bank3_open_0_0_; 
wire u2_u0__abc_73914_auto_rtlil_cc_1942_NotGate_71538; 
wire u2_u0__abc_73914_new_n136_; 
wire u2_u0__abc_73914_new_n137_; 
wire u2_u0__abc_73914_new_n138_; 
wire u2_u0__abc_73914_new_n139_; 
wire u2_u0__abc_73914_new_n140_; 
wire u2_u0__abc_73914_new_n141_; 
wire u2_u0__abc_73914_new_n143_; 
wire u2_u0__abc_73914_new_n144_; 
wire u2_u0__abc_73914_new_n146_; 
wire u2_u0__abc_73914_new_n147_; 
wire u2_u0__abc_73914_new_n149_; 
wire u2_u0__abc_73914_new_n150_; 
wire u2_u0__abc_73914_new_n152_; 
wire u2_u0__abc_73914_new_n153_; 
wire u2_u0__abc_73914_new_n155_; 
wire u2_u0__abc_73914_new_n156_; 
wire u2_u0__abc_73914_new_n158_; 
wire u2_u0__abc_73914_new_n159_; 
wire u2_u0__abc_73914_new_n161_; 
wire u2_u0__abc_73914_new_n162_; 
wire u2_u0__abc_73914_new_n164_; 
wire u2_u0__abc_73914_new_n165_; 
wire u2_u0__abc_73914_new_n167_; 
wire u2_u0__abc_73914_new_n168_; 
wire u2_u0__abc_73914_new_n170_; 
wire u2_u0__abc_73914_new_n171_; 
wire u2_u0__abc_73914_new_n173_; 
wire u2_u0__abc_73914_new_n174_; 
wire u2_u0__abc_73914_new_n176_; 
wire u2_u0__abc_73914_new_n177_; 
wire u2_u0__abc_73914_new_n179_; 
wire u2_u0__abc_73914_new_n180_; 
wire u2_u0__abc_73914_new_n181_; 
wire u2_u0__abc_73914_new_n182_; 
wire u2_u0__abc_73914_new_n184_; 
wire u2_u0__abc_73914_new_n186_; 
wire u2_u0__abc_73914_new_n188_; 
wire u2_u0__abc_73914_new_n190_; 
wire u2_u0__abc_73914_new_n192_; 
wire u2_u0__abc_73914_new_n194_; 
wire u2_u0__abc_73914_new_n196_; 
wire u2_u0__abc_73914_new_n198_; 
wire u2_u0__abc_73914_new_n200_; 
wire u2_u0__abc_73914_new_n202_; 
wire u2_u0__abc_73914_new_n204_; 
wire u2_u0__abc_73914_new_n206_; 
wire u2_u0__abc_73914_new_n208_; 
wire u2_u0__abc_73914_new_n209_; 
wire u2_u0__abc_73914_new_n210_; 
wire u2_u0__abc_73914_new_n211_; 
wire u2_u0__abc_73914_new_n213_; 
wire u2_u0__abc_73914_new_n215_; 
wire u2_u0__abc_73914_new_n217_; 
wire u2_u0__abc_73914_new_n219_; 
wire u2_u0__abc_73914_new_n221_; 
wire u2_u0__abc_73914_new_n223_; 
wire u2_u0__abc_73914_new_n225_; 
wire u2_u0__abc_73914_new_n227_; 
wire u2_u0__abc_73914_new_n229_; 
wire u2_u0__abc_73914_new_n231_; 
wire u2_u0__abc_73914_new_n233_; 
wire u2_u0__abc_73914_new_n235_; 
wire u2_u0__abc_73914_new_n237_; 
wire u2_u0__abc_73914_new_n238_; 
wire u2_u0__abc_73914_new_n239_; 
wire u2_u0__abc_73914_new_n240_; 
wire u2_u0__abc_73914_new_n242_; 
wire u2_u0__abc_73914_new_n244_; 
wire u2_u0__abc_73914_new_n246_; 
wire u2_u0__abc_73914_new_n248_; 
wire u2_u0__abc_73914_new_n250_; 
wire u2_u0__abc_73914_new_n252_; 
wire u2_u0__abc_73914_new_n254_; 
wire u2_u0__abc_73914_new_n256_; 
wire u2_u0__abc_73914_new_n258_; 
wire u2_u0__abc_73914_new_n260_; 
wire u2_u0__abc_73914_new_n262_; 
wire u2_u0__abc_73914_new_n264_; 
wire u2_u0__abc_73914_new_n266_; 
wire u2_u0__abc_73914_new_n267_; 
wire u2_u0__abc_73914_new_n268_; 
wire u2_u0__abc_73914_new_n269_; 
wire u2_u0__abc_73914_new_n270_; 
wire u2_u0__abc_73914_new_n271_; 
wire u2_u0__abc_73914_new_n272_; 
wire u2_u0__abc_73914_new_n273_; 
wire u2_u0__abc_73914_new_n274_; 
wire u2_u0__abc_73914_new_n275_; 
wire u2_u0__abc_73914_new_n276_; 
wire u2_u0__abc_73914_new_n277_; 
wire u2_u0__abc_73914_new_n278_; 
wire u2_u0__abc_73914_new_n279_; 
wire u2_u0__abc_73914_new_n280_; 
wire u2_u0__abc_73914_new_n281_; 
wire u2_u0__abc_73914_new_n282_; 
wire u2_u0__abc_73914_new_n283_; 
wire u2_u0__abc_73914_new_n284_; 
wire u2_u0__abc_73914_new_n285_; 
wire u2_u0__abc_73914_new_n286_; 
wire u2_u0__abc_73914_new_n287_; 
wire u2_u0__abc_73914_new_n288_; 
wire u2_u0__abc_73914_new_n289_; 
wire u2_u0__abc_73914_new_n290_; 
wire u2_u0__abc_73914_new_n291_; 
wire u2_u0__abc_73914_new_n292_; 
wire u2_u0__abc_73914_new_n293_; 
wire u2_u0__abc_73914_new_n294_; 
wire u2_u0__abc_73914_new_n295_; 
wire u2_u0__abc_73914_new_n296_; 
wire u2_u0__abc_73914_new_n297_; 
wire u2_u0__abc_73914_new_n298_; 
wire u2_u0__abc_73914_new_n299_; 
wire u2_u0__abc_73914_new_n300_; 
wire u2_u0__abc_73914_new_n301_; 
wire u2_u0__abc_73914_new_n302_; 
wire u2_u0__abc_73914_new_n303_; 
wire u2_u0__abc_73914_new_n304_; 
wire u2_u0__abc_73914_new_n305_; 
wire u2_u0__abc_73914_new_n306_; 
wire u2_u0__abc_73914_new_n307_; 
wire u2_u0__abc_73914_new_n308_; 
wire u2_u0__abc_73914_new_n309_; 
wire u2_u0__abc_73914_new_n310_; 
wire u2_u0__abc_73914_new_n311_; 
wire u2_u0__abc_73914_new_n312_; 
wire u2_u0__abc_73914_new_n313_; 
wire u2_u0__abc_73914_new_n314_; 
wire u2_u0__abc_73914_new_n315_; 
wire u2_u0__abc_73914_new_n316_; 
wire u2_u0__abc_73914_new_n317_; 
wire u2_u0__abc_73914_new_n318_; 
wire u2_u0__abc_73914_new_n319_; 
wire u2_u0__abc_73914_new_n320_; 
wire u2_u0__abc_73914_new_n321_; 
wire u2_u0__abc_73914_new_n322_; 
wire u2_u0__abc_73914_new_n323_; 
wire u2_u0__abc_73914_new_n324_; 
wire u2_u0__abc_73914_new_n325_; 
wire u2_u0__abc_73914_new_n326_; 
wire u2_u0__abc_73914_new_n327_; 
wire u2_u0__abc_73914_new_n328_; 
wire u2_u0__abc_73914_new_n329_; 
wire u2_u0__abc_73914_new_n330_; 
wire u2_u0__abc_73914_new_n331_; 
wire u2_u0__abc_73914_new_n332_; 
wire u2_u0__abc_73914_new_n333_; 
wire u2_u0__abc_73914_new_n334_; 
wire u2_u0__abc_73914_new_n335_; 
wire u2_u0__abc_73914_new_n336_; 
wire u2_u0__abc_73914_new_n337_; 
wire u2_u0__abc_73914_new_n338_; 
wire u2_u0__abc_73914_new_n339_; 
wire u2_u0__abc_73914_new_n340_; 
wire u2_u0__abc_73914_new_n341_; 
wire u2_u0__abc_73914_new_n342_; 
wire u2_u0__abc_73914_new_n343_; 
wire u2_u0__abc_73914_new_n344_; 
wire u2_u0__abc_73914_new_n345_; 
wire u2_u0__abc_73914_new_n346_; 
wire u2_u0__abc_73914_new_n347_; 
wire u2_u0__abc_73914_new_n348_; 
wire u2_u0__abc_73914_new_n349_; 
wire u2_u0__abc_73914_new_n350_; 
wire u2_u0__abc_73914_new_n351_; 
wire u2_u0__abc_73914_new_n352_; 
wire u2_u0__abc_73914_new_n353_; 
wire u2_u0__abc_73914_new_n354_; 
wire u2_u0__abc_73914_new_n355_; 
wire u2_u0__abc_73914_new_n356_; 
wire u2_u0__abc_73914_new_n357_; 
wire u2_u0__abc_73914_new_n358_; 
wire u2_u0__abc_73914_new_n359_; 
wire u2_u0__abc_73914_new_n360_; 
wire u2_u0__abc_73914_new_n361_; 
wire u2_u0__abc_73914_new_n362_; 
wire u2_u0__abc_73914_new_n363_; 
wire u2_u0__abc_73914_new_n364_; 
wire u2_u0__abc_73914_new_n365_; 
wire u2_u0__abc_73914_new_n366_; 
wire u2_u0__abc_73914_new_n367_; 
wire u2_u0__abc_73914_new_n368_; 
wire u2_u0__abc_73914_new_n369_; 
wire u2_u0__abc_73914_new_n370_; 
wire u2_u0__abc_73914_new_n371_; 
wire u2_u0__abc_73914_new_n372_; 
wire u2_u0__abc_73914_new_n373_; 
wire u2_u0__abc_73914_new_n374_; 
wire u2_u0__abc_73914_new_n375_; 
wire u2_u0__abc_73914_new_n376_; 
wire u2_u0__abc_73914_new_n377_; 
wire u2_u0__abc_73914_new_n378_; 
wire u2_u0__abc_73914_new_n379_; 
wire u2_u0__abc_73914_new_n380_; 
wire u2_u0__abc_73914_new_n381_; 
wire u2_u0__abc_73914_new_n382_; 
wire u2_u0__abc_73914_new_n383_; 
wire u2_u0__abc_73914_new_n384_; 
wire u2_u0__abc_73914_new_n385_; 
wire u2_u0__abc_73914_new_n386_; 
wire u2_u0__abc_73914_new_n387_; 
wire u2_u0__abc_73914_new_n388_; 
wire u2_u0__abc_73914_new_n389_; 
wire u2_u0__abc_73914_new_n390_; 
wire u2_u0__abc_73914_new_n391_; 
wire u2_u0__abc_73914_new_n392_; 
wire u2_u0__abc_73914_new_n393_; 
wire u2_u0__abc_73914_new_n394_; 
wire u2_u0__abc_73914_new_n395_; 
wire u2_u0__abc_73914_new_n396_; 
wire u2_u0__abc_73914_new_n398_; 
wire u2_u0__abc_73914_new_n399_; 
wire u2_u0__abc_73914_new_n400_; 
wire u2_u0__abc_73914_new_n401_; 
wire u2_u0__abc_73914_new_n402_; 
wire u2_u0__abc_73914_new_n404_; 
wire u2_u0__abc_73914_new_n405_; 
wire u2_u0__abc_73914_new_n406_; 
wire u2_u0__abc_73914_new_n407_; 
wire u2_u0__abc_73914_new_n409_; 
wire u2_u0__abc_73914_new_n410_; 
wire u2_u0__abc_73914_new_n411_; 
wire u2_u0__abc_73914_new_n415_; 
wire u2_u0__abc_73914_new_n416_; 
wire u2_u0__abc_73914_new_n418_; 
wire u2_u0__abc_73914_new_n419_; 
wire u2_u0_b0_last_row_0_; 
wire u2_u0_b0_last_row_10_; 
wire u2_u0_b0_last_row_11_; 
wire u2_u0_b0_last_row_12_; 
wire u2_u0_b0_last_row_1_; 
wire u2_u0_b0_last_row_2_; 
wire u2_u0_b0_last_row_3_; 
wire u2_u0_b0_last_row_4_; 
wire u2_u0_b0_last_row_5_; 
wire u2_u0_b0_last_row_6_; 
wire u2_u0_b0_last_row_7_; 
wire u2_u0_b0_last_row_8_; 
wire u2_u0_b0_last_row_9_; 
wire u2_u0_b1_last_row_0_; 
wire u2_u0_b1_last_row_10_; 
wire u2_u0_b1_last_row_11_; 
wire u2_u0_b1_last_row_12_; 
wire u2_u0_b1_last_row_1_; 
wire u2_u0_b1_last_row_2_; 
wire u2_u0_b1_last_row_3_; 
wire u2_u0_b1_last_row_4_; 
wire u2_u0_b1_last_row_5_; 
wire u2_u0_b1_last_row_6_; 
wire u2_u0_b1_last_row_7_; 
wire u2_u0_b1_last_row_8_; 
wire u2_u0_b1_last_row_9_; 
wire u2_u0_b2_last_row_0_; 
wire u2_u0_b2_last_row_10_; 
wire u2_u0_b2_last_row_11_; 
wire u2_u0_b2_last_row_12_; 
wire u2_u0_b2_last_row_1_; 
wire u2_u0_b2_last_row_2_; 
wire u2_u0_b2_last_row_3_; 
wire u2_u0_b2_last_row_4_; 
wire u2_u0_b2_last_row_5_; 
wire u2_u0_b2_last_row_6_; 
wire u2_u0_b2_last_row_7_; 
wire u2_u0_b2_last_row_8_; 
wire u2_u0_b2_last_row_9_; 
wire u2_u0_b3_last_row_0_; 
wire u2_u0_b3_last_row_10_; 
wire u2_u0_b3_last_row_11_; 
wire u2_u0_b3_last_row_12_; 
wire u2_u0_b3_last_row_1_; 
wire u2_u0_b3_last_row_2_; 
wire u2_u0_b3_last_row_3_; 
wire u2_u0_b3_last_row_4_; 
wire u2_u0_b3_last_row_5_; 
wire u2_u0_b3_last_row_6_; 
wire u2_u0_b3_last_row_7_; 
wire u2_u0_b3_last_row_8_; 
wire u2_u0_b3_last_row_9_; 
wire u2_u0_bank0_open; 
wire u2_u0_bank1_open; 
wire u2_u0_bank2_open; 
wire u2_u0_bank3_open; 
wire u2_u1__0b0_last_row_12_0__0_; 
wire u2_u1__0b0_last_row_12_0__10_; 
wire u2_u1__0b0_last_row_12_0__11_; 
wire u2_u1__0b0_last_row_12_0__12_; 
wire u2_u1__0b0_last_row_12_0__1_; 
wire u2_u1__0b0_last_row_12_0__2_; 
wire u2_u1__0b0_last_row_12_0__3_; 
wire u2_u1__0b0_last_row_12_0__4_; 
wire u2_u1__0b0_last_row_12_0__5_; 
wire u2_u1__0b0_last_row_12_0__6_; 
wire u2_u1__0b0_last_row_12_0__7_; 
wire u2_u1__0b0_last_row_12_0__8_; 
wire u2_u1__0b0_last_row_12_0__9_; 
wire u2_u1__0b1_last_row_12_0__0_; 
wire u2_u1__0b1_last_row_12_0__10_; 
wire u2_u1__0b1_last_row_12_0__11_; 
wire u2_u1__0b1_last_row_12_0__12_; 
wire u2_u1__0b1_last_row_12_0__1_; 
wire u2_u1__0b1_last_row_12_0__2_; 
wire u2_u1__0b1_last_row_12_0__3_; 
wire u2_u1__0b1_last_row_12_0__4_; 
wire u2_u1__0b1_last_row_12_0__5_; 
wire u2_u1__0b1_last_row_12_0__6_; 
wire u2_u1__0b1_last_row_12_0__7_; 
wire u2_u1__0b1_last_row_12_0__8_; 
wire u2_u1__0b1_last_row_12_0__9_; 
wire u2_u1__0b2_last_row_12_0__0_; 
wire u2_u1__0b2_last_row_12_0__10_; 
wire u2_u1__0b2_last_row_12_0__11_; 
wire u2_u1__0b2_last_row_12_0__12_; 
wire u2_u1__0b2_last_row_12_0__1_; 
wire u2_u1__0b2_last_row_12_0__2_; 
wire u2_u1__0b2_last_row_12_0__3_; 
wire u2_u1__0b2_last_row_12_0__4_; 
wire u2_u1__0b2_last_row_12_0__5_; 
wire u2_u1__0b2_last_row_12_0__6_; 
wire u2_u1__0b2_last_row_12_0__7_; 
wire u2_u1__0b2_last_row_12_0__8_; 
wire u2_u1__0b2_last_row_12_0__9_; 
wire u2_u1__0b3_last_row_12_0__0_; 
wire u2_u1__0b3_last_row_12_0__10_; 
wire u2_u1__0b3_last_row_12_0__11_; 
wire u2_u1__0b3_last_row_12_0__12_; 
wire u2_u1__0b3_last_row_12_0__1_; 
wire u2_u1__0b3_last_row_12_0__2_; 
wire u2_u1__0b3_last_row_12_0__3_; 
wire u2_u1__0b3_last_row_12_0__4_; 
wire u2_u1__0b3_last_row_12_0__5_; 
wire u2_u1__0b3_last_row_12_0__6_; 
wire u2_u1__0b3_last_row_12_0__7_; 
wire u2_u1__0b3_last_row_12_0__8_; 
wire u2_u1__0b3_last_row_12_0__9_; 
wire u2_u1__0bank0_open_0_0_; 
wire u2_u1__0bank1_open_0_0_; 
wire u2_u1__0bank2_open_0_0_; 
wire u2_u1__0bank3_open_0_0_; 
wire u2_u1__abc_73914_auto_rtlil_cc_1942_NotGate_71538; 
wire u2_u1__abc_73914_new_n136_; 
wire u2_u1__abc_73914_new_n137_; 
wire u2_u1__abc_73914_new_n138_; 
wire u2_u1__abc_73914_new_n139_; 
wire u2_u1__abc_73914_new_n140_; 
wire u2_u1__abc_73914_new_n141_; 
wire u2_u1__abc_73914_new_n143_; 
wire u2_u1__abc_73914_new_n144_; 
wire u2_u1__abc_73914_new_n146_; 
wire u2_u1__abc_73914_new_n147_; 
wire u2_u1__abc_73914_new_n149_; 
wire u2_u1__abc_73914_new_n150_; 
wire u2_u1__abc_73914_new_n152_; 
wire u2_u1__abc_73914_new_n153_; 
wire u2_u1__abc_73914_new_n155_; 
wire u2_u1__abc_73914_new_n156_; 
wire u2_u1__abc_73914_new_n158_; 
wire u2_u1__abc_73914_new_n159_; 
wire u2_u1__abc_73914_new_n161_; 
wire u2_u1__abc_73914_new_n162_; 
wire u2_u1__abc_73914_new_n164_; 
wire u2_u1__abc_73914_new_n165_; 
wire u2_u1__abc_73914_new_n167_; 
wire u2_u1__abc_73914_new_n168_; 
wire u2_u1__abc_73914_new_n170_; 
wire u2_u1__abc_73914_new_n171_; 
wire u2_u1__abc_73914_new_n173_; 
wire u2_u1__abc_73914_new_n174_; 
wire u2_u1__abc_73914_new_n176_; 
wire u2_u1__abc_73914_new_n177_; 
wire u2_u1__abc_73914_new_n179_; 
wire u2_u1__abc_73914_new_n180_; 
wire u2_u1__abc_73914_new_n181_; 
wire u2_u1__abc_73914_new_n182_; 
wire u2_u1__abc_73914_new_n184_; 
wire u2_u1__abc_73914_new_n186_; 
wire u2_u1__abc_73914_new_n188_; 
wire u2_u1__abc_73914_new_n190_; 
wire u2_u1__abc_73914_new_n192_; 
wire u2_u1__abc_73914_new_n194_; 
wire u2_u1__abc_73914_new_n196_; 
wire u2_u1__abc_73914_new_n198_; 
wire u2_u1__abc_73914_new_n200_; 
wire u2_u1__abc_73914_new_n202_; 
wire u2_u1__abc_73914_new_n204_; 
wire u2_u1__abc_73914_new_n206_; 
wire u2_u1__abc_73914_new_n208_; 
wire u2_u1__abc_73914_new_n209_; 
wire u2_u1__abc_73914_new_n210_; 
wire u2_u1__abc_73914_new_n211_; 
wire u2_u1__abc_73914_new_n213_; 
wire u2_u1__abc_73914_new_n215_; 
wire u2_u1__abc_73914_new_n217_; 
wire u2_u1__abc_73914_new_n219_; 
wire u2_u1__abc_73914_new_n221_; 
wire u2_u1__abc_73914_new_n223_; 
wire u2_u1__abc_73914_new_n225_; 
wire u2_u1__abc_73914_new_n227_; 
wire u2_u1__abc_73914_new_n229_; 
wire u2_u1__abc_73914_new_n231_; 
wire u2_u1__abc_73914_new_n233_; 
wire u2_u1__abc_73914_new_n235_; 
wire u2_u1__abc_73914_new_n237_; 
wire u2_u1__abc_73914_new_n238_; 
wire u2_u1__abc_73914_new_n239_; 
wire u2_u1__abc_73914_new_n240_; 
wire u2_u1__abc_73914_new_n242_; 
wire u2_u1__abc_73914_new_n244_; 
wire u2_u1__abc_73914_new_n246_; 
wire u2_u1__abc_73914_new_n248_; 
wire u2_u1__abc_73914_new_n250_; 
wire u2_u1__abc_73914_new_n252_; 
wire u2_u1__abc_73914_new_n254_; 
wire u2_u1__abc_73914_new_n256_; 
wire u2_u1__abc_73914_new_n258_; 
wire u2_u1__abc_73914_new_n260_; 
wire u2_u1__abc_73914_new_n262_; 
wire u2_u1__abc_73914_new_n264_; 
wire u2_u1__abc_73914_new_n266_; 
wire u2_u1__abc_73914_new_n267_; 
wire u2_u1__abc_73914_new_n268_; 
wire u2_u1__abc_73914_new_n269_; 
wire u2_u1__abc_73914_new_n270_; 
wire u2_u1__abc_73914_new_n271_; 
wire u2_u1__abc_73914_new_n272_; 
wire u2_u1__abc_73914_new_n273_; 
wire u2_u1__abc_73914_new_n274_; 
wire u2_u1__abc_73914_new_n275_; 
wire u2_u1__abc_73914_new_n276_; 
wire u2_u1__abc_73914_new_n277_; 
wire u2_u1__abc_73914_new_n278_; 
wire u2_u1__abc_73914_new_n279_; 
wire u2_u1__abc_73914_new_n280_; 
wire u2_u1__abc_73914_new_n281_; 
wire u2_u1__abc_73914_new_n282_; 
wire u2_u1__abc_73914_new_n283_; 
wire u2_u1__abc_73914_new_n284_; 
wire u2_u1__abc_73914_new_n285_; 
wire u2_u1__abc_73914_new_n286_; 
wire u2_u1__abc_73914_new_n287_; 
wire u2_u1__abc_73914_new_n288_; 
wire u2_u1__abc_73914_new_n289_; 
wire u2_u1__abc_73914_new_n290_; 
wire u2_u1__abc_73914_new_n291_; 
wire u2_u1__abc_73914_new_n292_; 
wire u2_u1__abc_73914_new_n293_; 
wire u2_u1__abc_73914_new_n294_; 
wire u2_u1__abc_73914_new_n295_; 
wire u2_u1__abc_73914_new_n296_; 
wire u2_u1__abc_73914_new_n297_; 
wire u2_u1__abc_73914_new_n298_; 
wire u2_u1__abc_73914_new_n299_; 
wire u2_u1__abc_73914_new_n300_; 
wire u2_u1__abc_73914_new_n301_; 
wire u2_u1__abc_73914_new_n302_; 
wire u2_u1__abc_73914_new_n303_; 
wire u2_u1__abc_73914_new_n304_; 
wire u2_u1__abc_73914_new_n305_; 
wire u2_u1__abc_73914_new_n306_; 
wire u2_u1__abc_73914_new_n307_; 
wire u2_u1__abc_73914_new_n308_; 
wire u2_u1__abc_73914_new_n309_; 
wire u2_u1__abc_73914_new_n310_; 
wire u2_u1__abc_73914_new_n311_; 
wire u2_u1__abc_73914_new_n312_; 
wire u2_u1__abc_73914_new_n313_; 
wire u2_u1__abc_73914_new_n314_; 
wire u2_u1__abc_73914_new_n315_; 
wire u2_u1__abc_73914_new_n316_; 
wire u2_u1__abc_73914_new_n317_; 
wire u2_u1__abc_73914_new_n318_; 
wire u2_u1__abc_73914_new_n319_; 
wire u2_u1__abc_73914_new_n320_; 
wire u2_u1__abc_73914_new_n321_; 
wire u2_u1__abc_73914_new_n322_; 
wire u2_u1__abc_73914_new_n323_; 
wire u2_u1__abc_73914_new_n324_; 
wire u2_u1__abc_73914_new_n325_; 
wire u2_u1__abc_73914_new_n326_; 
wire u2_u1__abc_73914_new_n327_; 
wire u2_u1__abc_73914_new_n328_; 
wire u2_u1__abc_73914_new_n329_; 
wire u2_u1__abc_73914_new_n330_; 
wire u2_u1__abc_73914_new_n331_; 
wire u2_u1__abc_73914_new_n332_; 
wire u2_u1__abc_73914_new_n333_; 
wire u2_u1__abc_73914_new_n334_; 
wire u2_u1__abc_73914_new_n335_; 
wire u2_u1__abc_73914_new_n336_; 
wire u2_u1__abc_73914_new_n337_; 
wire u2_u1__abc_73914_new_n338_; 
wire u2_u1__abc_73914_new_n339_; 
wire u2_u1__abc_73914_new_n340_; 
wire u2_u1__abc_73914_new_n341_; 
wire u2_u1__abc_73914_new_n342_; 
wire u2_u1__abc_73914_new_n343_; 
wire u2_u1__abc_73914_new_n344_; 
wire u2_u1__abc_73914_new_n345_; 
wire u2_u1__abc_73914_new_n346_; 
wire u2_u1__abc_73914_new_n347_; 
wire u2_u1__abc_73914_new_n348_; 
wire u2_u1__abc_73914_new_n349_; 
wire u2_u1__abc_73914_new_n350_; 
wire u2_u1__abc_73914_new_n351_; 
wire u2_u1__abc_73914_new_n352_; 
wire u2_u1__abc_73914_new_n353_; 
wire u2_u1__abc_73914_new_n354_; 
wire u2_u1__abc_73914_new_n355_; 
wire u2_u1__abc_73914_new_n356_; 
wire u2_u1__abc_73914_new_n357_; 
wire u2_u1__abc_73914_new_n358_; 
wire u2_u1__abc_73914_new_n359_; 
wire u2_u1__abc_73914_new_n360_; 
wire u2_u1__abc_73914_new_n361_; 
wire u2_u1__abc_73914_new_n362_; 
wire u2_u1__abc_73914_new_n363_; 
wire u2_u1__abc_73914_new_n364_; 
wire u2_u1__abc_73914_new_n365_; 
wire u2_u1__abc_73914_new_n366_; 
wire u2_u1__abc_73914_new_n367_; 
wire u2_u1__abc_73914_new_n368_; 
wire u2_u1__abc_73914_new_n369_; 
wire u2_u1__abc_73914_new_n370_; 
wire u2_u1__abc_73914_new_n371_; 
wire u2_u1__abc_73914_new_n372_; 
wire u2_u1__abc_73914_new_n373_; 
wire u2_u1__abc_73914_new_n374_; 
wire u2_u1__abc_73914_new_n375_; 
wire u2_u1__abc_73914_new_n376_; 
wire u2_u1__abc_73914_new_n377_; 
wire u2_u1__abc_73914_new_n378_; 
wire u2_u1__abc_73914_new_n379_; 
wire u2_u1__abc_73914_new_n380_; 
wire u2_u1__abc_73914_new_n381_; 
wire u2_u1__abc_73914_new_n382_; 
wire u2_u1__abc_73914_new_n383_; 
wire u2_u1__abc_73914_new_n384_; 
wire u2_u1__abc_73914_new_n385_; 
wire u2_u1__abc_73914_new_n386_; 
wire u2_u1__abc_73914_new_n387_; 
wire u2_u1__abc_73914_new_n388_; 
wire u2_u1__abc_73914_new_n389_; 
wire u2_u1__abc_73914_new_n390_; 
wire u2_u1__abc_73914_new_n391_; 
wire u2_u1__abc_73914_new_n392_; 
wire u2_u1__abc_73914_new_n393_; 
wire u2_u1__abc_73914_new_n394_; 
wire u2_u1__abc_73914_new_n395_; 
wire u2_u1__abc_73914_new_n396_; 
wire u2_u1__abc_73914_new_n398_; 
wire u2_u1__abc_73914_new_n399_; 
wire u2_u1__abc_73914_new_n400_; 
wire u2_u1__abc_73914_new_n401_; 
wire u2_u1__abc_73914_new_n402_; 
wire u2_u1__abc_73914_new_n404_; 
wire u2_u1__abc_73914_new_n405_; 
wire u2_u1__abc_73914_new_n406_; 
wire u2_u1__abc_73914_new_n407_; 
wire u2_u1__abc_73914_new_n409_; 
wire u2_u1__abc_73914_new_n410_; 
wire u2_u1__abc_73914_new_n411_; 
wire u2_u1__abc_73914_new_n415_; 
wire u2_u1__abc_73914_new_n416_; 
wire u2_u1__abc_73914_new_n418_; 
wire u2_u1__abc_73914_new_n419_; 
wire u2_u1_b0_last_row_0_; 
wire u2_u1_b0_last_row_10_; 
wire u2_u1_b0_last_row_11_; 
wire u2_u1_b0_last_row_12_; 
wire u2_u1_b0_last_row_1_; 
wire u2_u1_b0_last_row_2_; 
wire u2_u1_b0_last_row_3_; 
wire u2_u1_b0_last_row_4_; 
wire u2_u1_b0_last_row_5_; 
wire u2_u1_b0_last_row_6_; 
wire u2_u1_b0_last_row_7_; 
wire u2_u1_b0_last_row_8_; 
wire u2_u1_b0_last_row_9_; 
wire u2_u1_b1_last_row_0_; 
wire u2_u1_b1_last_row_10_; 
wire u2_u1_b1_last_row_11_; 
wire u2_u1_b1_last_row_12_; 
wire u2_u1_b1_last_row_1_; 
wire u2_u1_b1_last_row_2_; 
wire u2_u1_b1_last_row_3_; 
wire u2_u1_b1_last_row_4_; 
wire u2_u1_b1_last_row_5_; 
wire u2_u1_b1_last_row_6_; 
wire u2_u1_b1_last_row_7_; 
wire u2_u1_b1_last_row_8_; 
wire u2_u1_b1_last_row_9_; 
wire u2_u1_b2_last_row_0_; 
wire u2_u1_b2_last_row_10_; 
wire u2_u1_b2_last_row_11_; 
wire u2_u1_b2_last_row_12_; 
wire u2_u1_b2_last_row_1_; 
wire u2_u1_b2_last_row_2_; 
wire u2_u1_b2_last_row_3_; 
wire u2_u1_b2_last_row_4_; 
wire u2_u1_b2_last_row_5_; 
wire u2_u1_b2_last_row_6_; 
wire u2_u1_b2_last_row_7_; 
wire u2_u1_b2_last_row_8_; 
wire u2_u1_b2_last_row_9_; 
wire u2_u1_b3_last_row_0_; 
wire u2_u1_b3_last_row_10_; 
wire u2_u1_b3_last_row_11_; 
wire u2_u1_b3_last_row_12_; 
wire u2_u1_b3_last_row_1_; 
wire u2_u1_b3_last_row_2_; 
wire u2_u1_b3_last_row_3_; 
wire u2_u1_b3_last_row_4_; 
wire u2_u1_b3_last_row_5_; 
wire u2_u1_b3_last_row_6_; 
wire u2_u1_b3_last_row_7_; 
wire u2_u1_b3_last_row_8_; 
wire u2_u1_b3_last_row_9_; 
wire u2_u1_bank0_open; 
wire u2_u1_bank1_open; 
wire u2_u1_bank2_open; 
wire u2_u1_bank3_open; 
wire u3__0byte0_7_0__0_; 
wire u3__0byte0_7_0__1_; 
wire u3__0byte0_7_0__2_; 
wire u3__0byte0_7_0__3_; 
wire u3__0byte0_7_0__4_; 
wire u3__0byte0_7_0__5_; 
wire u3__0byte0_7_0__6_; 
wire u3__0byte0_7_0__7_; 
wire u3__0byte1_7_0__0_; 
wire u3__0byte1_7_0__1_; 
wire u3__0byte1_7_0__2_; 
wire u3__0byte1_7_0__3_; 
wire u3__0byte1_7_0__4_; 
wire u3__0byte1_7_0__5_; 
wire u3__0byte1_7_0__6_; 
wire u3__0byte1_7_0__7_; 
wire u3__0byte2_7_0__0_; 
wire u3__0byte2_7_0__1_; 
wire u3__0byte2_7_0__2_; 
wire u3__0byte2_7_0__3_; 
wire u3__0byte2_7_0__4_; 
wire u3__0byte2_7_0__5_; 
wire u3__0byte2_7_0__6_; 
wire u3__0byte2_7_0__7_; 
wire u3__0mc_data_o_31_0__0_; 
wire u3__0mc_data_o_31_0__10_; 
wire u3__0mc_data_o_31_0__11_; 
wire u3__0mc_data_o_31_0__12_; 
wire u3__0mc_data_o_31_0__13_; 
wire u3__0mc_data_o_31_0__14_; 
wire u3__0mc_data_o_31_0__15_; 
wire u3__0mc_data_o_31_0__16_; 
wire u3__0mc_data_o_31_0__17_; 
wire u3__0mc_data_o_31_0__18_; 
wire u3__0mc_data_o_31_0__19_; 
wire u3__0mc_data_o_31_0__1_; 
wire u3__0mc_data_o_31_0__20_; 
wire u3__0mc_data_o_31_0__21_; 
wire u3__0mc_data_o_31_0__22_; 
wire u3__0mc_data_o_31_0__23_; 
wire u3__0mc_data_o_31_0__24_; 
wire u3__0mc_data_o_31_0__25_; 
wire u3__0mc_data_o_31_0__26_; 
wire u3__0mc_data_o_31_0__27_; 
wire u3__0mc_data_o_31_0__28_; 
wire u3__0mc_data_o_31_0__29_; 
wire u3__0mc_data_o_31_0__2_; 
wire u3__0mc_data_o_31_0__30_; 
wire u3__0mc_data_o_31_0__31_; 
wire u3__0mc_data_o_31_0__3_; 
wire u3__0mc_data_o_31_0__4_; 
wire u3__0mc_data_o_31_0__5_; 
wire u3__0mc_data_o_31_0__6_; 
wire u3__0mc_data_o_31_0__7_; 
wire u3__0mc_data_o_31_0__8_; 
wire u3__0mc_data_o_31_0__9_; 
wire u3__0mc_dp_o_3_0__0_; 
wire u3__0mc_dp_o_3_0__1_; 
wire u3__0mc_dp_o_3_0__2_; 
wire u3__0mc_dp_o_3_0__3_; 
wire u3__abc_73372_new_n275_; 
wire u3__abc_73372_new_n276_; 
wire u3__abc_73372_new_n277_; 
wire u3__abc_73372_new_n278_; 
wire u3__abc_73372_new_n279_; 
wire u3__abc_73372_new_n280_; 
wire u3__abc_73372_new_n281_; 
wire u3__abc_73372_new_n282_; 
wire u3__abc_73372_new_n283_; 
wire u3__abc_73372_new_n284_; 
wire u3__abc_73372_new_n285_; 
wire u3__abc_73372_new_n286_; 
wire u3__abc_73372_new_n288_; 
wire u3__abc_73372_new_n289_; 
wire u3__abc_73372_new_n290_; 
wire u3__abc_73372_new_n291_; 
wire u3__abc_73372_new_n292_; 
wire u3__abc_73372_new_n293_; 
wire u3__abc_73372_new_n294_; 
wire u3__abc_73372_new_n295_; 
wire u3__abc_73372_new_n297_; 
wire u3__abc_73372_new_n298_; 
wire u3__abc_73372_new_n299_; 
wire u3__abc_73372_new_n300_; 
wire u3__abc_73372_new_n301_; 
wire u3__abc_73372_new_n302_; 
wire u3__abc_73372_new_n303_; 
wire u3__abc_73372_new_n304_; 
wire u3__abc_73372_new_n306_; 
wire u3__abc_73372_new_n307_; 
wire u3__abc_73372_new_n308_; 
wire u3__abc_73372_new_n309_; 
wire u3__abc_73372_new_n310_; 
wire u3__abc_73372_new_n311_; 
wire u3__abc_73372_new_n312_; 
wire u3__abc_73372_new_n313_; 
wire u3__abc_73372_new_n315_; 
wire u3__abc_73372_new_n316_; 
wire u3__abc_73372_new_n318_; 
wire u3__abc_73372_new_n319_; 
wire u3__abc_73372_new_n321_; 
wire u3__abc_73372_new_n322_; 
wire u3__abc_73372_new_n324_; 
wire u3__abc_73372_new_n325_; 
wire u3__abc_73372_new_n327_; 
wire u3__abc_73372_new_n328_; 
wire u3__abc_73372_new_n330_; 
wire u3__abc_73372_new_n331_; 
wire u3__abc_73372_new_n333_; 
wire u3__abc_73372_new_n334_; 
wire u3__abc_73372_new_n336_; 
wire u3__abc_73372_new_n337_; 
wire u3__abc_73372_new_n339_; 
wire u3__abc_73372_new_n340_; 
wire u3__abc_73372_new_n341_; 
wire u3__abc_73372_new_n342_; 
wire u3__abc_73372_new_n343_; 
wire u3__abc_73372_new_n344_; 
wire u3__abc_73372_new_n345_; 
wire u3__abc_73372_new_n346_; 
wire u3__abc_73372_new_n347_; 
wire u3__abc_73372_new_n348_; 
wire u3__abc_73372_new_n349_; 
wire u3__abc_73372_new_n351_; 
wire u3__abc_73372_new_n352_; 
wire u3__abc_73372_new_n353_; 
wire u3__abc_73372_new_n354_; 
wire u3__abc_73372_new_n356_; 
wire u3__abc_73372_new_n357_; 
wire u3__abc_73372_new_n358_; 
wire u3__abc_73372_new_n359_; 
wire u3__abc_73372_new_n361_; 
wire u3__abc_73372_new_n362_; 
wire u3__abc_73372_new_n363_; 
wire u3__abc_73372_new_n364_; 
wire u3__abc_73372_new_n366_; 
wire u3__abc_73372_new_n367_; 
wire u3__abc_73372_new_n368_; 
wire u3__abc_73372_new_n369_; 
wire u3__abc_73372_new_n371_; 
wire u3__abc_73372_new_n372_; 
wire u3__abc_73372_new_n373_; 
wire u3__abc_73372_new_n374_; 
wire u3__abc_73372_new_n376_; 
wire u3__abc_73372_new_n377_; 
wire u3__abc_73372_new_n378_; 
wire u3__abc_73372_new_n379_; 
wire u3__abc_73372_new_n381_; 
wire u3__abc_73372_new_n382_; 
wire u3__abc_73372_new_n383_; 
wire u3__abc_73372_new_n384_; 
wire u3__abc_73372_new_n386_; 
wire u3__abc_73372_new_n388_; 
wire u3__abc_73372_new_n390_; 
wire u3__abc_73372_new_n392_; 
wire u3__abc_73372_new_n394_; 
wire u3__abc_73372_new_n396_; 
wire u3__abc_73372_new_n398_; 
wire u3__abc_73372_new_n400_; 
wire u3__abc_73372_new_n402_; 
wire u3__abc_73372_new_n403_; 
wire u3__abc_73372_new_n405_; 
wire u3__abc_73372_new_n406_; 
wire u3__abc_73372_new_n408_; 
wire u3__abc_73372_new_n409_; 
wire u3__abc_73372_new_n411_; 
wire u3__abc_73372_new_n412_; 
wire u3__abc_73372_new_n414_; 
wire u3__abc_73372_new_n415_; 
wire u3__abc_73372_new_n417_; 
wire u3__abc_73372_new_n418_; 
wire u3__abc_73372_new_n420_; 
wire u3__abc_73372_new_n421_; 
wire u3__abc_73372_new_n423_; 
wire u3__abc_73372_new_n424_; 
wire u3__abc_73372_new_n426_; 
wire u3__abc_73372_new_n427_; 
wire u3__abc_73372_new_n429_; 
wire u3__abc_73372_new_n430_; 
wire u3__abc_73372_new_n432_; 
wire u3__abc_73372_new_n433_; 
wire u3__abc_73372_new_n435_; 
wire u3__abc_73372_new_n436_; 
wire u3__abc_73372_new_n438_; 
wire u3__abc_73372_new_n439_; 
wire u3__abc_73372_new_n441_; 
wire u3__abc_73372_new_n442_; 
wire u3__abc_73372_new_n444_; 
wire u3__abc_73372_new_n445_; 
wire u3__abc_73372_new_n447_; 
wire u3__abc_73372_new_n448_; 
wire u3__abc_73372_new_n450_; 
wire u3__abc_73372_new_n451_; 
wire u3__abc_73372_new_n453_; 
wire u3__abc_73372_new_n454_; 
wire u3__abc_73372_new_n456_; 
wire u3__abc_73372_new_n457_; 
wire u3__abc_73372_new_n459_; 
wire u3__abc_73372_new_n460_; 
wire u3__abc_73372_new_n462_; 
wire u3__abc_73372_new_n463_; 
wire u3__abc_73372_new_n465_; 
wire u3__abc_73372_new_n466_; 
wire u3__abc_73372_new_n468_; 
wire u3__abc_73372_new_n469_; 
wire u3__abc_73372_new_n471_; 
wire u3__abc_73372_new_n472_; 
wire u3__abc_73372_new_n474_; 
wire u3__abc_73372_new_n475_; 
wire u3__abc_73372_new_n477_; 
wire u3__abc_73372_new_n478_; 
wire u3__abc_73372_new_n480_; 
wire u3__abc_73372_new_n481_; 
wire u3__abc_73372_new_n483_; 
wire u3__abc_73372_new_n484_; 
wire u3__abc_73372_new_n486_; 
wire u3__abc_73372_new_n487_; 
wire u3__abc_73372_new_n489_; 
wire u3__abc_73372_new_n490_; 
wire u3__abc_73372_new_n492_; 
wire u3__abc_73372_new_n493_; 
wire u3__abc_73372_new_n495_; 
wire u3__abc_73372_new_n496_; 
wire u3__abc_73372_new_n498_; 
wire u3__abc_73372_new_n499_; 
wire u3__abc_73372_new_n500_; 
wire u3__abc_73372_new_n502_; 
wire u3__abc_73372_new_n503_; 
wire u3__abc_73372_new_n504_; 
wire u3__abc_73372_new_n506_; 
wire u3__abc_73372_new_n507_; 
wire u3__abc_73372_new_n508_; 
wire u3__abc_73372_new_n510_; 
wire u3__abc_73372_new_n511_; 
wire u3__abc_73372_new_n512_; 
wire u3__abc_73372_new_n514_; 
wire u3__abc_73372_new_n515_; 
wire u3__abc_73372_new_n516_; 
wire u3__abc_73372_new_n518_; 
wire u3__abc_73372_new_n519_; 
wire u3__abc_73372_new_n520_; 
wire u3__abc_73372_new_n522_; 
wire u3__abc_73372_new_n523_; 
wire u3__abc_73372_new_n524_; 
wire u3__abc_73372_new_n526_; 
wire u3__abc_73372_new_n527_; 
wire u3__abc_73372_new_n528_; 
wire u3__abc_73372_new_n530_; 
wire u3__abc_73372_new_n531_; 
wire u3__abc_73372_new_n532_; 
wire u3__abc_73372_new_n534_; 
wire u3__abc_73372_new_n535_; 
wire u3__abc_73372_new_n536_; 
wire u3__abc_73372_new_n538_; 
wire u3__abc_73372_new_n539_; 
wire u3__abc_73372_new_n540_; 
wire u3__abc_73372_new_n542_; 
wire u3__abc_73372_new_n543_; 
wire u3__abc_73372_new_n544_; 
wire u3__abc_73372_new_n546_; 
wire u3__abc_73372_new_n547_; 
wire u3__abc_73372_new_n548_; 
wire u3__abc_73372_new_n550_; 
wire u3__abc_73372_new_n551_; 
wire u3__abc_73372_new_n552_; 
wire u3__abc_73372_new_n554_; 
wire u3__abc_73372_new_n555_; 
wire u3__abc_73372_new_n556_; 
wire u3__abc_73372_new_n558_; 
wire u3__abc_73372_new_n559_; 
wire u3__abc_73372_new_n560_; 
wire u3__abc_73372_new_n562_; 
wire u3__abc_73372_new_n563_; 
wire u3__abc_73372_new_n564_; 
wire u3__abc_73372_new_n566_; 
wire u3__abc_73372_new_n567_; 
wire u3__abc_73372_new_n568_; 
wire u3__abc_73372_new_n570_; 
wire u3__abc_73372_new_n571_; 
wire u3__abc_73372_new_n572_; 
wire u3__abc_73372_new_n574_; 
wire u3__abc_73372_new_n575_; 
wire u3__abc_73372_new_n576_; 
wire u3__abc_73372_new_n578_; 
wire u3__abc_73372_new_n579_; 
wire u3__abc_73372_new_n580_; 
wire u3__abc_73372_new_n582_; 
wire u3__abc_73372_new_n583_; 
wire u3__abc_73372_new_n584_; 
wire u3__abc_73372_new_n586_; 
wire u3__abc_73372_new_n587_; 
wire u3__abc_73372_new_n588_; 
wire u3__abc_73372_new_n590_; 
wire u3__abc_73372_new_n591_; 
wire u3__abc_73372_new_n592_; 
wire u3__abc_73372_new_n594_; 
wire u3__abc_73372_new_n595_; 
wire u3__abc_73372_new_n596_; 
wire u3__abc_73372_new_n598_; 
wire u3__abc_73372_new_n599_; 
wire u3__abc_73372_new_n600_; 
wire u3__abc_73372_new_n602_; 
wire u3__abc_73372_new_n603_; 
wire u3__abc_73372_new_n604_; 
wire u3__abc_73372_new_n606_; 
wire u3__abc_73372_new_n607_; 
wire u3__abc_73372_new_n608_; 
wire u3__abc_73372_new_n610_; 
wire u3__abc_73372_new_n611_; 
wire u3__abc_73372_new_n612_; 
wire u3__abc_73372_new_n614_; 
wire u3__abc_73372_new_n615_; 
wire u3__abc_73372_new_n616_; 
wire u3__abc_73372_new_n618_; 
wire u3__abc_73372_new_n619_; 
wire u3__abc_73372_new_n620_; 
wire u3__abc_73372_new_n622_; 
wire u3__abc_73372_new_n623_; 
wire u3__abc_73372_new_n624_; 
wire u3__abc_73372_new_n626_; 
wire u3__abc_73372_new_n627_; 
wire u3__abc_73372_new_n630_; 
wire u3__abc_73372_new_n631_; 
wire u3__abc_73372_new_n632_; 
wire u3__abc_73372_new_n633_; 
wire u3__abc_73372_new_n634_; 
wire u3__abc_73372_new_n635_; 
wire u3__abc_73372_new_n636_; 
wire u3__abc_73372_new_n637_; 
wire u3__abc_73372_new_n638_; 
wire u3__abc_73372_new_n639_; 
wire u3__abc_73372_new_n640_; 
wire u3__abc_73372_new_n641_; 
wire u3__abc_73372_new_n642_; 
wire u3__abc_73372_new_n643_; 
wire u3__abc_73372_new_n644_; 
wire u3__abc_73372_new_n645_; 
wire u3__abc_73372_new_n646_; 
wire u3__abc_73372_new_n647_; 
wire u3__abc_73372_new_n648_; 
wire u3__abc_73372_new_n649_; 
wire u3__abc_73372_new_n650_; 
wire u3__abc_73372_new_n651_; 
wire u3__abc_73372_new_n652_; 
wire u3__abc_73372_new_n653_; 
wire u3__abc_73372_new_n654_; 
wire u3__abc_73372_new_n655_; 
wire u3__abc_73372_new_n656_; 
wire u3__abc_73372_new_n657_; 
wire u3__abc_73372_new_n658_; 
wire u3__abc_73372_new_n659_; 
wire u3__abc_73372_new_n660_; 
wire u3__abc_73372_new_n661_; 
wire u3__abc_73372_new_n662_; 
wire u3__abc_73372_new_n663_; 
wire u3__abc_73372_new_n664_; 
wire u3__abc_73372_new_n665_; 
wire u3__abc_73372_new_n666_; 
wire u3__abc_73372_new_n667_; 
wire u3__abc_73372_new_n668_; 
wire u3__abc_73372_new_n669_; 
wire u3__abc_73372_new_n670_; 
wire u3__abc_73372_new_n671_; 
wire u3__abc_73372_new_n672_; 
wire u3__abc_73372_new_n673_; 
wire u3__abc_73372_new_n674_; 
wire u3__abc_73372_new_n675_; 
wire u3__abc_73372_new_n676_; 
wire u3__abc_73372_new_n677_; 
wire u3__abc_73372_new_n678_; 
wire u3__abc_73372_new_n679_; 
wire u3__abc_73372_new_n680_; 
wire u3__abc_73372_new_n681_; 
wire u3__abc_73372_new_n682_; 
wire u3__abc_73372_new_n683_; 
wire u3__abc_73372_new_n684_; 
wire u3__abc_73372_new_n685_; 
wire u3__abc_73372_new_n686_; 
wire u3__abc_73372_new_n687_; 
wire u3__abc_73372_new_n688_; 
wire u3__abc_73372_new_n689_; 
wire u3__abc_73372_new_n690_; 
wire u3__abc_73372_new_n691_; 
wire u3__abc_73372_new_n692_; 
wire u3__abc_73372_new_n693_; 
wire u3__abc_73372_new_n694_; 
wire u3__abc_73372_new_n695_; 
wire u3__abc_73372_new_n696_; 
wire u3__abc_73372_new_n697_; 
wire u3__abc_73372_new_n698_; 
wire u3__abc_73372_new_n699_; 
wire u3__abc_73372_new_n700_; 
wire u3__abc_73372_new_n701_; 
wire u3__abc_73372_new_n702_; 
wire u3__abc_73372_new_n703_; 
wire u3__abc_73372_new_n704_; 
wire u3__abc_73372_new_n705_; 
wire u3__abc_73372_new_n706_; 
wire u3__abc_73372_new_n707_; 
wire u3__abc_73372_new_n708_; 
wire u3__abc_73372_new_n709_; 
wire u3__abc_73372_new_n710_; 
wire u3__abc_73372_new_n711_; 
wire u3__abc_73372_new_n712_; 
wire u3__abc_73372_new_n713_; 
wire u3__abc_73372_new_n714_; 
wire u3__abc_73372_new_n715_; 
wire u3__abc_73372_new_n716_; 
wire u3__abc_73372_new_n717_; 
wire u3__abc_73372_new_n718_; 
wire u3__abc_73372_new_n719_; 
wire u3__abc_73372_new_n720_; 
wire u3__abc_73372_new_n721_; 
wire u3__abc_73372_new_n722_; 
wire u3__abc_73372_new_n723_; 
wire u3__abc_73372_new_n724_; 
wire u3__abc_73372_new_n725_; 
wire u3__abc_73372_new_n726_; 
wire u3__abc_73372_new_n727_; 
wire u3__abc_73372_new_n728_; 
wire u3__abc_73372_new_n729_; 
wire u3_byte0_0_; 
wire u3_byte0_1_; 
wire u3_byte0_2_; 
wire u3_byte0_3_; 
wire u3_byte0_4_; 
wire u3_byte0_5_; 
wire u3_byte0_6_; 
wire u3_byte0_7_; 
wire u3_byte1_0_; 
wire u3_byte1_1_; 
wire u3_byte1_2_; 
wire u3_byte1_3_; 
wire u3_byte1_4_; 
wire u3_byte1_5_; 
wire u3_byte1_6_; 
wire u3_byte1_7_; 
wire u3_byte2_0_; 
wire u3_byte2_1_; 
wire u3_byte2_2_; 
wire u3_byte2_3_; 
wire u3_byte2_4_; 
wire u3_byte2_5_; 
wire u3_byte2_6_; 
wire u3_byte2_7_; 
wire u3_pen; 
wire u3_rd_fifo_clr; 
wire u3_rd_fifo_out_0_; 
wire u3_rd_fifo_out_10_; 
wire u3_rd_fifo_out_11_; 
wire u3_rd_fifo_out_12_; 
wire u3_rd_fifo_out_13_; 
wire u3_rd_fifo_out_14_; 
wire u3_rd_fifo_out_15_; 
wire u3_rd_fifo_out_16_; 
wire u3_rd_fifo_out_17_; 
wire u3_rd_fifo_out_18_; 
wire u3_rd_fifo_out_19_; 
wire u3_rd_fifo_out_1_; 
wire u3_rd_fifo_out_20_; 
wire u3_rd_fifo_out_21_; 
wire u3_rd_fifo_out_22_; 
wire u3_rd_fifo_out_23_; 
wire u3_rd_fifo_out_24_; 
wire u3_rd_fifo_out_25_; 
wire u3_rd_fifo_out_26_; 
wire u3_rd_fifo_out_27_; 
wire u3_rd_fifo_out_28_; 
wire u3_rd_fifo_out_29_; 
wire u3_rd_fifo_out_2_; 
wire u3_rd_fifo_out_30_; 
wire u3_rd_fifo_out_31_; 
wire u3_rd_fifo_out_32_; 
wire u3_rd_fifo_out_33_; 
wire u3_rd_fifo_out_34_; 
wire u3_rd_fifo_out_35_; 
wire u3_rd_fifo_out_3_; 
wire u3_rd_fifo_out_4_; 
wire u3_rd_fifo_out_5_; 
wire u3_rd_fifo_out_6_; 
wire u3_rd_fifo_out_7_; 
wire u3_rd_fifo_out_8_; 
wire u3_rd_fifo_out_9_; 
wire u3_re; 
wire u3_u0__0r0_35_0__0_; 
wire u3_u0__0r0_35_0__10_; 
wire u3_u0__0r0_35_0__11_; 
wire u3_u0__0r0_35_0__12_; 
wire u3_u0__0r0_35_0__13_; 
wire u3_u0__0r0_35_0__14_; 
wire u3_u0__0r0_35_0__15_; 
wire u3_u0__0r0_35_0__16_; 
wire u3_u0__0r0_35_0__17_; 
wire u3_u0__0r0_35_0__18_; 
wire u3_u0__0r0_35_0__19_; 
wire u3_u0__0r0_35_0__1_; 
wire u3_u0__0r0_35_0__20_; 
wire u3_u0__0r0_35_0__21_; 
wire u3_u0__0r0_35_0__22_; 
wire u3_u0__0r0_35_0__23_; 
wire u3_u0__0r0_35_0__24_; 
wire u3_u0__0r0_35_0__25_; 
wire u3_u0__0r0_35_0__26_; 
wire u3_u0__0r0_35_0__27_; 
wire u3_u0__0r0_35_0__28_; 
wire u3_u0__0r0_35_0__29_; 
wire u3_u0__0r0_35_0__2_; 
wire u3_u0__0r0_35_0__30_; 
wire u3_u0__0r0_35_0__31_; 
wire u3_u0__0r0_35_0__32_; 
wire u3_u0__0r0_35_0__33_; 
wire u3_u0__0r0_35_0__34_; 
wire u3_u0__0r0_35_0__35_; 
wire u3_u0__0r0_35_0__3_; 
wire u3_u0__0r0_35_0__4_; 
wire u3_u0__0r0_35_0__5_; 
wire u3_u0__0r0_35_0__6_; 
wire u3_u0__0r0_35_0__7_; 
wire u3_u0__0r0_35_0__8_; 
wire u3_u0__0r0_35_0__9_; 
wire u3_u0__0r1_35_0__0_; 
wire u3_u0__0r1_35_0__10_; 
wire u3_u0__0r1_35_0__11_; 
wire u3_u0__0r1_35_0__12_; 
wire u3_u0__0r1_35_0__13_; 
wire u3_u0__0r1_35_0__14_; 
wire u3_u0__0r1_35_0__15_; 
wire u3_u0__0r1_35_0__16_; 
wire u3_u0__0r1_35_0__17_; 
wire u3_u0__0r1_35_0__18_; 
wire u3_u0__0r1_35_0__19_; 
wire u3_u0__0r1_35_0__1_; 
wire u3_u0__0r1_35_0__20_; 
wire u3_u0__0r1_35_0__21_; 
wire u3_u0__0r1_35_0__22_; 
wire u3_u0__0r1_35_0__23_; 
wire u3_u0__0r1_35_0__24_; 
wire u3_u0__0r1_35_0__25_; 
wire u3_u0__0r1_35_0__26_; 
wire u3_u0__0r1_35_0__27_; 
wire u3_u0__0r1_35_0__28_; 
wire u3_u0__0r1_35_0__29_; 
wire u3_u0__0r1_35_0__2_; 
wire u3_u0__0r1_35_0__30_; 
wire u3_u0__0r1_35_0__31_; 
wire u3_u0__0r1_35_0__32_; 
wire u3_u0__0r1_35_0__33_; 
wire u3_u0__0r1_35_0__34_; 
wire u3_u0__0r1_35_0__35_; 
wire u3_u0__0r1_35_0__3_; 
wire u3_u0__0r1_35_0__4_; 
wire u3_u0__0r1_35_0__5_; 
wire u3_u0__0r1_35_0__6_; 
wire u3_u0__0r1_35_0__7_; 
wire u3_u0__0r1_35_0__8_; 
wire u3_u0__0r1_35_0__9_; 
wire u3_u0__0r2_35_0__0_; 
wire u3_u0__0r2_35_0__10_; 
wire u3_u0__0r2_35_0__11_; 
wire u3_u0__0r2_35_0__12_; 
wire u3_u0__0r2_35_0__13_; 
wire u3_u0__0r2_35_0__14_; 
wire u3_u0__0r2_35_0__15_; 
wire u3_u0__0r2_35_0__16_; 
wire u3_u0__0r2_35_0__17_; 
wire u3_u0__0r2_35_0__18_; 
wire u3_u0__0r2_35_0__19_; 
wire u3_u0__0r2_35_0__1_; 
wire u3_u0__0r2_35_0__20_; 
wire u3_u0__0r2_35_0__21_; 
wire u3_u0__0r2_35_0__22_; 
wire u3_u0__0r2_35_0__23_; 
wire u3_u0__0r2_35_0__24_; 
wire u3_u0__0r2_35_0__25_; 
wire u3_u0__0r2_35_0__26_; 
wire u3_u0__0r2_35_0__27_; 
wire u3_u0__0r2_35_0__28_; 
wire u3_u0__0r2_35_0__29_; 
wire u3_u0__0r2_35_0__2_; 
wire u3_u0__0r2_35_0__30_; 
wire u3_u0__0r2_35_0__31_; 
wire u3_u0__0r2_35_0__32_; 
wire u3_u0__0r2_35_0__33_; 
wire u3_u0__0r2_35_0__34_; 
wire u3_u0__0r2_35_0__35_; 
wire u3_u0__0r2_35_0__3_; 
wire u3_u0__0r2_35_0__4_; 
wire u3_u0__0r2_35_0__5_; 
wire u3_u0__0r2_35_0__6_; 
wire u3_u0__0r2_35_0__7_; 
wire u3_u0__0r2_35_0__8_; 
wire u3_u0__0r2_35_0__9_; 
wire u3_u0__0r3_35_0__0_; 
wire u3_u0__0r3_35_0__10_; 
wire u3_u0__0r3_35_0__11_; 
wire u3_u0__0r3_35_0__12_; 
wire u3_u0__0r3_35_0__13_; 
wire u3_u0__0r3_35_0__14_; 
wire u3_u0__0r3_35_0__15_; 
wire u3_u0__0r3_35_0__16_; 
wire u3_u0__0r3_35_0__17_; 
wire u3_u0__0r3_35_0__18_; 
wire u3_u0__0r3_35_0__19_; 
wire u3_u0__0r3_35_0__1_; 
wire u3_u0__0r3_35_0__20_; 
wire u3_u0__0r3_35_0__21_; 
wire u3_u0__0r3_35_0__22_; 
wire u3_u0__0r3_35_0__23_; 
wire u3_u0__0r3_35_0__24_; 
wire u3_u0__0r3_35_0__25_; 
wire u3_u0__0r3_35_0__26_; 
wire u3_u0__0r3_35_0__27_; 
wire u3_u0__0r3_35_0__28_; 
wire u3_u0__0r3_35_0__29_; 
wire u3_u0__0r3_35_0__2_; 
wire u3_u0__0r3_35_0__30_; 
wire u3_u0__0r3_35_0__31_; 
wire u3_u0__0r3_35_0__32_; 
wire u3_u0__0r3_35_0__33_; 
wire u3_u0__0r3_35_0__34_; 
wire u3_u0__0r3_35_0__35_; 
wire u3_u0__0r3_35_0__3_; 
wire u3_u0__0r3_35_0__4_; 
wire u3_u0__0r3_35_0__5_; 
wire u3_u0__0r3_35_0__6_; 
wire u3_u0__0r3_35_0__7_; 
wire u3_u0__0r3_35_0__8_; 
wire u3_u0__0r3_35_0__9_; 
wire u3_u0__0rd_adr_3_0__0_; 
wire u3_u0__0rd_adr_3_0__1_; 
wire u3_u0__0rd_adr_3_0__2_; 
wire u3_u0__0rd_adr_3_0__3_; 
wire u3_u0__0wr_adr_3_0__0_; 
wire u3_u0__0wr_adr_3_0__1_; 
wire u3_u0__0wr_adr_3_0__2_; 
wire u3_u0__0wr_adr_3_0__3_; 
wire u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546; 
wire u3_u0__abc_74260_new_n382_; 
wire u3_u0__abc_74260_new_n383_; 
wire u3_u0__abc_74260_new_n384_; 
wire u3_u0__abc_74260_new_n386_; 
wire u3_u0__abc_74260_new_n387_; 
wire u3_u0__abc_74260_new_n389_; 
wire u3_u0__abc_74260_new_n390_; 
wire u3_u0__abc_74260_new_n392_; 
wire u3_u0__abc_74260_new_n393_; 
wire u3_u0__abc_74260_new_n395_; 
wire u3_u0__abc_74260_new_n396_; 
wire u3_u0__abc_74260_new_n398_; 
wire u3_u0__abc_74260_new_n399_; 
wire u3_u0__abc_74260_new_n401_; 
wire u3_u0__abc_74260_new_n402_; 
wire u3_u0__abc_74260_new_n404_; 
wire u3_u0__abc_74260_new_n405_; 
wire u3_u0__abc_74260_new_n407_; 
wire u3_u0__abc_74260_new_n408_; 
wire u3_u0__abc_74260_new_n410_; 
wire u3_u0__abc_74260_new_n411_; 
wire u3_u0__abc_74260_new_n413_; 
wire u3_u0__abc_74260_new_n414_; 
wire u3_u0__abc_74260_new_n416_; 
wire u3_u0__abc_74260_new_n417_; 
wire u3_u0__abc_74260_new_n419_; 
wire u3_u0__abc_74260_new_n420_; 
wire u3_u0__abc_74260_new_n422_; 
wire u3_u0__abc_74260_new_n423_; 
wire u3_u0__abc_74260_new_n425_; 
wire u3_u0__abc_74260_new_n426_; 
wire u3_u0__abc_74260_new_n428_; 
wire u3_u0__abc_74260_new_n429_; 
wire u3_u0__abc_74260_new_n431_; 
wire u3_u0__abc_74260_new_n432_; 
wire u3_u0__abc_74260_new_n434_; 
wire u3_u0__abc_74260_new_n435_; 
wire u3_u0__abc_74260_new_n437_; 
wire u3_u0__abc_74260_new_n438_; 
wire u3_u0__abc_74260_new_n440_; 
wire u3_u0__abc_74260_new_n441_; 
wire u3_u0__abc_74260_new_n443_; 
wire u3_u0__abc_74260_new_n444_; 
wire u3_u0__abc_74260_new_n446_; 
wire u3_u0__abc_74260_new_n447_; 
wire u3_u0__abc_74260_new_n449_; 
wire u3_u0__abc_74260_new_n450_; 
wire u3_u0__abc_74260_new_n452_; 
wire u3_u0__abc_74260_new_n453_; 
wire u3_u0__abc_74260_new_n455_; 
wire u3_u0__abc_74260_new_n456_; 
wire u3_u0__abc_74260_new_n458_; 
wire u3_u0__abc_74260_new_n459_; 
wire u3_u0__abc_74260_new_n461_; 
wire u3_u0__abc_74260_new_n462_; 
wire u3_u0__abc_74260_new_n464_; 
wire u3_u0__abc_74260_new_n465_; 
wire u3_u0__abc_74260_new_n467_; 
wire u3_u0__abc_74260_new_n468_; 
wire u3_u0__abc_74260_new_n470_; 
wire u3_u0__abc_74260_new_n471_; 
wire u3_u0__abc_74260_new_n473_; 
wire u3_u0__abc_74260_new_n474_; 
wire u3_u0__abc_74260_new_n476_; 
wire u3_u0__abc_74260_new_n477_; 
wire u3_u0__abc_74260_new_n479_; 
wire u3_u0__abc_74260_new_n480_; 
wire u3_u0__abc_74260_new_n482_; 
wire u3_u0__abc_74260_new_n483_; 
wire u3_u0__abc_74260_new_n485_; 
wire u3_u0__abc_74260_new_n486_; 
wire u3_u0__abc_74260_new_n488_; 
wire u3_u0__abc_74260_new_n489_; 
wire u3_u0__abc_74260_new_n491_; 
wire u3_u0__abc_74260_new_n492_; 
wire u3_u0__abc_74260_new_n494_; 
wire u3_u0__abc_74260_new_n496_; 
wire u3_u0__abc_74260_new_n498_; 
wire u3_u0__abc_74260_new_n500_; 
wire u3_u0__abc_74260_new_n502_; 
wire u3_u0__abc_74260_new_n504_; 
wire u3_u0__abc_74260_new_n506_; 
wire u3_u0__abc_74260_new_n508_; 
wire u3_u0__abc_74260_new_n510_; 
wire u3_u0__abc_74260_new_n512_; 
wire u3_u0__abc_74260_new_n514_; 
wire u3_u0__abc_74260_new_n516_; 
wire u3_u0__abc_74260_new_n518_; 
wire u3_u0__abc_74260_new_n520_; 
wire u3_u0__abc_74260_new_n522_; 
wire u3_u0__abc_74260_new_n524_; 
wire u3_u0__abc_74260_new_n526_; 
wire u3_u0__abc_74260_new_n528_; 
wire u3_u0__abc_74260_new_n530_; 
wire u3_u0__abc_74260_new_n532_; 
wire u3_u0__abc_74260_new_n534_; 
wire u3_u0__abc_74260_new_n536_; 
wire u3_u0__abc_74260_new_n538_; 
wire u3_u0__abc_74260_new_n540_; 
wire u3_u0__abc_74260_new_n542_; 
wire u3_u0__abc_74260_new_n544_; 
wire u3_u0__abc_74260_new_n546_; 
wire u3_u0__abc_74260_new_n548_; 
wire u3_u0__abc_74260_new_n550_; 
wire u3_u0__abc_74260_new_n552_; 
wire u3_u0__abc_74260_new_n554_; 
wire u3_u0__abc_74260_new_n556_; 
wire u3_u0__abc_74260_new_n558_; 
wire u3_u0__abc_74260_new_n560_; 
wire u3_u0__abc_74260_new_n562_; 
wire u3_u0__abc_74260_new_n564_; 
wire u3_u0__abc_74260_new_n565_; 
wire u3_u0__abc_74260_new_n567_; 
wire u3_u0__abc_74260_new_n569_; 
wire u3_u0__abc_74260_new_n571_; 
wire u3_u0__abc_74260_new_n573_; 
wire u3_u0__abc_74260_new_n575_; 
wire u3_u0__abc_74260_new_n577_; 
wire u3_u0__abc_74260_new_n579_; 
wire u3_u0__abc_74260_new_n581_; 
wire u3_u0__abc_74260_new_n583_; 
wire u3_u0__abc_74260_new_n585_; 
wire u3_u0__abc_74260_new_n587_; 
wire u3_u0__abc_74260_new_n589_; 
wire u3_u0__abc_74260_new_n591_; 
wire u3_u0__abc_74260_new_n593_; 
wire u3_u0__abc_74260_new_n595_; 
wire u3_u0__abc_74260_new_n597_; 
wire u3_u0__abc_74260_new_n599_; 
wire u3_u0__abc_74260_new_n601_; 
wire u3_u0__abc_74260_new_n603_; 
wire u3_u0__abc_74260_new_n605_; 
wire u3_u0__abc_74260_new_n607_; 
wire u3_u0__abc_74260_new_n609_; 
wire u3_u0__abc_74260_new_n611_; 
wire u3_u0__abc_74260_new_n613_; 
wire u3_u0__abc_74260_new_n615_; 
wire u3_u0__abc_74260_new_n617_; 
wire u3_u0__abc_74260_new_n619_; 
wire u3_u0__abc_74260_new_n621_; 
wire u3_u0__abc_74260_new_n623_; 
wire u3_u0__abc_74260_new_n625_; 
wire u3_u0__abc_74260_new_n627_; 
wire u3_u0__abc_74260_new_n629_; 
wire u3_u0__abc_74260_new_n631_; 
wire u3_u0__abc_74260_new_n633_; 
wire u3_u0__abc_74260_new_n635_; 
wire u3_u0__abc_74260_new_n637_; 
wire u3_u0__abc_74260_new_n638_; 
wire u3_u0__abc_74260_new_n640_; 
wire u3_u0__abc_74260_new_n641_; 
wire u3_u0__abc_74260_new_n642_; 
wire u3_u0__abc_74260_new_n643_; 
wire u3_u0__abc_74260_new_n645_; 
wire u3_u0__abc_74260_new_n646_; 
wire u3_u0__abc_74260_new_n648_; 
wire u3_u0__abc_74260_new_n649_; 
wire u3_u0__abc_74260_new_n651_; 
wire u3_u0__abc_74260_new_n652_; 
wire u3_u0__abc_74260_new_n654_; 
wire u3_u0__abc_74260_new_n655_; 
wire u3_u0__abc_74260_new_n656_; 
wire u3_u0__abc_74260_new_n658_; 
wire u3_u0__abc_74260_new_n660_; 
wire u3_u0__abc_74260_new_n662_; 
wire u3_u0__abc_74260_new_n664_; 
wire u3_u0__abc_74260_new_n666_; 
wire u3_u0__abc_74260_new_n668_; 
wire u3_u0__abc_74260_new_n670_; 
wire u3_u0__abc_74260_new_n672_; 
wire u3_u0__abc_74260_new_n674_; 
wire u3_u0__abc_74260_new_n676_; 
wire u3_u0__abc_74260_new_n678_; 
wire u3_u0__abc_74260_new_n680_; 
wire u3_u0__abc_74260_new_n682_; 
wire u3_u0__abc_74260_new_n684_; 
wire u3_u0__abc_74260_new_n686_; 
wire u3_u0__abc_74260_new_n688_; 
wire u3_u0__abc_74260_new_n690_; 
wire u3_u0__abc_74260_new_n692_; 
wire u3_u0__abc_74260_new_n694_; 
wire u3_u0__abc_74260_new_n696_; 
wire u3_u0__abc_74260_new_n698_; 
wire u3_u0__abc_74260_new_n700_; 
wire u3_u0__abc_74260_new_n702_; 
wire u3_u0__abc_74260_new_n704_; 
wire u3_u0__abc_74260_new_n706_; 
wire u3_u0__abc_74260_new_n708_; 
wire u3_u0__abc_74260_new_n710_; 
wire u3_u0__abc_74260_new_n712_; 
wire u3_u0__abc_74260_new_n714_; 
wire u3_u0__abc_74260_new_n716_; 
wire u3_u0__abc_74260_new_n718_; 
wire u3_u0__abc_74260_new_n720_; 
wire u3_u0__abc_74260_new_n722_; 
wire u3_u0__abc_74260_new_n724_; 
wire u3_u0__abc_74260_new_n726_; 
wire u3_u0__abc_74260_new_n728_; 
wire u3_u0__abc_74260_new_n730_; 
wire u3_u0__abc_74260_new_n732_; 
wire u3_u0__abc_74260_new_n734_; 
wire u3_u0__abc_74260_new_n735_; 
wire u3_u0__abc_74260_new_n736_; 
wire u3_u0__abc_74260_new_n737_; 
wire u3_u0__abc_74260_new_n738_; 
wire u3_u0__abc_74260_new_n739_; 
wire u3_u0__abc_74260_new_n740_; 
wire u3_u0__abc_74260_new_n741_; 
wire u3_u0__abc_74260_new_n742_; 
wire u3_u0__abc_74260_new_n743_; 
wire u3_u0__abc_74260_new_n744_; 
wire u3_u0__abc_74260_new_n745_; 
wire u3_u0__abc_74260_new_n746_; 
wire u3_u0__abc_74260_new_n747_; 
wire u3_u0__abc_74260_new_n748_; 
wire u3_u0__abc_74260_new_n750_; 
wire u3_u0__abc_74260_new_n751_; 
wire u3_u0__abc_74260_new_n752_; 
wire u3_u0__abc_74260_new_n754_; 
wire u3_u0__abc_74260_new_n755_; 
wire u3_u0__abc_74260_new_n756_; 
wire u3_u0__abc_74260_new_n758_; 
wire u3_u0__abc_74260_new_n759_; 
wire u3_u0__abc_74260_new_n760_; 
wire u3_u0__abc_74260_new_n762_; 
wire u3_u0__abc_74260_new_n763_; 
wire u3_u0__abc_74260_new_n764_; 
wire u3_u0__abc_74260_new_n766_; 
wire u3_u0__abc_74260_new_n767_; 
wire u3_u0__abc_74260_new_n768_; 
wire u3_u0__abc_74260_new_n770_; 
wire u3_u0__abc_74260_new_n771_; 
wire u3_u0__abc_74260_new_n772_; 
wire u3_u0__abc_74260_new_n774_; 
wire u3_u0__abc_74260_new_n775_; 
wire u3_u0__abc_74260_new_n776_; 
wire u3_u0__abc_74260_new_n778_; 
wire u3_u0__abc_74260_new_n779_; 
wire u3_u0__abc_74260_new_n780_; 
wire u3_u0__abc_74260_new_n782_; 
wire u3_u0__abc_74260_new_n783_; 
wire u3_u0__abc_74260_new_n784_; 
wire u3_u0__abc_74260_new_n786_; 
wire u3_u0__abc_74260_new_n787_; 
wire u3_u0__abc_74260_new_n788_; 
wire u3_u0__abc_74260_new_n790_; 
wire u3_u0__abc_74260_new_n791_; 
wire u3_u0__abc_74260_new_n792_; 
wire u3_u0__abc_74260_new_n794_; 
wire u3_u0__abc_74260_new_n795_; 
wire u3_u0__abc_74260_new_n796_; 
wire u3_u0__abc_74260_new_n798_; 
wire u3_u0__abc_74260_new_n799_; 
wire u3_u0__abc_74260_new_n800_; 
wire u3_u0__abc_74260_new_n802_; 
wire u3_u0__abc_74260_new_n803_; 
wire u3_u0__abc_74260_new_n804_; 
wire u3_u0__abc_74260_new_n806_; 
wire u3_u0__abc_74260_new_n807_; 
wire u3_u0__abc_74260_new_n808_; 
wire u3_u0__abc_74260_new_n810_; 
wire u3_u0__abc_74260_new_n811_; 
wire u3_u0__abc_74260_new_n812_; 
wire u3_u0__abc_74260_new_n814_; 
wire u3_u0__abc_74260_new_n815_; 
wire u3_u0__abc_74260_new_n816_; 
wire u3_u0__abc_74260_new_n818_; 
wire u3_u0__abc_74260_new_n819_; 
wire u3_u0__abc_74260_new_n820_; 
wire u3_u0__abc_74260_new_n822_; 
wire u3_u0__abc_74260_new_n823_; 
wire u3_u0__abc_74260_new_n824_; 
wire u3_u0__abc_74260_new_n826_; 
wire u3_u0__abc_74260_new_n827_; 
wire u3_u0__abc_74260_new_n828_; 
wire u3_u0__abc_74260_new_n830_; 
wire u3_u0__abc_74260_new_n831_; 
wire u3_u0__abc_74260_new_n832_; 
wire u3_u0__abc_74260_new_n834_; 
wire u3_u0__abc_74260_new_n835_; 
wire u3_u0__abc_74260_new_n836_; 
wire u3_u0__abc_74260_new_n838_; 
wire u3_u0__abc_74260_new_n839_; 
wire u3_u0__abc_74260_new_n840_; 
wire u3_u0__abc_74260_new_n842_; 
wire u3_u0__abc_74260_new_n843_; 
wire u3_u0__abc_74260_new_n844_; 
wire u3_u0__abc_74260_new_n846_; 
wire u3_u0__abc_74260_new_n847_; 
wire u3_u0__abc_74260_new_n848_; 
wire u3_u0__abc_74260_new_n850_; 
wire u3_u0__abc_74260_new_n851_; 
wire u3_u0__abc_74260_new_n852_; 
wire u3_u0__abc_74260_new_n854_; 
wire u3_u0__abc_74260_new_n855_; 
wire u3_u0__abc_74260_new_n856_; 
wire u3_u0__abc_74260_new_n858_; 
wire u3_u0__abc_74260_new_n859_; 
wire u3_u0__abc_74260_new_n860_; 
wire u3_u0__abc_74260_new_n862_; 
wire u3_u0__abc_74260_new_n863_; 
wire u3_u0__abc_74260_new_n864_; 
wire u3_u0__abc_74260_new_n866_; 
wire u3_u0__abc_74260_new_n867_; 
wire u3_u0__abc_74260_new_n868_; 
wire u3_u0__abc_74260_new_n870_; 
wire u3_u0__abc_74260_new_n871_; 
wire u3_u0__abc_74260_new_n872_; 
wire u3_u0__abc_74260_new_n874_; 
wire u3_u0__abc_74260_new_n875_; 
wire u3_u0__abc_74260_new_n876_; 
wire u3_u0__abc_74260_new_n878_; 
wire u3_u0__abc_74260_new_n879_; 
wire u3_u0__abc_74260_new_n880_; 
wire u3_u0__abc_74260_new_n882_; 
wire u3_u0__abc_74260_new_n883_; 
wire u3_u0__abc_74260_new_n884_; 
wire u3_u0__abc_74260_new_n886_; 
wire u3_u0__abc_74260_new_n887_; 
wire u3_u0__abc_74260_new_n888_; 
wire u3_u0_r0_0_; 
wire u3_u0_r0_10_; 
wire u3_u0_r0_11_; 
wire u3_u0_r0_12_; 
wire u3_u0_r0_13_; 
wire u3_u0_r0_14_; 
wire u3_u0_r0_15_; 
wire u3_u0_r0_16_; 
wire u3_u0_r0_17_; 
wire u3_u0_r0_18_; 
wire u3_u0_r0_19_; 
wire u3_u0_r0_1_; 
wire u3_u0_r0_20_; 
wire u3_u0_r0_21_; 
wire u3_u0_r0_22_; 
wire u3_u0_r0_23_; 
wire u3_u0_r0_24_; 
wire u3_u0_r0_25_; 
wire u3_u0_r0_26_; 
wire u3_u0_r0_27_; 
wire u3_u0_r0_28_; 
wire u3_u0_r0_29_; 
wire u3_u0_r0_2_; 
wire u3_u0_r0_30_; 
wire u3_u0_r0_31_; 
wire u3_u0_r0_32_; 
wire u3_u0_r0_33_; 
wire u3_u0_r0_34_; 
wire u3_u0_r0_35_; 
wire u3_u0_r0_3_; 
wire u3_u0_r0_4_; 
wire u3_u0_r0_5_; 
wire u3_u0_r0_6_; 
wire u3_u0_r0_7_; 
wire u3_u0_r0_8_; 
wire u3_u0_r0_9_; 
wire u3_u0_r1_0_; 
wire u3_u0_r1_10_; 
wire u3_u0_r1_11_; 
wire u3_u0_r1_12_; 
wire u3_u0_r1_13_; 
wire u3_u0_r1_14_; 
wire u3_u0_r1_15_; 
wire u3_u0_r1_16_; 
wire u3_u0_r1_17_; 
wire u3_u0_r1_18_; 
wire u3_u0_r1_19_; 
wire u3_u0_r1_1_; 
wire u3_u0_r1_20_; 
wire u3_u0_r1_21_; 
wire u3_u0_r1_22_; 
wire u3_u0_r1_23_; 
wire u3_u0_r1_24_; 
wire u3_u0_r1_25_; 
wire u3_u0_r1_26_; 
wire u3_u0_r1_27_; 
wire u3_u0_r1_28_; 
wire u3_u0_r1_29_; 
wire u3_u0_r1_2_; 
wire u3_u0_r1_30_; 
wire u3_u0_r1_31_; 
wire u3_u0_r1_32_; 
wire u3_u0_r1_33_; 
wire u3_u0_r1_34_; 
wire u3_u0_r1_35_; 
wire u3_u0_r1_3_; 
wire u3_u0_r1_4_; 
wire u3_u0_r1_5_; 
wire u3_u0_r1_6_; 
wire u3_u0_r1_7_; 
wire u3_u0_r1_8_; 
wire u3_u0_r1_9_; 
wire u3_u0_r2_0_; 
wire u3_u0_r2_10_; 
wire u3_u0_r2_11_; 
wire u3_u0_r2_12_; 
wire u3_u0_r2_13_; 
wire u3_u0_r2_14_; 
wire u3_u0_r2_15_; 
wire u3_u0_r2_16_; 
wire u3_u0_r2_17_; 
wire u3_u0_r2_18_; 
wire u3_u0_r2_19_; 
wire u3_u0_r2_1_; 
wire u3_u0_r2_20_; 
wire u3_u0_r2_21_; 
wire u3_u0_r2_22_; 
wire u3_u0_r2_23_; 
wire u3_u0_r2_24_; 
wire u3_u0_r2_25_; 
wire u3_u0_r2_26_; 
wire u3_u0_r2_27_; 
wire u3_u0_r2_28_; 
wire u3_u0_r2_29_; 
wire u3_u0_r2_2_; 
wire u3_u0_r2_30_; 
wire u3_u0_r2_31_; 
wire u3_u0_r2_32_; 
wire u3_u0_r2_33_; 
wire u3_u0_r2_34_; 
wire u3_u0_r2_35_; 
wire u3_u0_r2_3_; 
wire u3_u0_r2_4_; 
wire u3_u0_r2_5_; 
wire u3_u0_r2_6_; 
wire u3_u0_r2_7_; 
wire u3_u0_r2_8_; 
wire u3_u0_r2_9_; 
wire u3_u0_r3_0_; 
wire u3_u0_r3_10_; 
wire u3_u0_r3_11_; 
wire u3_u0_r3_12_; 
wire u3_u0_r3_13_; 
wire u3_u0_r3_14_; 
wire u3_u0_r3_15_; 
wire u3_u0_r3_16_; 
wire u3_u0_r3_17_; 
wire u3_u0_r3_18_; 
wire u3_u0_r3_19_; 
wire u3_u0_r3_1_; 
wire u3_u0_r3_20_; 
wire u3_u0_r3_21_; 
wire u3_u0_r3_22_; 
wire u3_u0_r3_23_; 
wire u3_u0_r3_24_; 
wire u3_u0_r3_25_; 
wire u3_u0_r3_26_; 
wire u3_u0_r3_27_; 
wire u3_u0_r3_28_; 
wire u3_u0_r3_29_; 
wire u3_u0_r3_2_; 
wire u3_u0_r3_30_; 
wire u3_u0_r3_31_; 
wire u3_u0_r3_32_; 
wire u3_u0_r3_33_; 
wire u3_u0_r3_34_; 
wire u3_u0_r3_35_; 
wire u3_u0_r3_3_; 
wire u3_u0_r3_4_; 
wire u3_u0_r3_5_; 
wire u3_u0_r3_6_; 
wire u3_u0_r3_7_; 
wire u3_u0_r3_8_; 
wire u3_u0_r3_9_; 
wire u3_u0_rd_adr_0_; 
wire u3_u0_rd_adr_1_; 
wire u3_u0_rd_adr_2_; 
wire u3_u0_rd_adr_3_; 
wire u3_u0_wr_adr_0_; 
wire u3_u0_wr_adr_1_; 
wire u3_u0_wr_adr_2_; 
wire u3_u0_wr_adr_3_; 
wire u3_wb_read_go; 
wire u4__0ps_cnt_7_0__0_; 
wire u4__0ps_cnt_7_0__1_; 
wire u4__0ps_cnt_7_0__2_; 
wire u4__0ps_cnt_7_0__3_; 
wire u4__0ps_cnt_7_0__4_; 
wire u4__0ps_cnt_7_0__5_; 
wire u4__0ps_cnt_7_0__6_; 
wire u4__0ps_cnt_7_0__7_; 
wire u4__0rfr_clr_0_0_; 
wire u4__0rfr_cnt_7_0__0_; 
wire u4__0rfr_cnt_7_0__1_; 
wire u4__0rfr_cnt_7_0__2_; 
wire u4__0rfr_cnt_7_0__3_; 
wire u4__0rfr_cnt_7_0__4_; 
wire u4__0rfr_cnt_7_0__5_; 
wire u4__0rfr_cnt_7_0__6_; 
wire u4__0rfr_cnt_7_0__7_; 
wire u4__0rfr_early_0_0_; 
wire u4__0rfr_en_0_0_; 
wire u4__0rfr_req_0_0_; 
wire u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562; 
wire u4__abc_74770_new_n101_; 
wire u4__abc_74770_new_n102_; 
wire u4__abc_74770_new_n103_; 
wire u4__abc_74770_new_n104_; 
wire u4__abc_74770_new_n106_; 
wire u4__abc_74770_new_n107_; 
wire u4__abc_74770_new_n108_; 
wire u4__abc_74770_new_n110_; 
wire u4__abc_74770_new_n111_; 
wire u4__abc_74770_new_n112_; 
wire u4__abc_74770_new_n113_; 
wire u4__abc_74770_new_n115_; 
wire u4__abc_74770_new_n117_; 
wire u4__abc_74770_new_n118_; 
wire u4__abc_74770_new_n119_; 
wire u4__abc_74770_new_n121_; 
wire u4__abc_74770_new_n122_; 
wire u4__abc_74770_new_n123_; 
wire u4__abc_74770_new_n124_; 
wire u4__abc_74770_new_n125_; 
wire u4__abc_74770_new_n127_; 
wire u4__abc_74770_new_n128_; 
wire u4__abc_74770_new_n129_; 
wire u4__abc_74770_new_n130_; 
wire u4__abc_74770_new_n131_; 
wire u4__abc_74770_new_n132_; 
wire u4__abc_74770_new_n134_; 
wire u4__abc_74770_new_n135_; 
wire u4__abc_74770_new_n136_; 
wire u4__abc_74770_new_n137_; 
wire u4__abc_74770_new_n139_; 
wire u4__abc_74770_new_n140_; 
wire u4__abc_74770_new_n141_; 
wire u4__abc_74770_new_n142_; 
wire u4__abc_74770_new_n144_; 
wire u4__abc_74770_new_n145_; 
wire u4__abc_74770_new_n147_; 
wire u4__abc_74770_new_n148_; 
wire u4__abc_74770_new_n149_; 
wire u4__abc_74770_new_n151_; 
wire u4__abc_74770_new_n152_; 
wire u4__abc_74770_new_n154_; 
wire u4__abc_74770_new_n155_; 
wire u4__abc_74770_new_n156_; 
wire u4__abc_74770_new_n157_; 
wire u4__abc_74770_new_n158_; 
wire u4__abc_74770_new_n159_; 
wire u4__abc_74770_new_n160_; 
wire u4__abc_74770_new_n162_; 
wire u4__abc_74770_new_n163_; 
wire u4__abc_74770_new_n165_; 
wire u4__abc_74770_new_n166_; 
wire u4__abc_74770_new_n167_; 
wire u4__abc_74770_new_n168_; 
wire u4__abc_74770_new_n169_; 
wire u4__abc_74770_new_n170_; 
wire u4__abc_74770_new_n172_; 
wire u4__abc_74770_new_n173_; 
wire u4__abc_74770_new_n174_; 
wire u4__abc_74770_new_n175_; 
wire u4__abc_74770_new_n176_; 
wire u4__abc_74770_new_n177_; 
wire u4__abc_74770_new_n178_; 
wire u4__abc_74770_new_n179_; 
wire u4__abc_74770_new_n180_; 
wire u4__abc_74770_new_n181_; 
wire u4__abc_74770_new_n182_; 
wire u4__abc_74770_new_n183_; 
wire u4__abc_74770_new_n184_; 
wire u4__abc_74770_new_n185_; 
wire u4__abc_74770_new_n65_; 
wire u4__abc_74770_new_n66_; 
wire u4__abc_74770_new_n67_; 
wire u4__abc_74770_new_n68_; 
wire u4__abc_74770_new_n69_; 
wire u4__abc_74770_new_n71_; 
wire u4__abc_74770_new_n72_; 
wire u4__abc_74770_new_n73_; 
wire u4__abc_74770_new_n74_; 
wire u4__abc_74770_new_n75_; 
wire u4__abc_74770_new_n76_; 
wire u4__abc_74770_new_n77_; 
wire u4__abc_74770_new_n78_; 
wire u4__abc_74770_new_n79_; 
wire u4__abc_74770_new_n80_; 
wire u4__abc_74770_new_n81_; 
wire u4__abc_74770_new_n82_; 
wire u4__abc_74770_new_n83_; 
wire u4__abc_74770_new_n84_; 
wire u4__abc_74770_new_n85_; 
wire u4__abc_74770_new_n86_; 
wire u4__abc_74770_new_n87_; 
wire u4__abc_74770_new_n88_; 
wire u4__abc_74770_new_n89_; 
wire u4__abc_74770_new_n91_; 
wire u4__abc_74770_new_n93_; 
wire u4__abc_74770_new_n94_; 
wire u4__abc_74770_new_n95_; 
wire u4__abc_74770_new_n97_; 
wire u4__abc_74770_new_n98_; 
wire u4__abc_74770_new_n99_; 
wire u4_ps_cnt_0_; 
wire u4_ps_cnt_1_; 
wire u4_ps_cnt_2_; 
wire u4_ps_cnt_3_; 
wire u4_ps_cnt_4_; 
wire u4_ps_cnt_5_; 
wire u4_ps_cnt_6_; 
wire u4_ps_cnt_7_; 
wire u4_ps_cnt_clr; 
wire u4_rfr_ce; 
wire u4_rfr_clr; 
wire u4_rfr_cnt_0_; 
wire u4_rfr_cnt_1_; 
wire u4_rfr_cnt_2_; 
wire u4_rfr_cnt_3_; 
wire u4_rfr_cnt_4_; 
wire u4_rfr_cnt_5_; 
wire u4_rfr_cnt_6_; 
wire u4_rfr_cnt_7_; 
wire u4_rfr_early; 
wire u4_rfr_en; 
wire u5__0ack_cnt_3_0__0_; 
wire u5__0ack_cnt_3_0__1_; 
wire u5__0ack_cnt_3_0__2_; 
wire u5__0ack_cnt_3_0__3_; 
wire u5__0ap_en_0_0_; 
wire u5__0burst_act_rd_0_0_; 
wire u5__0burst_cnt_10_0__0_; 
wire u5__0burst_cnt_10_0__10_; 
wire u5__0burst_cnt_10_0__1_; 
wire u5__0burst_cnt_10_0__2_; 
wire u5__0burst_cnt_10_0__3_; 
wire u5__0burst_cnt_10_0__4_; 
wire u5__0burst_cnt_10_0__5_; 
wire u5__0burst_cnt_10_0__6_; 
wire u5__0burst_cnt_10_0__7_; 
wire u5__0burst_cnt_10_0__8_; 
wire u5__0burst_cnt_10_0__9_; 
wire u5__0cke__0_0_; 
wire u5__0cmd_asserted2_0_0_; 
wire u5__0cmd_asserted_0_0_; 
wire u5__0data_oe_0_0_; 
wire u5__0ir_cnt_3_0__0_; 
wire u5__0ir_cnt_3_0__1_; 
wire u5__0ir_cnt_3_0__2_; 
wire u5__0ir_cnt_3_0__3_; 
wire u5__0ir_cnt_done_0_0_; 
wire u5__0lookup_ready1_0_0_; 
wire u5__0lookup_ready2_0_0_; 
wire u5__0mc_adv_r1_0_0_; 
wire u5__0mc_adv_r_0_0_; 
wire u5__0mc_le_0_0_; 
wire u5__0no_wb_cycle_0_0_; 
wire u5__0oe__0_0_; 
wire u5__0susp_sel_r_0_0_; 
wire u5__0timer2_8_0__0_; 
wire u5__0timer2_8_0__1_; 
wire u5__0timer2_8_0__2_; 
wire u5__0timer2_8_0__3_; 
wire u5__0timer2_8_0__4_; 
wire u5__0timer2_8_0__5_; 
wire u5__0timer2_8_0__6_; 
wire u5__0timer2_8_0__7_; 
wire u5__0timer2_8_0__8_; 
wire u5__0timer_7_0__0_; 
wire u5__0timer_7_0__1_; 
wire u5__0timer_7_0__2_; 
wire u5__0timer_7_0__3_; 
wire u5__0timer_7_0__4_; 
wire u5__0timer_7_0__5_; 
wire u5__0timer_7_0__6_; 
wire u5__0timer_7_0__7_; 
wire u5__0tmr2_done_0_0_; 
wire u5__0wb_cycle_0_0_; 
wire u5__0wb_stb_first_0_0_; 
wire u5__0wr_cycle_0_0_; 
wire u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962; 
wire u5__abc_78290_auto_rtlil_cc_1942_NotGate_72182; 
wire u5__abc_78290_new_n1000_; 
wire u5__abc_78290_new_n1001_; 
wire u5__abc_78290_new_n1002_; 
wire u5__abc_78290_new_n1003_; 
wire u5__abc_78290_new_n1004_; 
wire u5__abc_78290_new_n1005_; 
wire u5__abc_78290_new_n1006_; 
wire u5__abc_78290_new_n1007_; 
wire u5__abc_78290_new_n1008_; 
wire u5__abc_78290_new_n1009_; 
wire u5__abc_78290_new_n1010_; 
wire u5__abc_78290_new_n1011_; 
wire u5__abc_78290_new_n1012_; 
wire u5__abc_78290_new_n1013_; 
wire u5__abc_78290_new_n1014_; 
wire u5__abc_78290_new_n1015_; 
wire u5__abc_78290_new_n1016_; 
wire u5__abc_78290_new_n1017_; 
wire u5__abc_78290_new_n1018_; 
wire u5__abc_78290_new_n1019_; 
wire u5__abc_78290_new_n1020_; 
wire u5__abc_78290_new_n1021_; 
wire u5__abc_78290_new_n1022_; 
wire u5__abc_78290_new_n1023_; 
wire u5__abc_78290_new_n1024_; 
wire u5__abc_78290_new_n1025_; 
wire u5__abc_78290_new_n1026_; 
wire u5__abc_78290_new_n1027_; 
wire u5__abc_78290_new_n1028_; 
wire u5__abc_78290_new_n1029_; 
wire u5__abc_78290_new_n1030_; 
wire u5__abc_78290_new_n1031_; 
wire u5__abc_78290_new_n1032_; 
wire u5__abc_78290_new_n1033_; 
wire u5__abc_78290_new_n1034_; 
wire u5__abc_78290_new_n1035_; 
wire u5__abc_78290_new_n1036_; 
wire u5__abc_78290_new_n1038_; 
wire u5__abc_78290_new_n1039_; 
wire u5__abc_78290_new_n1040_; 
wire u5__abc_78290_new_n1041_; 
wire u5__abc_78290_new_n1042_; 
wire u5__abc_78290_new_n1043_; 
wire u5__abc_78290_new_n1044_; 
wire u5__abc_78290_new_n1045_; 
wire u5__abc_78290_new_n1046_; 
wire u5__abc_78290_new_n1047_; 
wire u5__abc_78290_new_n1048_; 
wire u5__abc_78290_new_n1049_; 
wire u5__abc_78290_new_n1050_; 
wire u5__abc_78290_new_n1051_; 
wire u5__abc_78290_new_n1052_; 
wire u5__abc_78290_new_n1053_; 
wire u5__abc_78290_new_n1054_; 
wire u5__abc_78290_new_n1055_; 
wire u5__abc_78290_new_n1056_; 
wire u5__abc_78290_new_n1057_; 
wire u5__abc_78290_new_n1058_; 
wire u5__abc_78290_new_n1059_; 
wire u5__abc_78290_new_n1060_; 
wire u5__abc_78290_new_n1061_; 
wire u5__abc_78290_new_n1062_; 
wire u5__abc_78290_new_n1063_; 
wire u5__abc_78290_new_n1064_; 
wire u5__abc_78290_new_n1065_; 
wire u5__abc_78290_new_n1066_; 
wire u5__abc_78290_new_n1067_; 
wire u5__abc_78290_new_n1068_; 
wire u5__abc_78290_new_n1069_; 
wire u5__abc_78290_new_n1070_; 
wire u5__abc_78290_new_n1071_; 
wire u5__abc_78290_new_n1072_; 
wire u5__abc_78290_new_n1073_; 
wire u5__abc_78290_new_n1074_; 
wire u5__abc_78290_new_n1075_; 
wire u5__abc_78290_new_n1076_; 
wire u5__abc_78290_new_n1077_; 
wire u5__abc_78290_new_n1078_; 
wire u5__abc_78290_new_n1079_; 
wire u5__abc_78290_new_n1080_; 
wire u5__abc_78290_new_n1081_; 
wire u5__abc_78290_new_n1082_; 
wire u5__abc_78290_new_n1083_; 
wire u5__abc_78290_new_n1084_; 
wire u5__abc_78290_new_n1085_; 
wire u5__abc_78290_new_n1086_; 
wire u5__abc_78290_new_n1087_; 
wire u5__abc_78290_new_n1088_; 
wire u5__abc_78290_new_n1089_; 
wire u5__abc_78290_new_n1090_; 
wire u5__abc_78290_new_n1091_; 
wire u5__abc_78290_new_n1092_; 
wire u5__abc_78290_new_n1093_; 
wire u5__abc_78290_new_n1094_; 
wire u5__abc_78290_new_n1095_; 
wire u5__abc_78290_new_n1096_; 
wire u5__abc_78290_new_n1097_; 
wire u5__abc_78290_new_n1098_; 
wire u5__abc_78290_new_n1099_; 
wire u5__abc_78290_new_n1100_; 
wire u5__abc_78290_new_n1101_; 
wire u5__abc_78290_new_n1102_; 
wire u5__abc_78290_new_n1103_; 
wire u5__abc_78290_new_n1104_; 
wire u5__abc_78290_new_n1105_; 
wire u5__abc_78290_new_n1106_; 
wire u5__abc_78290_new_n1107_; 
wire u5__abc_78290_new_n1108_; 
wire u5__abc_78290_new_n1109_; 
wire u5__abc_78290_new_n1110_; 
wire u5__abc_78290_new_n1111_; 
wire u5__abc_78290_new_n1112_; 
wire u5__abc_78290_new_n1113_; 
wire u5__abc_78290_new_n1114_; 
wire u5__abc_78290_new_n1115_; 
wire u5__abc_78290_new_n1116_; 
wire u5__abc_78290_new_n1117_; 
wire u5__abc_78290_new_n1118_; 
wire u5__abc_78290_new_n1119_; 
wire u5__abc_78290_new_n1120_; 
wire u5__abc_78290_new_n1121_; 
wire u5__abc_78290_new_n1122_; 
wire u5__abc_78290_new_n1123_; 
wire u5__abc_78290_new_n1124_; 
wire u5__abc_78290_new_n1125_; 
wire u5__abc_78290_new_n1126_; 
wire u5__abc_78290_new_n1127_; 
wire u5__abc_78290_new_n1128_; 
wire u5__abc_78290_new_n1129_; 
wire u5__abc_78290_new_n1130_; 
wire u5__abc_78290_new_n1131_; 
wire u5__abc_78290_new_n1132_; 
wire u5__abc_78290_new_n1133_; 
wire u5__abc_78290_new_n1134_; 
wire u5__abc_78290_new_n1135_; 
wire u5__abc_78290_new_n1136_; 
wire u5__abc_78290_new_n1137_; 
wire u5__abc_78290_new_n1138_; 
wire u5__abc_78290_new_n1139_; 
wire u5__abc_78290_new_n1140_; 
wire u5__abc_78290_new_n1141_; 
wire u5__abc_78290_new_n1142_; 
wire u5__abc_78290_new_n1143_; 
wire u5__abc_78290_new_n1144_; 
wire u5__abc_78290_new_n1145_; 
wire u5__abc_78290_new_n1146_; 
wire u5__abc_78290_new_n1147_; 
wire u5__abc_78290_new_n1148_; 
wire u5__abc_78290_new_n1149_; 
wire u5__abc_78290_new_n1150_; 
wire u5__abc_78290_new_n1151_; 
wire u5__abc_78290_new_n1152_; 
wire u5__abc_78290_new_n1153_; 
wire u5__abc_78290_new_n1154_; 
wire u5__abc_78290_new_n1155_; 
wire u5__abc_78290_new_n1156_; 
wire u5__abc_78290_new_n1157_; 
wire u5__abc_78290_new_n1158_; 
wire u5__abc_78290_new_n1159_; 
wire u5__abc_78290_new_n1160_; 
wire u5__abc_78290_new_n1161_; 
wire u5__abc_78290_new_n1162_; 
wire u5__abc_78290_new_n1163_; 
wire u5__abc_78290_new_n1164_; 
wire u5__abc_78290_new_n1165_; 
wire u5__abc_78290_new_n1166_; 
wire u5__abc_78290_new_n1167_; 
wire u5__abc_78290_new_n1168_; 
wire u5__abc_78290_new_n1169_; 
wire u5__abc_78290_new_n1170_; 
wire u5__abc_78290_new_n1171_; 
wire u5__abc_78290_new_n1172_; 
wire u5__abc_78290_new_n1173_; 
wire u5__abc_78290_new_n1174_; 
wire u5__abc_78290_new_n1175_; 
wire u5__abc_78290_new_n1176_; 
wire u5__abc_78290_new_n1177_; 
wire u5__abc_78290_new_n1178_; 
wire u5__abc_78290_new_n1179_; 
wire u5__abc_78290_new_n1180_; 
wire u5__abc_78290_new_n1181_; 
wire u5__abc_78290_new_n1182_; 
wire u5__abc_78290_new_n1183_; 
wire u5__abc_78290_new_n1184_; 
wire u5__abc_78290_new_n1185_; 
wire u5__abc_78290_new_n1186_; 
wire u5__abc_78290_new_n1187_; 
wire u5__abc_78290_new_n1188_; 
wire u5__abc_78290_new_n1189_; 
wire u5__abc_78290_new_n1190_; 
wire u5__abc_78290_new_n1191_; 
wire u5__abc_78290_new_n1192_; 
wire u5__abc_78290_new_n1193_; 
wire u5__abc_78290_new_n1194_; 
wire u5__abc_78290_new_n1195_; 
wire u5__abc_78290_new_n1196_; 
wire u5__abc_78290_new_n1197_; 
wire u5__abc_78290_new_n1198_; 
wire u5__abc_78290_new_n1199_; 
wire u5__abc_78290_new_n1200_; 
wire u5__abc_78290_new_n1201_; 
wire u5__abc_78290_new_n1202_; 
wire u5__abc_78290_new_n1203_; 
wire u5__abc_78290_new_n1204_; 
wire u5__abc_78290_new_n1205_; 
wire u5__abc_78290_new_n1206_; 
wire u5__abc_78290_new_n1207_; 
wire u5__abc_78290_new_n1208_; 
wire u5__abc_78290_new_n1209_; 
wire u5__abc_78290_new_n1210_; 
wire u5__abc_78290_new_n1211_; 
wire u5__abc_78290_new_n1212_; 
wire u5__abc_78290_new_n1213_; 
wire u5__abc_78290_new_n1214_; 
wire u5__abc_78290_new_n1215_; 
wire u5__abc_78290_new_n1216_; 
wire u5__abc_78290_new_n1217_; 
wire u5__abc_78290_new_n1218_; 
wire u5__abc_78290_new_n1219_; 
wire u5__abc_78290_new_n1220_; 
wire u5__abc_78290_new_n1221_; 
wire u5__abc_78290_new_n1222_; 
wire u5__abc_78290_new_n1223_; 
wire u5__abc_78290_new_n1224_; 
wire u5__abc_78290_new_n1225_; 
wire u5__abc_78290_new_n1226_; 
wire u5__abc_78290_new_n1227_; 
wire u5__abc_78290_new_n1228_; 
wire u5__abc_78290_new_n1229_; 
wire u5__abc_78290_new_n1230_; 
wire u5__abc_78290_new_n1231_; 
wire u5__abc_78290_new_n1232_; 
wire u5__abc_78290_new_n1233_; 
wire u5__abc_78290_new_n1234_; 
wire u5__abc_78290_new_n1235_; 
wire u5__abc_78290_new_n1236_; 
wire u5__abc_78290_new_n1237_; 
wire u5__abc_78290_new_n1238_; 
wire u5__abc_78290_new_n1239_; 
wire u5__abc_78290_new_n1240_; 
wire u5__abc_78290_new_n1241_; 
wire u5__abc_78290_new_n1242_; 
wire u5__abc_78290_new_n1243_; 
wire u5__abc_78290_new_n1244_; 
wire u5__abc_78290_new_n1245_; 
wire u5__abc_78290_new_n1246_; 
wire u5__abc_78290_new_n1247_; 
wire u5__abc_78290_new_n1248_; 
wire u5__abc_78290_new_n1249_; 
wire u5__abc_78290_new_n1250_; 
wire u5__abc_78290_new_n1251_; 
wire u5__abc_78290_new_n1252_; 
wire u5__abc_78290_new_n1253_; 
wire u5__abc_78290_new_n1254_; 
wire u5__abc_78290_new_n1255_; 
wire u5__abc_78290_new_n1256_; 
wire u5__abc_78290_new_n1257_; 
wire u5__abc_78290_new_n1258_; 
wire u5__abc_78290_new_n1259_; 
wire u5__abc_78290_new_n1260_; 
wire u5__abc_78290_new_n1261_; 
wire u5__abc_78290_new_n1262_; 
wire u5__abc_78290_new_n1263_; 
wire u5__abc_78290_new_n1264_; 
wire u5__abc_78290_new_n1265_; 
wire u5__abc_78290_new_n1266_; 
wire u5__abc_78290_new_n1267_; 
wire u5__abc_78290_new_n1268_; 
wire u5__abc_78290_new_n1269_; 
wire u5__abc_78290_new_n1270_; 
wire u5__abc_78290_new_n1271_; 
wire u5__abc_78290_new_n1272_; 
wire u5__abc_78290_new_n1273_; 
wire u5__abc_78290_new_n1274_; 
wire u5__abc_78290_new_n1275_; 
wire u5__abc_78290_new_n1276_; 
wire u5__abc_78290_new_n1277_; 
wire u5__abc_78290_new_n1278_; 
wire u5__abc_78290_new_n1279_; 
wire u5__abc_78290_new_n1280_; 
wire u5__abc_78290_new_n1281_; 
wire u5__abc_78290_new_n1282_; 
wire u5__abc_78290_new_n1283_; 
wire u5__abc_78290_new_n1284_; 
wire u5__abc_78290_new_n1285_; 
wire u5__abc_78290_new_n1286_; 
wire u5__abc_78290_new_n1287_; 
wire u5__abc_78290_new_n1288_; 
wire u5__abc_78290_new_n1289_; 
wire u5__abc_78290_new_n1290_; 
wire u5__abc_78290_new_n1291_; 
wire u5__abc_78290_new_n1292_; 
wire u5__abc_78290_new_n1293_; 
wire u5__abc_78290_new_n1294_; 
wire u5__abc_78290_new_n1295_; 
wire u5__abc_78290_new_n1296_; 
wire u5__abc_78290_new_n1297_; 
wire u5__abc_78290_new_n1298_; 
wire u5__abc_78290_new_n1299_; 
wire u5__abc_78290_new_n1300_; 
wire u5__abc_78290_new_n1301_; 
wire u5__abc_78290_new_n1302_; 
wire u5__abc_78290_new_n1303_; 
wire u5__abc_78290_new_n1304_; 
wire u5__abc_78290_new_n1305_; 
wire u5__abc_78290_new_n1306_; 
wire u5__abc_78290_new_n1307_; 
wire u5__abc_78290_new_n1308_; 
wire u5__abc_78290_new_n1309_; 
wire u5__abc_78290_new_n1310_; 
wire u5__abc_78290_new_n1311_; 
wire u5__abc_78290_new_n1312_; 
wire u5__abc_78290_new_n1313_; 
wire u5__abc_78290_new_n1314_; 
wire u5__abc_78290_new_n1315_; 
wire u5__abc_78290_new_n1316_; 
wire u5__abc_78290_new_n1317_; 
wire u5__abc_78290_new_n1318_; 
wire u5__abc_78290_new_n1319_; 
wire u5__abc_78290_new_n1320_; 
wire u5__abc_78290_new_n1321_; 
wire u5__abc_78290_new_n1322_; 
wire u5__abc_78290_new_n1323_; 
wire u5__abc_78290_new_n1324_; 
wire u5__abc_78290_new_n1325_; 
wire u5__abc_78290_new_n1326_; 
wire u5__abc_78290_new_n1327_; 
wire u5__abc_78290_new_n1328_; 
wire u5__abc_78290_new_n1329_; 
wire u5__abc_78290_new_n1330_; 
wire u5__abc_78290_new_n1331_; 
wire u5__abc_78290_new_n1332_; 
wire u5__abc_78290_new_n1333_; 
wire u5__abc_78290_new_n1334_; 
wire u5__abc_78290_new_n1335_; 
wire u5__abc_78290_new_n1336_; 
wire u5__abc_78290_new_n1337_; 
wire u5__abc_78290_new_n1338_; 
wire u5__abc_78290_new_n1339_; 
wire u5__abc_78290_new_n1340_; 
wire u5__abc_78290_new_n1341_; 
wire u5__abc_78290_new_n1342_; 
wire u5__abc_78290_new_n1343_; 
wire u5__abc_78290_new_n1344_; 
wire u5__abc_78290_new_n1345_; 
wire u5__abc_78290_new_n1346_; 
wire u5__abc_78290_new_n1347_; 
wire u5__abc_78290_new_n1348_; 
wire u5__abc_78290_new_n1349_; 
wire u5__abc_78290_new_n1350_; 
wire u5__abc_78290_new_n1351_; 
wire u5__abc_78290_new_n1352_; 
wire u5__abc_78290_new_n1353_; 
wire u5__abc_78290_new_n1354_; 
wire u5__abc_78290_new_n1355_; 
wire u5__abc_78290_new_n1356_; 
wire u5__abc_78290_new_n1357_; 
wire u5__abc_78290_new_n1358_; 
wire u5__abc_78290_new_n1359_; 
wire u5__abc_78290_new_n1360_; 
wire u5__abc_78290_new_n1361_; 
wire u5__abc_78290_new_n1362_; 
wire u5__abc_78290_new_n1363_; 
wire u5__abc_78290_new_n1364_; 
wire u5__abc_78290_new_n1365_; 
wire u5__abc_78290_new_n1366_; 
wire u5__abc_78290_new_n1367_; 
wire u5__abc_78290_new_n1368_; 
wire u5__abc_78290_new_n1369_; 
wire u5__abc_78290_new_n1370_; 
wire u5__abc_78290_new_n1371_; 
wire u5__abc_78290_new_n1372_; 
wire u5__abc_78290_new_n1373_; 
wire u5__abc_78290_new_n1374_; 
wire u5__abc_78290_new_n1375_; 
wire u5__abc_78290_new_n1376_; 
wire u5__abc_78290_new_n1377_; 
wire u5__abc_78290_new_n1378_; 
wire u5__abc_78290_new_n1379_; 
wire u5__abc_78290_new_n1380_; 
wire u5__abc_78290_new_n1381_; 
wire u5__abc_78290_new_n1382_; 
wire u5__abc_78290_new_n1383_; 
wire u5__abc_78290_new_n1384_; 
wire u5__abc_78290_new_n1385_; 
wire u5__abc_78290_new_n1386_; 
wire u5__abc_78290_new_n1387_; 
wire u5__abc_78290_new_n1388_; 
wire u5__abc_78290_new_n1389_; 
wire u5__abc_78290_new_n1390_; 
wire u5__abc_78290_new_n1391_; 
wire u5__abc_78290_new_n1392_; 
wire u5__abc_78290_new_n1393_; 
wire u5__abc_78290_new_n1394_; 
wire u5__abc_78290_new_n1395_; 
wire u5__abc_78290_new_n1396_; 
wire u5__abc_78290_new_n1397_; 
wire u5__abc_78290_new_n1398_; 
wire u5__abc_78290_new_n1399_; 
wire u5__abc_78290_new_n1400_; 
wire u5__abc_78290_new_n1401_; 
wire u5__abc_78290_new_n1402_; 
wire u5__abc_78290_new_n1403_; 
wire u5__abc_78290_new_n1404_; 
wire u5__abc_78290_new_n1405_; 
wire u5__abc_78290_new_n1406_; 
wire u5__abc_78290_new_n1407_; 
wire u5__abc_78290_new_n1408_; 
wire u5__abc_78290_new_n1409_; 
wire u5__abc_78290_new_n1410_; 
wire u5__abc_78290_new_n1411_; 
wire u5__abc_78290_new_n1412_; 
wire u5__abc_78290_new_n1413_; 
wire u5__abc_78290_new_n1414_; 
wire u5__abc_78290_new_n1415_; 
wire u5__abc_78290_new_n1416_; 
wire u5__abc_78290_new_n1417_; 
wire u5__abc_78290_new_n1418_; 
wire u5__abc_78290_new_n1419_; 
wire u5__abc_78290_new_n1420_; 
wire u5__abc_78290_new_n1421_; 
wire u5__abc_78290_new_n1422_; 
wire u5__abc_78290_new_n1423_; 
wire u5__abc_78290_new_n1424_; 
wire u5__abc_78290_new_n1425_; 
wire u5__abc_78290_new_n1426_; 
wire u5__abc_78290_new_n1428_; 
wire u5__abc_78290_new_n1429_; 
wire u5__abc_78290_new_n1430_; 
wire u5__abc_78290_new_n1432_; 
wire u5__abc_78290_new_n1433_; 
wire u5__abc_78290_new_n1434_; 
wire u5__abc_78290_new_n1435_; 
wire u5__abc_78290_new_n1436_; 
wire u5__abc_78290_new_n1437_; 
wire u5__abc_78290_new_n1438_; 
wire u5__abc_78290_new_n1439_; 
wire u5__abc_78290_new_n1440_; 
wire u5__abc_78290_new_n1441_; 
wire u5__abc_78290_new_n1442_; 
wire u5__abc_78290_new_n1443_; 
wire u5__abc_78290_new_n1444_; 
wire u5__abc_78290_new_n1445_; 
wire u5__abc_78290_new_n1446_; 
wire u5__abc_78290_new_n1447_; 
wire u5__abc_78290_new_n1448_; 
wire u5__abc_78290_new_n1449_; 
wire u5__abc_78290_new_n1451_; 
wire u5__abc_78290_new_n1452_; 
wire u5__abc_78290_new_n1454_; 
wire u5__abc_78290_new_n1455_; 
wire u5__abc_78290_new_n1456_; 
wire u5__abc_78290_new_n1457_; 
wire u5__abc_78290_new_n1458_; 
wire u5__abc_78290_new_n1459_; 
wire u5__abc_78290_new_n1460_; 
wire u5__abc_78290_new_n1461_; 
wire u5__abc_78290_new_n1462_; 
wire u5__abc_78290_new_n1463_; 
wire u5__abc_78290_new_n1465_; 
wire u5__abc_78290_new_n1466_; 
wire u5__abc_78290_new_n1468_; 
wire u5__abc_78290_new_n1469_; 
wire u5__abc_78290_new_n1470_; 
wire u5__abc_78290_new_n1471_; 
wire u5__abc_78290_new_n1472_; 
wire u5__abc_78290_new_n1473_; 
wire u5__abc_78290_new_n1474_; 
wire u5__abc_78290_new_n1475_; 
wire u5__abc_78290_new_n1476_; 
wire u5__abc_78290_new_n1477_; 
wire u5__abc_78290_new_n1478_; 
wire u5__abc_78290_new_n1479_; 
wire u5__abc_78290_new_n1480_; 
wire u5__abc_78290_new_n1481_; 
wire u5__abc_78290_new_n1482_; 
wire u5__abc_78290_new_n1483_; 
wire u5__abc_78290_new_n1484_; 
wire u5__abc_78290_new_n1485_; 
wire u5__abc_78290_new_n1486_; 
wire u5__abc_78290_new_n1487_; 
wire u5__abc_78290_new_n1488_; 
wire u5__abc_78290_new_n1489_; 
wire u5__abc_78290_new_n1490_; 
wire u5__abc_78290_new_n1491_; 
wire u5__abc_78290_new_n1492_; 
wire u5__abc_78290_new_n1493_; 
wire u5__abc_78290_new_n1494_; 
wire u5__abc_78290_new_n1495_; 
wire u5__abc_78290_new_n1496_; 
wire u5__abc_78290_new_n1497_; 
wire u5__abc_78290_new_n1498_; 
wire u5__abc_78290_new_n1499_; 
wire u5__abc_78290_new_n1500_; 
wire u5__abc_78290_new_n1501_; 
wire u5__abc_78290_new_n1502_; 
wire u5__abc_78290_new_n1503_; 
wire u5__abc_78290_new_n1504_; 
wire u5__abc_78290_new_n1505_; 
wire u5__abc_78290_new_n1506_; 
wire u5__abc_78290_new_n1507_; 
wire u5__abc_78290_new_n1508_; 
wire u5__abc_78290_new_n1510_; 
wire u5__abc_78290_new_n1512_; 
wire u5__abc_78290_new_n1513_; 
wire u5__abc_78290_new_n1514_; 
wire u5__abc_78290_new_n1515_; 
wire u5__abc_78290_new_n1516_; 
wire u5__abc_78290_new_n1517_; 
wire u5__abc_78290_new_n1518_; 
wire u5__abc_78290_new_n1519_; 
wire u5__abc_78290_new_n1520_; 
wire u5__abc_78290_new_n1522_; 
wire u5__abc_78290_new_n1523_; 
wire u5__abc_78290_new_n1525_; 
wire u5__abc_78290_new_n1526_; 
wire u5__abc_78290_new_n1527_; 
wire u5__abc_78290_new_n1528_; 
wire u5__abc_78290_new_n1529_; 
wire u5__abc_78290_new_n1530_; 
wire u5__abc_78290_new_n1531_; 
wire u5__abc_78290_new_n1532_; 
wire u5__abc_78290_new_n1533_; 
wire u5__abc_78290_new_n1534_; 
wire u5__abc_78290_new_n1535_; 
wire u5__abc_78290_new_n1536_; 
wire u5__abc_78290_new_n1537_; 
wire u5__abc_78290_new_n1538_; 
wire u5__abc_78290_new_n1539_; 
wire u5__abc_78290_new_n1540_; 
wire u5__abc_78290_new_n1541_; 
wire u5__abc_78290_new_n1542_; 
wire u5__abc_78290_new_n1543_; 
wire u5__abc_78290_new_n1544_; 
wire u5__abc_78290_new_n1545_; 
wire u5__abc_78290_new_n1546_; 
wire u5__abc_78290_new_n1547_; 
wire u5__abc_78290_new_n1548_; 
wire u5__abc_78290_new_n1549_; 
wire u5__abc_78290_new_n1550_; 
wire u5__abc_78290_new_n1551_; 
wire u5__abc_78290_new_n1552_; 
wire u5__abc_78290_new_n1553_; 
wire u5__abc_78290_new_n1554_; 
wire u5__abc_78290_new_n1555_; 
wire u5__abc_78290_new_n1556_; 
wire u5__abc_78290_new_n1557_; 
wire u5__abc_78290_new_n1558_; 
wire u5__abc_78290_new_n1559_; 
wire u5__abc_78290_new_n1560_; 
wire u5__abc_78290_new_n1561_; 
wire u5__abc_78290_new_n1562_; 
wire u5__abc_78290_new_n1563_; 
wire u5__abc_78290_new_n1564_; 
wire u5__abc_78290_new_n1565_; 
wire u5__abc_78290_new_n1566_; 
wire u5__abc_78290_new_n1567_; 
wire u5__abc_78290_new_n1568_; 
wire u5__abc_78290_new_n1570_; 
wire u5__abc_78290_new_n1571_; 
wire u5__abc_78290_new_n1572_; 
wire u5__abc_78290_new_n1573_; 
wire u5__abc_78290_new_n1574_; 
wire u5__abc_78290_new_n1575_; 
wire u5__abc_78290_new_n1576_; 
wire u5__abc_78290_new_n1577_; 
wire u5__abc_78290_new_n1578_; 
wire u5__abc_78290_new_n1579_; 
wire u5__abc_78290_new_n1580_; 
wire u5__abc_78290_new_n1581_; 
wire u5__abc_78290_new_n1582_; 
wire u5__abc_78290_new_n1583_; 
wire u5__abc_78290_new_n1584_; 
wire u5__abc_78290_new_n1585_; 
wire u5__abc_78290_new_n1587_; 
wire u5__abc_78290_new_n1588_; 
wire u5__abc_78290_new_n1589_; 
wire u5__abc_78290_new_n1590_; 
wire u5__abc_78290_new_n1591_; 
wire u5__abc_78290_new_n1593_; 
wire u5__abc_78290_new_n1594_; 
wire u5__abc_78290_new_n1595_; 
wire u5__abc_78290_new_n1596_; 
wire u5__abc_78290_new_n1597_; 
wire u5__abc_78290_new_n1598_; 
wire u5__abc_78290_new_n1599_; 
wire u5__abc_78290_new_n1600_; 
wire u5__abc_78290_new_n1601_; 
wire u5__abc_78290_new_n1602_; 
wire u5__abc_78290_new_n1603_; 
wire u5__abc_78290_new_n1604_; 
wire u5__abc_78290_new_n1605_; 
wire u5__abc_78290_new_n1606_; 
wire u5__abc_78290_new_n1607_; 
wire u5__abc_78290_new_n1608_; 
wire u5__abc_78290_new_n1609_; 
wire u5__abc_78290_new_n1610_; 
wire u5__abc_78290_new_n1611_; 
wire u5__abc_78290_new_n1612_; 
wire u5__abc_78290_new_n1613_; 
wire u5__abc_78290_new_n1614_; 
wire u5__abc_78290_new_n1615_; 
wire u5__abc_78290_new_n1616_; 
wire u5__abc_78290_new_n1617_; 
wire u5__abc_78290_new_n1618_; 
wire u5__abc_78290_new_n1619_; 
wire u5__abc_78290_new_n1620_; 
wire u5__abc_78290_new_n1621_; 
wire u5__abc_78290_new_n1622_; 
wire u5__abc_78290_new_n1623_; 
wire u5__abc_78290_new_n1624_; 
wire u5__abc_78290_new_n1625_; 
wire u5__abc_78290_new_n1626_; 
wire u5__abc_78290_new_n1627_; 
wire u5__abc_78290_new_n1629_; 
wire u5__abc_78290_new_n1631_; 
wire u5__abc_78290_new_n1632_; 
wire u5__abc_78290_new_n1633_; 
wire u5__abc_78290_new_n1634_; 
wire u5__abc_78290_new_n1636_; 
wire u5__abc_78290_new_n1637_; 
wire u5__abc_78290_new_n1638_; 
wire u5__abc_78290_new_n1639_; 
wire u5__abc_78290_new_n1640_; 
wire u5__abc_78290_new_n1641_; 
wire u5__abc_78290_new_n1642_; 
wire u5__abc_78290_new_n1643_; 
wire u5__abc_78290_new_n1644_; 
wire u5__abc_78290_new_n1645_; 
wire u5__abc_78290_new_n1646_; 
wire u5__abc_78290_new_n1647_; 
wire u5__abc_78290_new_n1648_; 
wire u5__abc_78290_new_n1649_; 
wire u5__abc_78290_new_n1650_; 
wire u5__abc_78290_new_n1651_; 
wire u5__abc_78290_new_n1652_; 
wire u5__abc_78290_new_n1653_; 
wire u5__abc_78290_new_n1654_; 
wire u5__abc_78290_new_n1655_; 
wire u5__abc_78290_new_n1656_; 
wire u5__abc_78290_new_n1657_; 
wire u5__abc_78290_new_n1658_; 
wire u5__abc_78290_new_n1659_; 
wire u5__abc_78290_new_n1660_; 
wire u5__abc_78290_new_n1661_; 
wire u5__abc_78290_new_n1662_; 
wire u5__abc_78290_new_n1663_; 
wire u5__abc_78290_new_n1664_; 
wire u5__abc_78290_new_n1665_; 
wire u5__abc_78290_new_n1666_; 
wire u5__abc_78290_new_n1667_; 
wire u5__abc_78290_new_n1668_; 
wire u5__abc_78290_new_n1669_; 
wire u5__abc_78290_new_n1670_; 
wire u5__abc_78290_new_n1672_; 
wire u5__abc_78290_new_n1673_; 
wire u5__abc_78290_new_n1674_; 
wire u5__abc_78290_new_n1675_; 
wire u5__abc_78290_new_n1676_; 
wire u5__abc_78290_new_n1677_; 
wire u5__abc_78290_new_n1679_; 
wire u5__abc_78290_new_n1680_; 
wire u5__abc_78290_new_n1681_; 
wire u5__abc_78290_new_n1682_; 
wire u5__abc_78290_new_n1683_; 
wire u5__abc_78290_new_n1685_; 
wire u5__abc_78290_new_n1686_; 
wire u5__abc_78290_new_n1687_; 
wire u5__abc_78290_new_n1688_; 
wire u5__abc_78290_new_n1689_; 
wire u5__abc_78290_new_n1690_; 
wire u5__abc_78290_new_n1692_; 
wire u5__abc_78290_new_n1693_; 
wire u5__abc_78290_new_n1694_; 
wire u5__abc_78290_new_n1695_; 
wire u5__abc_78290_new_n1696_; 
wire u5__abc_78290_new_n1697_; 
wire u5__abc_78290_new_n1699_; 
wire u5__abc_78290_new_n1700_; 
wire u5__abc_78290_new_n1701_; 
wire u5__abc_78290_new_n1702_; 
wire u5__abc_78290_new_n1703_; 
wire u5__abc_78290_new_n1705_; 
wire u5__abc_78290_new_n1706_; 
wire u5__abc_78290_new_n1707_; 
wire u5__abc_78290_new_n1708_; 
wire u5__abc_78290_new_n1709_; 
wire u5__abc_78290_new_n1711_; 
wire u5__abc_78290_new_n1712_; 
wire u5__abc_78290_new_n1713_; 
wire u5__abc_78290_new_n1714_; 
wire u5__abc_78290_new_n1715_; 
wire u5__abc_78290_new_n1716_; 
wire u5__abc_78290_new_n1717_; 
wire u5__abc_78290_new_n1718_; 
wire u5__abc_78290_new_n1719_; 
wire u5__abc_78290_new_n1720_; 
wire u5__abc_78290_new_n1721_; 
wire u5__abc_78290_new_n1722_; 
wire u5__abc_78290_new_n1723_; 
wire u5__abc_78290_new_n1724_; 
wire u5__abc_78290_new_n1725_; 
wire u5__abc_78290_new_n1726_; 
wire u5__abc_78290_new_n1727_; 
wire u5__abc_78290_new_n1728_; 
wire u5__abc_78290_new_n1729_; 
wire u5__abc_78290_new_n1730_; 
wire u5__abc_78290_new_n1731_; 
wire u5__abc_78290_new_n1732_; 
wire u5__abc_78290_new_n1733_; 
wire u5__abc_78290_new_n1734_; 
wire u5__abc_78290_new_n1735_; 
wire u5__abc_78290_new_n1736_; 
wire u5__abc_78290_new_n1737_; 
wire u5__abc_78290_new_n1738_; 
wire u5__abc_78290_new_n1739_; 
wire u5__abc_78290_new_n1740_; 
wire u5__abc_78290_new_n1741_; 
wire u5__abc_78290_new_n1742_; 
wire u5__abc_78290_new_n1743_; 
wire u5__abc_78290_new_n1744_; 
wire u5__abc_78290_new_n1745_; 
wire u5__abc_78290_new_n1746_; 
wire u5__abc_78290_new_n1747_; 
wire u5__abc_78290_new_n1748_; 
wire u5__abc_78290_new_n1749_; 
wire u5__abc_78290_new_n1750_; 
wire u5__abc_78290_new_n1751_; 
wire u5__abc_78290_new_n1752_; 
wire u5__abc_78290_new_n1753_; 
wire u5__abc_78290_new_n1754_; 
wire u5__abc_78290_new_n1755_; 
wire u5__abc_78290_new_n1756_; 
wire u5__abc_78290_new_n1757_; 
wire u5__abc_78290_new_n1758_; 
wire u5__abc_78290_new_n1759_; 
wire u5__abc_78290_new_n1760_; 
wire u5__abc_78290_new_n1761_; 
wire u5__abc_78290_new_n1762_; 
wire u5__abc_78290_new_n1763_; 
wire u5__abc_78290_new_n1764_; 
wire u5__abc_78290_new_n1765_; 
wire u5__abc_78290_new_n1766_; 
wire u5__abc_78290_new_n1767_; 
wire u5__abc_78290_new_n1768_; 
wire u5__abc_78290_new_n1769_; 
wire u5__abc_78290_new_n1770_; 
wire u5__abc_78290_new_n1771_; 
wire u5__abc_78290_new_n1772_; 
wire u5__abc_78290_new_n1773_; 
wire u5__abc_78290_new_n1774_; 
wire u5__abc_78290_new_n1775_; 
wire u5__abc_78290_new_n1776_; 
wire u5__abc_78290_new_n1777_; 
wire u5__abc_78290_new_n1778_; 
wire u5__abc_78290_new_n1779_; 
wire u5__abc_78290_new_n1780_; 
wire u5__abc_78290_new_n1781_; 
wire u5__abc_78290_new_n1782_; 
wire u5__abc_78290_new_n1783_; 
wire u5__abc_78290_new_n1784_; 
wire u5__abc_78290_new_n1785_; 
wire u5__abc_78290_new_n1786_; 
wire u5__abc_78290_new_n1787_; 
wire u5__abc_78290_new_n1788_; 
wire u5__abc_78290_new_n1789_; 
wire u5__abc_78290_new_n1790_; 
wire u5__abc_78290_new_n1791_; 
wire u5__abc_78290_new_n1792_; 
wire u5__abc_78290_new_n1793_; 
wire u5__abc_78290_new_n1794_; 
wire u5__abc_78290_new_n1795_; 
wire u5__abc_78290_new_n1796_; 
wire u5__abc_78290_new_n1797_; 
wire u5__abc_78290_new_n1798_; 
wire u5__abc_78290_new_n1799_; 
wire u5__abc_78290_new_n1800_; 
wire u5__abc_78290_new_n1801_; 
wire u5__abc_78290_new_n1802_; 
wire u5__abc_78290_new_n1803_; 
wire u5__abc_78290_new_n1804_; 
wire u5__abc_78290_new_n1805_; 
wire u5__abc_78290_new_n1806_; 
wire u5__abc_78290_new_n1807_; 
wire u5__abc_78290_new_n1808_; 
wire u5__abc_78290_new_n1809_; 
wire u5__abc_78290_new_n1810_; 
wire u5__abc_78290_new_n1811_; 
wire u5__abc_78290_new_n1812_; 
wire u5__abc_78290_new_n1813_; 
wire u5__abc_78290_new_n1814_; 
wire u5__abc_78290_new_n1815_; 
wire u5__abc_78290_new_n1816_; 
wire u5__abc_78290_new_n1817_; 
wire u5__abc_78290_new_n1818_; 
wire u5__abc_78290_new_n1819_; 
wire u5__abc_78290_new_n1820_; 
wire u5__abc_78290_new_n1821_; 
wire u5__abc_78290_new_n1822_; 
wire u5__abc_78290_new_n1823_; 
wire u5__abc_78290_new_n1824_; 
wire u5__abc_78290_new_n1825_; 
wire u5__abc_78290_new_n1826_; 
wire u5__abc_78290_new_n1827_; 
wire u5__abc_78290_new_n1828_; 
wire u5__abc_78290_new_n1829_; 
wire u5__abc_78290_new_n1830_; 
wire u5__abc_78290_new_n1831_; 
wire u5__abc_78290_new_n1832_; 
wire u5__abc_78290_new_n1833_; 
wire u5__abc_78290_new_n1834_; 
wire u5__abc_78290_new_n1835_; 
wire u5__abc_78290_new_n1836_; 
wire u5__abc_78290_new_n1837_; 
wire u5__abc_78290_new_n1838_; 
wire u5__abc_78290_new_n1839_; 
wire u5__abc_78290_new_n1840_; 
wire u5__abc_78290_new_n1841_; 
wire u5__abc_78290_new_n1842_; 
wire u5__abc_78290_new_n1843_; 
wire u5__abc_78290_new_n1844_; 
wire u5__abc_78290_new_n1845_; 
wire u5__abc_78290_new_n1846_; 
wire u5__abc_78290_new_n1847_; 
wire u5__abc_78290_new_n1848_; 
wire u5__abc_78290_new_n1849_; 
wire u5__abc_78290_new_n1850_; 
wire u5__abc_78290_new_n1851_; 
wire u5__abc_78290_new_n1852_; 
wire u5__abc_78290_new_n1853_; 
wire u5__abc_78290_new_n1854_; 
wire u5__abc_78290_new_n1855_; 
wire u5__abc_78290_new_n1856_; 
wire u5__abc_78290_new_n1857_; 
wire u5__abc_78290_new_n1858_; 
wire u5__abc_78290_new_n1859_; 
wire u5__abc_78290_new_n1860_; 
wire u5__abc_78290_new_n1861_; 
wire u5__abc_78290_new_n1862_; 
wire u5__abc_78290_new_n1863_; 
wire u5__abc_78290_new_n1864_; 
wire u5__abc_78290_new_n1865_; 
wire u5__abc_78290_new_n1866_; 
wire u5__abc_78290_new_n1867_; 
wire u5__abc_78290_new_n1868_; 
wire u5__abc_78290_new_n1869_; 
wire u5__abc_78290_new_n1870_; 
wire u5__abc_78290_new_n1871_; 
wire u5__abc_78290_new_n1872_; 
wire u5__abc_78290_new_n1873_; 
wire u5__abc_78290_new_n1874_; 
wire u5__abc_78290_new_n1875_; 
wire u5__abc_78290_new_n1876_; 
wire u5__abc_78290_new_n1877_; 
wire u5__abc_78290_new_n1878_; 
wire u5__abc_78290_new_n1879_; 
wire u5__abc_78290_new_n1880_; 
wire u5__abc_78290_new_n1881_; 
wire u5__abc_78290_new_n1882_; 
wire u5__abc_78290_new_n1883_; 
wire u5__abc_78290_new_n1884_; 
wire u5__abc_78290_new_n1885_; 
wire u5__abc_78290_new_n1886_; 
wire u5__abc_78290_new_n1887_; 
wire u5__abc_78290_new_n1888_; 
wire u5__abc_78290_new_n1889_; 
wire u5__abc_78290_new_n1890_; 
wire u5__abc_78290_new_n1891_; 
wire u5__abc_78290_new_n1892_; 
wire u5__abc_78290_new_n1893_; 
wire u5__abc_78290_new_n1894_; 
wire u5__abc_78290_new_n1895_; 
wire u5__abc_78290_new_n1896_; 
wire u5__abc_78290_new_n1897_; 
wire u5__abc_78290_new_n1898_; 
wire u5__abc_78290_new_n1899_; 
wire u5__abc_78290_new_n1900_; 
wire u5__abc_78290_new_n1901_; 
wire u5__abc_78290_new_n1902_; 
wire u5__abc_78290_new_n1903_; 
wire u5__abc_78290_new_n1904_; 
wire u5__abc_78290_new_n1905_; 
wire u5__abc_78290_new_n1906_; 
wire u5__abc_78290_new_n1907_; 
wire u5__abc_78290_new_n1908_; 
wire u5__abc_78290_new_n1909_; 
wire u5__abc_78290_new_n1910_; 
wire u5__abc_78290_new_n1911_; 
wire u5__abc_78290_new_n1912_; 
wire u5__abc_78290_new_n1913_; 
wire u5__abc_78290_new_n1914_; 
wire u5__abc_78290_new_n1915_; 
wire u5__abc_78290_new_n1916_; 
wire u5__abc_78290_new_n1917_; 
wire u5__abc_78290_new_n1918_; 
wire u5__abc_78290_new_n1919_; 
wire u5__abc_78290_new_n1920_; 
wire u5__abc_78290_new_n1921_; 
wire u5__abc_78290_new_n1922_; 
wire u5__abc_78290_new_n1923_; 
wire u5__abc_78290_new_n1924_; 
wire u5__abc_78290_new_n1925_; 
wire u5__abc_78290_new_n1926_; 
wire u5__abc_78290_new_n1927_; 
wire u5__abc_78290_new_n1928_; 
wire u5__abc_78290_new_n1929_; 
wire u5__abc_78290_new_n1930_; 
wire u5__abc_78290_new_n1931_; 
wire u5__abc_78290_new_n1932_; 
wire u5__abc_78290_new_n1933_; 
wire u5__abc_78290_new_n1934_; 
wire u5__abc_78290_new_n1935_; 
wire u5__abc_78290_new_n1936_; 
wire u5__abc_78290_new_n1937_; 
wire u5__abc_78290_new_n1938_; 
wire u5__abc_78290_new_n1939_; 
wire u5__abc_78290_new_n1940_; 
wire u5__abc_78290_new_n1941_; 
wire u5__abc_78290_new_n1942_; 
wire u5__abc_78290_new_n1943_; 
wire u5__abc_78290_new_n1944_; 
wire u5__abc_78290_new_n1945_; 
wire u5__abc_78290_new_n1946_; 
wire u5__abc_78290_new_n1947_; 
wire u5__abc_78290_new_n1948_; 
wire u5__abc_78290_new_n1949_; 
wire u5__abc_78290_new_n1950_; 
wire u5__abc_78290_new_n1951_; 
wire u5__abc_78290_new_n1952_; 
wire u5__abc_78290_new_n1953_; 
wire u5__abc_78290_new_n1954_; 
wire u5__abc_78290_new_n1955_; 
wire u5__abc_78290_new_n1956_; 
wire u5__abc_78290_new_n1957_; 
wire u5__abc_78290_new_n1959_; 
wire u5__abc_78290_new_n1960_; 
wire u5__abc_78290_new_n1961_; 
wire u5__abc_78290_new_n1962_; 
wire u5__abc_78290_new_n1963_; 
wire u5__abc_78290_new_n1964_; 
wire u5__abc_78290_new_n1965_; 
wire u5__abc_78290_new_n1967_; 
wire u5__abc_78290_new_n1968_; 
wire u5__abc_78290_new_n1969_; 
wire u5__abc_78290_new_n1970_; 
wire u5__abc_78290_new_n1971_; 
wire u5__abc_78290_new_n1972_; 
wire u5__abc_78290_new_n1973_; 
wire u5__abc_78290_new_n1975_; 
wire u5__abc_78290_new_n1976_; 
wire u5__abc_78290_new_n1977_; 
wire u5__abc_78290_new_n1978_; 
wire u5__abc_78290_new_n1979_; 
wire u5__abc_78290_new_n1980_; 
wire u5__abc_78290_new_n1982_; 
wire u5__abc_78290_new_n1983_; 
wire u5__abc_78290_new_n1984_; 
wire u5__abc_78290_new_n1985_; 
wire u5__abc_78290_new_n1986_; 
wire u5__abc_78290_new_n1987_; 
wire u5__abc_78290_new_n1988_; 
wire u5__abc_78290_new_n1989_; 
wire u5__abc_78290_new_n1990_; 
wire u5__abc_78290_new_n1991_; 
wire u5__abc_78290_new_n1992_; 
wire u5__abc_78290_new_n1993_; 
wire u5__abc_78290_new_n1994_; 
wire u5__abc_78290_new_n1995_; 
wire u5__abc_78290_new_n1996_; 
wire u5__abc_78290_new_n1997_; 
wire u5__abc_78290_new_n1998_; 
wire u5__abc_78290_new_n1999_; 
wire u5__abc_78290_new_n2000_; 
wire u5__abc_78290_new_n2001_; 
wire u5__abc_78290_new_n2002_; 
wire u5__abc_78290_new_n2003_; 
wire u5__abc_78290_new_n2004_; 
wire u5__abc_78290_new_n2005_; 
wire u5__abc_78290_new_n2006_; 
wire u5__abc_78290_new_n2007_; 
wire u5__abc_78290_new_n2008_; 
wire u5__abc_78290_new_n2009_; 
wire u5__abc_78290_new_n2010_; 
wire u5__abc_78290_new_n2011_; 
wire u5__abc_78290_new_n2013_; 
wire u5__abc_78290_new_n2015_; 
wire u5__abc_78290_new_n2016_; 
wire u5__abc_78290_new_n2017_; 
wire u5__abc_78290_new_n2018_; 
wire u5__abc_78290_new_n2020_; 
wire u5__abc_78290_new_n2021_; 
wire u5__abc_78290_new_n2023_; 
wire u5__abc_78290_new_n2024_; 
wire u5__abc_78290_new_n2025_; 
wire u5__abc_78290_new_n2026_; 
wire u5__abc_78290_new_n2027_; 
wire u5__abc_78290_new_n2028_; 
wire u5__abc_78290_new_n2029_; 
wire u5__abc_78290_new_n2030_; 
wire u5__abc_78290_new_n2031_; 
wire u5__abc_78290_new_n2032_; 
wire u5__abc_78290_new_n2033_; 
wire u5__abc_78290_new_n2034_; 
wire u5__abc_78290_new_n2035_; 
wire u5__abc_78290_new_n2036_; 
wire u5__abc_78290_new_n2037_; 
wire u5__abc_78290_new_n2038_; 
wire u5__abc_78290_new_n2039_; 
wire u5__abc_78290_new_n2040_; 
wire u5__abc_78290_new_n2041_; 
wire u5__abc_78290_new_n2042_; 
wire u5__abc_78290_new_n2043_; 
wire u5__abc_78290_new_n2044_; 
wire u5__abc_78290_new_n2045_; 
wire u5__abc_78290_new_n2046_; 
wire u5__abc_78290_new_n2047_; 
wire u5__abc_78290_new_n2048_; 
wire u5__abc_78290_new_n2049_; 
wire u5__abc_78290_new_n2050_; 
wire u5__abc_78290_new_n2051_; 
wire u5__abc_78290_new_n2052_; 
wire u5__abc_78290_new_n2053_; 
wire u5__abc_78290_new_n2054_; 
wire u5__abc_78290_new_n2055_; 
wire u5__abc_78290_new_n2056_; 
wire u5__abc_78290_new_n2057_; 
wire u5__abc_78290_new_n2058_; 
wire u5__abc_78290_new_n2059_; 
wire u5__abc_78290_new_n2060_; 
wire u5__abc_78290_new_n2061_; 
wire u5__abc_78290_new_n2062_; 
wire u5__abc_78290_new_n2063_; 
wire u5__abc_78290_new_n2064_; 
wire u5__abc_78290_new_n2065_; 
wire u5__abc_78290_new_n2066_; 
wire u5__abc_78290_new_n2067_; 
wire u5__abc_78290_new_n2068_; 
wire u5__abc_78290_new_n2069_; 
wire u5__abc_78290_new_n2070_; 
wire u5__abc_78290_new_n2071_; 
wire u5__abc_78290_new_n2072_; 
wire u5__abc_78290_new_n2073_; 
wire u5__abc_78290_new_n2074_; 
wire u5__abc_78290_new_n2075_; 
wire u5__abc_78290_new_n2076_; 
wire u5__abc_78290_new_n2077_; 
wire u5__abc_78290_new_n2078_; 
wire u5__abc_78290_new_n2079_; 
wire u5__abc_78290_new_n2080_; 
wire u5__abc_78290_new_n2081_; 
wire u5__abc_78290_new_n2082_; 
wire u5__abc_78290_new_n2083_; 
wire u5__abc_78290_new_n2084_; 
wire u5__abc_78290_new_n2085_; 
wire u5__abc_78290_new_n2086_; 
wire u5__abc_78290_new_n2087_; 
wire u5__abc_78290_new_n2088_; 
wire u5__abc_78290_new_n2089_; 
wire u5__abc_78290_new_n2090_; 
wire u5__abc_78290_new_n2091_; 
wire u5__abc_78290_new_n2092_; 
wire u5__abc_78290_new_n2093_; 
wire u5__abc_78290_new_n2094_; 
wire u5__abc_78290_new_n2095_; 
wire u5__abc_78290_new_n2096_; 
wire u5__abc_78290_new_n2097_; 
wire u5__abc_78290_new_n2098_; 
wire u5__abc_78290_new_n2099_; 
wire u5__abc_78290_new_n2100_; 
wire u5__abc_78290_new_n2101_; 
wire u5__abc_78290_new_n2102_; 
wire u5__abc_78290_new_n2103_; 
wire u5__abc_78290_new_n2104_; 
wire u5__abc_78290_new_n2105_; 
wire u5__abc_78290_new_n2106_; 
wire u5__abc_78290_new_n2107_; 
wire u5__abc_78290_new_n2108_; 
wire u5__abc_78290_new_n2109_; 
wire u5__abc_78290_new_n2110_; 
wire u5__abc_78290_new_n2111_; 
wire u5__abc_78290_new_n2112_; 
wire u5__abc_78290_new_n2113_; 
wire u5__abc_78290_new_n2114_; 
wire u5__abc_78290_new_n2115_; 
wire u5__abc_78290_new_n2116_; 
wire u5__abc_78290_new_n2117_; 
wire u5__abc_78290_new_n2118_; 
wire u5__abc_78290_new_n2119_; 
wire u5__abc_78290_new_n2120_; 
wire u5__abc_78290_new_n2121_; 
wire u5__abc_78290_new_n2122_; 
wire u5__abc_78290_new_n2123_; 
wire u5__abc_78290_new_n2124_; 
wire u5__abc_78290_new_n2125_; 
wire u5__abc_78290_new_n2126_; 
wire u5__abc_78290_new_n2127_; 
wire u5__abc_78290_new_n2128_; 
wire u5__abc_78290_new_n2129_; 
wire u5__abc_78290_new_n2130_; 
wire u5__abc_78290_new_n2131_; 
wire u5__abc_78290_new_n2132_; 
wire u5__abc_78290_new_n2133_; 
wire u5__abc_78290_new_n2134_; 
wire u5__abc_78290_new_n2135_; 
wire u5__abc_78290_new_n2136_; 
wire u5__abc_78290_new_n2137_; 
wire u5__abc_78290_new_n2138_; 
wire u5__abc_78290_new_n2139_; 
wire u5__abc_78290_new_n2140_; 
wire u5__abc_78290_new_n2141_; 
wire u5__abc_78290_new_n2142_; 
wire u5__abc_78290_new_n2143_; 
wire u5__abc_78290_new_n2144_; 
wire u5__abc_78290_new_n2145_; 
wire u5__abc_78290_new_n2146_; 
wire u5__abc_78290_new_n2147_; 
wire u5__abc_78290_new_n2148_; 
wire u5__abc_78290_new_n2149_; 
wire u5__abc_78290_new_n2150_; 
wire u5__abc_78290_new_n2151_; 
wire u5__abc_78290_new_n2152_; 
wire u5__abc_78290_new_n2153_; 
wire u5__abc_78290_new_n2154_; 
wire u5__abc_78290_new_n2155_; 
wire u5__abc_78290_new_n2156_; 
wire u5__abc_78290_new_n2157_; 
wire u5__abc_78290_new_n2158_; 
wire u5__abc_78290_new_n2159_; 
wire u5__abc_78290_new_n2160_; 
wire u5__abc_78290_new_n2161_; 
wire u5__abc_78290_new_n2162_; 
wire u5__abc_78290_new_n2163_; 
wire u5__abc_78290_new_n2164_; 
wire u5__abc_78290_new_n2165_; 
wire u5__abc_78290_new_n2166_; 
wire u5__abc_78290_new_n2167_; 
wire u5__abc_78290_new_n2168_; 
wire u5__abc_78290_new_n2169_; 
wire u5__abc_78290_new_n2170_; 
wire u5__abc_78290_new_n2171_; 
wire u5__abc_78290_new_n2172_; 
wire u5__abc_78290_new_n2173_; 
wire u5__abc_78290_new_n2174_; 
wire u5__abc_78290_new_n2175_; 
wire u5__abc_78290_new_n2176_; 
wire u5__abc_78290_new_n2177_; 
wire u5__abc_78290_new_n2178_; 
wire u5__abc_78290_new_n2179_; 
wire u5__abc_78290_new_n2180_; 
wire u5__abc_78290_new_n2181_; 
wire u5__abc_78290_new_n2182_; 
wire u5__abc_78290_new_n2183_; 
wire u5__abc_78290_new_n2184_; 
wire u5__abc_78290_new_n2185_; 
wire u5__abc_78290_new_n2186_; 
wire u5__abc_78290_new_n2187_; 
wire u5__abc_78290_new_n2188_; 
wire u5__abc_78290_new_n2189_; 
wire u5__abc_78290_new_n2190_; 
wire u5__abc_78290_new_n2191_; 
wire u5__abc_78290_new_n2192_; 
wire u5__abc_78290_new_n2193_; 
wire u5__abc_78290_new_n2194_; 
wire u5__abc_78290_new_n2195_; 
wire u5__abc_78290_new_n2196_; 
wire u5__abc_78290_new_n2197_; 
wire u5__abc_78290_new_n2198_; 
wire u5__abc_78290_new_n2199_; 
wire u5__abc_78290_new_n2200_; 
wire u5__abc_78290_new_n2201_; 
wire u5__abc_78290_new_n2202_; 
wire u5__abc_78290_new_n2203_; 
wire u5__abc_78290_new_n2204_; 
wire u5__abc_78290_new_n2205_; 
wire u5__abc_78290_new_n2206_; 
wire u5__abc_78290_new_n2207_; 
wire u5__abc_78290_new_n2208_; 
wire u5__abc_78290_new_n2209_; 
wire u5__abc_78290_new_n2210_; 
wire u5__abc_78290_new_n2211_; 
wire u5__abc_78290_new_n2212_; 
wire u5__abc_78290_new_n2213_; 
wire u5__abc_78290_new_n2214_; 
wire u5__abc_78290_new_n2215_; 
wire u5__abc_78290_new_n2216_; 
wire u5__abc_78290_new_n2217_; 
wire u5__abc_78290_new_n2218_; 
wire u5__abc_78290_new_n2219_; 
wire u5__abc_78290_new_n2220_; 
wire u5__abc_78290_new_n2221_; 
wire u5__abc_78290_new_n2222_; 
wire u5__abc_78290_new_n2223_; 
wire u5__abc_78290_new_n2224_; 
wire u5__abc_78290_new_n2225_; 
wire u5__abc_78290_new_n2226_; 
wire u5__abc_78290_new_n2227_; 
wire u5__abc_78290_new_n2228_; 
wire u5__abc_78290_new_n2230_; 
wire u5__abc_78290_new_n2231_; 
wire u5__abc_78290_new_n2232_; 
wire u5__abc_78290_new_n2233_; 
wire u5__abc_78290_new_n2234_; 
wire u5__abc_78290_new_n2235_; 
wire u5__abc_78290_new_n2236_; 
wire u5__abc_78290_new_n2237_; 
wire u5__abc_78290_new_n2238_; 
wire u5__abc_78290_new_n2239_; 
wire u5__abc_78290_new_n2240_; 
wire u5__abc_78290_new_n2241_; 
wire u5__abc_78290_new_n2242_; 
wire u5__abc_78290_new_n2243_; 
wire u5__abc_78290_new_n2244_; 
wire u5__abc_78290_new_n2245_; 
wire u5__abc_78290_new_n2246_; 
wire u5__abc_78290_new_n2247_; 
wire u5__abc_78290_new_n2248_; 
wire u5__abc_78290_new_n2249_; 
wire u5__abc_78290_new_n2250_; 
wire u5__abc_78290_new_n2251_; 
wire u5__abc_78290_new_n2252_; 
wire u5__abc_78290_new_n2253_; 
wire u5__abc_78290_new_n2254_; 
wire u5__abc_78290_new_n2255_; 
wire u5__abc_78290_new_n2256_; 
wire u5__abc_78290_new_n2257_; 
wire u5__abc_78290_new_n2258_; 
wire u5__abc_78290_new_n2259_; 
wire u5__abc_78290_new_n2260_; 
wire u5__abc_78290_new_n2261_; 
wire u5__abc_78290_new_n2263_; 
wire u5__abc_78290_new_n2264_; 
wire u5__abc_78290_new_n2265_; 
wire u5__abc_78290_new_n2266_; 
wire u5__abc_78290_new_n2267_; 
wire u5__abc_78290_new_n2268_; 
wire u5__abc_78290_new_n2269_; 
wire u5__abc_78290_new_n2270_; 
wire u5__abc_78290_new_n2271_; 
wire u5__abc_78290_new_n2272_; 
wire u5__abc_78290_new_n2273_; 
wire u5__abc_78290_new_n2274_; 
wire u5__abc_78290_new_n2275_; 
wire u5__abc_78290_new_n2276_; 
wire u5__abc_78290_new_n2277_; 
wire u5__abc_78290_new_n2278_; 
wire u5__abc_78290_new_n2279_; 
wire u5__abc_78290_new_n2280_; 
wire u5__abc_78290_new_n2281_; 
wire u5__abc_78290_new_n2282_; 
wire u5__abc_78290_new_n2283_; 
wire u5__abc_78290_new_n2284_; 
wire u5__abc_78290_new_n2285_; 
wire u5__abc_78290_new_n2286_; 
wire u5__abc_78290_new_n2287_; 
wire u5__abc_78290_new_n2288_; 
wire u5__abc_78290_new_n2289_; 
wire u5__abc_78290_new_n2290_; 
wire u5__abc_78290_new_n2291_; 
wire u5__abc_78290_new_n2292_; 
wire u5__abc_78290_new_n2293_; 
wire u5__abc_78290_new_n2294_; 
wire u5__abc_78290_new_n2295_; 
wire u5__abc_78290_new_n2296_; 
wire u5__abc_78290_new_n2297_; 
wire u5__abc_78290_new_n2298_; 
wire u5__abc_78290_new_n2299_; 
wire u5__abc_78290_new_n2300_; 
wire u5__abc_78290_new_n2301_; 
wire u5__abc_78290_new_n2302_; 
wire u5__abc_78290_new_n2303_; 
wire u5__abc_78290_new_n2304_; 
wire u5__abc_78290_new_n2305_; 
wire u5__abc_78290_new_n2306_; 
wire u5__abc_78290_new_n2308_; 
wire u5__abc_78290_new_n2309_; 
wire u5__abc_78290_new_n2310_; 
wire u5__abc_78290_new_n2311_; 
wire u5__abc_78290_new_n2312_; 
wire u5__abc_78290_new_n2313_; 
wire u5__abc_78290_new_n2314_; 
wire u5__abc_78290_new_n2315_; 
wire u5__abc_78290_new_n2316_; 
wire u5__abc_78290_new_n2317_; 
wire u5__abc_78290_new_n2318_; 
wire u5__abc_78290_new_n2319_; 
wire u5__abc_78290_new_n2320_; 
wire u5__abc_78290_new_n2321_; 
wire u5__abc_78290_new_n2322_; 
wire u5__abc_78290_new_n2323_; 
wire u5__abc_78290_new_n2324_; 
wire u5__abc_78290_new_n2325_; 
wire u5__abc_78290_new_n2326_; 
wire u5__abc_78290_new_n2327_; 
wire u5__abc_78290_new_n2329_; 
wire u5__abc_78290_new_n2330_; 
wire u5__abc_78290_new_n2331_; 
wire u5__abc_78290_new_n2332_; 
wire u5__abc_78290_new_n2333_; 
wire u5__abc_78290_new_n2334_; 
wire u5__abc_78290_new_n2335_; 
wire u5__abc_78290_new_n2336_; 
wire u5__abc_78290_new_n2337_; 
wire u5__abc_78290_new_n2338_; 
wire u5__abc_78290_new_n2339_; 
wire u5__abc_78290_new_n2340_; 
wire u5__abc_78290_new_n2341_; 
wire u5__abc_78290_new_n2342_; 
wire u5__abc_78290_new_n2343_; 
wire u5__abc_78290_new_n2344_; 
wire u5__abc_78290_new_n2345_; 
wire u5__abc_78290_new_n2346_; 
wire u5__abc_78290_new_n2348_; 
wire u5__abc_78290_new_n2349_; 
wire u5__abc_78290_new_n2350_; 
wire u5__abc_78290_new_n2351_; 
wire u5__abc_78290_new_n2352_; 
wire u5__abc_78290_new_n2353_; 
wire u5__abc_78290_new_n2354_; 
wire u5__abc_78290_new_n2356_; 
wire u5__abc_78290_new_n2357_; 
wire u5__abc_78290_new_n2358_; 
wire u5__abc_78290_new_n2359_; 
wire u5__abc_78290_new_n2360_; 
wire u5__abc_78290_new_n2361_; 
wire u5__abc_78290_new_n2363_; 
wire u5__abc_78290_new_n2364_; 
wire u5__abc_78290_new_n2365_; 
wire u5__abc_78290_new_n2367_; 
wire u5__abc_78290_new_n2368_; 
wire u5__abc_78290_new_n2369_; 
wire u5__abc_78290_new_n2370_; 
wire u5__abc_78290_new_n2371_; 
wire u5__abc_78290_new_n2372_; 
wire u5__abc_78290_new_n2373_; 
wire u5__abc_78290_new_n2374_; 
wire u5__abc_78290_new_n2375_; 
wire u5__abc_78290_new_n2376_; 
wire u5__abc_78290_new_n2377_; 
wire u5__abc_78290_new_n2378_; 
wire u5__abc_78290_new_n2379_; 
wire u5__abc_78290_new_n2380_; 
wire u5__abc_78290_new_n2381_; 
wire u5__abc_78290_new_n2382_; 
wire u5__abc_78290_new_n2383_; 
wire u5__abc_78290_new_n2384_; 
wire u5__abc_78290_new_n2385_; 
wire u5__abc_78290_new_n2386_; 
wire u5__abc_78290_new_n2387_; 
wire u5__abc_78290_new_n2388_; 
wire u5__abc_78290_new_n2389_; 
wire u5__abc_78290_new_n2390_; 
wire u5__abc_78290_new_n2391_; 
wire u5__abc_78290_new_n2392_; 
wire u5__abc_78290_new_n2393_; 
wire u5__abc_78290_new_n2394_; 
wire u5__abc_78290_new_n2395_; 
wire u5__abc_78290_new_n2396_; 
wire u5__abc_78290_new_n2397_; 
wire u5__abc_78290_new_n2398_; 
wire u5__abc_78290_new_n2399_; 
wire u5__abc_78290_new_n2400_; 
wire u5__abc_78290_new_n2401_; 
wire u5__abc_78290_new_n2402_; 
wire u5__abc_78290_new_n2403_; 
wire u5__abc_78290_new_n2404_; 
wire u5__abc_78290_new_n2405_; 
wire u5__abc_78290_new_n2406_; 
wire u5__abc_78290_new_n2407_; 
wire u5__abc_78290_new_n2408_; 
wire u5__abc_78290_new_n2409_; 
wire u5__abc_78290_new_n2410_; 
wire u5__abc_78290_new_n2411_; 
wire u5__abc_78290_new_n2412_; 
wire u5__abc_78290_new_n2413_; 
wire u5__abc_78290_new_n2414_; 
wire u5__abc_78290_new_n2415_; 
wire u5__abc_78290_new_n2416_; 
wire u5__abc_78290_new_n2417_; 
wire u5__abc_78290_new_n2418_; 
wire u5__abc_78290_new_n2419_; 
wire u5__abc_78290_new_n2420_; 
wire u5__abc_78290_new_n2421_; 
wire u5__abc_78290_new_n2422_; 
wire u5__abc_78290_new_n2423_; 
wire u5__abc_78290_new_n2424_; 
wire u5__abc_78290_new_n2425_; 
wire u5__abc_78290_new_n2426_; 
wire u5__abc_78290_new_n2427_; 
wire u5__abc_78290_new_n2428_; 
wire u5__abc_78290_new_n2429_; 
wire u5__abc_78290_new_n2430_; 
wire u5__abc_78290_new_n2431_; 
wire u5__abc_78290_new_n2433_; 
wire u5__abc_78290_new_n2434_; 
wire u5__abc_78290_new_n2435_; 
wire u5__abc_78290_new_n2436_; 
wire u5__abc_78290_new_n2437_; 
wire u5__abc_78290_new_n2438_; 
wire u5__abc_78290_new_n2439_; 
wire u5__abc_78290_new_n2440_; 
wire u5__abc_78290_new_n2441_; 
wire u5__abc_78290_new_n2442_; 
wire u5__abc_78290_new_n2443_; 
wire u5__abc_78290_new_n2444_; 
wire u5__abc_78290_new_n2445_; 
wire u5__abc_78290_new_n2446_; 
wire u5__abc_78290_new_n2447_; 
wire u5__abc_78290_new_n2448_; 
wire u5__abc_78290_new_n2449_; 
wire u5__abc_78290_new_n2450_; 
wire u5__abc_78290_new_n2451_; 
wire u5__abc_78290_new_n2452_; 
wire u5__abc_78290_new_n2453_; 
wire u5__abc_78290_new_n2454_; 
wire u5__abc_78290_new_n2455_; 
wire u5__abc_78290_new_n2456_; 
wire u5__abc_78290_new_n2457_; 
wire u5__abc_78290_new_n2458_; 
wire u5__abc_78290_new_n2459_; 
wire u5__abc_78290_new_n2460_; 
wire u5__abc_78290_new_n2461_; 
wire u5__abc_78290_new_n2462_; 
wire u5__abc_78290_new_n2464_; 
wire u5__abc_78290_new_n2465_; 
wire u5__abc_78290_new_n2466_; 
wire u5__abc_78290_new_n2467_; 
wire u5__abc_78290_new_n2468_; 
wire u5__abc_78290_new_n2469_; 
wire u5__abc_78290_new_n2470_; 
wire u5__abc_78290_new_n2471_; 
wire u5__abc_78290_new_n2472_; 
wire u5__abc_78290_new_n2473_; 
wire u5__abc_78290_new_n2474_; 
wire u5__abc_78290_new_n2475_; 
wire u5__abc_78290_new_n2476_; 
wire u5__abc_78290_new_n2477_; 
wire u5__abc_78290_new_n2478_; 
wire u5__abc_78290_new_n2479_; 
wire u5__abc_78290_new_n2480_; 
wire u5__abc_78290_new_n2481_; 
wire u5__abc_78290_new_n2483_; 
wire u5__abc_78290_new_n2484_; 
wire u5__abc_78290_new_n2485_; 
wire u5__abc_78290_new_n2486_; 
wire u5__abc_78290_new_n2487_; 
wire u5__abc_78290_new_n2488_; 
wire u5__abc_78290_new_n2489_; 
wire u5__abc_78290_new_n2490_; 
wire u5__abc_78290_new_n2491_; 
wire u5__abc_78290_new_n2492_; 
wire u5__abc_78290_new_n2493_; 
wire u5__abc_78290_new_n2494_; 
wire u5__abc_78290_new_n2495_; 
wire u5__abc_78290_new_n2497_; 
wire u5__abc_78290_new_n2498_; 
wire u5__abc_78290_new_n2499_; 
wire u5__abc_78290_new_n2500_; 
wire u5__abc_78290_new_n2501_; 
wire u5__abc_78290_new_n2502_; 
wire u5__abc_78290_new_n2503_; 
wire u5__abc_78290_new_n2504_; 
wire u5__abc_78290_new_n2505_; 
wire u5__abc_78290_new_n2506_; 
wire u5__abc_78290_new_n2507_; 
wire u5__abc_78290_new_n2508_; 
wire u5__abc_78290_new_n2510_; 
wire u5__abc_78290_new_n2511_; 
wire u5__abc_78290_new_n2512_; 
wire u5__abc_78290_new_n2513_; 
wire u5__abc_78290_new_n2514_; 
wire u5__abc_78290_new_n2515_; 
wire u5__abc_78290_new_n2516_; 
wire u5__abc_78290_new_n2517_; 
wire u5__abc_78290_new_n2518_; 
wire u5__abc_78290_new_n2520_; 
wire u5__abc_78290_new_n2521_; 
wire u5__abc_78290_new_n2522_; 
wire u5__abc_78290_new_n2523_; 
wire u5__abc_78290_new_n2524_; 
wire u5__abc_78290_new_n2526_; 
wire u5__abc_78290_new_n2527_; 
wire u5__abc_78290_new_n2528_; 
wire u5__abc_78290_new_n2529_; 
wire u5__abc_78290_new_n2531_; 
wire u5__abc_78290_new_n2532_; 
wire u5__abc_78290_new_n2534_; 
wire u5__abc_78290_new_n2535_; 
wire u5__abc_78290_new_n2536_; 
wire u5__abc_78290_new_n2537_; 
wire u5__abc_78290_new_n2538_; 
wire u5__abc_78290_new_n2539_; 
wire u5__abc_78290_new_n2541_; 
wire u5__abc_78290_new_n2542_; 
wire u5__abc_78290_new_n2543_; 
wire u5__abc_78290_new_n2544_; 
wire u5__abc_78290_new_n2545_; 
wire u5__abc_78290_new_n2546_; 
wire u5__abc_78290_new_n2548_; 
wire u5__abc_78290_new_n2549_; 
wire u5__abc_78290_new_n2550_; 
wire u5__abc_78290_new_n2551_; 
wire u5__abc_78290_new_n2553_; 
wire u5__abc_78290_new_n2554_; 
wire u5__abc_78290_new_n2555_; 
wire u5__abc_78290_new_n2556_; 
wire u5__abc_78290_new_n2558_; 
wire u5__abc_78290_new_n2560_; 
wire u5__abc_78290_new_n2562_; 
wire u5__abc_78290_new_n2563_; 
wire u5__abc_78290_new_n2565_; 
wire u5__abc_78290_new_n2566_; 
wire u5__abc_78290_new_n2567_; 
wire u5__abc_78290_new_n2568_; 
wire u5__abc_78290_new_n2569_; 
wire u5__abc_78290_new_n2570_; 
wire u5__abc_78290_new_n2571_; 
wire u5__abc_78290_new_n2572_; 
wire u5__abc_78290_new_n2574_; 
wire u5__abc_78290_new_n2576_; 
wire u5__abc_78290_new_n2577_; 
wire u5__abc_78290_new_n2578_; 
wire u5__abc_78290_new_n2579_; 
wire u5__abc_78290_new_n2580_; 
wire u5__abc_78290_new_n2581_; 
wire u5__abc_78290_new_n2582_; 
wire u5__abc_78290_new_n2583_; 
wire u5__abc_78290_new_n2584_; 
wire u5__abc_78290_new_n2586_; 
wire u5__abc_78290_new_n2587_; 
wire u5__abc_78290_new_n2588_; 
wire u5__abc_78290_new_n2589_; 
wire u5__abc_78290_new_n2590_; 
wire u5__abc_78290_new_n2591_; 
wire u5__abc_78290_new_n2592_; 
wire u5__abc_78290_new_n2593_; 
wire u5__abc_78290_new_n2594_; 
wire u5__abc_78290_new_n2595_; 
wire u5__abc_78290_new_n2596_; 
wire u5__abc_78290_new_n2597_; 
wire u5__abc_78290_new_n2598_; 
wire u5__abc_78290_new_n2599_; 
wire u5__abc_78290_new_n2600_; 
wire u5__abc_78290_new_n2601_; 
wire u5__abc_78290_new_n2602_; 
wire u5__abc_78290_new_n2603_; 
wire u5__abc_78290_new_n2605_; 
wire u5__abc_78290_new_n2606_; 
wire u5__abc_78290_new_n2607_; 
wire u5__abc_78290_new_n2608_; 
wire u5__abc_78290_new_n2609_; 
wire u5__abc_78290_new_n2610_; 
wire u5__abc_78290_new_n2611_; 
wire u5__abc_78290_new_n2612_; 
wire u5__abc_78290_new_n2613_; 
wire u5__abc_78290_new_n2614_; 
wire u5__abc_78290_new_n2615_; 
wire u5__abc_78290_new_n2616_; 
wire u5__abc_78290_new_n2617_; 
wire u5__abc_78290_new_n2618_; 
wire u5__abc_78290_new_n2619_; 
wire u5__abc_78290_new_n2620_; 
wire u5__abc_78290_new_n2621_; 
wire u5__abc_78290_new_n2622_; 
wire u5__abc_78290_new_n2623_; 
wire u5__abc_78290_new_n2624_; 
wire u5__abc_78290_new_n2625_; 
wire u5__abc_78290_new_n2626_; 
wire u5__abc_78290_new_n2627_; 
wire u5__abc_78290_new_n2628_; 
wire u5__abc_78290_new_n2629_; 
wire u5__abc_78290_new_n2630_; 
wire u5__abc_78290_new_n2631_; 
wire u5__abc_78290_new_n2632_; 
wire u5__abc_78290_new_n2633_; 
wire u5__abc_78290_new_n2634_; 
wire u5__abc_78290_new_n2635_; 
wire u5__abc_78290_new_n2636_; 
wire u5__abc_78290_new_n2637_; 
wire u5__abc_78290_new_n2638_; 
wire u5__abc_78290_new_n2639_; 
wire u5__abc_78290_new_n2640_; 
wire u5__abc_78290_new_n2641_; 
wire u5__abc_78290_new_n2643_; 
wire u5__abc_78290_new_n2644_; 
wire u5__abc_78290_new_n2645_; 
wire u5__abc_78290_new_n2647_; 
wire u5__abc_78290_new_n2648_; 
wire u5__abc_78290_new_n2649_; 
wire u5__abc_78290_new_n2650_; 
wire u5__abc_78290_new_n2651_; 
wire u5__abc_78290_new_n2652_; 
wire u5__abc_78290_new_n2653_; 
wire u5__abc_78290_new_n2654_; 
wire u5__abc_78290_new_n2655_; 
wire u5__abc_78290_new_n2656_; 
wire u5__abc_78290_new_n2657_; 
wire u5__abc_78290_new_n2659_; 
wire u5__abc_78290_new_n2660_; 
wire u5__abc_78290_new_n2661_; 
wire u5__abc_78290_new_n2663_; 
wire u5__abc_78290_new_n2664_; 
wire u5__abc_78290_new_n2665_; 
wire u5__abc_78290_new_n2666_; 
wire u5__abc_78290_new_n2667_; 
wire u5__abc_78290_new_n2668_; 
wire u5__abc_78290_new_n2669_; 
wire u5__abc_78290_new_n2670_; 
wire u5__abc_78290_new_n2671_; 
wire u5__abc_78290_new_n2672_; 
wire u5__abc_78290_new_n2673_; 
wire u5__abc_78290_new_n2674_; 
wire u5__abc_78290_new_n2675_; 
wire u5__abc_78290_new_n2676_; 
wire u5__abc_78290_new_n2678_; 
wire u5__abc_78290_new_n2679_; 
wire u5__abc_78290_new_n2680_; 
wire u5__abc_78290_new_n2681_; 
wire u5__abc_78290_new_n2682_; 
wire u5__abc_78290_new_n2683_; 
wire u5__abc_78290_new_n2684_; 
wire u5__abc_78290_new_n2685_; 
wire u5__abc_78290_new_n2687_; 
wire u5__abc_78290_new_n2688_; 
wire u5__abc_78290_new_n2689_; 
wire u5__abc_78290_new_n2690_; 
wire u5__abc_78290_new_n2691_; 
wire u5__abc_78290_new_n2692_; 
wire u5__abc_78290_new_n2693_; 
wire u5__abc_78290_new_n2694_; 
wire u5__abc_78290_new_n2696_; 
wire u5__abc_78290_new_n2697_; 
wire u5__abc_78290_new_n2698_; 
wire u5__abc_78290_new_n2699_; 
wire u5__abc_78290_new_n2700_; 
wire u5__abc_78290_new_n2701_; 
wire u5__abc_78290_new_n2702_; 
wire u5__abc_78290_new_n2703_; 
wire u5__abc_78290_new_n2704_; 
wire u5__abc_78290_new_n2705_; 
wire u5__abc_78290_new_n2706_; 
wire u5__abc_78290_new_n2707_; 
wire u5__abc_78290_new_n2709_; 
wire u5__abc_78290_new_n2710_; 
wire u5__abc_78290_new_n2712_; 
wire u5__abc_78290_new_n2713_; 
wire u5__abc_78290_new_n2714_; 
wire u5__abc_78290_new_n2715_; 
wire u5__abc_78290_new_n2716_; 
wire u5__abc_78290_new_n2717_; 
wire u5__abc_78290_new_n2718_; 
wire u5__abc_78290_new_n2719_; 
wire u5__abc_78290_new_n2721_; 
wire u5__abc_78290_new_n2722_; 
wire u5__abc_78290_new_n2723_; 
wire u5__abc_78290_new_n2724_; 
wire u5__abc_78290_new_n2726_; 
wire u5__abc_78290_new_n2727_; 
wire u5__abc_78290_new_n2728_; 
wire u5__abc_78290_new_n2729_; 
wire u5__abc_78290_new_n2731_; 
wire u5__abc_78290_new_n2732_; 
wire u5__abc_78290_new_n2733_; 
wire u5__abc_78290_new_n2734_; 
wire u5__abc_78290_new_n2735_; 
wire u5__abc_78290_new_n2736_; 
wire u5__abc_78290_new_n2737_; 
wire u5__abc_78290_new_n2738_; 
wire u5__abc_78290_new_n2740_; 
wire u5__abc_78290_new_n2741_; 
wire u5__abc_78290_new_n2742_; 
wire u5__abc_78290_new_n2743_; 
wire u5__abc_78290_new_n2744_; 
wire u5__abc_78290_new_n2745_; 
wire u5__abc_78290_new_n2746_; 
wire u5__abc_78290_new_n2747_; 
wire u5__abc_78290_new_n2748_; 
wire u5__abc_78290_new_n2749_; 
wire u5__abc_78290_new_n2750_; 
wire u5__abc_78290_new_n2751_; 
wire u5__abc_78290_new_n2752_; 
wire u5__abc_78290_new_n2753_; 
wire u5__abc_78290_new_n2754_; 
wire u5__abc_78290_new_n2756_; 
wire u5__abc_78290_new_n2757_; 
wire u5__abc_78290_new_n2758_; 
wire u5__abc_78290_new_n2759_; 
wire u5__abc_78290_new_n2760_; 
wire u5__abc_78290_new_n2761_; 
wire u5__abc_78290_new_n2762_; 
wire u5__abc_78290_new_n2763_; 
wire u5__abc_78290_new_n2764_; 
wire u5__abc_78290_new_n2765_; 
wire u5__abc_78290_new_n2766_; 
wire u5__abc_78290_new_n2767_; 
wire u5__abc_78290_new_n2768_; 
wire u5__abc_78290_new_n2769_; 
wire u5__abc_78290_new_n2770_; 
wire u5__abc_78290_new_n2772_; 
wire u5__abc_78290_new_n2773_; 
wire u5__abc_78290_new_n2774_; 
wire u5__abc_78290_new_n2775_; 
wire u5__abc_78290_new_n2776_; 
wire u5__abc_78290_new_n2777_; 
wire u5__abc_78290_new_n2778_; 
wire u5__abc_78290_new_n2779_; 
wire u5__abc_78290_new_n2780_; 
wire u5__abc_78290_new_n2782_; 
wire u5__abc_78290_new_n2783_; 
wire u5__abc_78290_new_n2784_; 
wire u5__abc_78290_new_n2785_; 
wire u5__abc_78290_new_n2786_; 
wire u5__abc_78290_new_n2788_; 
wire u5__abc_78290_new_n2789_; 
wire u5__abc_78290_new_n2790_; 
wire u5__abc_78290_new_n2791_; 
wire u5__abc_78290_new_n2792_; 
wire u5__abc_78290_new_n2793_; 
wire u5__abc_78290_new_n2795_; 
wire u5__abc_78290_new_n2796_; 
wire u5__abc_78290_new_n2797_; 
wire u5__abc_78290_new_n2798_; 
wire u5__abc_78290_new_n2799_; 
wire u5__abc_78290_new_n2800_; 
wire u5__abc_78290_new_n2802_; 
wire u5__abc_78290_new_n2804_; 
wire u5__abc_78290_new_n2805_; 
wire u5__abc_78290_new_n2806_; 
wire u5__abc_78290_new_n2808_; 
wire u5__abc_78290_new_n2809_; 
wire u5__abc_78290_new_n2810_; 
wire u5__abc_78290_new_n2811_; 
wire u5__abc_78290_new_n2813_; 
wire u5__abc_78290_new_n2814_; 
wire u5__abc_78290_new_n2815_; 
wire u5__abc_78290_new_n2816_; 
wire u5__abc_78290_new_n2817_; 
wire u5__abc_78290_new_n2818_; 
wire u5__abc_78290_new_n2820_; 
wire u5__abc_78290_new_n2821_; 
wire u5__abc_78290_new_n2822_; 
wire u5__abc_78290_new_n2823_; 
wire u5__abc_78290_new_n2825_; 
wire u5__abc_78290_new_n2826_; 
wire u5__abc_78290_new_n2827_; 
wire u5__abc_78290_new_n2828_; 
wire u5__abc_78290_new_n2830_; 
wire u5__abc_78290_new_n2831_; 
wire u5__abc_78290_new_n2833_; 
wire u5__abc_78290_new_n2834_; 
wire u5__abc_78290_new_n2835_; 
wire u5__abc_78290_new_n2836_; 
wire u5__abc_78290_new_n2837_; 
wire u5__abc_78290_new_n2839_; 
wire u5__abc_78290_new_n2840_; 
wire u5__abc_78290_new_n2841_; 
wire u5__abc_78290_new_n2842_; 
wire u5__abc_78290_new_n2844_; 
wire u5__abc_78290_new_n2845_; 
wire u5__abc_78290_new_n2846_; 
wire u5__abc_78290_new_n2847_; 
wire u5__abc_78290_new_n2849_; 
wire u5__abc_78290_new_n2850_; 
wire u5__abc_78290_new_n2852_; 
wire u5__abc_78290_new_n2853_; 
wire u5__abc_78290_new_n2854_; 
wire u5__abc_78290_new_n2856_; 
wire u5__abc_78290_new_n2859_; 
wire u5__abc_78290_new_n2861_; 
wire u5__abc_78290_new_n2862_; 
wire u5__abc_78290_new_n2863_; 
wire u5__abc_78290_new_n2864_; 
wire u5__abc_78290_new_n2865_; 
wire u5__abc_78290_new_n2866_; 
wire u5__abc_78290_new_n2867_; 
wire u5__abc_78290_new_n2869_; 
wire u5__abc_78290_new_n2870_; 
wire u5__abc_78290_new_n2871_; 
wire u5__abc_78290_new_n2873_; 
wire u5__abc_78290_new_n2874_; 
wire u5__abc_78290_new_n2875_; 
wire u5__abc_78290_new_n2877_; 
wire u5__abc_78290_new_n2878_; 
wire u5__abc_78290_new_n2879_; 
wire u5__abc_78290_new_n2882_; 
wire u5__abc_78290_new_n2883_; 
wire u5__abc_78290_new_n2884_; 
wire u5__abc_78290_new_n2886_; 
wire u5__abc_78290_new_n2887_; 
wire u5__abc_78290_new_n2888_; 
wire u5__abc_78290_new_n2890_; 
wire u5__abc_78290_new_n2891_; 
wire u5__abc_78290_new_n2893_; 
wire u5__abc_78290_new_n2894_; 
wire u5__abc_78290_new_n2896_; 
wire u5__abc_78290_new_n2897_; 
wire u5__abc_78290_new_n2898_; 
wire u5__abc_78290_new_n2899_; 
wire u5__abc_78290_new_n2900_; 
wire u5__abc_78290_new_n2902_; 
wire u5__abc_78290_new_n2903_; 
wire u5__abc_78290_new_n2905_; 
wire u5__abc_78290_new_n2906_; 
wire u5__abc_78290_new_n2908_; 
wire u5__abc_78290_new_n2909_; 
wire u5__abc_78290_new_n2910_; 
wire u5__abc_78290_new_n2912_; 
wire u5__abc_78290_new_n2914_; 
wire u5__abc_78290_new_n2915_; 
wire u5__abc_78290_new_n2917_; 
wire u5__abc_78290_new_n2919_; 
wire u5__abc_78290_new_n2920_; 
wire u5__abc_78290_new_n2921_; 
wire u5__abc_78290_new_n2922_; 
wire u5__abc_78290_new_n2923_; 
wire u5__abc_78290_new_n2924_; 
wire u5__abc_78290_new_n2926_; 
wire u5__abc_78290_new_n2927_; 
wire u5__abc_78290_new_n2928_; 
wire u5__abc_78290_new_n2930_; 
wire u5__abc_78290_new_n2931_; 
wire u5__abc_78290_new_n2932_; 
wire u5__abc_78290_new_n2934_; 
wire u5__abc_78290_new_n2935_; 
wire u5__abc_78290_new_n2936_; 
wire u5__abc_78290_new_n2937_; 
wire u5__abc_78290_new_n2938_; 
wire u5__abc_78290_new_n2940_; 
wire u5__abc_78290_new_n2941_; 
wire u5__abc_78290_new_n2942_; 
wire u5__abc_78290_new_n2943_; 
wire u5__abc_78290_new_n2944_; 
wire u5__abc_78290_new_n2945_; 
wire u5__abc_78290_new_n2947_; 
wire u5__abc_78290_new_n2948_; 
wire u5__abc_78290_new_n2949_; 
wire u5__abc_78290_new_n2950_; 
wire u5__abc_78290_new_n2951_; 
wire u5__abc_78290_new_n2952_; 
wire u5__abc_78290_new_n2953_; 
wire u5__abc_78290_new_n2954_; 
wire u5__abc_78290_new_n2956_; 
wire u5__abc_78290_new_n2957_; 
wire u5__abc_78290_new_n2958_; 
wire u5__abc_78290_new_n2959_; 
wire u5__abc_78290_new_n2960_; 
wire u5__abc_78290_new_n2961_; 
wire u5__abc_78290_new_n2963_; 
wire u5__abc_78290_new_n2964_; 
wire u5__abc_78290_new_n2965_; 
wire u5__abc_78290_new_n2967_; 
wire u5__abc_78290_new_n2968_; 
wire u5__abc_78290_new_n2969_; 
wire u5__abc_78290_new_n2970_; 
wire u5__abc_78290_new_n2971_; 
wire u5__abc_78290_new_n2973_; 
wire u5__abc_78290_new_n2974_; 
wire u5__abc_78290_new_n2975_; 
wire u5__abc_78290_new_n2976_; 
wire u5__abc_78290_new_n2977_; 
wire u5__abc_78290_new_n2979_; 
wire u5__abc_78290_new_n2981_; 
wire u5__abc_78290_new_n2982_; 
wire u5__abc_78290_new_n2983_; 
wire u5__abc_78290_new_n2984_; 
wire u5__abc_78290_new_n2985_; 
wire u5__abc_78290_new_n2987_; 
wire u5__abc_78290_new_n2988_; 
wire u5__abc_78290_new_n2989_; 
wire u5__abc_78290_new_n2991_; 
wire u5__abc_78290_new_n2993_; 
wire u5__abc_78290_new_n2994_; 
wire u5__abc_78290_new_n2995_; 
wire u5__abc_78290_new_n2996_; 
wire u5__abc_78290_new_n2997_; 
wire u5__abc_78290_new_n2998_; 
wire u5__abc_78290_new_n2999_; 
wire u5__abc_78290_new_n3000_; 
wire u5__abc_78290_new_n3001_; 
wire u5__abc_78290_new_n3003_; 
wire u5__abc_78290_new_n3004_; 
wire u5__abc_78290_new_n3005_; 
wire u5__abc_78290_new_n3006_; 
wire u5__abc_78290_new_n3007_; 
wire u5__abc_78290_new_n3008_; 
wire u5__abc_78290_new_n3009_; 
wire u5__abc_78290_new_n3010_; 
wire u5__abc_78290_new_n3011_; 
wire u5__abc_78290_new_n3012_; 
wire u5__abc_78290_new_n3013_; 
wire u5__abc_78290_new_n3014_; 
wire u5__abc_78290_new_n3016_; 
wire u5__abc_78290_new_n3017_; 
wire u5__abc_78290_new_n3018_; 
wire u5__abc_78290_new_n3019_; 
wire u5__abc_78290_new_n3020_; 
wire u5__abc_78290_new_n3021_; 
wire u5__abc_78290_new_n3023_; 
wire u5__abc_78290_new_n3024_; 
wire u5__abc_78290_new_n3026_; 
wire u5__abc_78290_new_n3027_; 
wire u5__abc_78290_new_n3028_; 
wire u5__abc_78290_new_n3029_; 
wire u5__abc_78290_new_n3030_; 
wire u5__abc_78290_new_n3031_; 
wire u5__abc_78290_new_n3032_; 
wire u5__abc_78290_new_n3033_; 
wire u5__abc_78290_new_n3035_; 
wire u5__abc_78290_new_n3036_; 
wire u5__abc_78290_new_n3037_; 
wire u5__abc_78290_new_n3038_; 
wire u5__abc_78290_new_n3039_; 
wire u5__abc_78290_new_n3040_; 
wire u5__abc_78290_new_n3041_; 
wire u5__abc_78290_new_n3042_; 
wire u5__abc_78290_new_n3043_; 
wire u5__abc_78290_new_n3044_; 
wire u5__abc_78290_new_n3045_; 
wire u5__abc_78290_new_n3046_; 
wire u5__abc_78290_new_n3047_; 
wire u5__abc_78290_new_n3048_; 
wire u5__abc_78290_new_n3050_; 
wire u5__abc_78290_new_n3051_; 
wire u5__abc_78290_new_n3052_; 
wire u5__abc_78290_new_n3053_; 
wire u5__abc_78290_new_n3054_; 
wire u5__abc_78290_new_n3055_; 
wire u5__abc_78290_new_n3056_; 
wire u5__abc_78290_new_n3057_; 
wire u5__abc_78290_new_n3058_; 
wire u5__abc_78290_new_n3060_; 
wire u5__abc_78290_new_n3061_; 
wire u5__abc_78290_new_n3062_; 
wire u5__abc_78290_new_n3063_; 
wire u5__abc_78290_new_n3064_; 
wire u5__abc_78290_new_n3065_; 
wire u5__abc_78290_new_n3067_; 
wire u5__abc_78290_new_n3068_; 
wire u5__abc_78290_new_n3069_; 
wire u5__abc_78290_new_n3070_; 
wire u5__abc_78290_new_n3072_; 
wire u5__abc_78290_new_n3073_; 
wire u5__abc_78290_new_n3074_; 
wire u5__abc_78290_new_n3075_; 
wire u5__abc_78290_new_n3076_; 
wire u5__abc_78290_new_n3077_; 
wire u5__abc_78290_new_n3078_; 
wire u5__abc_78290_new_n3079_; 
wire u5__abc_78290_new_n3080_; 
wire u5__abc_78290_new_n3081_; 
wire u5__abc_78290_new_n3082_; 
wire u5__abc_78290_new_n3084_; 
wire u5__abc_78290_new_n3085_; 
wire u5__abc_78290_new_n3087_; 
wire u5__abc_78290_new_n3088_; 
wire u5__abc_78290_new_n3089_; 
wire u5__abc_78290_new_n3090_; 
wire u5__abc_78290_new_n3091_; 
wire u5__abc_78290_new_n3092_; 
wire u5__abc_78290_new_n3093_; 
wire u5__abc_78290_new_n3094_; 
wire u5__abc_78290_new_n3095_; 
wire u5__abc_78290_new_n3096_; 
wire u5__abc_78290_new_n3097_; 
wire u5__abc_78290_new_n3098_; 
wire u5__abc_78290_new_n3099_; 
wire u5__abc_78290_new_n3100_; 
wire u5__abc_78290_new_n3101_; 
wire u5__abc_78290_new_n3102_; 
wire u5__abc_78290_new_n3103_; 
wire u5__abc_78290_new_n3104_; 
wire u5__abc_78290_new_n3105_; 
wire u5__abc_78290_new_n3106_; 
wire u5__abc_78290_new_n3107_; 
wire u5__abc_78290_new_n3108_; 
wire u5__abc_78290_new_n3109_; 
wire u5__abc_78290_new_n3110_; 
wire u5__abc_78290_new_n3111_; 
wire u5__abc_78290_new_n3112_; 
wire u5__abc_78290_new_n3113_; 
wire u5__abc_78290_new_n3114_; 
wire u5__abc_78290_new_n3116_; 
wire u5__abc_78290_new_n3117_; 
wire u5__abc_78290_new_n3118_; 
wire u5__abc_78290_new_n3119_; 
wire u5__abc_78290_new_n3121_; 
wire u5__abc_78290_new_n3122_; 
wire u5__abc_78290_new_n3123_; 
wire u5__abc_78290_new_n3124_; 
wire u5__abc_78290_new_n3126_; 
wire u5__abc_78290_new_n3127_; 
wire u5__abc_78290_new_n3129_; 
wire u5__abc_78290_new_n3130_; 
wire u5__abc_78290_new_n3132_; 
wire u5__abc_78290_new_n3133_; 
wire u5__abc_78290_new_n3134_; 
wire u5__abc_78290_new_n3135_; 
wire u5__abc_78290_new_n3136_; 
wire u5__abc_78290_new_n3137_; 
wire u5__abc_78290_new_n3138_; 
wire u5__abc_78290_new_n3139_; 
wire u5__abc_78290_new_n3141_; 
wire u5__abc_78290_new_n3143_; 
wire u5__abc_78290_new_n3145_; 
wire u5__abc_78290_new_n3146_; 
wire u5__abc_78290_new_n3147_; 
wire u5__abc_78290_new_n3149_; 
wire u5__abc_78290_new_n3150_; 
wire u5__abc_78290_new_n3151_; 
wire u5__abc_78290_new_n3153_; 
wire u5__abc_78290_new_n3155_; 
wire u5__abc_78290_new_n3156_; 
wire u5__abc_78290_new_n3157_; 
wire u5__abc_78290_new_n366_; 
wire u5__abc_78290_new_n367_; 
wire u5__abc_78290_new_n368_; 
wire u5__abc_78290_new_n369_; 
wire u5__abc_78290_new_n370_; 
wire u5__abc_78290_new_n371_; 
wire u5__abc_78290_new_n372_; 
wire u5__abc_78290_new_n373_; 
wire u5__abc_78290_new_n374_; 
wire u5__abc_78290_new_n375_; 
wire u5__abc_78290_new_n376_; 
wire u5__abc_78290_new_n378_; 
wire u5__abc_78290_new_n379_; 
wire u5__abc_78290_new_n380_; 
wire u5__abc_78290_new_n381_; 
wire u5__abc_78290_new_n382_; 
wire u5__abc_78290_new_n383_; 
wire u5__abc_78290_new_n384_; 
wire u5__abc_78290_new_n385_; 
wire u5__abc_78290_new_n386_; 
wire u5__abc_78290_new_n387_; 
wire u5__abc_78290_new_n388_; 
wire u5__abc_78290_new_n389_; 
wire u5__abc_78290_new_n390_; 
wire u5__abc_78290_new_n391_; 
wire u5__abc_78290_new_n392_; 
wire u5__abc_78290_new_n393_; 
wire u5__abc_78290_new_n394_; 
wire u5__abc_78290_new_n395_; 
wire u5__abc_78290_new_n396_; 
wire u5__abc_78290_new_n397_; 
wire u5__abc_78290_new_n398_; 
wire u5__abc_78290_new_n399_; 
wire u5__abc_78290_new_n400_; 
wire u5__abc_78290_new_n401_; 
wire u5__abc_78290_new_n402_; 
wire u5__abc_78290_new_n403_; 
wire u5__abc_78290_new_n404_; 
wire u5__abc_78290_new_n405_; 
wire u5__abc_78290_new_n406_; 
wire u5__abc_78290_new_n407_; 
wire u5__abc_78290_new_n408_; 
wire u5__abc_78290_new_n409_; 
wire u5__abc_78290_new_n410_; 
wire u5__abc_78290_new_n411_; 
wire u5__abc_78290_new_n412_; 
wire u5__abc_78290_new_n413_; 
wire u5__abc_78290_new_n414_; 
wire u5__abc_78290_new_n415_; 
wire u5__abc_78290_new_n416_; 
wire u5__abc_78290_new_n417_; 
wire u5__abc_78290_new_n418_; 
wire u5__abc_78290_new_n419_; 
wire u5__abc_78290_new_n420_; 
wire u5__abc_78290_new_n421_; 
wire u5__abc_78290_new_n422_; 
wire u5__abc_78290_new_n423_; 
wire u5__abc_78290_new_n424_; 
wire u5__abc_78290_new_n425_; 
wire u5__abc_78290_new_n426_; 
wire u5__abc_78290_new_n427_; 
wire u5__abc_78290_new_n428_; 
wire u5__abc_78290_new_n429_; 
wire u5__abc_78290_new_n430_; 
wire u5__abc_78290_new_n431_; 
wire u5__abc_78290_new_n432_; 
wire u5__abc_78290_new_n433_; 
wire u5__abc_78290_new_n434_; 
wire u5__abc_78290_new_n435_; 
wire u5__abc_78290_new_n436_; 
wire u5__abc_78290_new_n437_; 
wire u5__abc_78290_new_n438_; 
wire u5__abc_78290_new_n439_; 
wire u5__abc_78290_new_n440_; 
wire u5__abc_78290_new_n441_; 
wire u5__abc_78290_new_n442_; 
wire u5__abc_78290_new_n443_; 
wire u5__abc_78290_new_n444_; 
wire u5__abc_78290_new_n445_; 
wire u5__abc_78290_new_n446_; 
wire u5__abc_78290_new_n447_; 
wire u5__abc_78290_new_n448_; 
wire u5__abc_78290_new_n449_; 
wire u5__abc_78290_new_n450_; 
wire u5__abc_78290_new_n451_; 
wire u5__abc_78290_new_n452_; 
wire u5__abc_78290_new_n453_; 
wire u5__abc_78290_new_n454_; 
wire u5__abc_78290_new_n455_; 
wire u5__abc_78290_new_n456_; 
wire u5__abc_78290_new_n457_; 
wire u5__abc_78290_new_n458_; 
wire u5__abc_78290_new_n459_; 
wire u5__abc_78290_new_n460_; 
wire u5__abc_78290_new_n461_; 
wire u5__abc_78290_new_n462_; 
wire u5__abc_78290_new_n463_; 
wire u5__abc_78290_new_n464_; 
wire u5__abc_78290_new_n465_; 
wire u5__abc_78290_new_n466_; 
wire u5__abc_78290_new_n467_; 
wire u5__abc_78290_new_n468_; 
wire u5__abc_78290_new_n469_; 
wire u5__abc_78290_new_n470_; 
wire u5__abc_78290_new_n471_; 
wire u5__abc_78290_new_n472_; 
wire u5__abc_78290_new_n473_; 
wire u5__abc_78290_new_n474_; 
wire u5__abc_78290_new_n475_; 
wire u5__abc_78290_new_n476_; 
wire u5__abc_78290_new_n477_; 
wire u5__abc_78290_new_n478_; 
wire u5__abc_78290_new_n479_; 
wire u5__abc_78290_new_n480_; 
wire u5__abc_78290_new_n481_; 
wire u5__abc_78290_new_n482_; 
wire u5__abc_78290_new_n483_; 
wire u5__abc_78290_new_n484_; 
wire u5__abc_78290_new_n486_; 
wire u5__abc_78290_new_n487_; 
wire u5__abc_78290_new_n488_; 
wire u5__abc_78290_new_n489_; 
wire u5__abc_78290_new_n490_; 
wire u5__abc_78290_new_n491_; 
wire u5__abc_78290_new_n492_; 
wire u5__abc_78290_new_n493_; 
wire u5__abc_78290_new_n494_; 
wire u5__abc_78290_new_n495_; 
wire u5__abc_78290_new_n496_; 
wire u5__abc_78290_new_n497_; 
wire u5__abc_78290_new_n498_; 
wire u5__abc_78290_new_n499_; 
wire u5__abc_78290_new_n500_; 
wire u5__abc_78290_new_n501_; 
wire u5__abc_78290_new_n502_; 
wire u5__abc_78290_new_n503_; 
wire u5__abc_78290_new_n504_; 
wire u5__abc_78290_new_n505_; 
wire u5__abc_78290_new_n506_; 
wire u5__abc_78290_new_n507_; 
wire u5__abc_78290_new_n508_; 
wire u5__abc_78290_new_n509_; 
wire u5__abc_78290_new_n510_; 
wire u5__abc_78290_new_n511_; 
wire u5__abc_78290_new_n512_; 
wire u5__abc_78290_new_n513_; 
wire u5__abc_78290_new_n514_; 
wire u5__abc_78290_new_n515_; 
wire u5__abc_78290_new_n516_; 
wire u5__abc_78290_new_n517_; 
wire u5__abc_78290_new_n518_; 
wire u5__abc_78290_new_n519_; 
wire u5__abc_78290_new_n520_; 
wire u5__abc_78290_new_n521_; 
wire u5__abc_78290_new_n522_; 
wire u5__abc_78290_new_n523_; 
wire u5__abc_78290_new_n524_; 
wire u5__abc_78290_new_n525_; 
wire u5__abc_78290_new_n526_; 
wire u5__abc_78290_new_n527_; 
wire u5__abc_78290_new_n528_; 
wire u5__abc_78290_new_n529_; 
wire u5__abc_78290_new_n530_; 
wire u5__abc_78290_new_n531_; 
wire u5__abc_78290_new_n532_; 
wire u5__abc_78290_new_n533_; 
wire u5__abc_78290_new_n534_; 
wire u5__abc_78290_new_n535_; 
wire u5__abc_78290_new_n536_; 
wire u5__abc_78290_new_n537_; 
wire u5__abc_78290_new_n538_; 
wire u5__abc_78290_new_n539_; 
wire u5__abc_78290_new_n540_; 
wire u5__abc_78290_new_n541_; 
wire u5__abc_78290_new_n542_; 
wire u5__abc_78290_new_n543_; 
wire u5__abc_78290_new_n544_; 
wire u5__abc_78290_new_n545_; 
wire u5__abc_78290_new_n546_; 
wire u5__abc_78290_new_n547_; 
wire u5__abc_78290_new_n548_; 
wire u5__abc_78290_new_n549_; 
wire u5__abc_78290_new_n550_; 
wire u5__abc_78290_new_n551_; 
wire u5__abc_78290_new_n552_; 
wire u5__abc_78290_new_n553_; 
wire u5__abc_78290_new_n554_; 
wire u5__abc_78290_new_n555_; 
wire u5__abc_78290_new_n556_; 
wire u5__abc_78290_new_n557_; 
wire u5__abc_78290_new_n558_; 
wire u5__abc_78290_new_n559_; 
wire u5__abc_78290_new_n560_; 
wire u5__abc_78290_new_n561_; 
wire u5__abc_78290_new_n562_; 
wire u5__abc_78290_new_n563_; 
wire u5__abc_78290_new_n564_; 
wire u5__abc_78290_new_n565_; 
wire u5__abc_78290_new_n566_; 
wire u5__abc_78290_new_n567_; 
wire u5__abc_78290_new_n568_; 
wire u5__abc_78290_new_n569_; 
wire u5__abc_78290_new_n570_; 
wire u5__abc_78290_new_n571_; 
wire u5__abc_78290_new_n572_; 
wire u5__abc_78290_new_n573_; 
wire u5__abc_78290_new_n574_; 
wire u5__abc_78290_new_n575_; 
wire u5__abc_78290_new_n576_; 
wire u5__abc_78290_new_n577_; 
wire u5__abc_78290_new_n578_; 
wire u5__abc_78290_new_n579_; 
wire u5__abc_78290_new_n580_; 
wire u5__abc_78290_new_n581_; 
wire u5__abc_78290_new_n582_; 
wire u5__abc_78290_new_n583_; 
wire u5__abc_78290_new_n584_; 
wire u5__abc_78290_new_n585_; 
wire u5__abc_78290_new_n586_; 
wire u5__abc_78290_new_n587_; 
wire u5__abc_78290_new_n588_; 
wire u5__abc_78290_new_n589_; 
wire u5__abc_78290_new_n590_; 
wire u5__abc_78290_new_n591_; 
wire u5__abc_78290_new_n592_; 
wire u5__abc_78290_new_n593_; 
wire u5__abc_78290_new_n594_; 
wire u5__abc_78290_new_n595_; 
wire u5__abc_78290_new_n596_; 
wire u5__abc_78290_new_n597_; 
wire u5__abc_78290_new_n598_; 
wire u5__abc_78290_new_n599_; 
wire u5__abc_78290_new_n600_; 
wire u5__abc_78290_new_n601_; 
wire u5__abc_78290_new_n602_; 
wire u5__abc_78290_new_n603_; 
wire u5__abc_78290_new_n604_; 
wire u5__abc_78290_new_n605_; 
wire u5__abc_78290_new_n606_; 
wire u5__abc_78290_new_n607_; 
wire u5__abc_78290_new_n608_; 
wire u5__abc_78290_new_n609_; 
wire u5__abc_78290_new_n610_; 
wire u5__abc_78290_new_n611_; 
wire u5__abc_78290_new_n612_; 
wire u5__abc_78290_new_n613_; 
wire u5__abc_78290_new_n614_; 
wire u5__abc_78290_new_n615_; 
wire u5__abc_78290_new_n616_; 
wire u5__abc_78290_new_n617_; 
wire u5__abc_78290_new_n618_; 
wire u5__abc_78290_new_n619_; 
wire u5__abc_78290_new_n620_; 
wire u5__abc_78290_new_n621_; 
wire u5__abc_78290_new_n622_; 
wire u5__abc_78290_new_n623_; 
wire u5__abc_78290_new_n624_; 
wire u5__abc_78290_new_n625_; 
wire u5__abc_78290_new_n626_; 
wire u5__abc_78290_new_n627_; 
wire u5__abc_78290_new_n628_; 
wire u5__abc_78290_new_n629_; 
wire u5__abc_78290_new_n630_; 
wire u5__abc_78290_new_n631_; 
wire u5__abc_78290_new_n632_; 
wire u5__abc_78290_new_n633_; 
wire u5__abc_78290_new_n634_; 
wire u5__abc_78290_new_n635_; 
wire u5__abc_78290_new_n636_; 
wire u5__abc_78290_new_n637_; 
wire u5__abc_78290_new_n638_; 
wire u5__abc_78290_new_n639_; 
wire u5__abc_78290_new_n640_; 
wire u5__abc_78290_new_n641_; 
wire u5__abc_78290_new_n642_; 
wire u5__abc_78290_new_n643_; 
wire u5__abc_78290_new_n644_; 
wire u5__abc_78290_new_n645_; 
wire u5__abc_78290_new_n646_; 
wire u5__abc_78290_new_n647_; 
wire u5__abc_78290_new_n648_; 
wire u5__abc_78290_new_n649_; 
wire u5__abc_78290_new_n650_; 
wire u5__abc_78290_new_n651_; 
wire u5__abc_78290_new_n652_; 
wire u5__abc_78290_new_n653_; 
wire u5__abc_78290_new_n654_; 
wire u5__abc_78290_new_n655_; 
wire u5__abc_78290_new_n656_; 
wire u5__abc_78290_new_n657_; 
wire u5__abc_78290_new_n658_; 
wire u5__abc_78290_new_n659_; 
wire u5__abc_78290_new_n660_; 
wire u5__abc_78290_new_n661_; 
wire u5__abc_78290_new_n662_; 
wire u5__abc_78290_new_n663_; 
wire u5__abc_78290_new_n664_; 
wire u5__abc_78290_new_n665_; 
wire u5__abc_78290_new_n666_; 
wire u5__abc_78290_new_n667_; 
wire u5__abc_78290_new_n668_; 
wire u5__abc_78290_new_n669_; 
wire u5__abc_78290_new_n670_; 
wire u5__abc_78290_new_n671_; 
wire u5__abc_78290_new_n672_; 
wire u5__abc_78290_new_n673_; 
wire u5__abc_78290_new_n674_; 
wire u5__abc_78290_new_n675_; 
wire u5__abc_78290_new_n676_; 
wire u5__abc_78290_new_n677_; 
wire u5__abc_78290_new_n678_; 
wire u5__abc_78290_new_n679_; 
wire u5__abc_78290_new_n680_; 
wire u5__abc_78290_new_n681_; 
wire u5__abc_78290_new_n682_; 
wire u5__abc_78290_new_n683_; 
wire u5__abc_78290_new_n684_; 
wire u5__abc_78290_new_n685_; 
wire u5__abc_78290_new_n686_; 
wire u5__abc_78290_new_n687_; 
wire u5__abc_78290_new_n688_; 
wire u5__abc_78290_new_n689_; 
wire u5__abc_78290_new_n690_; 
wire u5__abc_78290_new_n691_; 
wire u5__abc_78290_new_n692_; 
wire u5__abc_78290_new_n693_; 
wire u5__abc_78290_new_n694_; 
wire u5__abc_78290_new_n695_; 
wire u5__abc_78290_new_n696_; 
wire u5__abc_78290_new_n697_; 
wire u5__abc_78290_new_n698_; 
wire u5__abc_78290_new_n699_; 
wire u5__abc_78290_new_n700_; 
wire u5__abc_78290_new_n701_; 
wire u5__abc_78290_new_n702_; 
wire u5__abc_78290_new_n703_; 
wire u5__abc_78290_new_n704_; 
wire u5__abc_78290_new_n705_; 
wire u5__abc_78290_new_n706_; 
wire u5__abc_78290_new_n707_; 
wire u5__abc_78290_new_n708_; 
wire u5__abc_78290_new_n709_; 
wire u5__abc_78290_new_n710_; 
wire u5__abc_78290_new_n711_; 
wire u5__abc_78290_new_n712_; 
wire u5__abc_78290_new_n713_; 
wire u5__abc_78290_new_n714_; 
wire u5__abc_78290_new_n715_; 
wire u5__abc_78290_new_n716_; 
wire u5__abc_78290_new_n717_; 
wire u5__abc_78290_new_n718_; 
wire u5__abc_78290_new_n719_; 
wire u5__abc_78290_new_n720_; 
wire u5__abc_78290_new_n721_; 
wire u5__abc_78290_new_n722_; 
wire u5__abc_78290_new_n723_; 
wire u5__abc_78290_new_n724_; 
wire u5__abc_78290_new_n725_; 
wire u5__abc_78290_new_n726_; 
wire u5__abc_78290_new_n727_; 
wire u5__abc_78290_new_n728_; 
wire u5__abc_78290_new_n729_; 
wire u5__abc_78290_new_n730_; 
wire u5__abc_78290_new_n731_; 
wire u5__abc_78290_new_n732_; 
wire u5__abc_78290_new_n733_; 
wire u5__abc_78290_new_n734_; 
wire u5__abc_78290_new_n735_; 
wire u5__abc_78290_new_n736_; 
wire u5__abc_78290_new_n737_; 
wire u5__abc_78290_new_n738_; 
wire u5__abc_78290_new_n739_; 
wire u5__abc_78290_new_n740_; 
wire u5__abc_78290_new_n741_; 
wire u5__abc_78290_new_n742_; 
wire u5__abc_78290_new_n743_; 
wire u5__abc_78290_new_n744_; 
wire u5__abc_78290_new_n745_; 
wire u5__abc_78290_new_n746_; 
wire u5__abc_78290_new_n747_; 
wire u5__abc_78290_new_n748_; 
wire u5__abc_78290_new_n749_; 
wire u5__abc_78290_new_n750_; 
wire u5__abc_78290_new_n751_; 
wire u5__abc_78290_new_n752_; 
wire u5__abc_78290_new_n753_; 
wire u5__abc_78290_new_n754_; 
wire u5__abc_78290_new_n755_; 
wire u5__abc_78290_new_n756_; 
wire u5__abc_78290_new_n757_; 
wire u5__abc_78290_new_n758_; 
wire u5__abc_78290_new_n759_; 
wire u5__abc_78290_new_n760_; 
wire u5__abc_78290_new_n761_; 
wire u5__abc_78290_new_n762_; 
wire u5__abc_78290_new_n763_; 
wire u5__abc_78290_new_n764_; 
wire u5__abc_78290_new_n765_; 
wire u5__abc_78290_new_n766_; 
wire u5__abc_78290_new_n767_; 
wire u5__abc_78290_new_n768_; 
wire u5__abc_78290_new_n769_; 
wire u5__abc_78290_new_n770_; 
wire u5__abc_78290_new_n771_; 
wire u5__abc_78290_new_n772_; 
wire u5__abc_78290_new_n773_; 
wire u5__abc_78290_new_n774_; 
wire u5__abc_78290_new_n775_; 
wire u5__abc_78290_new_n776_; 
wire u5__abc_78290_new_n777_; 
wire u5__abc_78290_new_n778_; 
wire u5__abc_78290_new_n779_; 
wire u5__abc_78290_new_n780_; 
wire u5__abc_78290_new_n781_; 
wire u5__abc_78290_new_n782_; 
wire u5__abc_78290_new_n783_; 
wire u5__abc_78290_new_n784_; 
wire u5__abc_78290_new_n785_; 
wire u5__abc_78290_new_n786_; 
wire u5__abc_78290_new_n787_; 
wire u5__abc_78290_new_n788_; 
wire u5__abc_78290_new_n789_; 
wire u5__abc_78290_new_n790_; 
wire u5__abc_78290_new_n791_; 
wire u5__abc_78290_new_n792_; 
wire u5__abc_78290_new_n793_; 
wire u5__abc_78290_new_n794_; 
wire u5__abc_78290_new_n795_; 
wire u5__abc_78290_new_n796_; 
wire u5__abc_78290_new_n797_; 
wire u5__abc_78290_new_n798_; 
wire u5__abc_78290_new_n799_; 
wire u5__abc_78290_new_n800_; 
wire u5__abc_78290_new_n801_; 
wire u5__abc_78290_new_n802_; 
wire u5__abc_78290_new_n803_; 
wire u5__abc_78290_new_n804_; 
wire u5__abc_78290_new_n805_; 
wire u5__abc_78290_new_n806_; 
wire u5__abc_78290_new_n807_; 
wire u5__abc_78290_new_n808_; 
wire u5__abc_78290_new_n809_; 
wire u5__abc_78290_new_n810_; 
wire u5__abc_78290_new_n811_; 
wire u5__abc_78290_new_n812_; 
wire u5__abc_78290_new_n813_; 
wire u5__abc_78290_new_n814_; 
wire u5__abc_78290_new_n815_; 
wire u5__abc_78290_new_n816_; 
wire u5__abc_78290_new_n817_; 
wire u5__abc_78290_new_n818_; 
wire u5__abc_78290_new_n819_; 
wire u5__abc_78290_new_n820_; 
wire u5__abc_78290_new_n821_; 
wire u5__abc_78290_new_n822_; 
wire u5__abc_78290_new_n823_; 
wire u5__abc_78290_new_n824_; 
wire u5__abc_78290_new_n825_; 
wire u5__abc_78290_new_n826_; 
wire u5__abc_78290_new_n827_; 
wire u5__abc_78290_new_n828_; 
wire u5__abc_78290_new_n829_; 
wire u5__abc_78290_new_n830_; 
wire u5__abc_78290_new_n831_; 
wire u5__abc_78290_new_n832_; 
wire u5__abc_78290_new_n833_; 
wire u5__abc_78290_new_n834_; 
wire u5__abc_78290_new_n835_; 
wire u5__abc_78290_new_n836_; 
wire u5__abc_78290_new_n837_; 
wire u5__abc_78290_new_n838_; 
wire u5__abc_78290_new_n839_; 
wire u5__abc_78290_new_n840_; 
wire u5__abc_78290_new_n841_; 
wire u5__abc_78290_new_n842_; 
wire u5__abc_78290_new_n843_; 
wire u5__abc_78290_new_n844_; 
wire u5__abc_78290_new_n845_; 
wire u5__abc_78290_new_n846_; 
wire u5__abc_78290_new_n847_; 
wire u5__abc_78290_new_n848_; 
wire u5__abc_78290_new_n849_; 
wire u5__abc_78290_new_n850_; 
wire u5__abc_78290_new_n851_; 
wire u5__abc_78290_new_n852_; 
wire u5__abc_78290_new_n853_; 
wire u5__abc_78290_new_n854_; 
wire u5__abc_78290_new_n855_; 
wire u5__abc_78290_new_n856_; 
wire u5__abc_78290_new_n857_; 
wire u5__abc_78290_new_n858_; 
wire u5__abc_78290_new_n859_; 
wire u5__abc_78290_new_n860_; 
wire u5__abc_78290_new_n861_; 
wire u5__abc_78290_new_n862_; 
wire u5__abc_78290_new_n863_; 
wire u5__abc_78290_new_n864_; 
wire u5__abc_78290_new_n865_; 
wire u5__abc_78290_new_n866_; 
wire u5__abc_78290_new_n867_; 
wire u5__abc_78290_new_n868_; 
wire u5__abc_78290_new_n869_; 
wire u5__abc_78290_new_n870_; 
wire u5__abc_78290_new_n871_; 
wire u5__abc_78290_new_n872_; 
wire u5__abc_78290_new_n873_; 
wire u5__abc_78290_new_n874_; 
wire u5__abc_78290_new_n875_; 
wire u5__abc_78290_new_n876_; 
wire u5__abc_78290_new_n877_; 
wire u5__abc_78290_new_n878_; 
wire u5__abc_78290_new_n879_; 
wire u5__abc_78290_new_n880_; 
wire u5__abc_78290_new_n881_; 
wire u5__abc_78290_new_n882_; 
wire u5__abc_78290_new_n883_; 
wire u5__abc_78290_new_n884_; 
wire u5__abc_78290_new_n885_; 
wire u5__abc_78290_new_n886_; 
wire u5__abc_78290_new_n887_; 
wire u5__abc_78290_new_n888_; 
wire u5__abc_78290_new_n889_; 
wire u5__abc_78290_new_n890_; 
wire u5__abc_78290_new_n891_; 
wire u5__abc_78290_new_n892_; 
wire u5__abc_78290_new_n893_; 
wire u5__abc_78290_new_n894_; 
wire u5__abc_78290_new_n895_; 
wire u5__abc_78290_new_n896_; 
wire u5__abc_78290_new_n897_; 
wire u5__abc_78290_new_n898_; 
wire u5__abc_78290_new_n899_; 
wire u5__abc_78290_new_n900_; 
wire u5__abc_78290_new_n901_; 
wire u5__abc_78290_new_n902_; 
wire u5__abc_78290_new_n903_; 
wire u5__abc_78290_new_n904_; 
wire u5__abc_78290_new_n905_; 
wire u5__abc_78290_new_n906_; 
wire u5__abc_78290_new_n907_; 
wire u5__abc_78290_new_n908_; 
wire u5__abc_78290_new_n909_; 
wire u5__abc_78290_new_n910_; 
wire u5__abc_78290_new_n911_; 
wire u5__abc_78290_new_n912_; 
wire u5__abc_78290_new_n913_; 
wire u5__abc_78290_new_n914_; 
wire u5__abc_78290_new_n915_; 
wire u5__abc_78290_new_n916_; 
wire u5__abc_78290_new_n917_; 
wire u5__abc_78290_new_n918_; 
wire u5__abc_78290_new_n919_; 
wire u5__abc_78290_new_n920_; 
wire u5__abc_78290_new_n921_; 
wire u5__abc_78290_new_n922_; 
wire u5__abc_78290_new_n923_; 
wire u5__abc_78290_new_n924_; 
wire u5__abc_78290_new_n925_; 
wire u5__abc_78290_new_n926_; 
wire u5__abc_78290_new_n927_; 
wire u5__abc_78290_new_n928_; 
wire u5__abc_78290_new_n929_; 
wire u5__abc_78290_new_n930_; 
wire u5__abc_78290_new_n931_; 
wire u5__abc_78290_new_n932_; 
wire u5__abc_78290_new_n933_; 
wire u5__abc_78290_new_n934_; 
wire u5__abc_78290_new_n935_; 
wire u5__abc_78290_new_n936_; 
wire u5__abc_78290_new_n937_; 
wire u5__abc_78290_new_n938_; 
wire u5__abc_78290_new_n939_; 
wire u5__abc_78290_new_n940_; 
wire u5__abc_78290_new_n941_; 
wire u5__abc_78290_new_n942_; 
wire u5__abc_78290_new_n943_; 
wire u5__abc_78290_new_n944_; 
wire u5__abc_78290_new_n945_; 
wire u5__abc_78290_new_n946_; 
wire u5__abc_78290_new_n947_; 
wire u5__abc_78290_new_n948_; 
wire u5__abc_78290_new_n949_; 
wire u5__abc_78290_new_n950_; 
wire u5__abc_78290_new_n951_; 
wire u5__abc_78290_new_n952_; 
wire u5__abc_78290_new_n953_; 
wire u5__abc_78290_new_n954_; 
wire u5__abc_78290_new_n955_; 
wire u5__abc_78290_new_n956_; 
wire u5__abc_78290_new_n957_; 
wire u5__abc_78290_new_n958_; 
wire u5__abc_78290_new_n961_; 
wire u5__abc_78290_new_n962_; 
wire u5__abc_78290_new_n963_; 
wire u5__abc_78290_new_n964_; 
wire u5__abc_78290_new_n965_; 
wire u5__abc_78290_new_n966_; 
wire u5__abc_78290_new_n967_; 
wire u5__abc_78290_new_n969_; 
wire u5__abc_78290_new_n970_; 
wire u5__abc_78290_new_n971_; 
wire u5__abc_78290_new_n974_; 
wire u5__abc_78290_new_n975_; 
wire u5__abc_78290_new_n976_; 
wire u5__abc_78290_new_n977_; 
wire u5__abc_78290_new_n978_; 
wire u5__abc_78290_new_n979_; 
wire u5__abc_78290_new_n980_; 
wire u5__abc_78290_new_n981_; 
wire u5__abc_78290_new_n982_; 
wire u5__abc_78290_new_n983_; 
wire u5__abc_78290_new_n984_; 
wire u5__abc_78290_new_n985_; 
wire u5__abc_78290_new_n986_; 
wire u5__abc_78290_new_n987_; 
wire u5__abc_78290_new_n988_; 
wire u5__abc_78290_new_n989_; 
wire u5__abc_78290_new_n990_; 
wire u5__abc_78290_new_n991_; 
wire u5__abc_78290_new_n992_; 
wire u5__abc_78290_new_n993_; 
wire u5__abc_78290_new_n994_; 
wire u5__abc_78290_new_n995_; 
wire u5__abc_78290_new_n996_; 
wire u5__abc_78290_new_n997_; 
wire u5__abc_78290_new_n998_; 
wire u5__abc_78290_new_n999_; 
wire u5_ack_cnt_0_; 
wire u5_ack_cnt_1_; 
wire u5_ack_cnt_2_; 
wire u5_ack_cnt_3_; 
wire u5_ap_en; 
wire u5_burst_act_rd; 
wire u5_burst_cnt_0_; 
wire u5_burst_cnt_10_; 
wire u5_burst_cnt_1_; 
wire u5_burst_cnt_2_; 
wire u5_burst_cnt_3_; 
wire u5_burst_cnt_4_; 
wire u5_burst_cnt_5_; 
wire u5_burst_cnt_6_; 
wire u5_burst_cnt_7_; 
wire u5_burst_cnt_8_; 
wire u5_burst_cnt_9_; 
wire u5_cke_d; 
wire u5_cke_o_del; 
wire u5_cke_o_r1; 
wire u5_cke_o_r2; 
wire u5_cke_r; 
wire u5_cmd_0_; 
wire u5_cmd_1_; 
wire u5_cmd_2_; 
wire u5_cmd_3_; 
wire u5_cmd_a10_r; 
wire u5_cmd_asserted; 
wire u5_cmd_asserted2; 
wire u5_cmd_del_0_; 
wire u5_cmd_del_1_; 
wire u5_cmd_del_2_; 
wire u5_cmd_del_3_; 
wire u5_cmd_r_0_; 
wire u5_cmd_r_1_; 
wire u5_cmd_r_2_; 
wire u5_cmd_r_3_; 
wire u5_cnt; 
wire u5_cnt_next; 
wire u5_cs_le_r; 
wire u5_cs_le_r1; 
wire u5_data_oe_d; 
wire u5_data_oe_r; 
wire u5_data_oe_r2; 
wire u5_dv_r; 
wire u5_ir_cnt_0_; 
wire u5_ir_cnt_1_; 
wire u5_ir_cnt_2_; 
wire u5_ir_cnt_3_; 
wire u5_ir_cnt_done; 
wire u5_kro; 
wire u5_lmr_ack_d; 
wire u5_lookup_ready1; 
wire u5_lookup_ready2; 
wire u5_mc_adv_r; 
wire u5_mc_adv_r1; 
wire u5_mc_c_oe_d; 
wire u5_mc_le; 
wire u5_mem_ack_r; 
wire u5_next_state_0_; 
wire u5_next_state_10_; 
wire u5_next_state_11_; 
wire u5_next_state_12_; 
wire u5_next_state_13_; 
wire u5_next_state_14_; 
wire u5_next_state_15_; 
wire u5_next_state_16_; 
wire u5_next_state_17_; 
wire u5_next_state_18_; 
wire u5_next_state_19_; 
wire u5_next_state_1_; 
wire u5_next_state_20_; 
wire u5_next_state_21_; 
wire u5_next_state_22_; 
wire u5_next_state_23_; 
wire u5_next_state_24_; 
wire u5_next_state_25_; 
wire u5_next_state_26_; 
wire u5_next_state_27_; 
wire u5_next_state_28_; 
wire u5_next_state_29_; 
wire u5_next_state_2_; 
wire u5_next_state_30_; 
wire u5_next_state_31_; 
wire u5_next_state_32_; 
wire u5_next_state_33_; 
wire u5_next_state_34_; 
wire u5_next_state_35_; 
wire u5_next_state_36_; 
wire u5_next_state_37_; 
wire u5_next_state_38_; 
wire u5_next_state_39_; 
wire u5_next_state_3_; 
wire u5_next_state_40_; 
wire u5_next_state_41_; 
wire u5_next_state_42_; 
wire u5_next_state_43_; 
wire u5_next_state_44_; 
wire u5_next_state_45_; 
wire u5_next_state_46_; 
wire u5_next_state_47_; 
wire u5_next_state_48_; 
wire u5_next_state_49_; 
wire u5_next_state_4_; 
wire u5_next_state_50_; 
wire u5_next_state_51_; 
wire u5_next_state_52_; 
wire u5_next_state_53_; 
wire u5_next_state_54_; 
wire u5_next_state_55_; 
wire u5_next_state_56_; 
wire u5_next_state_57_; 
wire u5_next_state_58_; 
wire u5_next_state_59_; 
wire u5_next_state_5_; 
wire u5_next_state_60_; 
wire u5_next_state_61_; 
wire u5_next_state_62_; 
wire u5_next_state_63_; 
wire u5_next_state_64_; 
wire u5_next_state_65_; 
wire u5_next_state_6_; 
wire u5_next_state_7_; 
wire u5_next_state_8_; 
wire u5_next_state_9_; 
wire u5_no_wb_cycle; 
wire u5_pack_le0_d; 
wire u5_pack_le1_d; 
wire u5_pack_le2_d; 
wire u5_resume_req_r; 
wire u5_rfr_ack_d; 
wire u5_rsts; 
wire u5_state_0_; 
wire u5_state_10_; 
wire u5_state_11_; 
wire u5_state_12_; 
wire u5_state_13_; 
wire u5_state_14_; 
wire u5_state_15_; 
wire u5_state_16_; 
wire u5_state_17_; 
wire u5_state_18_; 
wire u5_state_19_; 
wire u5_state_1_; 
wire u5_state_20_; 
wire u5_state_21_; 
wire u5_state_22_; 
wire u5_state_23_; 
wire u5_state_24_; 
wire u5_state_25_; 
wire u5_state_26_; 
wire u5_state_27_; 
wire u5_state_28_; 
wire u5_state_29_; 
wire u5_state_2_; 
wire u5_state_30_; 
wire u5_state_31_; 
wire u5_state_32_; 
wire u5_state_33_; 
wire u5_state_34_; 
wire u5_state_35_; 
wire u5_state_36_; 
wire u5_state_37_; 
wire u5_state_38_; 
wire u5_state_39_; 
wire u5_state_3_; 
wire u5_state_40_; 
wire u5_state_41_; 
wire u5_state_42_; 
wire u5_state_43_; 
wire u5_state_44_; 
wire u5_state_45_; 
wire u5_state_46_; 
wire u5_state_47_; 
wire u5_state_48_; 
wire u5_state_49_; 
wire u5_state_4_; 
wire u5_state_50_; 
wire u5_state_51_; 
wire u5_state_52_; 
wire u5_state_53_; 
wire u5_state_54_; 
wire u5_state_55_; 
wire u5_state_56_; 
wire u5_state_57_; 
wire u5_state_58_; 
wire u5_state_59_; 
wire u5_state_5_; 
wire u5_state_60_; 
wire u5_state_61_; 
wire u5_state_62_; 
wire u5_state_63_; 
wire u5_state_64_; 
wire u5_state_65_; 
wire u5_state_6_; 
wire u5_state_7_; 
wire u5_state_8_; 
wire u5_state_9_; 
wire u5_susp_req_r; 
wire u5_suspended_d; 
wire u5_timer2_0_; 
wire u5_timer2_1_; 
wire u5_timer2_2_; 
wire u5_timer2_3_; 
wire u5_timer2_4_; 
wire u5_timer2_5_; 
wire u5_timer2_6_; 
wire u5_timer2_7_; 
wire u5_timer2_8_; 
wire u5_timer_0_; 
wire u5_timer_1_; 
wire u5_timer_2_; 
wire u5_timer_3_; 
wire u5_timer_4_; 
wire u5_timer_5_; 
wire u5_timer_6_; 
wire u5_timer_7_; 
wire u5_timer_is_zero; 
wire u5_tmr2_done; 
wire u5_tmr_done; 
wire u5_wb_cycle; 
wire u5_wb_first; 
wire u5_wb_stb_first; 
wire u5_wb_wait; 
wire u5_wb_wait_r; 
wire u5_wb_wait_r2; 
wire u5_wb_write_go_r; 
wire u5_we_; 
wire u6__0read_go_r1_0_0_; 
wire u6__0read_go_r_0_0_; 
wire u6__0rmw_en_0_0_; 
wire u6__0rmw_r_0_0_; 
wire u6__0wb_ack_o_0_0_; 
wire u6__0wb_data_o_31_0__0_; 
wire u6__0wb_data_o_31_0__10_; 
wire u6__0wb_data_o_31_0__11_; 
wire u6__0wb_data_o_31_0__12_; 
wire u6__0wb_data_o_31_0__13_; 
wire u6__0wb_data_o_31_0__14_; 
wire u6__0wb_data_o_31_0__15_; 
wire u6__0wb_data_o_31_0__16_; 
wire u6__0wb_data_o_31_0__17_; 
wire u6__0wb_data_o_31_0__18_; 
wire u6__0wb_data_o_31_0__19_; 
wire u6__0wb_data_o_31_0__1_; 
wire u6__0wb_data_o_31_0__20_; 
wire u6__0wb_data_o_31_0__21_; 
wire u6__0wb_data_o_31_0__22_; 
wire u6__0wb_data_o_31_0__23_; 
wire u6__0wb_data_o_31_0__24_; 
wire u6__0wb_data_o_31_0__25_; 
wire u6__0wb_data_o_31_0__26_; 
wire u6__0wb_data_o_31_0__27_; 
wire u6__0wb_data_o_31_0__28_; 
wire u6__0wb_data_o_31_0__29_; 
wire u6__0wb_data_o_31_0__2_; 
wire u6__0wb_data_o_31_0__30_; 
wire u6__0wb_data_o_31_0__31_; 
wire u6__0wb_data_o_31_0__3_; 
wire u6__0wb_data_o_31_0__4_; 
wire u6__0wb_data_o_31_0__5_; 
wire u6__0wb_data_o_31_0__6_; 
wire u6__0wb_data_o_31_0__7_; 
wire u6__0wb_data_o_31_0__8_; 
wire u6__0wb_data_o_31_0__9_; 
wire u6__0wb_err_0_0_; 
wire u6__0wb_first_r_0_0_; 
wire u6__0wr_hold_0_0_; 
wire u6__0write_go_r1_0_0_; 
wire u6__0write_go_r_0_0_; 
wire u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188; 
wire u6__abc_81318_new_n133_; 
wire u6__abc_81318_new_n134_; 
wire u6__abc_81318_new_n135_; 
wire u6__abc_81318_new_n136_; 
wire u6__abc_81318_new_n137_; 
wire u6__abc_81318_new_n138_; 
wire u6__abc_81318_new_n139_; 
wire u6__abc_81318_new_n140_; 
wire u6__abc_81318_new_n141_; 
wire u6__abc_81318_new_n142_; 
wire u6__abc_81318_new_n143_; 
wire u6__abc_81318_new_n144_; 
wire u6__abc_81318_new_n146_; 
wire u6__abc_81318_new_n147_; 
wire u6__abc_81318_new_n149_; 
wire u6__abc_81318_new_n150_; 
wire u6__abc_81318_new_n152_; 
wire u6__abc_81318_new_n153_; 
wire u6__abc_81318_new_n155_; 
wire u6__abc_81318_new_n156_; 
wire u6__abc_81318_new_n158_; 
wire u6__abc_81318_new_n159_; 
wire u6__abc_81318_new_n161_; 
wire u6__abc_81318_new_n162_; 
wire u6__abc_81318_new_n164_; 
wire u6__abc_81318_new_n165_; 
wire u6__abc_81318_new_n167_; 
wire u6__abc_81318_new_n168_; 
wire u6__abc_81318_new_n170_; 
wire u6__abc_81318_new_n171_; 
wire u6__abc_81318_new_n173_; 
wire u6__abc_81318_new_n174_; 
wire u6__abc_81318_new_n176_; 
wire u6__abc_81318_new_n177_; 
wire u6__abc_81318_new_n179_; 
wire u6__abc_81318_new_n180_; 
wire u6__abc_81318_new_n182_; 
wire u6__abc_81318_new_n183_; 
wire u6__abc_81318_new_n185_; 
wire u6__abc_81318_new_n186_; 
wire u6__abc_81318_new_n188_; 
wire u6__abc_81318_new_n189_; 
wire u6__abc_81318_new_n191_; 
wire u6__abc_81318_new_n192_; 
wire u6__abc_81318_new_n194_; 
wire u6__abc_81318_new_n195_; 
wire u6__abc_81318_new_n197_; 
wire u6__abc_81318_new_n198_; 
wire u6__abc_81318_new_n200_; 
wire u6__abc_81318_new_n201_; 
wire u6__abc_81318_new_n203_; 
wire u6__abc_81318_new_n204_; 
wire u6__abc_81318_new_n206_; 
wire u6__abc_81318_new_n207_; 
wire u6__abc_81318_new_n209_; 
wire u6__abc_81318_new_n210_; 
wire u6__abc_81318_new_n212_; 
wire u6__abc_81318_new_n213_; 
wire u6__abc_81318_new_n215_; 
wire u6__abc_81318_new_n216_; 
wire u6__abc_81318_new_n218_; 
wire u6__abc_81318_new_n219_; 
wire u6__abc_81318_new_n221_; 
wire u6__abc_81318_new_n222_; 
wire u6__abc_81318_new_n224_; 
wire u6__abc_81318_new_n225_; 
wire u6__abc_81318_new_n227_; 
wire u6__abc_81318_new_n228_; 
wire u6__abc_81318_new_n230_; 
wire u6__abc_81318_new_n231_; 
wire u6__abc_81318_new_n233_; 
wire u6__abc_81318_new_n234_; 
wire u6__abc_81318_new_n236_; 
wire u6__abc_81318_new_n237_; 
wire u6__abc_81318_new_n239_; 
wire u6__abc_81318_new_n240_; 
wire u6__abc_81318_new_n242_; 
wire u6__abc_81318_new_n243_; 
wire u6__abc_81318_new_n245_; 
wire u6__abc_81318_new_n247_; 
wire u6__abc_81318_new_n248_; 
wire u6__abc_81318_new_n249_; 
wire u6__abc_81318_new_n250_; 
wire u6__abc_81318_new_n251_; 
wire u6__abc_81318_new_n252_; 
wire u6__abc_81318_new_n253_; 
wire u6__abc_81318_new_n254_; 
wire u6__abc_81318_new_n255_; 
wire u6__abc_81318_new_n256_; 
wire u6__abc_81318_new_n258_; 
wire u6__abc_81318_new_n260_; 
wire u6__abc_81318_new_n262_; 
wire u6__abc_81318_new_n263_; 
wire u6__abc_81318_new_n265_; 
wire u6__abc_81318_new_n267_; 
wire u6__abc_81318_new_n269_; 
wire u6__abc_81318_new_n270_; 
wire u6__abc_81318_new_n271_; 
wire u6__abc_81318_new_n273_; 
wire u6__abc_81318_new_n275_; 
wire u6_read_go_r; 
wire u6_read_go_r1; 
wire u6_rmw_en; 
wire u6_rmw_r; 
wire u6_wb_first_r; 
wire u6_write_go_r; 
wire u6_write_go_r1; 
wire u7__0mc_adsc__0_0_; 
wire u7__0mc_adv__0_0_; 
wire u7__0mc_cs__0_0_; 
wire u7__0mc_cs__1_1_; 
wire u7__0mc_cs__2_2_; 
wire u7__0mc_cs__3_3_; 
wire u7__0mc_cs__4_4_; 
wire u7__0mc_cs__5_5_; 
wire u7__0mc_cs__6_6_; 
wire u7__0mc_cs__7_7_; 
wire u7__0mc_data_oe_0_0_; 
wire u7__0mc_dqm_3_0__0_; 
wire u7__0mc_dqm_3_0__1_; 
wire u7__0mc_dqm_3_0__2_; 
wire u7__0mc_dqm_3_0__3_; 
wire u7__0mc_dqm_r_3_0__0_; 
wire u7__0mc_dqm_r_3_0__1_; 
wire u7__0mc_dqm_r_3_0__2_; 
wire u7__0mc_dqm_r_3_0__3_; 
wire u7__0mc_oe__0_0_; 
wire u7__0mc_rp_0_0_; 
wire u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518; 
wire u7__abc_73829_new_n100_; 
wire u7__abc_73829_new_n101_; 
wire u7__abc_73829_new_n102_; 
wire u7__abc_73829_new_n103_; 
wire u7__abc_73829_new_n104_; 
wire u7__abc_73829_new_n105_; 
wire u7__abc_73829_new_n106_; 
wire u7__abc_73829_new_n107_; 
wire u7__abc_73829_new_n108_; 
wire u7__abc_73829_new_n110_; 
wire u7__abc_73829_new_n111_; 
wire u7__abc_73829_new_n112_; 
wire u7__abc_73829_new_n113_; 
wire u7__abc_73829_new_n114_; 
wire u7__abc_73829_new_n116_; 
wire u7__abc_73829_new_n117_; 
wire u7__abc_73829_new_n118_; 
wire u7__abc_73829_new_n119_; 
wire u7__abc_73829_new_n120_; 
wire u7__abc_73829_new_n122_; 
wire u7__abc_73829_new_n123_; 
wire u7__abc_73829_new_n124_; 
wire u7__abc_73829_new_n125_; 
wire u7__abc_73829_new_n126_; 
wire u7__abc_73829_new_n128_; 
wire u7__abc_73829_new_n129_; 
wire u7__abc_73829_new_n130_; 
wire u7__abc_73829_new_n131_; 
wire u7__abc_73829_new_n132_; 
wire u7__abc_73829_new_n134_; 
wire u7__abc_73829_new_n135_; 
wire u7__abc_73829_new_n136_; 
wire u7__abc_73829_new_n137_; 
wire u7__abc_73829_new_n138_; 
wire u7__abc_73829_new_n140_; 
wire u7__abc_73829_new_n141_; 
wire u7__abc_73829_new_n142_; 
wire u7__abc_73829_new_n143_; 
wire u7__abc_73829_new_n144_; 
wire u7__abc_73829_new_n146_; 
wire u7__abc_73829_new_n147_; 
wire u7__abc_73829_new_n148_; 
wire u7__abc_73829_new_n149_; 
wire u7__abc_73829_new_n150_; 
wire u7__abc_73829_new_n155_; 
wire u7__abc_73829_new_n75_; 
wire u7__abc_73829_new_n76_; 
wire u7__abc_73829_new_n77_; 
wire u7__abc_73829_new_n78_; 
wire u7__abc_73829_new_n79_; 
wire u7__abc_73829_new_n81_; 
wire u7__abc_73829_new_n83_; 
wire u7__abc_73829_new_n85_; 
wire u7__abc_73829_new_n87_; 
wire u7__abc_73829_new_n88_; 
wire u7__abc_73829_new_n89_; 
wire u7__abc_73829_new_n91_; 
wire u7__abc_73829_new_n92_; 
wire u7__abc_73829_new_n94_; 
wire u7__abc_73829_new_n95_; 
wire u7__abc_73829_new_n97_; 
wire u7__abc_73829_new_n98_; 
wire u7_mc_dqm_r2_0_; 
wire u7_mc_dqm_r2_1_; 
wire u7_mc_dqm_r2_2_; 
wire u7_mc_dqm_r2_3_; 
wire u7_mc_dqm_r_0_; 
wire u7_mc_dqm_r_1_; 
wire u7_mc_dqm_r_2_; 
wire u7_mc_dqm_r_3_; 
output wb_ack_o;
input \wb_addr_i[0] ;
input \wb_addr_i[10] ;
input \wb_addr_i[11] ;
input \wb_addr_i[12] ;
input \wb_addr_i[13] ;
input \wb_addr_i[14] ;
input \wb_addr_i[15] ;
input \wb_addr_i[16] ;
input \wb_addr_i[17] ;
input \wb_addr_i[18] ;
input \wb_addr_i[19] ;
input \wb_addr_i[1] ;
input \wb_addr_i[20] ;
input \wb_addr_i[21] ;
input \wb_addr_i[22] ;
input \wb_addr_i[23] ;
input \wb_addr_i[24] ;
input \wb_addr_i[25] ;
input \wb_addr_i[26] ;
input \wb_addr_i[27] ;
input \wb_addr_i[28] ;
input \wb_addr_i[29] ;
input \wb_addr_i[2] ;
input \wb_addr_i[30] ;
input \wb_addr_i[31] ;
input \wb_addr_i[3] ;
input \wb_addr_i[4] ;
input \wb_addr_i[5] ;
input \wb_addr_i[6] ;
input \wb_addr_i[7] ;
input \wb_addr_i[8] ;
input \wb_addr_i[9] ;
input wb_cyc_i;
input \wb_data_i[0] ;
input \wb_data_i[10] ;
input \wb_data_i[11] ;
input \wb_data_i[12] ;
input \wb_data_i[13] ;
input \wb_data_i[14] ;
input \wb_data_i[15] ;
input \wb_data_i[16] ;
input \wb_data_i[17] ;
input \wb_data_i[18] ;
input \wb_data_i[19] ;
input \wb_data_i[1] ;
input \wb_data_i[20] ;
input \wb_data_i[21] ;
input \wb_data_i[22] ;
input \wb_data_i[23] ;
input \wb_data_i[24] ;
input \wb_data_i[25] ;
input \wb_data_i[26] ;
input \wb_data_i[27] ;
input \wb_data_i[28] ;
input \wb_data_i[29] ;
input \wb_data_i[2] ;
input \wb_data_i[30] ;
input \wb_data_i[31] ;
input \wb_data_i[3] ;
input \wb_data_i[4] ;
input \wb_data_i[5] ;
input \wb_data_i[6] ;
input \wb_data_i[7] ;
input \wb_data_i[8] ;
input \wb_data_i[9] ;
output \wb_data_o[0] ;
output \wb_data_o[10] ;
output \wb_data_o[11] ;
output \wb_data_o[12] ;
output \wb_data_o[13] ;
output \wb_data_o[14] ;
output \wb_data_o[15] ;
output \wb_data_o[16] ;
output \wb_data_o[17] ;
output \wb_data_o[18] ;
output \wb_data_o[19] ;
output \wb_data_o[1] ;
output \wb_data_o[20] ;
output \wb_data_o[21] ;
output \wb_data_o[22] ;
output \wb_data_o[23] ;
output \wb_data_o[24] ;
output \wb_data_o[25] ;
output \wb_data_o[26] ;
output \wb_data_o[27] ;
output \wb_data_o[28] ;
output \wb_data_o[29] ;
output \wb_data_o[2] ;
output \wb_data_o[30] ;
output \wb_data_o[31] ;
output \wb_data_o[3] ;
output \wb_data_o[4] ;
output \wb_data_o[5] ;
output \wb_data_o[6] ;
output \wb_data_o[7] ;
output \wb_data_o[8] ;
output \wb_data_o[9] ;
output wb_err_o;
input \wb_sel_i[0] ;
input \wb_sel_i[1] ;
input \wb_sel_i[2] ;
input \wb_sel_i[3] ;
input wb_stb_i;
input wb_we_i;
AND2X2 AND2X2_1 ( .A(wb_stb_i), .B(wb_cyc_i), .Y(u0__abc_74894_new_n1154_));
AND2X2 AND2X2_10 ( .A(u0__abc_74894_new_n3728_), .B(u0__abc_74894_new_n3769_), .Y(u0__abc_74894_new_n3770_));
AND2X2 AND2X2_100 ( .A(u5__abc_78290_new_n393_), .B(u5__abc_78290_new_n394_), .Y(u5__abc_78290_new_n395_));
AND2X2 AND2X2_101 ( .A(u5__abc_78290_new_n396_), .B(u5__abc_78290_new_n397_), .Y(u5__abc_78290_new_n398_));
AND2X2 AND2X2_102 ( .A(u5__abc_78290_new_n400_), .B(u5__abc_78290_new_n401_), .Y(u5__abc_78290_new_n402_));
AND2X2 AND2X2_103 ( .A(u5__abc_78290_new_n403_), .B(u5__abc_78290_new_n404_), .Y(u5__abc_78290_new_n405_));
AND2X2 AND2X2_104 ( .A(u5__abc_78290_new_n409_), .B(u5__abc_78290_new_n410_), .Y(u5__abc_78290_new_n411_));
AND2X2 AND2X2_105 ( .A(u5__abc_78290_new_n412_), .B(u5__abc_78290_new_n413_), .Y(u5__abc_78290_new_n414_));
AND2X2 AND2X2_106 ( .A(u5__abc_78290_new_n416_), .B(u5__abc_78290_new_n417_), .Y(u5__abc_78290_new_n418_));
AND2X2 AND2X2_107 ( .A(u5__abc_78290_new_n419_), .B(u5__abc_78290_new_n420_), .Y(u5__abc_78290_new_n421_));
AND2X2 AND2X2_108 ( .A(u5__abc_78290_new_n434_), .B(u5__abc_78290_new_n435_), .Y(u5__abc_78290_new_n473_));
AND2X2 AND2X2_109 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n479_), .Y(u5__abc_78290_new_n480_));
AND2X2 AND2X2_11 ( .A(u0__abc_74894_new_n3881_), .B(u0__abc_74894_new_n3882_), .Y(u0__abc_74894_new_n3883_));
AND2X2 AND2X2_110 ( .A(u5__abc_78290_new_n493_), .B(u5__abc_78290_new_n413_), .Y(u5__abc_78290_new_n494_));
AND2X2 AND2X2_111 ( .A(u5__abc_78290_new_n438_), .B(u5__abc_78290_new_n451_), .Y(u5__abc_78290_new_n499_));
AND2X2 AND2X2_112 ( .A(u5__abc_78290_new_n517_), .B(u5__abc_78290_new_n514_), .Y(u5__abc_78290_new_n518_));
AND2X2 AND2X2_113 ( .A(u5__abc_78290_new_n431_), .B(u5__abc_78290_new_n545_), .Y(u5__abc_78290_new_n546_));
AND2X2 AND2X2_114 ( .A(u5__abc_78290_new_n553_), .B(u5__abc_78290_new_n547_), .Y(u5__abc_78290_new_n554_));
AND2X2 AND2X2_115 ( .A(u5__abc_78290_new_n427_), .B(u5__abc_78290_new_n429_), .Y(u5__abc_78290_new_n562_));
AND2X2 AND2X2_116 ( .A(u5__abc_78290_new_n424_), .B(u5__abc_78290_new_n425_), .Y(u5__abc_78290_new_n588_));
AND2X2 AND2X2_117 ( .A(u5__abc_78290_new_n427_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n589_));
AND2X2 AND2X2_118 ( .A(u5__abc_78290_new_n580_), .B(u5__abc_78290_new_n609_), .Y(u5__abc_78290_new_n610_));
AND2X2 AND2X2_119 ( .A(u5__abc_78290_new_n416_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n626_));
AND2X2 AND2X2_12 ( .A(u0__abc_74894_new_n4004_), .B(u0__abc_74894_new_n4007_), .Y(u0__abc_74894_new_n4008_));
AND2X2 AND2X2_120 ( .A(u5__abc_78290_new_n428_), .B(u5_state_8_), .Y(u5__abc_78290_new_n725_));
AND2X2 AND2X2_121 ( .A(u5__abc_78290_new_n412_), .B(u5__abc_78290_new_n726_), .Y(u5__abc_78290_new_n727_));
AND2X2 AND2X2_122 ( .A(u5__abc_78290_new_n736_), .B(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n737_));
AND2X2 AND2X2_123 ( .A(u5__abc_78290_new_n428_), .B(u5_state_9_), .Y(u5__abc_78290_new_n740_));
AND2X2 AND2X2_124 ( .A(u5__abc_78290_new_n412_), .B(u5__abc_78290_new_n741_), .Y(u5__abc_78290_new_n742_));
AND2X2 AND2X2_125 ( .A(u5__abc_78290_new_n447_), .B(u5__abc_78290_new_n409_), .Y(u5__abc_78290_new_n750_));
AND2X2 AND2X2_126 ( .A(u5__abc_78290_new_n826_), .B(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n827_));
AND2X2 AND2X2_127 ( .A(u5__abc_78290_new_n832_), .B(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n833_));
AND2X2 AND2X2_128 ( .A(u5__abc_78290_new_n810_), .B(u5__abc_78290_new_n836_), .Y(u5__abc_78290_new_n837_));
AND2X2 AND2X2_129 ( .A(u5__abc_78290_new_n884_), .B(u5__abc_78290_new_n845_), .Y(u5__abc_78290_new_n885_));
AND2X2 AND2X2_13 ( .A(u0__abc_74894_new_n4026_), .B(u0__abc_74894_new_n4029_), .Y(u0__abc_74894_new_n4030_));
AND2X2 AND2X2_130 ( .A(u5__abc_78290_new_n428_), .B(u5_state_11_), .Y(u5__abc_78290_new_n889_));
AND2X2 AND2X2_131 ( .A(u5__abc_78290_new_n413_), .B(u5__abc_78290_new_n757_), .Y(u5__abc_78290_new_n890_));
AND2X2 AND2X2_132 ( .A(u5__abc_78290_new_n772_), .B(u5__abc_78290_new_n416_), .Y(u5__abc_78290_new_n1020_));
AND2X2 AND2X2_133 ( .A(u5__abc_78290_new_n628_), .B(u5__abc_78290_new_n416_), .Y(u5__abc_78290_new_n1024_));
AND2X2 AND2X2_134 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n1079_), .Y(u5__abc_78290_new_n1085_));
AND2X2 AND2X2_135 ( .A(u5__abc_78290_new_n1102_), .B(u5__abc_78290_new_n1096_), .Y(u5__abc_78290_new_n1103_));
AND2X2 AND2X2_136 ( .A(u5__abc_78290_new_n1166_), .B(u5__abc_78290_new_n1157_), .Y(u5__abc_78290_new_n1167_));
AND2X2 AND2X2_137 ( .A(u5__abc_78290_new_n1194_), .B(u5__abc_78290_new_n499_), .Y(u5__abc_78290_new_n1195_));
AND2X2 AND2X2_138 ( .A(u5__abc_78290_new_n1204_), .B(u5__abc_78290_new_n1207_), .Y(u5__abc_78290_new_n1208_));
AND2X2 AND2X2_139 ( .A(u5__abc_78290_new_n1201_), .B(u5__abc_78290_new_n1208_), .Y(u5__abc_78290_new_n1209_));
AND2X2 AND2X2_14 ( .A(u0__abc_74894_new_n4045_), .B(u0__abc_74894_new_n4041_), .Y(u0__abc_74894_new_n4046_));
AND2X2 AND2X2_140 ( .A(u5__abc_78290_new_n1239_), .B(u5__abc_78290_new_n484_), .Y(u5__abc_78290_new_n1240_));
AND2X2 AND2X2_141 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n566_), .Y(u5__abc_78290_new_n1304_));
AND2X2 AND2X2_142 ( .A(u5__abc_78290_new_n480_), .B(u5__abc_78290_new_n1304_), .Y(u5__abc_78290_new_n1305_));
AND2X2 AND2X2_143 ( .A(u5__abc_78290_new_n1327_), .B(u5__abc_78290_new_n1328_), .Y(u5__abc_78290_new_n1329_));
AND2X2 AND2X2_144 ( .A(u5__abc_78290_new_n1240_), .B(u5__abc_78290_new_n1062_), .Y(u5__abc_78290_new_n1367_));
AND2X2 AND2X2_145 ( .A(u5__abc_78290_new_n1373_), .B(u5__abc_78290_new_n1378_), .Y(u5__abc_78290_new_n1379_));
AND2X2 AND2X2_146 ( .A(u5__abc_78290_new_n1440_), .B(u5__abc_78290_new_n1444_), .Y(u5__abc_78290_new_n1445_));
AND2X2 AND2X2_147 ( .A(u5__abc_78290_new_n1469_), .B(mc_c_oe_d), .Y(u5__abc_78290_new_n1470_));
AND2X2 AND2X2_148 ( .A(u5__abc_78290_new_n1204_), .B(u5__abc_78290_new_n1491_), .Y(u5__abc_78290_new_n1492_));
AND2X2 AND2X2_149 ( .A(u5__abc_78290_new_n1549_), .B(u5__abc_78290_new_n1538_), .Y(u5__abc_78290_new_n1550_));
AND2X2 AND2X2_15 ( .A(u0__abc_74894_new_n4055_), .B(u0__abc_74894_new_n4058_), .Y(u0__abc_74894_new_n4059_));
AND2X2 AND2X2_150 ( .A(u5__abc_78290_new_n1497_), .B(u5__abc_78290_new_n1552_), .Y(u5__abc_78290_new_n1553_));
AND2X2 AND2X2_151 ( .A(u5__abc_78290_new_n1610_), .B(u1_wr_cycle), .Y(u5__abc_78290_new_n1611_));
AND2X2 AND2X2_152 ( .A(u5__abc_78290_new_n1624_), .B(u5__abc_78290_new_n1617_), .Y(u5__abc_78290_new_n1625_));
AND2X2 AND2X2_153 ( .A(u5__abc_78290_new_n1660_), .B(u5__abc_78290_new_n1661_), .Y(u5__abc_78290_new_n1662_));
AND2X2 AND2X2_154 ( .A(u5__abc_78290_new_n1665_), .B(u5__abc_78290_new_n1664_), .Y(u5__abc_78290_new_n1666_));
AND2X2 AND2X2_155 ( .A(u5__abc_78290_new_n1675_), .B(1'h0), .Y(u5__abc_78290_new_n1676_));
AND2X2 AND2X2_156 ( .A(u5__abc_78290_new_n1675_), .B(1'h0), .Y(u5__abc_78290_new_n1702_));
AND2X2 AND2X2_157 ( .A(u5__abc_78290_new_n1675_), .B(1'h0), .Y(u5__abc_78290_new_n1708_));
AND2X2 AND2X2_158 ( .A(u5__abc_78290_new_n1734_), .B(u5__abc_78290_new_n450_), .Y(u5__abc_78290_new_n1735_));
AND2X2 AND2X2_159 ( .A(u5__abc_78290_new_n591_), .B(u5__abc_78290_new_n427_), .Y(u5__abc_78290_new_n1738_));
AND2X2 AND2X2_16 ( .A(u0__abc_74894_new_n4087_), .B(u0__abc_74894_new_n4083_), .Y(u0__abc_74894_new_n4088_));
AND2X2 AND2X2_160 ( .A(u5__abc_78290_new_n1740_), .B(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n1741_));
AND2X2 AND2X2_161 ( .A(u5__abc_78290_new_n604_), .B(u5__abc_78290_new_n429_), .Y(u5__abc_78290_new_n1748_));
AND2X2 AND2X2_162 ( .A(u5__abc_78290_new_n1763_), .B(u5__abc_78290_new_n450_), .Y(u5__abc_78290_new_n1764_));
AND2X2 AND2X2_163 ( .A(u5__abc_78290_new_n1237_), .B(u5__abc_78290_new_n465_), .Y(u5__abc_78290_new_n1766_));
AND2X2 AND2X2_164 ( .A(u5__abc_78290_new_n1218_), .B(u5__abc_78290_new_n465_), .Y(u5__abc_78290_new_n1770_));
AND2X2 AND2X2_165 ( .A(u5__abc_78290_new_n1773_), .B(u5__abc_78290_new_n453_), .Y(u5__abc_78290_new_n1774_));
AND2X2 AND2X2_166 ( .A(u5__abc_78290_new_n1230_), .B(u5__abc_78290_new_n410_), .Y(u5__abc_78290_new_n1782_));
AND2X2 AND2X2_167 ( .A(u5__abc_78290_new_n1308_), .B(u5__abc_78290_new_n419_), .Y(u5__abc_78290_new_n1791_));
AND2X2 AND2X2_168 ( .A(u5__abc_78290_new_n1793_), .B(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n1794_));
AND2X2 AND2X2_169 ( .A(u5__abc_78290_new_n1279_), .B(u5__abc_78290_new_n413_), .Y(u5__abc_78290_new_n1797_));
AND2X2 AND2X2_17 ( .A(u0__abc_74894_new_n4097_), .B(u0__abc_74894_new_n4100_), .Y(u0__abc_74894_new_n4101_));
AND2X2 AND2X2_170 ( .A(u5__abc_78290_new_n1264_), .B(u5__abc_78290_new_n412_), .Y(u5__abc_78290_new_n1803_));
AND2X2 AND2X2_171 ( .A(u5__abc_78290_new_n1269_), .B(u5__abc_78290_new_n410_), .Y(u5__abc_78290_new_n1807_));
AND2X2 AND2X2_172 ( .A(u5__abc_78290_new_n1259_), .B(u5__abc_78290_new_n412_), .Y(u5__abc_78290_new_n1817_));
AND2X2 AND2X2_173 ( .A(u5__abc_78290_new_n1288_), .B(u5__abc_78290_new_n417_), .Y(u5__abc_78290_new_n1822_));
AND2X2 AND2X2_174 ( .A(u5__abc_78290_new_n1285_), .B(u5__abc_78290_new_n417_), .Y(u5__abc_78290_new_n1825_));
AND2X2 AND2X2_175 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n1837_), .Y(u5__abc_78290_new_n1838_));
AND2X2 AND2X2_176 ( .A(u5__abc_78290_new_n1140_), .B(u5__abc_78290_new_n388_), .Y(u5__abc_78290_new_n1844_));
AND2X2 AND2X2_177 ( .A(u5__abc_78290_new_n1846_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1847_));
AND2X2 AND2X2_178 ( .A(u5__abc_78290_new_n1855_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1856_));
AND2X2 AND2X2_179 ( .A(u5__abc_78290_new_n1119_), .B(u5__abc_78290_new_n465_), .Y(u5__abc_78290_new_n1860_));
AND2X2 AND2X2_18 ( .A(u0__abc_74894_new_n4109_), .B(u0__abc_74894_new_n4105_), .Y(u0__abc_74894_new_n4110_));
AND2X2 AND2X2_180 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n1874_), .Y(u5__abc_78290_new_n1875_));
AND2X2 AND2X2_181 ( .A(u5__abc_78290_new_n1885_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1886_));
AND2X2 AND2X2_182 ( .A(u5__abc_78290_new_n1056_), .B(u5__abc_78290_new_n420_), .Y(u5__abc_78290_new_n1909_));
AND2X2 AND2X2_183 ( .A(u5__abc_78290_new_n1911_), .B(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n1912_));
AND2X2 AND2X2_184 ( .A(u5__abc_78290_new_n1913_), .B(u5__abc_78290_new_n1904_), .Y(u5__abc_78290_new_n1914_));
AND2X2 AND2X2_185 ( .A(u5__abc_78290_new_n1924_), .B(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n1925_));
AND2X2 AND2X2_186 ( .A(u5__abc_78290_new_n1100_), .B(u5__abc_78290_new_n382_), .Y(u5__abc_78290_new_n1927_));
AND2X2 AND2X2_187 ( .A(u5__abc_78290_new_n1106_), .B(u5__abc_78290_new_n381_), .Y(u5__abc_78290_new_n1931_));
AND2X2 AND2X2_188 ( .A(u5__abc_78290_new_n1110_), .B(u5__abc_78290_new_n386_), .Y(u5__abc_78290_new_n1943_));
AND2X2 AND2X2_189 ( .A(u5__abc_78290_new_n1945_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1946_));
AND2X2 AND2X2_19 ( .A(u0__abc_74894_new_n4119_), .B(u0__abc_74894_new_n4122_), .Y(u0__abc_74894_new_n4123_));
AND2X2 AND2X2_190 ( .A(u5__abc_78290_new_n1675_), .B(1'h0), .Y(u5__abc_78290_new_n1956_));
AND2X2 AND2X2_191 ( .A(u5__abc_78290_new_n1675_), .B(page_size_8_), .Y(u5__abc_78290_new_n1964_));
AND2X2 AND2X2_192 ( .A(u5__abc_78290_new_n1675_), .B(page_size_9_), .Y(u5__abc_78290_new_n1972_));
AND2X2 AND2X2_193 ( .A(u5__abc_78290_new_n1675_), .B(page_size_10_), .Y(u5__abc_78290_new_n1979_));
AND2X2 AND2X2_194 ( .A(u5__abc_78290_new_n1985_), .B(u5__abc_78290_new_n1984_), .Y(u5__abc_78290_new_n1986_));
AND2X2 AND2X2_195 ( .A(u5__abc_78290_new_n2001_), .B(u5__abc_78290_new_n1187_), .Y(u5__abc_78290_new_n2002_));
AND2X2 AND2X2_196 ( .A(u5__abc_78290_new_n2015_), .B(u5_ir_cnt_2_), .Y(u5__abc_78290_new_n2016_));
AND2X2 AND2X2_197 ( .A(u5__abc_78290_new_n2025_), .B(u5__abc_78290_new_n1544_), .Y(u5__abc_78290_new_n2026_));
AND2X2 AND2X2_198 ( .A(u5__abc_78290_new_n1240_), .B(u5__abc_78290_new_n1984_), .Y(u5__abc_78290_new_n2028_));
AND2X2 AND2X2_199 ( .A(u5__abc_78290_new_n798_), .B(u5__abc_78290_new_n2050_), .Y(u5__abc_78290_new_n2051_));
AND2X2 AND2X2_2 ( .A(u0__abc_74894_new_n3710_), .B(u0__abc_74894_new_n3705_), .Y(u0__abc_74894_new_n3711_));
AND2X2 AND2X2_20 ( .A(u0__abc_74894_new_n4134_), .B(u0__abc_74894_new_n4137_), .Y(u0__abc_74894_new_n4138_));
AND2X2 AND2X2_200 ( .A(u5__abc_78290_new_n521_), .B(u5__abc_78290_new_n511_), .Y(u5__abc_78290_new_n2058_));
AND2X2 AND2X2_201 ( .A(u5__abc_78290_new_n2088_), .B(u5__abc_78290_new_n2089_), .Y(u5__abc_78290_new_n2090_));
AND2X2 AND2X2_202 ( .A(u5__abc_78290_new_n2094_), .B(u5__abc_78290_new_n2090_), .Y(u5__abc_78290_new_n2095_));
AND2X2 AND2X2_203 ( .A(u5__abc_78290_new_n1539_), .B(u5__abc_78290_new_n419_), .Y(u5__abc_78290_new_n2098_));
AND2X2 AND2X2_204 ( .A(u5__abc_78290_new_n2117_), .B(u5__abc_78290_new_n2116_), .Y(u5__abc_78290_new_n2118_));
AND2X2 AND2X2_205 ( .A(u5__abc_78290_new_n2121_), .B(u5__abc_78290_new_n2118_), .Y(u5__abc_78290_new_n2122_));
AND2X2 AND2X2_206 ( .A(u5__abc_78290_new_n2129_), .B(u5__abc_78290_new_n2131_), .Y(u5__abc_78290_new_n2132_));
AND2X2 AND2X2_207 ( .A(u5__abc_78290_new_n837_), .B(u5__abc_78290_new_n2137_), .Y(u5__abc_78290_new_n2138_));
AND2X2 AND2X2_208 ( .A(u5__abc_78290_new_n612_), .B(u5__abc_78290_new_n997_), .Y(u5__abc_78290_new_n2139_));
AND2X2 AND2X2_209 ( .A(u5__abc_78290_new_n2139_), .B(u5__abc_78290_new_n2138_), .Y(u5__abc_78290_new_n2140_));
AND2X2 AND2X2_21 ( .A(u0__abc_74894_new_n4176_), .B(u0__abc_74894_new_n4179_), .Y(u0__abc_74894_new_n4180_));
AND2X2 AND2X2_210 ( .A(u5__abc_78290_new_n868_), .B(u5__abc_78290_new_n874_), .Y(u5__abc_78290_new_n2152_));
AND2X2 AND2X2_211 ( .A(u5__abc_78290_new_n2153_), .B(u5__abc_78290_new_n2152_), .Y(u5__abc_78290_new_n2154_));
AND2X2 AND2X2_212 ( .A(u5__abc_78290_new_n952_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n2155_));
AND2X2 AND2X2_213 ( .A(u5__abc_78290_new_n2025_), .B(u5__abc_78290_new_n2170_), .Y(u5__abc_78290_new_n2171_));
AND2X2 AND2X2_214 ( .A(u5__abc_78290_new_n2178_), .B(u5__abc_78290_new_n2186_), .Y(u5__abc_78290_new_n2187_));
AND2X2 AND2X2_215 ( .A(u5__abc_78290_new_n2191_), .B(u5__abc_78290_new_n1148_), .Y(u5__abc_78290_new_n2192_));
AND2X2 AND2X2_216 ( .A(u5__abc_78290_new_n2208_), .B(u5__abc_78290_new_n2205_), .Y(u5__abc_78290_new_n2209_));
AND2X2 AND2X2_217 ( .A(u5__abc_78290_new_n2235_), .B(u5__abc_78290_new_n2233_), .Y(u5__abc_78290_new_n2236_));
AND2X2 AND2X2_218 ( .A(u5__abc_78290_new_n2241_), .B(u5__abc_78290_new_n2242_), .Y(u5__abc_78290_new_n2243_));
AND2X2 AND2X2_219 ( .A(u5__abc_78290_new_n2280_), .B(u5__abc_78290_new_n2277_), .Y(u5__abc_78290_new_n2281_));
AND2X2 AND2X2_22 ( .A(u0__abc_74894_new_n3701_), .B(1'h0), .Y(u0__abc_74894_new_n4420_));
AND2X2 AND2X2_220 ( .A(u5__abc_78290_new_n580_), .B(u5__abc_78290_new_n1984_), .Y(u5__abc_78290_new_n2284_));
AND2X2 AND2X2_221 ( .A(u5__abc_78290_new_n2335_), .B(u5__abc_78290_new_n2034_), .Y(u5__abc_78290_new_n2336_));
AND2X2 AND2X2_222 ( .A(u5__abc_78290_new_n2342_), .B(u5_timer_5_), .Y(u5__abc_78290_new_n2349_));
AND2X2 AND2X2_223 ( .A(u5__abc_78290_new_n2336_), .B(u5__abc_78290_new_n2338_), .Y(u5__abc_78290_new_n2350_));
AND2X2 AND2X2_224 ( .A(u5__abc_78290_new_n648_), .B(u5__abc_78290_new_n659_), .Y(u5__abc_78290_new_n2372_));
AND2X2 AND2X2_225 ( .A(u5__abc_78290_new_n1567_), .B(u5__abc_78290_new_n2384_), .Y(u5__abc_78290_new_n2385_));
AND2X2 AND2X2_226 ( .A(u5__abc_78290_new_n1495_), .B(u5__abc_78290_new_n1297_), .Y(u5__abc_78290_new_n2386_));
AND2X2 AND2X2_227 ( .A(u5__abc_78290_new_n2416_), .B(u5__abc_78290_new_n2422_), .Y(u5__abc_78290_new_n2423_));
AND2X2 AND2X2_228 ( .A(u5__abc_78290_new_n2435_), .B(u5__abc_78290_new_n668_), .Y(u5__abc_78290_new_n2436_));
AND2X2 AND2X2_229 ( .A(u5__abc_78290_new_n2371_), .B(u5__abc_78290_new_n2436_), .Y(u5__abc_78290_new_n2437_));
AND2X2 AND2X2_23 ( .A(u0__abc_74894_new_n4444_), .B(1'h0), .Y(cs_need_rfr_2_));
AND2X2 AND2X2_230 ( .A(u5__abc_78290_new_n2047_), .B(u5__abc_78290_new_n2050_), .Y(u5__abc_78290_new_n2445_));
AND2X2 AND2X2_231 ( .A(u5__abc_78290_new_n2443_), .B(u5__abc_78290_new_n2449_), .Y(u5__abc_78290_new_n2450_));
AND2X2 AND2X2_232 ( .A(u5__abc_78290_new_n2457_), .B(u5__abc_78290_new_n2459_), .Y(u5__abc_78290_new_n2460_));
AND2X2 AND2X2_233 ( .A(u5__abc_78290_new_n1567_), .B(u5__abc_78290_new_n2388_), .Y(u5__abc_78290_new_n2467_));
AND2X2 AND2X2_234 ( .A(u5__abc_78290_new_n1567_), .B(u5__abc_78290_new_n2390_), .Y(u5__abc_78290_new_n2497_));
AND2X2 AND2X2_235 ( .A(u5__abc_78290_new_n2568_), .B(u5__abc_78290_new_n1349_), .Y(u5__abc_78290_new_n2569_));
AND2X2 AND2X2_236 ( .A(u5__abc_78290_new_n2632_), .B(u5__abc_78290_new_n2630_), .Y(u5__abc_78290_new_n2633_));
AND2X2 AND2X2_237 ( .A(u5__abc_78290_new_n2623_), .B(u5__abc_78290_new_n2633_), .Y(u5__abc_78290_new_n2634_));
AND2X2 AND2X2_238 ( .A(u5__abc_78290_new_n2713_), .B(u5__abc_78290_new_n2714_), .Y(u5__abc_78290_new_n2715_));
AND2X2 AND2X2_239 ( .A(u5__abc_78290_new_n2680_), .B(u5_state_32_), .Y(u5__abc_78290_new_n2853_));
AND2X2 AND2X2_24 ( .A(u0__abc_74894_new_n4450_), .B(1'h0), .Y(cs_need_rfr_4_));
AND2X2 AND2X2_240 ( .A(u5__abc_78290_new_n2861_), .B(u5_state_36_), .Y(u5__abc_78290_new_n2862_));
AND2X2 AND2X2_241 ( .A(u5__abc_78290_new_n1526_), .B(u5_tmr2_done), .Y(u5__abc_78290_new_n2883_));
AND2X2 AND2X2_242 ( .A(u5__abc_78290_new_n2948_), .B(u5__abc_78290_new_n2953_), .Y(u5__abc_78290_new_n2954_));
AND2X2 AND2X2_243 ( .A(u5__abc_78290_new_n2997_), .B(u5__abc_78290_new_n2998_), .Y(u5__abc_78290_new_n2999_));
AND2X2 AND2X2_244 ( .A(u5__abc_78290_new_n3001_), .B(u5__abc_78290_new_n2993_), .Y(u5_pack_le0_d));
AND2X2 AND2X2_245 ( .A(u5__abc_78290_new_n484_), .B(u5__abc_78290_new_n1222_), .Y(u5__abc_78290_new_n3029_));
AND2X2 AND2X2_246 ( .A(u5__abc_78290_new_n3031_), .B(u5__abc_78290_new_n3028_), .Y(u5__abc_78290_new_n3032_));
AND2X2 AND2X2_247 ( .A(u5__abc_78290_new_n2283_), .B(u5__abc_78290_new_n2024_), .Y(u5__abc_78290_new_n3056_));
AND2X2 AND2X2_248 ( .A(u5__abc_78290_new_n3062_), .B(u5__abc_78290_new_n2171_), .Y(u5__abc_78290_new_n3063_));
AND2X2 AND2X2_249 ( .A(u5__abc_78290_new_n3068_), .B(u5__abc_78290_new_n2278_), .Y(u5__abc_78290_new_n3069_));
AND2X2 AND2X2_25 ( .A(u0__abc_74894_new_n4459_), .B(1'h0), .Y(cs_need_rfr_7_));
AND2X2 AND2X2_250 ( .A(u5__abc_78290_new_n1377_), .B(u5_cmd_a10_r), .Y(u5__abc_78290_new_n3110_));
AND2X2 AND2X2_251 ( .A(u5__abc_78290_new_n3103_), .B(u5__abc_78290_new_n3113_), .Y(u5__abc_78290_new_n3114_));
AND2X2 AND2X2_252 ( .A(u5__abc_78290_new_n2381_), .B(u5__abc_78290_new_n3117_), .Y(u5__abc_78290_new_n3118_));
AND2X2 AND2X2_253 ( .A(u5__abc_78290_new_n3136_), .B(u5__abc_78290_new_n2283_), .Y(u5__abc_78290_new_n3137_));
AND2X2 AND2X2_26 ( .A(u0__abc_74894_new_n4467_), .B(u0__abc_74894_new_n4468_), .Y(u0__abc_74894_new_n4469_));
AND2X2 AND2X2_27 ( .A(u0_u0__abc_72207_new_n214_), .B(u0_u0_addr_r_4_), .Y(u0_u0__abc_72207_new_n319_));
AND2X2 AND2X2_28 ( .A(u0_csc0_21_), .B(\wb_addr_i[26] ), .Y(u0_u0__abc_72207_new_n435_));
AND2X2 AND2X2_29 ( .A(u0_csc0_19_), .B(\wb_addr_i[24] ), .Y(u0_u0__abc_72207_new_n437_));
AND2X2 AND2X2_3 ( .A(u0__abc_74894_new_n3712_), .B(u0__abc_74894_new_n3705_), .Y(u0__abc_74894_new_n3713_));
AND2X2 AND2X2_30 ( .A(u0_csc0_16_), .B(\wb_addr_i[21] ), .Y(u0_u0__abc_72207_new_n443_));
AND2X2 AND2X2_31 ( .A(u0_csc0_18_), .B(\wb_addr_i[23] ), .Y(u0_u0__abc_72207_new_n445_));
AND2X2 AND2X2_32 ( .A(u0_csc0_23_), .B(\wb_addr_i[28] ), .Y(u0_u0__abc_72207_new_n449_));
AND2X2 AND2X2_33 ( .A(u0_csc0_22_), .B(\wb_addr_i[27] ), .Y(u0_u0__abc_72207_new_n452_));
AND2X2 AND2X2_34 ( .A(u0_csc0_20_), .B(\wb_addr_i[25] ), .Y(u0_u0__abc_72207_new_n454_));
AND2X2 AND2X2_35 ( .A(u0_csc1_21_), .B(\wb_addr_i[26] ), .Y(u0_u1__abc_72470_new_n412_));
AND2X2 AND2X2_36 ( .A(u0_csc1_19_), .B(\wb_addr_i[24] ), .Y(u0_u1__abc_72470_new_n414_));
AND2X2 AND2X2_37 ( .A(u0_csc1_16_), .B(\wb_addr_i[21] ), .Y(u0_u1__abc_72470_new_n419_));
AND2X2 AND2X2_38 ( .A(u0_csc1_18_), .B(\wb_addr_i[23] ), .Y(u0_u1__abc_72470_new_n421_));
AND2X2 AND2X2_39 ( .A(u0_csc1_23_), .B(\wb_addr_i[28] ), .Y(u0_u1__abc_72470_new_n425_));
AND2X2 AND2X2_4 ( .A(\wb_addr_i[5] ), .B(\wb_addr_i[4] ), .Y(u0__abc_74894_new_n3718_));
AND2X2 AND2X2_40 ( .A(u0_csc1_22_), .B(\wb_addr_i[27] ), .Y(u0_u1__abc_72470_new_n428_));
AND2X2 AND2X2_41 ( .A(u0_csc1_20_), .B(\wb_addr_i[25] ), .Y(u0_u1__abc_72470_new_n430_));
AND2X2 AND2X2_42 ( .A(u1__abc_72801_new_n353_), .B(u1__abc_72801_new_n354_), .Y(u1__abc_72801_new_n355_));
AND2X2 AND2X2_43 ( .A(u1__abc_72801_new_n361_), .B(u1__abc_72801_new_n341_), .Y(u1__abc_72801_new_n362_));
AND2X2 AND2X2_44 ( .A(u1__abc_72801_new_n365_), .B(u1__abc_72801_new_n366_), .Y(u1__abc_72801_new_n367_));
AND2X2 AND2X2_45 ( .A(u1__abc_72801_new_n373_), .B(u1__abc_72801_new_n374_), .Y(u1__abc_72801_new_n375_));
AND2X2 AND2X2_46 ( .A(u1__abc_72801_new_n383_), .B(u1__abc_72801_new_n384_), .Y(u1__abc_72801_new_n385_));
AND2X2 AND2X2_47 ( .A(u1__abc_72801_new_n392_), .B(u1__abc_72801_new_n393_), .Y(u1__abc_72801_new_n394_));
AND2X2 AND2X2_48 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[2] ), .Y(u1__abc_72801_new_n506_));
AND2X2 AND2X2_49 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[3] ), .Y(u1__abc_72801_new_n511_));
AND2X2 AND2X2_5 ( .A(u0__abc_74894_new_n3688_), .B(u0__abc_74894_new_n3724_), .Y(u0__abc_74894_new_n3727_));
AND2X2 AND2X2_50 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[4] ), .Y(u1__abc_72801_new_n516_));
AND2X2 AND2X2_51 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[5] ), .Y(u1__abc_72801_new_n521_));
AND2X2 AND2X2_52 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[6] ), .Y(u1__abc_72801_new_n526_));
AND2X2 AND2X2_53 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[7] ), .Y(u1__abc_72801_new_n531_));
AND2X2 AND2X2_54 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[8] ), .Y(u1__abc_72801_new_n536_));
AND2X2 AND2X2_55 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[10] ), .Y(u1__abc_72801_new_n549_));
AND2X2 AND2X2_56 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[11] ), .Y(u1__abc_72801_new_n554_));
AND2X2 AND2X2_57 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[12] ), .Y(u1__abc_72801_new_n559_));
AND2X2 AND2X2_58 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[13] ), .Y(u1__abc_72801_new_n564_));
AND2X2 AND2X2_59 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[17] ), .Y(u1__abc_72801_new_n586_));
AND2X2 AND2X2_6 ( .A(u0__abc_74894_new_n3712_), .B(u0__abc_74894_new_n3718_), .Y(u0__abc_74894_new_n3741_));
AND2X2 AND2X2_60 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[18] ), .Y(u1__abc_72801_new_n592_));
AND2X2 AND2X2_61 ( .A(u1_u0__abc_72719_new_n67_), .B(u1_u0__abc_72719_new_n71_), .Y(u1_u0__0out_r_12_0__7_));
AND2X2 AND2X2_62 ( .A(u1_u0__abc_72719_new_n76_), .B(u1_u0__abc_72719_new_n78_), .Y(u1_u0__0out_r_12_0__9_));
AND2X2 AND2X2_63 ( .A(u1_u0__abc_72719_new_n86_), .B(u1_u0__abc_72719_new_n85_), .Y(u1_u0__0out_r_12_0__11_));
AND2X2 AND2X2_64 ( .A(u1_u0_inc_next), .B(u1_acs_addr_12_), .Y(u1_u0__abc_72719_new_n89_));
AND2X2 AND2X2_65 ( .A(u1_acs_addr_14_), .B(u1_acs_addr_15_), .Y(u1_u0__abc_72719_new_n96_));
AND2X2 AND2X2_66 ( .A(u1_u0__abc_72719_new_n95_), .B(u1_u0__abc_72719_new_n97_), .Y(u1_acs_addr_pl1_15_));
AND2X2 AND2X2_67 ( .A(u1_acs_addr_16_), .B(u1_acs_addr_17_), .Y(u1_u0__abc_72719_new_n113_));
AND2X2 AND2X2_68 ( .A(u1_acs_addr_18_), .B(u1_acs_addr_19_), .Y(u1_u0__abc_72719_new_n114_));
AND2X2 AND2X2_69 ( .A(u1_u0__abc_72719_new_n116_), .B(u1_u0__abc_72719_new_n111_), .Y(u1_acs_addr_pl1_20_));
AND2X2 AND2X2_7 ( .A(u0__abc_74894_new_n3706_), .B(u0__abc_74894_new_n3718_), .Y(u0__abc_74894_new_n3743_));
AND2X2 AND2X2_70 ( .A(u2__abc_74202_new_n100_), .B(u2__abc_74202_new_n101_), .Y(u2__abc_74202_new_n102_));
AND2X2 AND2X2_71 ( .A(u2__abc_74202_new_n103_), .B(u2__abc_74202_new_n104_), .Y(u2__abc_74202_new_n105_));
AND2X2 AND2X2_72 ( .A(u2__abc_74202_new_n107_), .B(u2__abc_74202_new_n108_), .Y(u2__abc_74202_new_n109_));
AND2X2 AND2X2_73 ( .A(u2__abc_74202_new_n110_), .B(u2__abc_74202_new_n111_), .Y(u2__abc_74202_new_n112_));
AND2X2 AND2X2_74 ( .A(u2_u0_b3_last_row_10_), .B(row_adr_10_), .Y(u2_u0__abc_73914_new_n285_));
AND2X2 AND2X2_75 ( .A(u2_u0_b3_last_row_3_), .B(row_adr_3_), .Y(u2_u0__abc_73914_new_n288_));
AND2X2 AND2X2_76 ( .A(row_adr_10_), .B(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_73914_new_n385_));
AND2X2 AND2X2_77 ( .A(row_adr_5_), .B(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_73914_new_n389_));
AND2X2 AND2X2_78 ( .A(u2_u1_b3_last_row_10_), .B(row_adr_10_), .Y(u2_u1__abc_73914_new_n285_));
AND2X2 AND2X2_79 ( .A(u2_u1_b3_last_row_3_), .B(row_adr_3_), .Y(u2_u1__abc_73914_new_n288_));
AND2X2 AND2X2_8 ( .A(u0__abc_74894_new_n3710_), .B(u0__abc_74894_new_n3718_), .Y(u0__abc_74894_new_n3745_));
AND2X2 AND2X2_80 ( .A(row_adr_10_), .B(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_73914_new_n385_));
AND2X2 AND2X2_81 ( .A(row_adr_5_), .B(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_73914_new_n389_));
AND2X2 AND2X2_82 ( .A(mem_ack_r), .B(u3_wb_read_go), .Y(u3_re));
AND2X2 AND2X2_83 ( .A(u3_rd_fifo_out_8_), .B(u3_rd_fifo_out_9_), .Y(u3__abc_73372_new_n636_));
AND2X2 AND2X2_84 ( .A(u3_rd_fifo_out_20_), .B(u3_rd_fifo_out_21_), .Y(u3__abc_73372_new_n665_));
AND2X2 AND2X2_85 ( .A(u3_rd_fifo_out_18_), .B(u3_rd_fifo_out_19_), .Y(u3__abc_73372_new_n672_));
AND2X2 AND2X2_86 ( .A(u3__abc_73372_new_n676_), .B(\wb_sel_i[2] ), .Y(u3__abc_73372_new_n677_));
AND2X2 AND2X2_87 ( .A(u3_rd_fifo_out_0_), .B(u3_rd_fifo_out_1_), .Y(u3__abc_73372_new_n685_));
AND2X2 AND2X2_88 ( .A(u3_rd_fifo_out_28_), .B(u3_rd_fifo_out_29_), .Y(u3__abc_73372_new_n715_));
AND2X2 AND2X2_89 ( .A(u3_rd_fifo_out_26_), .B(u3_rd_fifo_out_27_), .Y(u3__abc_73372_new_n722_));
AND2X2 AND2X2_9 ( .A(u0__abc_74894_new_n3706_), .B(u0__abc_74894_new_n3688_), .Y(u0__abc_74894_new_n3749_));
AND2X2 AND2X2_90 ( .A(u3__abc_73372_new_n726_), .B(\wb_sel_i[3] ), .Y(u3__abc_73372_new_n727_));
AND2X2 AND2X2_91 ( .A(u3_u0__abc_74260_new_n738_), .B(u3_u0__abc_74260_new_n737_), .Y(u3_u0__abc_74260_new_n742_));
AND2X2 AND2X2_92 ( .A(u4__abc_74770_new_n65_), .B(u4__abc_74770_new_n66_), .Y(u4__abc_74770_new_n67_));
AND2X2 AND2X2_93 ( .A(u4_rfr_ce), .B(u4_rfr_cnt_0_), .Y(u4__abc_74770_new_n93_));
AND2X2 AND2X2_94 ( .A(u4__abc_74770_new_n127_), .B(u4__abc_74770_new_n128_), .Y(u4__abc_74770_new_n129_));
AND2X2 AND2X2_95 ( .A(u4__0rfr_early_0_0_), .B(u4__abc_74770_new_n132_), .Y(u4_ps_cnt_clr));
AND2X2 AND2X2_96 ( .A(u5__abc_78290_new_n378_), .B(u5__abc_78290_new_n379_), .Y(u5__abc_78290_new_n380_));
AND2X2 AND2X2_97 ( .A(u5__abc_78290_new_n381_), .B(u5__abc_78290_new_n382_), .Y(u5__abc_78290_new_n383_));
AND2X2 AND2X2_98 ( .A(u5__abc_78290_new_n385_), .B(u5__abc_78290_new_n386_), .Y(u5__abc_78290_new_n387_));
AND2X2 AND2X2_99 ( .A(u5__abc_78290_new_n388_), .B(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n390_));
AOI21X1 AOI21X1_1 ( .A(_abc_81086_new_n464_), .B(_abc_81086_new_n463_), .C(_abc_81086_new_n465_), .Y(not_mem_cyc));
AOI21X1 AOI21X1_10 ( .A(u0__abc_74894_new_n1247_), .B(u0__abc_74894_new_n1248_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1249_));
AOI21X1 AOI21X1_100 ( .A(u0__abc_74894_new_n2645_), .B(u0__abc_74894_new_n2646_), .C(u0_cs1), .Y(u0__abc_74894_new_n2647_));
AOI21X1 AOI21X1_101 ( .A(u0__abc_74894_new_n1412_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2649_));
AOI21X1 AOI21X1_102 ( .A(u0__abc_74894_new_n2661_), .B(u0__abc_74894_new_n2662_), .C(u0_cs1), .Y(u0__abc_74894_new_n2663_));
AOI21X1 AOI21X1_103 ( .A(u0__abc_74894_new_n1432_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2665_));
AOI21X1 AOI21X1_104 ( .A(u0__abc_74894_new_n2677_), .B(u0__abc_74894_new_n2678_), .C(u0_cs1), .Y(u0__abc_74894_new_n2679_));
AOI21X1 AOI21X1_105 ( .A(u0__abc_74894_new_n1452_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2681_));
AOI21X1 AOI21X1_106 ( .A(u0__abc_74894_new_n2693_), .B(u0__abc_74894_new_n2694_), .C(u0_cs1), .Y(u0__abc_74894_new_n2695_));
AOI21X1 AOI21X1_107 ( .A(u0__abc_74894_new_n1472_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2697_));
AOI21X1 AOI21X1_108 ( .A(u0__abc_74894_new_n2709_), .B(u0__abc_74894_new_n2710_), .C(u0_cs1), .Y(u0__abc_74894_new_n2711_));
AOI21X1 AOI21X1_109 ( .A(u0__abc_74894_new_n1492_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2713_));
AOI21X1 AOI21X1_11 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1252_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1253_));
AOI21X1 AOI21X1_110 ( .A(u0__abc_74894_new_n2725_), .B(u0__abc_74894_new_n2726_), .C(u0_cs1), .Y(u0__abc_74894_new_n2727_));
AOI21X1 AOI21X1_111 ( .A(u0__abc_74894_new_n1512_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2729_));
AOI21X1 AOI21X1_112 ( .A(u0__abc_74894_new_n2741_), .B(u0__abc_74894_new_n2742_), .C(u0_cs1), .Y(u0__abc_74894_new_n2743_));
AOI21X1 AOI21X1_113 ( .A(u0__abc_74894_new_n1532_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2745_));
AOI21X1 AOI21X1_114 ( .A(u0__abc_74894_new_n2757_), .B(u0__abc_74894_new_n2758_), .C(u0_cs1), .Y(u0__abc_74894_new_n2759_));
AOI21X1 AOI21X1_115 ( .A(u0__abc_74894_new_n1552_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2761_));
AOI21X1 AOI21X1_116 ( .A(u0__abc_74894_new_n2773_), .B(u0__abc_74894_new_n2774_), .C(u0_cs1), .Y(u0__abc_74894_new_n2775_));
AOI21X1 AOI21X1_117 ( .A(u0__abc_74894_new_n1572_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2777_));
AOI21X1 AOI21X1_118 ( .A(u0__abc_74894_new_n2789_), .B(u0__abc_74894_new_n2790_), .C(u0_cs1), .Y(u0__abc_74894_new_n2791_));
AOI21X1 AOI21X1_119 ( .A(u0__abc_74894_new_n1592_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2793_));
AOI21X1 AOI21X1_12 ( .A(u0__abc_74894_new_n1267_), .B(u0__abc_74894_new_n1268_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1269_));
AOI21X1 AOI21X1_120 ( .A(u0__abc_74894_new_n2805_), .B(u0__abc_74894_new_n2806_), .C(u0_cs1), .Y(u0__abc_74894_new_n2807_));
AOI21X1 AOI21X1_121 ( .A(u0__abc_74894_new_n1612_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2809_));
AOI21X1 AOI21X1_122 ( .A(u0__abc_74894_new_n2821_), .B(u0__abc_74894_new_n2822_), .C(u0_cs1), .Y(u0__abc_74894_new_n2823_));
AOI21X1 AOI21X1_123 ( .A(u0__abc_74894_new_n1632_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2825_));
AOI21X1 AOI21X1_124 ( .A(u0__abc_74894_new_n2837_), .B(u0__abc_74894_new_n2838_), .C(u0_cs1), .Y(u0__abc_74894_new_n2839_));
AOI21X1 AOI21X1_125 ( .A(u0__abc_74894_new_n1652_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2841_));
AOI21X1 AOI21X1_126 ( .A(u0__abc_74894_new_n2853_), .B(u0__abc_74894_new_n2854_), .C(u0_cs1), .Y(u0__abc_74894_new_n2855_));
AOI21X1 AOI21X1_127 ( .A(u0__abc_74894_new_n1672_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2857_));
AOI21X1 AOI21X1_128 ( .A(u0__abc_74894_new_n2869_), .B(u0__abc_74894_new_n2870_), .C(u0_cs1), .Y(u0__abc_74894_new_n2871_));
AOI21X1 AOI21X1_129 ( .A(u0__abc_74894_new_n1692_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2873_));
AOI21X1 AOI21X1_13 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1272_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1273_));
AOI21X1 AOI21X1_130 ( .A(u0__abc_74894_new_n2885_), .B(u0__abc_74894_new_n2886_), .C(u0_cs1), .Y(u0__abc_74894_new_n2887_));
AOI21X1 AOI21X1_131 ( .A(u0__abc_74894_new_n1712_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2889_));
AOI21X1 AOI21X1_132 ( .A(u0__abc_74894_new_n2984_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2985_), .Y(u0__abc_74894_new_n2986_));
AOI21X1 AOI21X1_133 ( .A(u0__abc_74894_new_n3000_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3001_), .Y(u0__abc_74894_new_n3002_));
AOI21X1 AOI21X1_134 ( .A(u0__abc_74894_new_n3016_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3017_), .Y(u0__abc_74894_new_n3018_));
AOI21X1 AOI21X1_135 ( .A(u0__abc_74894_new_n3032_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3033_), .Y(u0__abc_74894_new_n3034_));
AOI21X1 AOI21X1_136 ( .A(u0__abc_74894_new_n3048_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3049_), .Y(u0__abc_74894_new_n3050_));
AOI21X1 AOI21X1_137 ( .A(u0__abc_74894_new_n3064_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3065_), .Y(u0__abc_74894_new_n3066_));
AOI21X1 AOI21X1_138 ( .A(u0__abc_74894_new_n3080_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3081_), .Y(u0__abc_74894_new_n3082_));
AOI21X1 AOI21X1_139 ( .A(u0__abc_74894_new_n3112_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3113_), .Y(u0__abc_74894_new_n3114_));
AOI21X1 AOI21X1_14 ( .A(u0__abc_74894_new_n1287_), .B(u0__abc_74894_new_n1288_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1289_));
AOI21X1 AOI21X1_140 ( .A(u0__abc_74894_new_n3128_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3129_), .Y(u0__abc_74894_new_n3130_));
AOI21X1 AOI21X1_141 ( .A(u0__abc_74894_new_n3144_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n3145_), .Y(u0__abc_74894_new_n3146_));
AOI21X1 AOI21X1_142 ( .A(u0__abc_74894_new_n2455_), .B(cs_le), .C(u0__abc_74894_new_n3479_), .Y(u0__0cs_7_0__0_));
AOI21X1 AOI21X1_143 ( .A(u0__abc_74894_new_n2454_), .B(cs_le), .C(u0__abc_74894_new_n3481_), .Y(u0__0cs_7_0__1_));
AOI21X1 AOI21X1_144 ( .A(u0__abc_74894_new_n2438_), .B(cs_le), .C(u0__abc_74894_new_n3483_), .Y(u0__0cs_7_0__2_));
AOI21X1 AOI21X1_145 ( .A(u0__abc_74894_new_n2440_), .B(cs_le), .C(u0__abc_74894_new_n3485_), .Y(u0__0cs_7_0__3_));
AOI21X1 AOI21X1_146 ( .A(u0__abc_74894_new_n2441_), .B(cs_le), .C(u0__abc_74894_new_n3487_), .Y(u0__0cs_7_0__4_));
AOI21X1 AOI21X1_147 ( .A(u0__abc_74894_new_n2443_), .B(cs_le), .C(u0__abc_74894_new_n3489_), .Y(u0__0cs_7_0__5_));
AOI21X1 AOI21X1_148 ( .A(u0__abc_74894_new_n2444_), .B(cs_le), .C(u0__abc_74894_new_n3491_), .Y(u0__0cs_7_0__6_));
AOI21X1 AOI21X1_149 ( .A(u0_csr_0_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n3739_), .Y(u0__abc_74894_new_n3740_));
AOI21X1 AOI21X1_15 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1292_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1293_));
AOI21X1 AOI21X1_150 ( .A(u0_csr_3_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n3819_), .Y(u0__abc_74894_new_n3820_));
AOI21X1 AOI21X1_151 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .C(u0__abc_74894_new_n3831_), .Y(u0__abc_74894_new_n3832_));
AOI21X1 AOI21X1_152 ( .A(u0_csr_5_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n3860_), .Y(u0__abc_74894_new_n3861_));
AOI21X1 AOI21X1_153 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .C(u0__abc_74894_new_n3872_), .Y(u0__abc_74894_new_n3873_));
AOI21X1 AOI21X1_154 ( .A(u0_csc1_7_), .B(u0__abc_74894_new_n3816_), .C(u0__abc_74894_new_n3890_), .Y(u0__abc_74894_new_n3891_));
AOI21X1 AOI21X1_155 ( .A(u0_tms1_7_), .B(u0__abc_74894_new_n3802_), .C(u0__abc_74894_new_n3895_), .Y(u0__abc_74894_new_n3896_));
AOI21X1 AOI21X1_156 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .C(u0__abc_74894_new_n3909_), .Y(u0__abc_74894_new_n3910_));
AOI21X1 AOI21X1_157 ( .A(u0_csc1_8_), .B(u0__abc_74894_new_n3816_), .C(u0__abc_74894_new_n3913_), .Y(u0__abc_74894_new_n3914_));
AOI21X1 AOI21X1_158 ( .A(u0_tms1_8_), .B(u0__abc_74894_new_n3802_), .C(u0__abc_74894_new_n3915_), .Y(u0__abc_74894_new_n3916_));
AOI21X1 AOI21X1_159 ( .A(ref_int_1_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n3936_), .Y(u0__abc_74894_new_n3937_));
AOI21X1 AOI21X1_16 ( .A(u0__abc_74894_new_n1307_), .B(u0__abc_74894_new_n1308_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1309_));
AOI21X1 AOI21X1_160 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .C(u0__abc_74894_new_n3948_), .Y(u0__abc_74894_new_n3949_));
AOI21X1 AOI21X1_161 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(u0__abc_74894_new_n4003_), .Y(u0__abc_74894_new_n4004_));
AOI21X1 AOI21X1_162 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .C(u0__abc_74894_new_n4006_), .Y(u0__abc_74894_new_n4007_));
AOI21X1 AOI21X1_163 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(u0__abc_74894_new_n4025_), .Y(u0__abc_74894_new_n4026_));
AOI21X1 AOI21X1_164 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .C(u0__abc_74894_new_n4028_), .Y(u0__abc_74894_new_n4029_));
AOI21X1 AOI21X1_165 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .C(u0__abc_74894_new_n4040_), .Y(u0__abc_74894_new_n4041_));
AOI21X1 AOI21X1_166 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(u0__abc_74894_new_n4050_), .Y(u0__abc_74894_new_n4051_));
AOI21X1 AOI21X1_167 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .C(u0__abc_74894_new_n4054_), .Y(u0__abc_74894_new_n4055_));
AOI21X1 AOI21X1_168 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(u0__abc_74894_new_n4057_), .Y(u0__abc_74894_new_n4058_));
AOI21X1 AOI21X1_169 ( .A(u0_csc1_16_), .B(u0__abc_74894_new_n3816_), .C(u0__abc_74894_new_n4069_), .Y(u0__abc_74894_new_n4070_));
AOI21X1 AOI21X1_17 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1312_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1313_));
AOI21X1 AOI21X1_170 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .C(u0__abc_74894_new_n4082_), .Y(u0__abc_74894_new_n4083_));
AOI21X1 AOI21X1_171 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(u0__abc_74894_new_n4092_), .Y(u0__abc_74894_new_n4093_));
AOI21X1 AOI21X1_172 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .C(u0__abc_74894_new_n4096_), .Y(u0__abc_74894_new_n4097_));
AOI21X1 AOI21X1_173 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(u0__abc_74894_new_n4099_), .Y(u0__abc_74894_new_n4100_));
AOI21X1 AOI21X1_174 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .C(u0__abc_74894_new_n4104_), .Y(u0__abc_74894_new_n4105_));
AOI21X1 AOI21X1_175 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(u0__abc_74894_new_n4114_), .Y(u0__abc_74894_new_n4115_));
AOI21X1 AOI21X1_176 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(u0__abc_74894_new_n4118_), .Y(u0__abc_74894_new_n4119_));
AOI21X1 AOI21X1_177 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .C(u0__abc_74894_new_n4121_), .Y(u0__abc_74894_new_n4122_));
AOI21X1 AOI21X1_178 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .C(u0__abc_74894_new_n4133_), .Y(u0__abc_74894_new_n4134_));
AOI21X1 AOI21X1_179 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(u0__abc_74894_new_n4136_), .Y(u0__abc_74894_new_n4137_));
AOI21X1 AOI21X1_18 ( .A(u0__abc_74894_new_n1327_), .B(u0__abc_74894_new_n1328_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1329_));
AOI21X1 AOI21X1_180 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(u0__abc_74894_new_n4175_), .Y(u0__abc_74894_new_n4176_));
AOI21X1 AOI21X1_181 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .C(u0__abc_74894_new_n4178_), .Y(u0__abc_74894_new_n4179_));
AOI21X1 AOI21X1_182 ( .A(u0_csc1_23_), .B(u0__abc_74894_new_n3816_), .C(u0__abc_74894_new_n4216_), .Y(u0__abc_74894_new_n4217_));
AOI21X1 AOI21X1_183 ( .A(rfr_ps_val_0_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n4240_), .Y(u0__abc_74894_new_n4241_));
AOI21X1 AOI21X1_184 ( .A(rfr_ps_val_1_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n4266_), .Y(u0__abc_74894_new_n4267_));
AOI21X1 AOI21X1_185 ( .A(rfr_ps_val_2_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n4292_), .Y(u0__abc_74894_new_n4293_));
AOI21X1 AOI21X1_186 ( .A(rfr_ps_val_3_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n4318_), .Y(u0__abc_74894_new_n4319_));
AOI21X1 AOI21X1_187 ( .A(rfr_ps_val_4_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n4345_), .Y(u0__abc_74894_new_n4346_));
AOI21X1 AOI21X1_188 ( .A(rfr_ps_val_5_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n4370_), .Y(u0__abc_74894_new_n4371_));
AOI21X1 AOI21X1_189 ( .A(rfr_ps_val_6_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n4394_), .Y(u0__abc_74894_new_n4395_));
AOI21X1 AOI21X1_19 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1332_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1333_));
AOI21X1 AOI21X1_190 ( .A(rfr_ps_val_7_), .B(u0__abc_74894_new_n3729_), .C(u0__abc_74894_new_n4418_), .Y(u0__abc_74894_new_n4419_));
AOI21X1 AOI21X1_191 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_0_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n223_));
AOI21X1 AOI21X1_192 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_1_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n226_));
AOI21X1 AOI21X1_193 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_2_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n229_));
AOI21X1 AOI21X1_194 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_3_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n232_));
AOI21X1 AOI21X1_195 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_4_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n235_));
AOI21X1 AOI21X1_196 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_5_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n238_));
AOI21X1 AOI21X1_197 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_6_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n241_));
AOI21X1 AOI21X1_198 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_7_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n244_));
AOI21X1 AOI21X1_199 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_8_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n247_));
AOI21X1 AOI21X1_2 ( .A(u0__abc_74894_new_n1167_), .B(u0__abc_74894_new_n1168_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1169_));
AOI21X1 AOI21X1_20 ( .A(u0__abc_74894_new_n1347_), .B(u0__abc_74894_new_n1348_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1349_));
AOI21X1 AOI21X1_200 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_9_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n250_));
AOI21X1 AOI21X1_201 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_10_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n253_));
AOI21X1 AOI21X1_202 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_11_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n256_));
AOI21X1 AOI21X1_203 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_12_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n259_));
AOI21X1 AOI21X1_204 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_13_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n262_));
AOI21X1 AOI21X1_205 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_14_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n265_));
AOI21X1 AOI21X1_206 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_15_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n268_));
AOI21X1 AOI21X1_207 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_16_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n271_));
AOI21X1 AOI21X1_208 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_17_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n274_));
AOI21X1 AOI21X1_209 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_18_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n277_));
AOI21X1 AOI21X1_21 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1352_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1353_));
AOI21X1 AOI21X1_210 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_19_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n280_));
AOI21X1 AOI21X1_211 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_20_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n283_));
AOI21X1 AOI21X1_212 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_21_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n286_));
AOI21X1 AOI21X1_213 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_22_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n289_));
AOI21X1 AOI21X1_214 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_23_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n292_));
AOI21X1 AOI21X1_215 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_24_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n295_));
AOI21X1 AOI21X1_216 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_25_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n298_));
AOI21X1 AOI21X1_217 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_26_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n301_));
AOI21X1 AOI21X1_218 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_27_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n304_));
AOI21X1 AOI21X1_219 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_28_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n307_));
AOI21X1 AOI21X1_22 ( .A(u0__abc_74894_new_n1367_), .B(u0__abc_74894_new_n1368_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1369_));
AOI21X1 AOI21X1_220 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_29_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n310_));
AOI21X1 AOI21X1_221 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_30_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n313_));
AOI21X1 AOI21X1_222 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_tms0_31_), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n316_));
AOI21X1 AOI21X1_223 ( .A(u0_u0__abc_72207_new_n219_), .B(u0_u0__abc_72207_new_n318_), .C(u0_csc0_1_), .Y(u0_u0__abc_72207_new_n333_));
AOI21X1 AOI21X1_224 ( .A(u0_u0__abc_72207_new_n219_), .B(u0_u0__abc_72207_new_n318_), .C(u0_csc0_2_), .Y(u0_u0__abc_72207_new_n337_));
AOI21X1 AOI21X1_225 ( .A(u0_u0__abc_72207_new_n206_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n340_), .Y(u0_u0__0csc_31_0__3_));
AOI21X1 AOI21X1_226 ( .A(u0_u0__abc_72207_new_n356_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n357_), .Y(u0_u0__0csc_31_0__6_));
AOI21X1 AOI21X1_227 ( .A(u0_u0__abc_72207_new_n359_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n360_), .Y(u0_u0__0csc_31_0__7_));
AOI21X1 AOI21X1_228 ( .A(u0_u0__abc_72207_new_n362_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n363_), .Y(u0_u0__0csc_31_0__8_));
AOI21X1 AOI21X1_229 ( .A(u0_u0__abc_72207_new_n365_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n366_), .Y(u0_u0__0csc_31_0__9_));
AOI21X1 AOI21X1_23 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1372_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1373_));
AOI21X1 AOI21X1_230 ( .A(u0_u0__abc_72207_new_n368_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n369_), .Y(u0_u0__0csc_31_0__10_));
AOI21X1 AOI21X1_231 ( .A(u0_u0__abc_72207_new_n371_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n372_), .Y(u0_u0__0csc_31_0__11_));
AOI21X1 AOI21X1_232 ( .A(u0_u0__abc_72207_new_n374_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n375_), .Y(u0_u0__0csc_31_0__12_));
AOI21X1 AOI21X1_233 ( .A(u0_u0__abc_72207_new_n377_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n378_), .Y(u0_u0__0csc_31_0__13_));
AOI21X1 AOI21X1_234 ( .A(u0_u0__abc_72207_new_n380_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n381_), .Y(u0_u0__0csc_31_0__14_));
AOI21X1 AOI21X1_235 ( .A(u0_u0__abc_72207_new_n383_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n384_), .Y(u0_u0__0csc_31_0__15_));
AOI21X1 AOI21X1_236 ( .A(u0_u0__abc_72207_new_n386_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n387_), .Y(u0_u0__0csc_31_0__16_));
AOI21X1 AOI21X1_237 ( .A(u0_u0__abc_72207_new_n389_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n390_), .Y(u0_u0__0csc_31_0__17_));
AOI21X1 AOI21X1_238 ( .A(u0_u0__abc_72207_new_n392_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n393_), .Y(u0_u0__0csc_31_0__18_));
AOI21X1 AOI21X1_239 ( .A(u0_u0__abc_72207_new_n395_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n396_), .Y(u0_u0__0csc_31_0__19_));
AOI21X1 AOI21X1_24 ( .A(u0__abc_74894_new_n1387_), .B(u0__abc_74894_new_n1388_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1389_));
AOI21X1 AOI21X1_240 ( .A(u0_u0__abc_72207_new_n398_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n399_), .Y(u0_u0__0csc_31_0__20_));
AOI21X1 AOI21X1_241 ( .A(u0_u0__abc_72207_new_n401_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n402_), .Y(u0_u0__0csc_31_0__21_));
AOI21X1 AOI21X1_242 ( .A(u0_u0__abc_72207_new_n404_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n405_), .Y(u0_u0__0csc_31_0__22_));
AOI21X1 AOI21X1_243 ( .A(u0_u0__abc_72207_new_n407_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n408_), .Y(u0_u0__0csc_31_0__23_));
AOI21X1 AOI21X1_244 ( .A(u0_u0__abc_72207_new_n410_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n411_), .Y(u0_u0__0csc_31_0__24_));
AOI21X1 AOI21X1_245 ( .A(u0_u0__abc_72207_new_n413_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n414_), .Y(u0_u0__0csc_31_0__25_));
AOI21X1 AOI21X1_246 ( .A(u0_u0__abc_72207_new_n416_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n417_), .Y(u0_u0__0csc_31_0__26_));
AOI21X1 AOI21X1_247 ( .A(u0_u0__abc_72207_new_n419_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n420_), .Y(u0_u0__0csc_31_0__27_));
AOI21X1 AOI21X1_248 ( .A(u0_u0__abc_72207_new_n422_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n423_), .Y(u0_u0__0csc_31_0__28_));
AOI21X1 AOI21X1_249 ( .A(u0_u0__abc_72207_new_n425_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n426_), .Y(u0_u0__0csc_31_0__29_));
AOI21X1 AOI21X1_25 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1392_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1393_));
AOI21X1 AOI21X1_250 ( .A(u0_u0__abc_72207_new_n428_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n429_), .Y(u0_u0__0csc_31_0__30_));
AOI21X1 AOI21X1_251 ( .A(u0_u0__abc_72207_new_n431_), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n432_), .Y(u0_u0__0csc_31_0__31_));
AOI21X1 AOI21X1_252 ( .A(u0_csc0_17_), .B(\wb_addr_i[22] ), .C(u0_u0__abc_72207_new_n441_), .Y(u0_u0__abc_72207_new_n442_));
AOI21X1 AOI21X1_253 ( .A(u0_csc0_8_), .B(wb_we_i), .C(u0_u0__abc_72207_new_n458_), .Y(u0_cs0));
AOI21X1 AOI21X1_254 ( .A(u0_u1__abc_72470_new_n219_), .B(u0_u1__abc_72470_new_n218_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__0_));
AOI21X1 AOI21X1_255 ( .A(u0_u1__abc_72470_new_n222_), .B(u0_u1__abc_72470_new_n221_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__1_));
AOI21X1 AOI21X1_256 ( .A(u0_u1__abc_72470_new_n225_), .B(u0_u1__abc_72470_new_n224_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__2_));
AOI21X1 AOI21X1_257 ( .A(u0_u1__abc_72470_new_n228_), .B(u0_u1__abc_72470_new_n227_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__3_));
AOI21X1 AOI21X1_258 ( .A(u0_u1__abc_72470_new_n231_), .B(u0_u1__abc_72470_new_n230_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__4_));
AOI21X1 AOI21X1_259 ( .A(u0_u1__abc_72470_new_n234_), .B(u0_u1__abc_72470_new_n233_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__5_));
AOI21X1 AOI21X1_26 ( .A(u0__abc_74894_new_n1407_), .B(u0__abc_74894_new_n1408_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1409_));
AOI21X1 AOI21X1_260 ( .A(u0_u1__abc_72470_new_n237_), .B(u0_u1__abc_72470_new_n236_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__6_));
AOI21X1 AOI21X1_261 ( .A(u0_u1__abc_72470_new_n240_), .B(u0_u1__abc_72470_new_n239_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__7_));
AOI21X1 AOI21X1_262 ( .A(u0_u1__abc_72470_new_n243_), .B(u0_u1__abc_72470_new_n242_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__8_));
AOI21X1 AOI21X1_263 ( .A(u0_u1__abc_72470_new_n246_), .B(u0_u1__abc_72470_new_n245_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__9_));
AOI21X1 AOI21X1_264 ( .A(u0_u1__abc_72470_new_n249_), .B(u0_u1__abc_72470_new_n248_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__10_));
AOI21X1 AOI21X1_265 ( .A(u0_u1__abc_72470_new_n252_), .B(u0_u1__abc_72470_new_n251_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__11_));
AOI21X1 AOI21X1_266 ( .A(u0_u1__abc_72470_new_n255_), .B(u0_u1__abc_72470_new_n254_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__12_));
AOI21X1 AOI21X1_267 ( .A(u0_u1__abc_72470_new_n258_), .B(u0_u1__abc_72470_new_n257_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__13_));
AOI21X1 AOI21X1_268 ( .A(u0_u1__abc_72470_new_n261_), .B(u0_u1__abc_72470_new_n260_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__14_));
AOI21X1 AOI21X1_269 ( .A(u0_u1__abc_72470_new_n264_), .B(u0_u1__abc_72470_new_n263_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__15_));
AOI21X1 AOI21X1_27 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1412_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1413_));
AOI21X1 AOI21X1_270 ( .A(u0_u1__abc_72470_new_n267_), .B(u0_u1__abc_72470_new_n266_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__16_));
AOI21X1 AOI21X1_271 ( .A(u0_u1__abc_72470_new_n270_), .B(u0_u1__abc_72470_new_n269_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__17_));
AOI21X1 AOI21X1_272 ( .A(u0_u1__abc_72470_new_n273_), .B(u0_u1__abc_72470_new_n272_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__18_));
AOI21X1 AOI21X1_273 ( .A(u0_u1__abc_72470_new_n276_), .B(u0_u1__abc_72470_new_n275_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__19_));
AOI21X1 AOI21X1_274 ( .A(u0_u1__abc_72470_new_n279_), .B(u0_u1__abc_72470_new_n278_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__20_));
AOI21X1 AOI21X1_275 ( .A(u0_u1__abc_72470_new_n282_), .B(u0_u1__abc_72470_new_n281_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__21_));
AOI21X1 AOI21X1_276 ( .A(u0_u1__abc_72470_new_n285_), .B(u0_u1__abc_72470_new_n284_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__22_));
AOI21X1 AOI21X1_277 ( .A(u0_u1__abc_72470_new_n288_), .B(u0_u1__abc_72470_new_n287_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__23_));
AOI21X1 AOI21X1_278 ( .A(u0_u1__abc_72470_new_n291_), .B(u0_u1__abc_72470_new_n290_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__24_));
AOI21X1 AOI21X1_279 ( .A(u0_u1__abc_72470_new_n294_), .B(u0_u1__abc_72470_new_n293_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__25_));
AOI21X1 AOI21X1_28 ( .A(u0__abc_74894_new_n1427_), .B(u0__abc_74894_new_n1428_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1429_));
AOI21X1 AOI21X1_280 ( .A(u0_u1__abc_72470_new_n297_), .B(u0_u1__abc_72470_new_n296_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__26_));
AOI21X1 AOI21X1_281 ( .A(u0_u1__abc_72470_new_n300_), .B(u0_u1__abc_72470_new_n299_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__27_));
AOI21X1 AOI21X1_282 ( .A(u0_u1__abc_72470_new_n303_), .B(u0_u1__abc_72470_new_n302_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__28_));
AOI21X1 AOI21X1_283 ( .A(u0_u1__abc_72470_new_n306_), .B(u0_u1__abc_72470_new_n305_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__29_));
AOI21X1 AOI21X1_284 ( .A(u0_u1__abc_72470_new_n309_), .B(u0_u1__abc_72470_new_n308_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__30_));
AOI21X1 AOI21X1_285 ( .A(u0_u1__abc_72470_new_n312_), .B(u0_u1__abc_72470_new_n311_), .C(u0_u1_rst_r2), .Y(u0_u1__0tms_31_0__31_));
AOI21X1 AOI21X1_286 ( .A(u0_u1__abc_72470_new_n316_), .B(u0_u1__abc_72470_new_n315_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__0_));
AOI21X1 AOI21X1_287 ( .A(u0_u1__abc_72470_new_n319_), .B(u0_u1__abc_72470_new_n318_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__1_));
AOI21X1 AOI21X1_288 ( .A(u0_u1__abc_72470_new_n322_), .B(u0_u1__abc_72470_new_n321_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__2_));
AOI21X1 AOI21X1_289 ( .A(u0_u1__abc_72470_new_n325_), .B(u0_u1__abc_72470_new_n324_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__3_));
AOI21X1 AOI21X1_29 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1432_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1433_));
AOI21X1 AOI21X1_290 ( .A(u0_u1__abc_72470_new_n328_), .B(u0_u1__abc_72470_new_n327_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__4_));
AOI21X1 AOI21X1_291 ( .A(u0_u1__abc_72470_new_n331_), .B(u0_u1__abc_72470_new_n330_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__5_));
AOI21X1 AOI21X1_292 ( .A(u0_u1__abc_72470_new_n334_), .B(u0_u1__abc_72470_new_n333_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__6_));
AOI21X1 AOI21X1_293 ( .A(u0_u1__abc_72470_new_n337_), .B(u0_u1__abc_72470_new_n336_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__7_));
AOI21X1 AOI21X1_294 ( .A(u0_u1__abc_72470_new_n340_), .B(u0_u1__abc_72470_new_n339_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__8_));
AOI21X1 AOI21X1_295 ( .A(u0_u1__abc_72470_new_n343_), .B(u0_u1__abc_72470_new_n342_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__9_));
AOI21X1 AOI21X1_296 ( .A(u0_u1__abc_72470_new_n346_), .B(u0_u1__abc_72470_new_n345_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__10_));
AOI21X1 AOI21X1_297 ( .A(u0_u1__abc_72470_new_n349_), .B(u0_u1__abc_72470_new_n348_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__11_));
AOI21X1 AOI21X1_298 ( .A(u0_u1__abc_72470_new_n352_), .B(u0_u1__abc_72470_new_n351_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__12_));
AOI21X1 AOI21X1_299 ( .A(u0_u1__abc_72470_new_n355_), .B(u0_u1__abc_72470_new_n354_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__13_));
AOI21X1 AOI21X1_3 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1172_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1173_));
AOI21X1 AOI21X1_30 ( .A(u0__abc_74894_new_n1447_), .B(u0__abc_74894_new_n1448_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1449_));
AOI21X1 AOI21X1_300 ( .A(u0_u1__abc_72470_new_n358_), .B(u0_u1__abc_72470_new_n357_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__14_));
AOI21X1 AOI21X1_301 ( .A(u0_u1__abc_72470_new_n361_), .B(u0_u1__abc_72470_new_n360_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__15_));
AOI21X1 AOI21X1_302 ( .A(u0_u1__abc_72470_new_n364_), .B(u0_u1__abc_72470_new_n363_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__16_));
AOI21X1 AOI21X1_303 ( .A(u0_u1__abc_72470_new_n367_), .B(u0_u1__abc_72470_new_n366_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__17_));
AOI21X1 AOI21X1_304 ( .A(u0_u1__abc_72470_new_n370_), .B(u0_u1__abc_72470_new_n369_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__18_));
AOI21X1 AOI21X1_305 ( .A(u0_u1__abc_72470_new_n373_), .B(u0_u1__abc_72470_new_n372_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__19_));
AOI21X1 AOI21X1_306 ( .A(u0_u1__abc_72470_new_n376_), .B(u0_u1__abc_72470_new_n375_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__20_));
AOI21X1 AOI21X1_307 ( .A(u0_u1__abc_72470_new_n379_), .B(u0_u1__abc_72470_new_n378_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__21_));
AOI21X1 AOI21X1_308 ( .A(u0_u1__abc_72470_new_n382_), .B(u0_u1__abc_72470_new_n381_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__22_));
AOI21X1 AOI21X1_309 ( .A(u0_u1__abc_72470_new_n385_), .B(u0_u1__abc_72470_new_n384_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__23_));
AOI21X1 AOI21X1_31 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1452_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1453_));
AOI21X1 AOI21X1_310 ( .A(u0_u1__abc_72470_new_n388_), .B(u0_u1__abc_72470_new_n387_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__24_));
AOI21X1 AOI21X1_311 ( .A(u0_u1__abc_72470_new_n391_), .B(u0_u1__abc_72470_new_n390_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__25_));
AOI21X1 AOI21X1_312 ( .A(u0_u1__abc_72470_new_n394_), .B(u0_u1__abc_72470_new_n393_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__26_));
AOI21X1 AOI21X1_313 ( .A(u0_u1__abc_72470_new_n397_), .B(u0_u1__abc_72470_new_n396_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__27_));
AOI21X1 AOI21X1_314 ( .A(u0_u1__abc_72470_new_n400_), .B(u0_u1__abc_72470_new_n399_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__28_));
AOI21X1 AOI21X1_315 ( .A(u0_u1__abc_72470_new_n403_), .B(u0_u1__abc_72470_new_n402_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__29_));
AOI21X1 AOI21X1_316 ( .A(u0_u1__abc_72470_new_n406_), .B(u0_u1__abc_72470_new_n405_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__30_));
AOI21X1 AOI21X1_317 ( .A(u0_u1__abc_72470_new_n409_), .B(u0_u1__abc_72470_new_n408_), .C(u0_u1_rst_r2), .Y(u0_u1__0csc_31_0__31_));
AOI21X1 AOI21X1_318 ( .A(u0_csc_mask_1_), .B(u0_u1__abc_72470_new_n418_), .C(u0_u1__abc_72470_new_n423_), .Y(u0_u1__abc_72470_new_n424_));
AOI21X1 AOI21X1_319 ( .A(u0_csc1_8_), .B(wb_we_i), .C(u0_u1__abc_72470_new_n434_), .Y(u0_cs1));
AOI21X1 AOI21X1_32 ( .A(u0__abc_74894_new_n1467_), .B(u0__abc_74894_new_n1468_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1469_));
AOI21X1 AOI21X1_320 ( .A(\wb_addr_i[22] ), .B(u1__abc_72801_new_n299_), .C(u1__abc_72801_new_n302_), .Y(u1__abc_72801_new_n303_));
AOI21X1 AOI21X1_321 ( .A(u1__abc_72801_new_n297_), .B(\wb_addr_i[25] ), .C(u1__abc_72801_new_n317_), .Y(u1__abc_72801_new_n318_));
AOI21X1 AOI21X1_322 ( .A(\wb_addr_i[22] ), .B(u1__abc_72801_new_n289_), .C(u1__abc_72801_new_n434_), .Y(u1__abc_72801_new_n435_));
AOI21X1 AOI21X1_323 ( .A(u1__abc_72801_new_n280_), .B(\wb_addr_i[1] ), .C(u1__abc_72801_new_n491_), .Y(u1__abc_72801_new_n494_));
AOI21X1 AOI21X1_324 ( .A(\wb_addr_i[0] ), .B(u1__abc_72801_new_n493_), .C(u1__abc_72801_new_n495_), .Y(u1__abc_72801_new_n496_));
AOI21X1 AOI21X1_325 ( .A(u1__abc_72801_new_n491_), .B(u1__abc_72801_new_n492_), .C(u1__abc_72801_new_n496_), .Y(u1__0acs_addr_23_0__0_));
AOI21X1 AOI21X1_326 ( .A(u1__abc_72801_new_n292_), .B(\wb_addr_i[16] ), .C(u1__abc_72801_new_n491_), .Y(u1__abc_72801_new_n569_));
AOI21X1 AOI21X1_327 ( .A(\wb_addr_i[14] ), .B(u1__abc_72801_new_n493_), .C(u1__abc_72801_new_n570_), .Y(u1__abc_72801_new_n571_));
AOI21X1 AOI21X1_328 ( .A(u1__abc_72801_new_n491_), .B(u1__abc_72801_new_n568_), .C(u1__abc_72801_new_n571_), .Y(u1__0acs_addr_23_0__14_));
AOI21X1 AOI21X1_329 ( .A(u1__abc_72801_new_n493_), .B(\wb_addr_i[20] ), .C(u1__abc_72801_new_n602_), .Y(u1__abc_72801_new_n603_));
AOI21X1 AOI21X1_33 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1472_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1473_));
AOI21X1 AOI21X1_330 ( .A(wb_stb_i), .B(u1__abc_72801_new_n460_), .C(u1__abc_72801_new_n620_), .Y(u1__0sram_addr_23_0__0_));
AOI21X1 AOI21X1_331 ( .A(wb_stb_i), .B(u1__abc_72801_new_n464_), .C(u1__abc_72801_new_n622_), .Y(u1__0sram_addr_23_0__1_));
AOI21X1 AOI21X1_332 ( .A(wb_stb_i), .B(u1__abc_72801_new_n467_), .C(u1__abc_72801_new_n624_), .Y(u1__0sram_addr_23_0__2_));
AOI21X1 AOI21X1_333 ( .A(wb_stb_i), .B(u1__abc_72801_new_n470_), .C(u1__abc_72801_new_n626_), .Y(u1__0sram_addr_23_0__3_));
AOI21X1 AOI21X1_334 ( .A(wb_stb_i), .B(u1__abc_72801_new_n473_), .C(u1__abc_72801_new_n628_), .Y(u1__0sram_addr_23_0__4_));
AOI21X1 AOI21X1_335 ( .A(wb_stb_i), .B(u1__abc_72801_new_n476_), .C(u1__abc_72801_new_n630_), .Y(u1__0sram_addr_23_0__5_));
AOI21X1 AOI21X1_336 ( .A(wb_stb_i), .B(u1__abc_72801_new_n479_), .C(u1__abc_72801_new_n632_), .Y(u1__0sram_addr_23_0__6_));
AOI21X1 AOI21X1_337 ( .A(wb_stb_i), .B(u1__abc_72801_new_n482_), .C(u1__abc_72801_new_n634_), .Y(u1__0sram_addr_23_0__7_));
AOI21X1 AOI21X1_338 ( .A(u1__abc_72801_new_n537_), .B(wb_stb_i), .C(u1__abc_72801_new_n636_), .Y(u1__0sram_addr_23_0__8_));
AOI21X1 AOI21X1_339 ( .A(u1__abc_72801_new_n543_), .B(wb_stb_i), .C(u1__abc_72801_new_n638_), .Y(u1__0sram_addr_23_0__9_));
AOI21X1 AOI21X1_34 ( .A(u0__abc_74894_new_n1487_), .B(u0__abc_74894_new_n1488_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1489_));
AOI21X1 AOI21X1_340 ( .A(u1__abc_72801_new_n277_), .B(wb_stb_i), .C(u1__abc_72801_new_n640_), .Y(u1__0sram_addr_23_0__10_));
AOI21X1 AOI21X1_341 ( .A(u1__abc_72801_new_n308_), .B(wb_stb_i), .C(u1__abc_72801_new_n642_), .Y(u1__0sram_addr_23_0__11_));
AOI21X1 AOI21X1_342 ( .A(u1__abc_72801_new_n324_), .B(wb_stb_i), .C(u1__abc_72801_new_n644_), .Y(u1__0sram_addr_23_0__12_));
AOI21X1 AOI21X1_343 ( .A(u1__abc_72801_new_n332_), .B(wb_stb_i), .C(u1__abc_72801_new_n646_), .Y(u1__0sram_addr_23_0__13_));
AOI21X1 AOI21X1_344 ( .A(u1__abc_72801_new_n399_), .B(wb_stb_i), .C(u1__abc_72801_new_n657_), .Y(u1__0sram_addr_23_0__17_));
AOI21X1 AOI21X1_345 ( .A(u1__abc_72801_new_n408_), .B(wb_stb_i), .C(u1__abc_72801_new_n659_), .Y(u1__0sram_addr_23_0__18_));
AOI21X1 AOI21X1_346 ( .A(u1__abc_72801_new_n300_), .B(wb_stb_i), .C(u1__abc_72801_new_n661_), .Y(u1__0sram_addr_23_0__19_));
AOI21X1 AOI21X1_347 ( .A(u1__abc_72801_new_n422_), .B(wb_stb_i), .C(u1__abc_72801_new_n663_), .Y(u1__0sram_addr_23_0__20_));
AOI21X1 AOI21X1_348 ( .A(u1__abc_72801_new_n423_), .B(wb_stb_i), .C(u1__abc_72801_new_n665_), .Y(u1__0sram_addr_23_0__21_));
AOI21X1 AOI21X1_349 ( .A(u1__abc_72801_new_n432_), .B(wb_stb_i), .C(u1__abc_72801_new_n667_), .Y(u1__0sram_addr_23_0__22_));
AOI21X1 AOI21X1_35 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1492_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1493_));
AOI21X1 AOI21X1_350 ( .A(u1__abc_72801_new_n287_), .B(wb_stb_i), .C(u1__abc_72801_new_n669_), .Y(u1__0sram_addr_23_0__23_));
AOI21X1 AOI21X1_351 ( .A(u1__abc_72801_new_n791_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n792_), .Y(mc_addr_d_15_));
AOI21X1 AOI21X1_352 ( .A(u1__abc_72801_new_n795_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n796_), .Y(mc_addr_d_16_));
AOI21X1 AOI21X1_353 ( .A(u1__abc_72801_new_n798_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n799_), .Y(mc_addr_d_17_));
AOI21X1 AOI21X1_354 ( .A(u1__abc_72801_new_n801_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n802_), .Y(mc_addr_d_18_));
AOI21X1 AOI21X1_355 ( .A(u1__abc_72801_new_n804_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n805_), .Y(mc_addr_d_19_));
AOI21X1 AOI21X1_356 ( .A(u1__abc_72801_new_n807_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n808_), .Y(mc_addr_d_20_));
AOI21X1 AOI21X1_357 ( .A(u1__abc_72801_new_n810_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n811_), .Y(mc_addr_d_21_));
AOI21X1 AOI21X1_358 ( .A(u1__abc_72801_new_n813_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n814_), .Y(mc_addr_d_22_));
AOI21X1 AOI21X1_359 ( .A(u1__abc_72801_new_n816_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n817_), .Y(mc_addr_d_23_));
AOI21X1 AOI21X1_36 ( .A(u0__abc_74894_new_n1507_), .B(u0__abc_74894_new_n1508_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1509_));
AOI21X1 AOI21X1_360 ( .A(u1__abc_72801_new_n825_), .B(u1__abc_72801_new_n672_), .C(rfr_ack), .Y(u1__abc_72801_new_n826_));
AOI21X1 AOI21X1_361 ( .A(u1_u0__abc_72719_new_n58_), .B(u1_acs_addr_4_), .C(u1_acs_addr_5_), .Y(u1_u0__abc_72719_new_n60_));
AOI21X1 AOI21X1_362 ( .A(u1_u0__abc_72719_new_n100_), .B(u1_acs_addr_16_), .C(u1_acs_addr_17_), .Y(u1_u0__abc_72719_new_n102_));
AOI21X1 AOI21X1_363 ( .A(u1_u0__abc_72719_new_n104_), .B(u1_acs_addr_18_), .C(u1_acs_addr_19_), .Y(u1_u0__abc_72719_new_n107_));
AOI21X1 AOI21X1_364 ( .A(u1_u0__abc_72719_new_n100_), .B(u1_u0__abc_72719_new_n109_), .C(u1_u0__abc_72719_new_n107_), .Y(u1_acs_addr_pl1_19_));
AOI21X1 AOI21X1_365 ( .A(u2_u0__abc_73914_new_n266_), .B(row_adr_8_), .C(u2_u0__abc_73914_new_n268_), .Y(u2_u0__abc_73914_new_n269_));
AOI21X1 AOI21X1_366 ( .A(u2_u0__abc_73914_new_n275_), .B(row_adr_1_), .C(u2_u0__abc_73914_new_n137_), .Y(u2_u0__abc_73914_new_n276_));
AOI21X1 AOI21X1_367 ( .A(u2_u0__abc_73914_new_n136_), .B(u2_u0_b1_last_row_0_), .C(u2_u0__abc_73914_new_n298_), .Y(u2_u0__abc_73914_new_n299_));
AOI21X1 AOI21X1_368 ( .A(u2_u0__abc_73914_new_n300_), .B(u2_u0__abc_73914_new_n301_), .C(u2_u0__abc_73914_new_n303_), .Y(u2_u0__abc_73914_new_n304_));
AOI21X1 AOI21X1_369 ( .A(u2_u0__abc_73914_new_n173_), .B(u2_u0_b1_last_row_11_), .C(u2_u0__abc_73914_new_n209_), .Y(u2_u0__abc_73914_new_n312_));
AOI21X1 AOI21X1_37 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1512_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1513_));
AOI21X1 AOI21X1_370 ( .A(u2_u0__abc_73914_new_n164_), .B(u2_u0_b0_last_row_8_), .C(u2_u0__abc_73914_new_n179_), .Y(u2_u0__abc_73914_new_n352_));
AOI21X1 AOI21X1_371 ( .A(u2_u0__abc_73914_new_n164_), .B(u2_u0_b2_last_row_8_), .C(u2_u0__abc_73914_new_n365_), .Y(u2_u0__abc_73914_new_n366_));
AOI21X1 AOI21X1_372 ( .A(u2_u0__abc_73914_new_n372_), .B(u2_u0__abc_73914_new_n373_), .C(u2_u0__abc_73914_new_n375_), .Y(u2_u0__abc_73914_new_n376_));
AOI21X1 AOI21X1_373 ( .A(u2_u0__abc_73914_new_n377_), .B(u2_u0__abc_73914_new_n378_), .C(u2_u0__abc_73914_new_n380_), .Y(u2_u0__abc_73914_new_n381_));
AOI21X1 AOI21X1_374 ( .A(u2_u1__abc_73914_new_n266_), .B(row_adr_8_), .C(u2_u1__abc_73914_new_n268_), .Y(u2_u1__abc_73914_new_n269_));
AOI21X1 AOI21X1_375 ( .A(u2_u1__abc_73914_new_n275_), .B(row_adr_1_), .C(u2_u1__abc_73914_new_n137_), .Y(u2_u1__abc_73914_new_n276_));
AOI21X1 AOI21X1_376 ( .A(u2_u1__abc_73914_new_n136_), .B(u2_u1_b1_last_row_0_), .C(u2_u1__abc_73914_new_n298_), .Y(u2_u1__abc_73914_new_n299_));
AOI21X1 AOI21X1_377 ( .A(u2_u1__abc_73914_new_n300_), .B(u2_u1__abc_73914_new_n301_), .C(u2_u1__abc_73914_new_n303_), .Y(u2_u1__abc_73914_new_n304_));
AOI21X1 AOI21X1_378 ( .A(u2_u1__abc_73914_new_n173_), .B(u2_u1_b1_last_row_11_), .C(u2_u1__abc_73914_new_n209_), .Y(u2_u1__abc_73914_new_n312_));
AOI21X1 AOI21X1_379 ( .A(u2_u1__abc_73914_new_n164_), .B(u2_u1_b0_last_row_8_), .C(u2_u1__abc_73914_new_n179_), .Y(u2_u1__abc_73914_new_n352_));
AOI21X1 AOI21X1_38 ( .A(u0__abc_74894_new_n1527_), .B(u0__abc_74894_new_n1528_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1529_));
AOI21X1 AOI21X1_380 ( .A(u2_u1__abc_73914_new_n164_), .B(u2_u1_b2_last_row_8_), .C(u2_u1__abc_73914_new_n365_), .Y(u2_u1__abc_73914_new_n366_));
AOI21X1 AOI21X1_381 ( .A(u2_u1__abc_73914_new_n372_), .B(u2_u1__abc_73914_new_n373_), .C(u2_u1__abc_73914_new_n375_), .Y(u2_u1__abc_73914_new_n376_));
AOI21X1 AOI21X1_382 ( .A(u2_u1__abc_73914_new_n377_), .B(u2_u1__abc_73914_new_n378_), .C(u2_u1__abc_73914_new_n380_), .Y(u2_u1__abc_73914_new_n381_));
AOI21X1 AOI21X1_383 ( .A(u3__abc_73372_new_n315_), .B(pack_le2), .C(u3__abc_73372_new_n316_), .Y(u3__0byte2_7_0__0_));
AOI21X1 AOI21X1_384 ( .A(pack_le2), .B(u3__abc_73372_new_n318_), .C(u3__abc_73372_new_n319_), .Y(u3__0byte2_7_0__1_));
AOI21X1 AOI21X1_385 ( .A(pack_le2), .B(u3__abc_73372_new_n321_), .C(u3__abc_73372_new_n322_), .Y(u3__0byte2_7_0__2_));
AOI21X1 AOI21X1_386 ( .A(pack_le2), .B(u3__abc_73372_new_n324_), .C(u3__abc_73372_new_n325_), .Y(u3__0byte2_7_0__3_));
AOI21X1 AOI21X1_387 ( .A(pack_le2), .B(u3__abc_73372_new_n327_), .C(u3__abc_73372_new_n328_), .Y(u3__0byte2_7_0__4_));
AOI21X1 AOI21X1_388 ( .A(pack_le2), .B(u3__abc_73372_new_n330_), .C(u3__abc_73372_new_n331_), .Y(u3__0byte2_7_0__5_));
AOI21X1 AOI21X1_389 ( .A(pack_le2), .B(u3__abc_73372_new_n333_), .C(u3__abc_73372_new_n334_), .Y(u3__0byte2_7_0__6_));
AOI21X1 AOI21X1_39 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1532_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1533_));
AOI21X1 AOI21X1_390 ( .A(pack_le2), .B(u3__abc_73372_new_n336_), .C(u3__abc_73372_new_n337_), .Y(u3__0byte2_7_0__7_));
AOI21X1 AOI21X1_391 ( .A(u3__abc_73372_new_n315_), .B(pack_le0), .C(u3__abc_73372_new_n386_), .Y(u3__0byte0_7_0__0_));
AOI21X1 AOI21X1_392 ( .A(u3__abc_73372_new_n318_), .B(pack_le0), .C(u3__abc_73372_new_n388_), .Y(u3__0byte0_7_0__1_));
AOI21X1 AOI21X1_393 ( .A(u3__abc_73372_new_n321_), .B(pack_le0), .C(u3__abc_73372_new_n390_), .Y(u3__0byte0_7_0__2_));
AOI21X1 AOI21X1_394 ( .A(u3__abc_73372_new_n324_), .B(pack_le0), .C(u3__abc_73372_new_n392_), .Y(u3__0byte0_7_0__3_));
AOI21X1 AOI21X1_395 ( .A(u3__abc_73372_new_n327_), .B(pack_le0), .C(u3__abc_73372_new_n394_), .Y(u3__0byte0_7_0__4_));
AOI21X1 AOI21X1_396 ( .A(u3__abc_73372_new_n330_), .B(pack_le0), .C(u3__abc_73372_new_n396_), .Y(u3__0byte0_7_0__5_));
AOI21X1 AOI21X1_397 ( .A(u3__abc_73372_new_n333_), .B(pack_le0), .C(u3__abc_73372_new_n398_), .Y(u3__0byte0_7_0__6_));
AOI21X1 AOI21X1_398 ( .A(u3__abc_73372_new_n336_), .B(pack_le0), .C(u3__abc_73372_new_n400_), .Y(u3__0byte0_7_0__7_));
AOI21X1 AOI21X1_399 ( .A(u3__abc_73372_new_n339_), .B(u3_byte2_0_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n564_));
AOI21X1 AOI21X1_4 ( .A(u0__abc_74894_new_n1187_), .B(u0__abc_74894_new_n1188_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1189_));
AOI21X1 AOI21X1_40 ( .A(u0__abc_74894_new_n1547_), .B(u0__abc_74894_new_n1548_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1549_));
AOI21X1 AOI21X1_400 ( .A(u3__abc_73372_new_n339_), .B(u3_byte2_1_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n568_));
AOI21X1 AOI21X1_401 ( .A(u3__abc_73372_new_n339_), .B(u3_byte2_2_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n572_));
AOI21X1 AOI21X1_402 ( .A(u3__abc_73372_new_n339_), .B(u3_byte2_3_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n576_));
AOI21X1 AOI21X1_403 ( .A(u3__abc_73372_new_n339_), .B(u3_byte2_4_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n580_));
AOI21X1 AOI21X1_404 ( .A(u3__abc_73372_new_n339_), .B(u3_byte2_5_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n584_));
AOI21X1 AOI21X1_405 ( .A(u3__abc_73372_new_n339_), .B(u3_byte2_6_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n588_));
AOI21X1 AOI21X1_406 ( .A(u3__abc_73372_new_n339_), .B(u3_byte2_7_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n592_));
AOI21X1 AOI21X1_407 ( .A(u3__abc_73372_new_n339_), .B(mc_data_ir_0_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n596_));
AOI21X1 AOI21X1_408 ( .A(u3__abc_73372_new_n339_), .B(mc_data_ir_1_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n600_));
AOI21X1 AOI21X1_409 ( .A(u3__abc_73372_new_n339_), .B(mc_data_ir_2_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n604_));
AOI21X1 AOI21X1_41 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1552_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1553_));
AOI21X1 AOI21X1_410 ( .A(u3__abc_73372_new_n339_), .B(mc_data_ir_3_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n608_));
AOI21X1 AOI21X1_411 ( .A(u3__abc_73372_new_n339_), .B(mc_data_ir_4_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n612_));
AOI21X1 AOI21X1_412 ( .A(u3__abc_73372_new_n339_), .B(mc_data_ir_5_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n616_));
AOI21X1 AOI21X1_413 ( .A(u3__abc_73372_new_n339_), .B(mc_data_ir_6_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n620_));
AOI21X1 AOI21X1_414 ( .A(u3__abc_73372_new_n339_), .B(mc_data_ir_7_), .C(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n624_));
AOI21X1 AOI21X1_415 ( .A(u3__abc_73372_new_n646_), .B(u3__abc_73372_new_n643_), .C(u3__abc_73372_new_n648_), .Y(u3__abc_73372_new_n649_));
AOI21X1 AOI21X1_416 ( .A(u3__abc_73372_new_n653_), .B(u3__abc_73372_new_n654_), .C(u3__abc_73372_new_n652_), .Y(u3__abc_73372_new_n655_));
AOI21X1 AOI21X1_417 ( .A(u3__abc_73372_new_n656_), .B(u3__abc_73372_new_n657_), .C(u3_rd_fifo_out_34_), .Y(u3__abc_73372_new_n658_));
AOI21X1 AOI21X1_418 ( .A(u3__abc_73372_new_n697_), .B(u3__abc_73372_new_n698_), .C(u3__abc_73372_new_n696_), .Y(u3__abc_73372_new_n699_));
AOI21X1 AOI21X1_419 ( .A(u3__abc_73372_new_n703_), .B(u3__abc_73372_new_n704_), .C(u3__abc_73372_new_n702_), .Y(u3__abc_73372_new_n705_));
AOI21X1 AOI21X1_42 ( .A(u0__abc_74894_new_n1567_), .B(u0__abc_74894_new_n1568_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1569_));
AOI21X1 AOI21X1_420 ( .A(u3__abc_73372_new_n706_), .B(u3__abc_73372_new_n707_), .C(u3_rd_fifo_out_35_), .Y(u3__abc_73372_new_n708_));
AOI21X1 AOI21X1_421 ( .A(u3__abc_73372_new_n678_), .B(u3__abc_73372_new_n728_), .C(u3__abc_73372_new_n729_), .Y(par_err));
AOI21X1 AOI21X1_422 ( .A(u3_u0_rd_adr_3_), .B(u3_re), .C(u3_rd_fifo_clr), .Y(u3_u0__abc_74260_new_n638_));
AOI21X1 AOI21X1_423 ( .A(u3_u0__abc_74260_new_n640_), .B(u3_u0__abc_74260_new_n641_), .C(u3_u0__abc_74260_new_n643_), .Y(u3_u0__0rd_adr_3_0__1_));
AOI21X1 AOI21X1_424 ( .A(u3_u0__abc_74260_new_n640_), .B(u3_u0__abc_74260_new_n645_), .C(u3_u0__abc_74260_new_n646_), .Y(u3_u0__0rd_adr_3_0__2_));
AOI21X1 AOI21X1_425 ( .A(u3_u0__abc_74260_new_n648_), .B(u3_u0__abc_74260_new_n640_), .C(u3_u0__abc_74260_new_n649_), .Y(u3_u0__0rd_adr_3_0__3_));
AOI21X1 AOI21X1_426 ( .A(dv), .B(u3_u0_wr_adr_3_), .C(u3_rd_fifo_clr), .Y(u3_u0__abc_74260_new_n652_));
AOI21X1 AOI21X1_427 ( .A(u3_u0_wr_adr_1_), .B(u3_u0__abc_74260_new_n654_), .C(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n656_));
AOI21X1 AOI21X1_428 ( .A(u3_u0__abc_74260_new_n658_), .B(u3_u0__abc_74260_new_n383_), .C(u3_rd_fifo_clr), .Y(u3_u0__0wr_adr_3_0__2_));
AOI21X1 AOI21X1_429 ( .A(u3_u0__abc_74260_new_n660_), .B(u3_u0__abc_74260_new_n564_), .C(u3_rd_fifo_clr), .Y(u3_u0__0wr_adr_3_0__3_));
AOI21X1 AOI21X1_43 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1572_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1573_));
AOI21X1 AOI21X1_430 ( .A(u3_u0__abc_74260_new_n382_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n662_), .Y(u3_u0__0r0_35_0__0_));
AOI21X1 AOI21X1_431 ( .A(u3_u0__abc_74260_new_n386_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n664_), .Y(u3_u0__0r0_35_0__1_));
AOI21X1 AOI21X1_432 ( .A(u3_u0__abc_74260_new_n389_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n666_), .Y(u3_u0__0r0_35_0__2_));
AOI21X1 AOI21X1_433 ( .A(u3_u0__abc_74260_new_n392_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n668_), .Y(u3_u0__0r0_35_0__3_));
AOI21X1 AOI21X1_434 ( .A(u3_u0__abc_74260_new_n395_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n670_), .Y(u3_u0__0r0_35_0__4_));
AOI21X1 AOI21X1_435 ( .A(u3_u0__abc_74260_new_n398_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n672_), .Y(u3_u0__0r0_35_0__5_));
AOI21X1 AOI21X1_436 ( .A(u3_u0__abc_74260_new_n401_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n674_), .Y(u3_u0__0r0_35_0__6_));
AOI21X1 AOI21X1_437 ( .A(u3_u0__abc_74260_new_n404_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n676_), .Y(u3_u0__0r0_35_0__7_));
AOI21X1 AOI21X1_438 ( .A(u3_u0__abc_74260_new_n407_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n678_), .Y(u3_u0__0r0_35_0__8_));
AOI21X1 AOI21X1_439 ( .A(u3_u0__abc_74260_new_n410_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n680_), .Y(u3_u0__0r0_35_0__9_));
AOI21X1 AOI21X1_44 ( .A(u0__abc_74894_new_n1587_), .B(u0__abc_74894_new_n1588_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1589_));
AOI21X1 AOI21X1_440 ( .A(u3_u0__abc_74260_new_n413_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n682_), .Y(u3_u0__0r0_35_0__10_));
AOI21X1 AOI21X1_441 ( .A(u3_u0__abc_74260_new_n416_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n684_), .Y(u3_u0__0r0_35_0__11_));
AOI21X1 AOI21X1_442 ( .A(u3_u0__abc_74260_new_n419_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n686_), .Y(u3_u0__0r0_35_0__12_));
AOI21X1 AOI21X1_443 ( .A(u3_u0__abc_74260_new_n422_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n688_), .Y(u3_u0__0r0_35_0__13_));
AOI21X1 AOI21X1_444 ( .A(u3_u0__abc_74260_new_n425_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n690_), .Y(u3_u0__0r0_35_0__14_));
AOI21X1 AOI21X1_445 ( .A(u3_u0__abc_74260_new_n428_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n692_), .Y(u3_u0__0r0_35_0__15_));
AOI21X1 AOI21X1_446 ( .A(u3_u0__abc_74260_new_n431_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n694_), .Y(u3_u0__0r0_35_0__16_));
AOI21X1 AOI21X1_447 ( .A(u3_u0__abc_74260_new_n434_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n696_), .Y(u3_u0__0r0_35_0__17_));
AOI21X1 AOI21X1_448 ( .A(u3_u0__abc_74260_new_n437_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n698_), .Y(u3_u0__0r0_35_0__18_));
AOI21X1 AOI21X1_449 ( .A(u3_u0__abc_74260_new_n440_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n700_), .Y(u3_u0__0r0_35_0__19_));
AOI21X1 AOI21X1_45 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1592_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1593_));
AOI21X1 AOI21X1_450 ( .A(u3_u0__abc_74260_new_n443_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n702_), .Y(u3_u0__0r0_35_0__20_));
AOI21X1 AOI21X1_451 ( .A(u3_u0__abc_74260_new_n446_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n704_), .Y(u3_u0__0r0_35_0__21_));
AOI21X1 AOI21X1_452 ( .A(u3_u0__abc_74260_new_n449_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n706_), .Y(u3_u0__0r0_35_0__22_));
AOI21X1 AOI21X1_453 ( .A(u3_u0__abc_74260_new_n452_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n708_), .Y(u3_u0__0r0_35_0__23_));
AOI21X1 AOI21X1_454 ( .A(u3_u0__abc_74260_new_n455_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n710_), .Y(u3_u0__0r0_35_0__24_));
AOI21X1 AOI21X1_455 ( .A(u3_u0__abc_74260_new_n458_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n712_), .Y(u3_u0__0r0_35_0__25_));
AOI21X1 AOI21X1_456 ( .A(u3_u0__abc_74260_new_n461_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n714_), .Y(u3_u0__0r0_35_0__26_));
AOI21X1 AOI21X1_457 ( .A(u3_u0__abc_74260_new_n464_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n716_), .Y(u3_u0__0r0_35_0__27_));
AOI21X1 AOI21X1_458 ( .A(u3_u0__abc_74260_new_n467_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n718_), .Y(u3_u0__0r0_35_0__28_));
AOI21X1 AOI21X1_459 ( .A(u3_u0__abc_74260_new_n470_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n720_), .Y(u3_u0__0r0_35_0__29_));
AOI21X1 AOI21X1_46 ( .A(u0__abc_74894_new_n1607_), .B(u0__abc_74894_new_n1608_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1609_));
AOI21X1 AOI21X1_460 ( .A(u3_u0__abc_74260_new_n473_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n722_), .Y(u3_u0__0r0_35_0__30_));
AOI21X1 AOI21X1_461 ( .A(u3_u0__abc_74260_new_n476_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n724_), .Y(u3_u0__0r0_35_0__31_));
AOI21X1 AOI21X1_462 ( .A(u3_u0__abc_74260_new_n479_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n726_), .Y(u3_u0__0r0_35_0__32_));
AOI21X1 AOI21X1_463 ( .A(u3_u0__abc_74260_new_n482_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n728_), .Y(u3_u0__0r0_35_0__33_));
AOI21X1 AOI21X1_464 ( .A(u3_u0__abc_74260_new_n485_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n730_), .Y(u3_u0__0r0_35_0__34_));
AOI21X1 AOI21X1_465 ( .A(u3_u0__abc_74260_new_n488_), .B(u3_u0__abc_74260_new_n655_), .C(u3_u0__abc_74260_new_n732_), .Y(u3_u0__0r0_35_0__35_));
AOI21X1 AOI21X1_466 ( .A(u4_rfr_ce), .B(u4__abc_74770_new_n107_), .C(u4__abc_74770_new_n108_), .Y(u4__0rfr_cnt_7_0__3_));
AOI21X1 AOI21X1_467 ( .A(u4__abc_74770_new_n107_), .B(u4_rfr_ce), .C(u4_rfr_cnt_4_), .Y(u4__abc_74770_new_n110_));
AOI21X1 AOI21X1_468 ( .A(u4_rfr_cnt_5_), .B(u4__abc_74770_new_n112_), .C(u4__abc_74770_new_n115_), .Y(u4__0rfr_cnt_7_0__5_));
AOI21X1 AOI21X1_469 ( .A(u4__abc_74770_new_n117_), .B(u4__abc_74770_new_n118_), .C(u4__abc_74770_new_n119_), .Y(u4__0rfr_cnt_7_0__6_));
AOI21X1 AOI21X1_47 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1612_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1613_));
AOI21X1 AOI21X1_470 ( .A(u4__abc_74770_new_n121_), .B(u4__abc_74770_new_n125_), .C(rfr_ack), .Y(u4__0rfr_cnt_7_0__7_));
AOI21X1 AOI21X1_471 ( .A(u4__0rfr_early_0_0_), .B(u4__abc_74770_new_n132_), .C(u4__abc_74770_new_n142_), .Y(u4__0ps_cnt_7_0__1_));
AOI21X1 AOI21X1_472 ( .A(u4__0rfr_early_0_0_), .B(u4__abc_74770_new_n132_), .C(u4__abc_74770_new_n149_), .Y(u4__0ps_cnt_7_0__3_));
AOI21X1 AOI21X1_473 ( .A(u4__0rfr_early_0_0_), .B(u4__abc_74770_new_n132_), .C(u4__abc_74770_new_n152_), .Y(u4__0ps_cnt_7_0__4_));
AOI21X1 AOI21X1_474 ( .A(u4__0rfr_early_0_0_), .B(u4__abc_74770_new_n132_), .C(u4__abc_74770_new_n160_), .Y(u4__0ps_cnt_7_0__5_));
AOI21X1 AOI21X1_475 ( .A(u4__0rfr_early_0_0_), .B(u4__abc_74770_new_n132_), .C(u4__abc_74770_new_n170_), .Y(u4__0ps_cnt_7_0__7_));
AOI21X1 AOI21X1_476 ( .A(u4_rfr_cnt_7_), .B(ref_int_1_), .C(u4__abc_74770_new_n174_), .Y(u4__abc_74770_new_n183_));
AOI21X1 AOI21X1_477 ( .A(u4__abc_74770_new_n180_), .B(u4__abc_74770_new_n185_), .C(u4__abc_74770_new_n172_), .Y(u4__0rfr_clr_0_0_));
AOI21X1 AOI21X1_478 ( .A(u5__abc_78290_new_n828_), .B(u5__abc_78290_new_n834_), .C(u5__abc_78290_new_n454_), .Y(u5__abc_78290_new_n835_));
AOI21X1 AOI21X1_479 ( .A(u5__abc_78290_new_n707_), .B(u5__abc_78290_new_n714_), .C(u5__abc_78290_new_n671_), .Y(u5__abc_78290_new_n991_));
AOI21X1 AOI21X1_48 ( .A(u0__abc_74894_new_n1627_), .B(u0__abc_74894_new_n1628_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1629_));
AOI21X1 AOI21X1_480 ( .A(u5__abc_78290_new_n730_), .B(u5__abc_78290_new_n745_), .C(u5__abc_78290_new_n454_), .Y(u5__abc_78290_new_n1003_));
AOI21X1 AOI21X1_481 ( .A(u5__abc_78290_new_n775_), .B(u5__abc_78290_new_n631_), .C(u5__abc_78290_new_n454_), .Y(u5__abc_78290_new_n1008_));
AOI21X1 AOI21X1_482 ( .A(u5__abc_78290_new_n578_), .B(u5__abc_78290_new_n1013_), .C(u5__abc_78290_new_n570_), .Y(u5__abc_78290_new_n1014_));
AOI21X1 AOI21X1_483 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n797_), .C(u5__abc_78290_new_n574_), .Y(u5__abc_78290_new_n1016_));
AOI21X1 AOI21X1_484 ( .A(u5__abc_78290_new_n1028_), .B(rfr_ack), .C(u5__abc_78290_new_n1035_), .Y(u5__abc_78290_new_n1036_));
AOI21X1 AOI21X1_485 ( .A(u5__abc_78290_new_n1120_), .B(u5__abc_78290_new_n1123_), .C(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1124_));
AOI21X1 AOI21X1_486 ( .A(u5__abc_78290_new_n1152_), .B(u5__abc_78290_new_n1155_), .C(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1156_));
AOI21X1 AOI21X1_487 ( .A(u5__abc_78290_new_n1171_), .B(u5__abc_78290_new_n1174_), .C(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1175_));
AOI21X1 AOI21X1_488 ( .A(u5__abc_78290_new_n1178_), .B(u5__abc_78290_new_n1181_), .C(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1182_));
AOI21X1 AOI21X1_489 ( .A(u5__abc_78290_new_n1188_), .B(u5__abc_78290_new_n1189_), .C(u5__abc_78290_new_n1014_), .Y(u5__abc_78290_new_n1190_));
AOI21X1 AOI21X1_49 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1632_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1633_));
AOI21X1 AOI21X1_490 ( .A(u5__abc_78290_new_n1085_), .B(u5__abc_78290_new_n1136_), .C(u5__abc_78290_new_n1358_), .Y(u5__abc_78290_new_n1359_));
AOI21X1 AOI21X1_491 ( .A(u5__abc_78290_new_n1155_), .B(u5__abc_78290_new_n1174_), .C(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1388_));
AOI21X1 AOI21X1_492 ( .A(u5__abc_78290_new_n1413_), .B(u5__abc_78290_new_n1419_), .C(u5__abc_78290_new_n1408_), .Y(u5__abc_78290_new_n1420_));
AOI21X1 AOI21X1_493 ( .A(u5__abc_78290_new_n1407_), .B(u5__abc_78290_new_n1420_), .C(u5__abc_78290_new_n1403_), .Y(u5__abc_78290_new_n1421_));
AOI21X1 AOI21X1_494 ( .A(u5__abc_78290_new_n1455_), .B(u5__abc_78290_new_n1456_), .C(u5__abc_78290_new_n1493_), .Y(u5__abc_78290_new_n1494_));
AOI21X1 AOI21X1_495 ( .A(u5__abc_78290_new_n1501_), .B(u5__abc_78290_new_n1273_), .C(u5__abc_78290_new_n1502_), .Y(u5__abc_78290_new_n1503_));
AOI21X1 AOI21X1_496 ( .A(u5__abc_78290_new_n1488_), .B(u5__abc_78290_new_n1515_), .C(u5__abc_78290_new_n1519_), .Y(u5__abc_78290_new_n1520_));
AOI21X1 AOI21X1_497 ( .A(u5__abc_78290_new_n1627_), .B(u5__abc_78290_new_n1605_), .C(u5__0no_wb_cycle_0_0_), .Y(mem_ack));
AOI21X1 AOI21X1_498 ( .A(wb_stb_i), .B(u5_wb_first), .C(u5_wb_stb_first), .Y(u5__abc_78290_new_n1629_));
AOI21X1 AOI21X1_499 ( .A(u5__abc_78290_new_n1361_), .B(u5__abc_78290_new_n1392_), .C(u5__abc_78290_new_n1442_), .Y(u5__abc_78290_new_n1639_));
AOI21X1 AOI21X1_5 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1192_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1193_));
AOI21X1 AOI21X1_50 ( .A(u0__abc_74894_new_n1647_), .B(u0__abc_74894_new_n1648_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1649_));
AOI21X1 AOI21X1_500 ( .A(u5__abc_78290_new_n1670_), .B(u5__abc_78290_new_n1663_), .C(u5__abc_78290_new_n1649_), .Y(u5__0burst_cnt_10_0__0_));
AOI21X1 AOI21X1_501 ( .A(u5__abc_78290_new_n1673_), .B(u5__abc_78290_new_n367_), .C(u5__abc_78290_new_n1318_), .Y(u5__abc_78290_new_n1674_));
AOI21X1 AOI21X1_502 ( .A(u5__abc_78290_new_n1672_), .B(u5__abc_78290_new_n1674_), .C(u5__abc_78290_new_n1677_), .Y(u5__0burst_cnt_10_0__1_));
AOI21X1 AOI21X1_503 ( .A(u5__abc_78290_new_n1673_), .B(u5__abc_78290_new_n367_), .C(u5__abc_78290_new_n366_), .Y(u5__abc_78290_new_n1680_));
AOI21X1 AOI21X1_504 ( .A(u5__abc_78290_new_n1679_), .B(u5__abc_78290_new_n1673_), .C(u5__abc_78290_new_n1680_), .Y(u5__abc_78290_new_n1681_));
AOI21X1 AOI21X1_505 ( .A(u5__abc_78290_new_n1654_), .B(1'h0), .C(u5__abc_78290_new_n1682_), .Y(u5__abc_78290_new_n1683_));
AOI21X1 AOI21X1_506 ( .A(u5__abc_78290_new_n1673_), .B(u5__abc_78290_new_n369_), .C(u5__abc_78290_new_n1318_), .Y(u5__abc_78290_new_n1686_));
AOI21X1 AOI21X1_507 ( .A(u5__abc_78290_new_n1686_), .B(u5__abc_78290_new_n1685_), .C(u5__abc_78290_new_n1690_), .Y(u5__0burst_cnt_10_0__3_));
AOI21X1 AOI21X1_508 ( .A(u5__abc_78290_new_n1673_), .B(u5__abc_78290_new_n369_), .C(u5__abc_78290_new_n1692_), .Y(u5__abc_78290_new_n1693_));
AOI21X1 AOI21X1_509 ( .A(u5__abc_78290_new_n1696_), .B(u5__abc_78290_new_n1697_), .C(u5__abc_78290_new_n1649_), .Y(u5__0burst_cnt_10_0__4_));
AOI21X1 AOI21X1_51 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1652_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1653_));
AOI21X1 AOI21X1_510 ( .A(u5__abc_78290_new_n1694_), .B(u5_burst_cnt_5_), .C(u5__abc_78290_new_n1318_), .Y(u5__abc_78290_new_n1701_));
AOI21X1 AOI21X1_511 ( .A(u5__abc_78290_new_n1700_), .B(u5__abc_78290_new_n1701_), .C(u5__abc_78290_new_n1703_), .Y(u5__0burst_cnt_10_0__5_));
AOI21X1 AOI21X1_512 ( .A(u5__abc_78290_new_n1707_), .B(u5__abc_78290_new_n1705_), .C(u5__abc_78290_new_n1709_), .Y(u5__0burst_cnt_10_0__6_));
AOI21X1 AOI21X1_513 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n1864_), .C(u5__abc_78290_new_n1862_), .Y(u5__abc_78290_new_n1865_));
AOI21X1 AOI21X1_514 ( .A(u5__abc_78290_new_n1160_), .B(u5__abc_78290_new_n1868_), .C(u5__abc_78290_new_n685_), .Y(u5__abc_78290_new_n1869_));
AOI21X1 AOI21X1_515 ( .A(u5__abc_78290_new_n1878_), .B(u5__abc_78290_new_n1879_), .C(u5__abc_78290_new_n685_), .Y(u5__abc_78290_new_n1880_));
AOI21X1 AOI21X1_516 ( .A(u5__abc_78290_new_n1899_), .B(u5__abc_78290_new_n1902_), .C(u5__abc_78290_new_n685_), .Y(u5__abc_78290_new_n1903_));
AOI21X1 AOI21X1_517 ( .A(u5__abc_78290_new_n1918_), .B(u5__abc_78290_new_n1921_), .C(u5__abc_78290_new_n685_), .Y(u5__abc_78290_new_n1922_));
AOI21X1 AOI21X1_518 ( .A(u5__abc_78290_new_n1933_), .B(u5__abc_78290_new_n1936_), .C(u5__abc_78290_new_n685_), .Y(u5__abc_78290_new_n1937_));
AOI21X1 AOI21X1_519 ( .A(u5__abc_78290_new_n1955_), .B(u5__abc_78290_new_n1952_), .C(u5__abc_78290_new_n1957_), .Y(u5__0burst_cnt_10_0__7_));
AOI21X1 AOI21X1_52 ( .A(u0__abc_74894_new_n1667_), .B(u0__abc_74894_new_n1668_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1669_));
AOI21X1 AOI21X1_520 ( .A(u5__abc_78290_new_n1962_), .B(u5__abc_78290_new_n1961_), .C(u5__abc_78290_new_n1318_), .Y(u5__abc_78290_new_n1963_));
AOI21X1 AOI21X1_521 ( .A(u5__abc_78290_new_n1963_), .B(u5__abc_78290_new_n1960_), .C(u5__abc_78290_new_n1965_), .Y(u5__0burst_cnt_10_0__8_));
AOI21X1 AOI21X1_522 ( .A(u5__abc_78290_new_n1971_), .B(u5__abc_78290_new_n1952_), .C(u5__abc_78290_new_n1973_), .Y(u5__0burst_cnt_10_0__9_));
AOI21X1 AOI21X1_523 ( .A(u5__abc_78290_new_n1978_), .B(u5__abc_78290_new_n1317_), .C(u5__abc_78290_new_n1980_), .Y(u5__0burst_cnt_10_0__10_));
AOI21X1 AOI21X1_524 ( .A(u5__abc_78290_new_n2004_), .B(u5__abc_78290_new_n2003_), .C(u5__abc_78290_new_n2011_), .Y(u5__0ir_cnt_3_0__0_));
AOI21X1 AOI21X1_525 ( .A(u5__abc_78290_new_n2003_), .B(u5_ir_cnt_1_), .C(u5__abc_78290_new_n2011_), .Y(u5__abc_78290_new_n2013_));
AOI21X1 AOI21X1_526 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n815_), .C(u5__abc_78290_new_n2052_), .Y(u5__abc_78290_new_n2053_));
AOI21X1 AOI21X1_527 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n791_), .C(u5__abc_78290_new_n574_), .Y(u5__abc_78290_new_n2061_));
AOI21X1 AOI21X1_528 ( .A(u5_mc_le), .B(u5_timer_0_), .C(u5__abc_78290_new_n2085_), .Y(u5__abc_78290_new_n2086_));
AOI21X1 AOI21X1_529 ( .A(u5__abc_78290_new_n2132_), .B(u5__abc_78290_new_n2034_), .C(u5__abc_78290_new_n2142_), .Y(u5__abc_78290_new_n2143_));
AOI21X1 AOI21X1_53 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1672_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1673_));
AOI21X1 AOI21X1_530 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n945_), .C(u5__abc_78290_new_n1433_), .Y(u5__abc_78290_new_n2160_));
AOI21X1 AOI21X1_531 ( .A(u5__abc_78290_new_n2189_), .B(u5__abc_78290_new_n2168_), .C(u5__abc_78290_new_n2211_), .Y(u5__abc_78290_new_n2212_));
AOI21X1 AOI21X1_532 ( .A(u5__abc_78290_new_n2243_), .B(u5__abc_78290_new_n2034_), .C(u5__abc_78290_new_n2246_), .Y(u5__abc_78290_new_n2247_));
AOI21X1 AOI21X1_533 ( .A(u5__abc_78290_new_n2249_), .B(u5__abc_78290_new_n2244_), .C(u5__abc_78290_new_n2251_), .Y(u5__abc_78290_new_n2252_));
AOI21X1 AOI21X1_534 ( .A(u5__abc_78290_new_n2252_), .B(u5__abc_78290_new_n2248_), .C(u5__abc_78290_new_n2141_), .Y(u5__abc_78290_new_n2253_));
AOI21X1 AOI21X1_535 ( .A(u5__abc_78290_new_n2189_), .B(u5__abc_78290_new_n2256_), .C(u5__abc_78290_new_n2211_), .Y(u5__abc_78290_new_n2257_));
AOI21X1 AOI21X1_536 ( .A(u5__abc_78290_new_n2252_), .B(u5__abc_78290_new_n2248_), .C(u5__abc_78290_new_n2251_), .Y(u5__abc_78290_new_n2272_));
AOI21X1 AOI21X1_537 ( .A(u5__abc_78290_new_n1472_), .B(u5__abc_78290_new_n2130_), .C(u5__abc_78290_new_n2033_), .Y(u5__abc_78290_new_n2275_));
AOI21X1 AOI21X1_538 ( .A(u5__abc_78290_new_n2291_), .B(u5__abc_78290_new_n2295_), .C(u5__abc_78290_new_n2293_), .Y(u5__abc_78290_new_n2296_));
AOI21X1 AOI21X1_539 ( .A(u5__abc_78290_new_n2033_), .B(u5__abc_78290_new_n2264_), .C(u5__abc_78290_new_n2140_), .Y(u5__abc_78290_new_n2299_));
AOI21X1 AOI21X1_54 ( .A(u0__abc_74894_new_n1687_), .B(u0__abc_74894_new_n1688_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1689_));
AOI21X1 AOI21X1_540 ( .A(u5__abc_78290_new_n2211_), .B(u5__abc_78290_new_n2304_), .C(u5__abc_78290_new_n2223_), .Y(u5__abc_78290_new_n2305_));
AOI21X1 AOI21X1_541 ( .A(u5__abc_78290_new_n2311_), .B(u5__abc_78290_new_n2309_), .C(u5__abc_78290_new_n2141_), .Y(u5__abc_78290_new_n2312_));
AOI21X1 AOI21X1_542 ( .A(u5__abc_78290_new_n2189_), .B(u5__abc_78290_new_n2323_), .C(u5__abc_78290_new_n2211_), .Y(u5__abc_78290_new_n2324_));
AOI21X1 AOI21X1_543 ( .A(u5__abc_78290_new_n2211_), .B(u5__abc_78290_new_n2326_), .C(u5__abc_78290_new_n2223_), .Y(u5__abc_78290_new_n2327_));
AOI21X1 AOI21X1_544 ( .A(u5__abc_78290_new_n1187_), .B(u5__abc_78290_new_n2290_), .C(u5__abc_78290_new_n2337_), .Y(u5__abc_78290_new_n2338_));
AOI21X1 AOI21X1_545 ( .A(u5__abc_78290_new_n2342_), .B(u5__abc_78290_new_n2343_), .C(u5__abc_78290_new_n2189_), .Y(u5__abc_78290_new_n2344_));
AOI21X1 AOI21X1_546 ( .A(u5__abc_78290_new_n2345_), .B(u5__abc_78290_new_n2346_), .C(u5__abc_78290_new_n2224_), .Y(u5__0timer_7_0__4_));
AOI21X1 AOI21X1_547 ( .A(u5__abc_78290_new_n2351_), .B(u5__abc_78290_new_n2188_), .C(u5__abc_78290_new_n2354_), .Y(u5__0timer_7_0__5_));
AOI21X1 AOI21X1_548 ( .A(u5__abc_78290_new_n2359_), .B(u5__abc_78290_new_n2188_), .C(u5__abc_78290_new_n2361_), .Y(u5__0timer_7_0__6_));
AOI21X1 AOI21X1_549 ( .A(u5__abc_78290_new_n2363_), .B(u5__abc_78290_new_n2188_), .C(u5__abc_78290_new_n2365_), .Y(u5__0timer_7_0__7_));
AOI21X1 AOI21X1_55 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1692_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1693_));
AOI21X1 AOI21X1_550 ( .A(u5__abc_78290_new_n2392_), .B(u5__abc_78290_new_n2407_), .C(u5__abc_78290_new_n2413_), .Y(u5__abc_78290_new_n2414_));
AOI21X1 AOI21X1_551 ( .A(u5__abc_78290_new_n2414_), .B(u5__abc_78290_new_n2391_), .C(u5__abc_78290_new_n2385_), .Y(u5__abc_78290_new_n2415_));
AOI21X1 AOI21X1_552 ( .A(u5__abc_78290_new_n2397_), .B(u5__abc_78290_new_n2452_), .C(u5__abc_78290_new_n2450_), .Y(u5__abc_78290_new_n2453_));
AOI21X1 AOI21X1_553 ( .A(u5__abc_78290_new_n2453_), .B(u5__abc_78290_new_n2407_), .C(u5__abc_78290_new_n2437_), .Y(u5__abc_78290_new_n2454_));
AOI21X1 AOI21X1_554 ( .A(u5__abc_78290_new_n2379_), .B(u5__abc_78290_new_n2244_), .C(u5__abc_78290_new_n2385_), .Y(u5__abc_78290_new_n2456_));
AOI21X1 AOI21X1_555 ( .A(u5__abc_78290_new_n2385_), .B(u5__abc_78290_new_n2268_), .C(u5__abc_78290_new_n2458_), .Y(u5__abc_78290_new_n2459_));
AOI21X1 AOI21X1_556 ( .A(u5__abc_78290_new_n2399_), .B(u5__abc_78290_new_n2470_), .C(u5__abc_78290_new_n2450_), .Y(u5__abc_78290_new_n2471_));
AOI21X1 AOI21X1_557 ( .A(u5__abc_78290_new_n2471_), .B(u5__abc_78290_new_n2407_), .C(u5__abc_78290_new_n2437_), .Y(u5__abc_78290_new_n2472_));
AOI21X1 AOI21X1_558 ( .A(u5__abc_78290_new_n2473_), .B(u5__abc_78290_new_n2468_), .C(u5__abc_78290_new_n2467_), .Y(u5__abc_78290_new_n2474_));
AOI21X1 AOI21X1_559 ( .A(u5__abc_78290_new_n2385_), .B(u5__abc_78290_new_n2433_), .C(u5__abc_78290_new_n2458_), .Y(u5__abc_78290_new_n2476_));
AOI21X1 AOI21X1_56 ( .A(u0__abc_74894_new_n1707_), .B(u0__abc_74894_new_n1708_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1709_));
AOI21X1 AOI21X1_560 ( .A(u5__abc_78290_new_n2487_), .B(u5__abc_78290_new_n2488_), .C(u5__abc_78290_new_n2450_), .Y(u5__abc_78290_new_n2489_));
AOI21X1 AOI21X1_561 ( .A(u5__abc_78290_new_n2489_), .B(u5__abc_78290_new_n2407_), .C(u5__abc_78290_new_n2437_), .Y(u5__abc_78290_new_n2490_));
AOI21X1 AOI21X1_562 ( .A(u5__abc_78290_new_n2379_), .B(u5__abc_78290_new_n2308_), .C(u5__abc_78290_new_n2385_), .Y(u5__abc_78290_new_n2493_));
AOI21X1 AOI21X1_563 ( .A(u5__abc_78290_new_n2492_), .B(u5__abc_78290_new_n2493_), .C(u5__abc_78290_new_n2494_), .Y(u5__abc_78290_new_n2495_));
AOI21X1 AOI21X1_564 ( .A(u5__abc_78290_new_n2500_), .B(u5__abc_78290_new_n2502_), .C(u5__abc_78290_new_n2497_), .Y(u5__abc_78290_new_n2503_));
AOI21X1 AOI21X1_565 ( .A(u5__abc_78290_new_n2379_), .B(u5__abc_78290_new_n2506_), .C(u5__abc_78290_new_n2385_), .Y(u5__abc_78290_new_n2507_));
AOI21X1 AOI21X1_566 ( .A(u5__abc_78290_new_n2500_), .B(u5__abc_78290_new_n2513_), .C(u5__abc_78290_new_n2497_), .Y(u5__abc_78290_new_n2514_));
AOI21X1 AOI21X1_567 ( .A(u5__abc_78290_new_n2514_), .B(u5__abc_78290_new_n2510_), .C(u5__abc_78290_new_n2467_), .Y(u5__abc_78290_new_n2515_));
AOI21X1 AOI21X1_568 ( .A(u5_ack_cnt_0_), .B(u5__abc_78290_new_n2537_), .C(u5__abc_78290_new_n2539_), .Y(u5__0ack_cnt_3_0__0_));
AOI21X1 AOI21X1_569 ( .A(u5__abc_78290_new_n2545_), .B(u5__abc_78290_new_n2534_), .C(u5__abc_78290_new_n2546_), .Y(u5__0ack_cnt_3_0__1_));
AOI21X1 AOI21X1_57 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1712_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1713_));
AOI21X1 AOI21X1_570 ( .A(u5__abc_78290_new_n2548_), .B(u5__abc_78290_new_n2550_), .C(u5__abc_78290_new_n2551_), .Y(u5__0ack_cnt_3_0__2_));
AOI21X1 AOI21X1_571 ( .A(u5__abc_78290_new_n2553_), .B(u5__abc_78290_new_n2534_), .C(u5__abc_78290_new_n2556_), .Y(u5__0ack_cnt_3_0__3_));
AOI21X1 AOI21X1_572 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n2566_), .C(u5__abc_78290_new_n2572_), .Y(mc_adv_d));
AOI21X1 AOI21X1_573 ( .A(u5__abc_78290_new_n2584_), .B(u5__abc_78290_new_n2576_), .C(u5__abc_78290_new_n787_), .Y(u5_next_state_0_));
AOI21X1 AOI21X1_574 ( .A(u5__abc_78290_new_n574_), .B(u5__abc_78290_new_n2602_), .C(u5__abc_78290_new_n2567_), .Y(u5__abc_78290_new_n2603_));
AOI21X1 AOI21X1_575 ( .A(u5__abc_78290_new_n2638_), .B(u5__abc_78290_new_n2640_), .C(u5__abc_78290_new_n2635_), .Y(u5__abc_78290_new_n2641_));
AOI21X1 AOI21X1_576 ( .A(u5__abc_78290_new_n1061_), .B(u5__abc_78290_new_n2644_), .C(u5__abc_78290_new_n1618_), .Y(u5__abc_78290_new_n2645_));
AOI21X1 AOI21X1_577 ( .A(u5__abc_78290_new_n1375_), .B(u5__abc_78290_new_n1554_), .C(u5__abc_78290_new_n2659_), .Y(u5__abc_78290_new_n2660_));
AOI21X1 AOI21X1_578 ( .A(u5__abc_78290_new_n733_), .B(u5__abc_78290_new_n1375_), .C(u5__abc_78290_new_n2673_), .Y(u5__abc_78290_new_n2674_));
AOI21X1 AOI21X1_579 ( .A(u5__abc_78290_new_n2653_), .B(u5__abc_78290_new_n2689_), .C(u5__abc_78290_new_n1335_), .Y(u5__abc_78290_new_n2690_));
AOI21X1 AOI21X1_58 ( .A(u0__abc_74894_new_n1828_), .B(u0__abc_74894_new_n1829_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1830_));
AOI21X1 AOI21X1_580 ( .A(u5__abc_78290_new_n1514_), .B(u5__abc_78290_new_n2687_), .C(u5__abc_78290_new_n1335_), .Y(u5__abc_78290_new_n2697_));
AOI21X1 AOI21X1_581 ( .A(u5__abc_78290_new_n1990_), .B(u5__abc_78290_new_n1257_), .C(u5__abc_78290_new_n2728_), .Y(u5__abc_78290_new_n2729_));
AOI21X1 AOI21X1_582 ( .A(u5__abc_78290_new_n829_), .B(u5__abc_78290_new_n1990_), .C(u5__abc_78290_new_n2732_), .Y(u5__abc_78290_new_n2733_));
AOI21X1 AOI21X1_583 ( .A(u5__abc_78290_new_n2750_), .B(u5__abc_78290_new_n2713_), .C(u5__abc_78290_new_n2748_), .Y(u5__abc_78290_new_n2751_));
AOI21X1 AOI21X1_584 ( .A(u5__abc_78290_new_n2753_), .B(u5__abc_78290_new_n2609_), .C(u5__abc_78290_new_n1418_), .Y(u5__abc_78290_new_n2754_));
AOI21X1 AOI21X1_585 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n2756_), .C(u5__abc_78290_new_n2639_), .Y(u5__abc_78290_new_n2757_));
AOI21X1 AOI21X1_586 ( .A(u5__abc_78290_new_n2624_), .B(u5_state_16_), .C(u5__abc_78290_new_n2628_), .Y(u5__abc_78290_new_n2761_));
AOI21X1 AOI21X1_587 ( .A(u5__abc_78290_new_n2631_), .B(u5__abc_78290_new_n2759_), .C(u5__abc_78290_new_n2762_), .Y(u5__abc_78290_new_n2763_));
AOI21X1 AOI21X1_588 ( .A(u5__abc_78290_new_n2731_), .B(u5__abc_78290_new_n2757_), .C(u5__abc_78290_new_n2764_), .Y(u5__abc_78290_new_n2765_));
AOI21X1 AOI21X1_589 ( .A(u5__abc_78290_new_n486_), .B(u5__abc_78290_new_n1410_), .C(u5__abc_78290_new_n1413_), .Y(u5__abc_78290_new_n2769_));
AOI21X1 AOI21X1_59 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1833_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1834_));
AOI21X1 AOI21X1_590 ( .A(u5__abc_78290_new_n2768_), .B(u5__abc_78290_new_n2769_), .C(u5__abc_78290_new_n1418_), .Y(u5__abc_78290_new_n2770_));
AOI21X1 AOI21X1_591 ( .A(u5__abc_78290_new_n603_), .B(u5__abc_78290_new_n1375_), .C(u5__abc_78290_new_n561_), .Y(u5__abc_78290_new_n2798_));
AOI21X1 AOI21X1_592 ( .A(u5__abc_78290_new_n2618_), .B(u5__abc_78290_new_n2799_), .C(u5__abc_78290_new_n2798_), .Y(u5__abc_78290_new_n2800_));
AOI21X1 AOI21X1_593 ( .A(u5__abc_78290_new_n2680_), .B(u5_state_21_), .C(init_req), .Y(u5__abc_78290_new_n2802_));
AOI21X1 AOI21X1_594 ( .A(u5__abc_78290_new_n582_), .B(u5__abc_78290_new_n1990_), .C(u5__abc_78290_new_n1207_), .Y(u5__abc_78290_new_n2821_));
AOI21X1 AOI21X1_595 ( .A(u5__abc_78290_new_n1197_), .B(u5__abc_78290_new_n2822_), .C(u5__abc_78290_new_n2821_), .Y(u5__abc_78290_new_n2823_));
AOI21X1 AOI21X1_596 ( .A(u5__abc_78290_new_n2788_), .B(u5_state_27_), .C(u5__abc_78290_new_n1339_), .Y(u5__abc_78290_new_n2831_));
AOI21X1 AOI21X1_597 ( .A(u5__abc_78290_new_n2783_), .B(u5__abc_78290_new_n2853_), .C(u5__abc_78290_new_n2052_), .Y(u5__abc_78290_new_n2854_));
AOI21X1 AOI21X1_598 ( .A(u5__abc_78290_new_n2620_), .B(mc_br_r), .C(u5__abc_78290_new_n1557_), .Y(u5__abc_78290_new_n2859_));
AOI21X1 AOI21X1_599 ( .A(u5__abc_78290_new_n1380_), .B(u5_tmr2_done), .C(u5_state_43_), .Y(u5__abc_78290_new_n2891_));
AOI21X1 AOI21X1_6 ( .A(u0__abc_74894_new_n1207_), .B(u0__abc_74894_new_n1208_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1209_));
AOI21X1 AOI21X1_60 ( .A(u0__abc_74894_new_n1848_), .B(u0__abc_74894_new_n1849_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1850_));
AOI21X1 AOI21X1_600 ( .A(u5__abc_78290_new_n2584_), .B(u5__abc_78290_new_n2890_), .C(u5__abc_78290_new_n2891_), .Y(u5_next_state_43_));
AOI21X1 AOI21X1_601 ( .A(u5__abc_78290_new_n1161_), .B(u5__abc_78290_new_n2902_), .C(u5__abc_78290_new_n1165_), .Y(u5__abc_78290_new_n2903_));
AOI21X1 AOI21X1_602 ( .A(u5__abc_78290_new_n2742_), .B(u5__abc_78290_new_n911_), .C(u5__abc_78290_new_n2697_), .Y(u5__abc_78290_new_n2941_));
AOI21X1 AOI21X1_603 ( .A(u5__abc_78290_new_n2922_), .B(u5__abc_78290_new_n2940_), .C(u5__abc_78290_new_n2944_), .Y(u5__abc_78290_new_n2945_));
AOI21X1 AOI21X1_604 ( .A(u5__abc_78290_new_n2745_), .B(u5__abc_78290_new_n909_), .C(u5__abc_78290_new_n2950_), .Y(u5__abc_78290_new_n2951_));
AOI21X1 AOI21X1_605 ( .A(u5__abc_78290_new_n2949_), .B(u5__abc_78290_new_n2951_), .C(u5__abc_78290_new_n2952_), .Y(u5__abc_78290_new_n2953_));
AOI21X1 AOI21X1_606 ( .A(u5__abc_78290_new_n2987_), .B(u5__abc_78290_new_n2988_), .C(u5__abc_78290_new_n1502_), .Y(u5__abc_78290_new_n2989_));
AOI21X1 AOI21X1_607 ( .A(u5__abc_78290_new_n489_), .B(u5__abc_78290_new_n2565_), .C(u5__abc_78290_new_n2991_), .Y(u5_next_state_65_));
AOI21X1 AOI21X1_608 ( .A(u5__abc_78290_new_n1273_), .B(u5__abc_78290_new_n3009_), .C(u5__abc_78290_new_n2835_), .Y(u5__abc_78290_new_n3010_));
AOI21X1 AOI21X1_609 ( .A(u5__abc_78290_new_n1061_), .B(u5__abc_78290_new_n2587_), .C(u5__abc_78290_new_n2567_), .Y(u5__abc_78290_new_n3040_));
AOI21X1 AOI21X1_61 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1853_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1854_));
AOI21X1 AOI21X1_610 ( .A(u5_wb_cycle), .B(u5__abc_78290_new_n3041_), .C(u5__abc_78290_new_n3047_), .Y(u5__abc_78290_new_n3048_));
AOI21X1 AOI21X1_611 ( .A(u5__abc_78290_new_n1262_), .B(u5__abc_78290_new_n1325_), .C(u5__abc_78290_new_n3105_), .Y(u5__abc_78290_new_n3106_));
AOI21X1 AOI21X1_612 ( .A(u5__abc_78290_new_n3107_), .B(u5__abc_78290_new_n3109_), .C(u5__abc_78290_new_n3112_), .Y(u5__abc_78290_new_n3113_));
AOI21X1 AOI21X1_613 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n1069_), .C(u5__abc_78290_new_n2190_), .Y(u5__abc_78290_new_n3126_));
AOI21X1 AOI21X1_614 ( .A(u5__abc_78290_new_n3135_), .B(u5__abc_78290_new_n3139_), .C(u5__abc_78290_new_n1416_), .Y(u5__0cke__0_0_));
AOI21X1 AOI21X1_615 ( .A(u6__abc_81318_new_n250_), .B(u6__abc_81318_new_n247_), .C(u6__abc_81318_new_n256_), .Y(u6__0read_go_r1_0_0_));
AOI21X1 AOI21X1_616 ( .A(u6__abc_81318_new_n263_), .B(u6__abc_81318_new_n262_), .C(u6__abc_81318_new_n136_), .Y(u6__0write_go_r1_0_0_));
AOI21X1 AOI21X1_617 ( .A(u6__abc_81318_new_n248_), .B(wb_stb_i), .C(u6__abc_81318_new_n265_), .Y(u6__0write_go_r_0_0_));
AOI21X1 AOI21X1_618 ( .A(u6__abc_81318_new_n260_), .B(u6__abc_81318_new_n267_), .C(u6__abc_81318_new_n275_), .Y(u5_wb_wait));
AOI21X1 AOI21X1_619 ( .A(u7__abc_73829_new_n107_), .B(u7__abc_73829_new_n105_), .C(u7__abc_73829_new_n106_), .Y(u7__abc_73829_new_n108_));
AOI21X1 AOI21X1_62 ( .A(u0__abc_74894_new_n1868_), .B(u0__abc_74894_new_n1869_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1870_));
AOI21X1 AOI21X1_620 ( .A(u7__abc_73829_new_n107_), .B(u7__abc_73829_new_n113_), .C(u7__abc_73829_new_n106_), .Y(u7__abc_73829_new_n114_));
AOI21X1 AOI21X1_621 ( .A(u7__abc_73829_new_n107_), .B(u7__abc_73829_new_n119_), .C(u7__abc_73829_new_n106_), .Y(u7__abc_73829_new_n120_));
AOI21X1 AOI21X1_622 ( .A(u7__abc_73829_new_n107_), .B(u7__abc_73829_new_n125_), .C(u7__abc_73829_new_n106_), .Y(u7__abc_73829_new_n126_));
AOI21X1 AOI21X1_623 ( .A(u7__abc_73829_new_n107_), .B(u7__abc_73829_new_n131_), .C(u7__abc_73829_new_n106_), .Y(u7__abc_73829_new_n132_));
AOI21X1 AOI21X1_624 ( .A(u7__abc_73829_new_n107_), .B(u7__abc_73829_new_n137_), .C(u7__abc_73829_new_n106_), .Y(u7__abc_73829_new_n138_));
AOI21X1 AOI21X1_625 ( .A(u7__abc_73829_new_n107_), .B(u7__abc_73829_new_n143_), .C(u7__abc_73829_new_n106_), .Y(u7__abc_73829_new_n144_));
AOI21X1 AOI21X1_626 ( .A(u7__abc_73829_new_n107_), .B(u7__abc_73829_new_n149_), .C(u7__abc_73829_new_n106_), .Y(u7__abc_73829_new_n150_));
AOI21X1 AOI21X1_63 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1873_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1874_));
AOI21X1 AOI21X1_64 ( .A(u0__abc_74894_new_n1888_), .B(u0__abc_74894_new_n1889_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1890_));
AOI21X1 AOI21X1_65 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1893_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1894_));
AOI21X1 AOI21X1_66 ( .A(u0__abc_74894_new_n1908_), .B(u0__abc_74894_new_n1909_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1910_));
AOI21X1 AOI21X1_67 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1913_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1914_));
AOI21X1 AOI21X1_68 ( .A(u0__abc_74894_new_n1928_), .B(u0__abc_74894_new_n1929_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1930_));
AOI21X1 AOI21X1_69 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1933_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1934_));
AOI21X1 AOI21X1_7 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1212_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1213_));
AOI21X1 AOI21X1_70 ( .A(u0__abc_74894_new_n1948_), .B(u0__abc_74894_new_n1949_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1950_));
AOI21X1 AOI21X1_71 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1953_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1954_));
AOI21X1 AOI21X1_72 ( .A(u0__abc_74894_new_n1988_), .B(u0__abc_74894_new_n1989_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1990_));
AOI21X1 AOI21X1_73 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1993_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1994_));
AOI21X1 AOI21X1_74 ( .A(u0__abc_74894_new_n2008_), .B(u0__abc_74894_new_n2009_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n2010_));
AOI21X1 AOI21X1_75 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n2013_), .C(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n2014_));
AOI21X1 AOI21X1_76 ( .A(u0__abc_74894_new_n2451_), .B(u0__abc_74894_new_n2452_), .C(u0_cs1), .Y(u0__abc_74894_new_n2453_));
AOI21X1 AOI21X1_77 ( .A(u0__abc_74894_new_n1172_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2457_));
AOI21X1 AOI21X1_78 ( .A(u0__abc_74894_new_n2469_), .B(u0__abc_74894_new_n2470_), .C(u0_cs1), .Y(u0__abc_74894_new_n2471_));
AOI21X1 AOI21X1_79 ( .A(u0__abc_74894_new_n1192_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2473_));
AOI21X1 AOI21X1_8 ( .A(u0__abc_74894_new_n1227_), .B(u0__abc_74894_new_n1228_), .C(spec_req_cs_1_), .Y(u0__abc_74894_new_n1229_));
AOI21X1 AOI21X1_80 ( .A(u0__abc_74894_new_n2485_), .B(u0__abc_74894_new_n2486_), .C(u0_cs1), .Y(u0__abc_74894_new_n2487_));
AOI21X1 AOI21X1_81 ( .A(u0__abc_74894_new_n1212_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2489_));
AOI21X1 AOI21X1_82 ( .A(u0__abc_74894_new_n2501_), .B(u0__abc_74894_new_n2502_), .C(u0_cs1), .Y(u0__abc_74894_new_n2503_));
AOI21X1 AOI21X1_83 ( .A(u0__abc_74894_new_n1232_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2505_));
AOI21X1 AOI21X1_84 ( .A(u0__abc_74894_new_n2517_), .B(u0__abc_74894_new_n2518_), .C(u0_cs1), .Y(u0__abc_74894_new_n2519_));
AOI21X1 AOI21X1_85 ( .A(u0__abc_74894_new_n1252_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2521_));
AOI21X1 AOI21X1_86 ( .A(u0__abc_74894_new_n2533_), .B(u0__abc_74894_new_n2534_), .C(u0_cs1), .Y(u0__abc_74894_new_n2535_));
AOI21X1 AOI21X1_87 ( .A(u0__abc_74894_new_n1272_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2537_));
AOI21X1 AOI21X1_88 ( .A(u0__abc_74894_new_n2549_), .B(u0__abc_74894_new_n2550_), .C(u0_cs1), .Y(u0__abc_74894_new_n2551_));
AOI21X1 AOI21X1_89 ( .A(u0__abc_74894_new_n1292_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2553_));
AOI21X1 AOI21X1_9 ( .A(spec_req_cs_0_), .B(u0__abc_74894_new_n1232_), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1233_));
AOI21X1 AOI21X1_90 ( .A(u0__abc_74894_new_n2565_), .B(u0__abc_74894_new_n2566_), .C(u0_cs1), .Y(u0__abc_74894_new_n2567_));
AOI21X1 AOI21X1_91 ( .A(u0__abc_74894_new_n1312_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2569_));
AOI21X1 AOI21X1_92 ( .A(u0__abc_74894_new_n2581_), .B(u0__abc_74894_new_n2582_), .C(u0_cs1), .Y(u0__abc_74894_new_n2583_));
AOI21X1 AOI21X1_93 ( .A(u0__abc_74894_new_n1332_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2585_));
AOI21X1 AOI21X1_94 ( .A(u0__abc_74894_new_n2597_), .B(u0__abc_74894_new_n2598_), .C(u0_cs1), .Y(u0__abc_74894_new_n2599_));
AOI21X1 AOI21X1_95 ( .A(u0__abc_74894_new_n1352_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2601_));
AOI21X1 AOI21X1_96 ( .A(u0__abc_74894_new_n2613_), .B(u0__abc_74894_new_n2614_), .C(u0_cs1), .Y(u0__abc_74894_new_n2615_));
AOI21X1 AOI21X1_97 ( .A(u0__abc_74894_new_n1372_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2617_));
AOI21X1 AOI21X1_98 ( .A(u0__abc_74894_new_n2629_), .B(u0__abc_74894_new_n2630_), .C(u0_cs1), .Y(u0__abc_74894_new_n2631_));
AOI21X1 AOI21X1_99 ( .A(u0__abc_74894_new_n1392_), .B(u0_cs0), .C(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2633_));
AOI22X1 AOI22X1_1 ( .A(u0__abc_74894_new_n3699_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3702_));
AOI22X1 AOI22X1_10 ( .A(u0__abc_74894_new_n3749_), .B(u0_csc_mask_1_), .C(\poc_o[1] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3772_));
AOI22X1 AOI22X1_100 ( .A(\wb_addr_i[11] ), .B(page_size_8_), .C(\wb_addr_i[12] ), .D(page_size_9_), .Y(u1__abc_72801_new_n309_));
AOI22X1 AOI22X1_101 ( .A(\wb_addr_i[12] ), .B(page_size_8_), .C(\wb_addr_i[13] ), .D(page_size_9_), .Y(u1__abc_72801_new_n325_));
AOI22X1 AOI22X1_102 ( .A(u1__abc_72801_new_n280_), .B(u1__abc_72801_new_n279_), .C(u1__abc_72801_new_n281_), .D(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n333_));
AOI22X1 AOI22X1_103 ( .A(u1__abc_72801_new_n292_), .B(u1__abc_72801_new_n279_), .C(u1__abc_72801_new_n280_), .D(u1__abc_72801_new_n335_), .Y(u1__abc_72801_new_n337_));
AOI22X1 AOI22X1_104 ( .A(\wb_addr_i[15] ), .B(u1__abc_72801_new_n340_), .C(\wb_addr_i[13] ), .D(page_size_8_), .Y(u1__abc_72801_new_n341_));
AOI22X1 AOI22X1_105 ( .A(\wb_addr_i[16] ), .B(u1__abc_72801_new_n340_), .C(\wb_addr_i[14] ), .D(page_size_8_), .Y(u1__abc_72801_new_n354_));
AOI22X1 AOI22X1_106 ( .A(\wb_addr_i[17] ), .B(u1__abc_72801_new_n340_), .C(\wb_addr_i[15] ), .D(page_size_8_), .Y(u1__abc_72801_new_n366_));
AOI22X1 AOI22X1_107 ( .A(\wb_addr_i[18] ), .B(u1__abc_72801_new_n340_), .C(\wb_addr_i[16] ), .D(page_size_8_), .Y(u1__abc_72801_new_n374_));
AOI22X1 AOI22X1_108 ( .A(\wb_addr_i[19] ), .B(u1__abc_72801_new_n340_), .C(\wb_addr_i[17] ), .D(page_size_8_), .Y(u1__abc_72801_new_n384_));
AOI22X1 AOI22X1_109 ( .A(\wb_addr_i[20] ), .B(u1__abc_72801_new_n340_), .C(\wb_addr_i[18] ), .D(page_size_8_), .Y(u1__abc_72801_new_n393_));
AOI22X1 AOI22X1_11 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_1_), .C(u0_tms0_1_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3774_));
AOI22X1 AOI22X1_110 ( .A(\wb_addr_i[19] ), .B(page_size_8_), .C(\wb_addr_i[20] ), .D(page_size_9_), .Y(u1__abc_72801_new_n403_));
AOI22X1 AOI22X1_111 ( .A(\wb_addr_i[20] ), .B(page_size_8_), .C(\wb_addr_i[21] ), .D(page_size_9_), .Y(u1__abc_72801_new_n413_));
AOI22X1 AOI22X1_112 ( .A(\wb_addr_i[22] ), .B(u1__abc_72801_new_n267_), .C(\wb_addr_i[21] ), .D(u1__abc_72801_new_n334_), .Y(u1__abc_72801_new_n421_));
AOI22X1 AOI22X1_113 ( .A(u1__abc_72801_new_n340_), .B(\wb_addr_i[24] ), .C(\wb_addr_i[23] ), .D(u1__abc_72801_new_n267_), .Y(u1__abc_72801_new_n436_));
AOI22X1 AOI22X1_114 ( .A(u1__abc_72801_new_n264_), .B(\wb_addr_i[23] ), .C(\wb_addr_i[22] ), .D(u1__abc_72801_new_n299_), .Y(u1__abc_72801_new_n437_));
AOI22X1 AOI22X1_115 ( .A(u1__abc_72801_new_n340_), .B(\wb_addr_i[26] ), .C(\wb_addr_i[25] ), .D(u1__abc_72801_new_n267_), .Y(u1__abc_72801_new_n454_));
AOI22X1 AOI22X1_116 ( .A(u1__abc_72801_new_n280_), .B(\wb_addr_i[16] ), .C(\wb_addr_i[17] ), .D(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n575_));
AOI22X1 AOI22X1_117 ( .A(u1__abc_72801_new_n280_), .B(\wb_addr_i[17] ), .C(\wb_addr_i[18] ), .D(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n581_));
AOI22X1 AOI22X1_118 ( .A(u1__abc_72801_new_n280_), .B(\wb_addr_i[20] ), .C(\wb_addr_i[21] ), .D(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n597_));
AOI22X1 AOI22X1_119 ( .A(u1__abc_72801_new_n280_), .B(\wb_addr_i[22] ), .C(\wb_addr_i[23] ), .D(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n606_));
AOI22X1 AOI22X1_12 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3778_));
AOI22X1 AOI22X1_120 ( .A(u1__abc_72801_new_n280_), .B(\wb_addr_i[23] ), .C(\wb_addr_i[24] ), .D(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n611_));
AOI22X1 AOI22X1_121 ( .A(u1__abc_72801_new_n280_), .B(\wb_addr_i[24] ), .C(\wb_addr_i[25] ), .D(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n616_));
AOI22X1 AOI22X1_122 ( .A(obct_cs_2_), .B(1'h0), .C(obct_cs_4_), .D(1'h0), .Y(u2__abc_74202_new_n100_));
AOI22X1 AOI22X1_123 ( .A(obct_cs_3_), .B(1'h0), .C(obct_cs_5_), .D(1'h0), .Y(u2__abc_74202_new_n101_));
AOI22X1 AOI22X1_124 ( .A(obct_cs_0_), .B(u2_bank_open_0), .C(obct_cs_1_), .D(u2_bank_open_1), .Y(u2__abc_74202_new_n103_));
AOI22X1 AOI22X1_125 ( .A(obct_cs_6_), .B(1'h0), .C(obct_cs_7_), .D(1'h0), .Y(u2__abc_74202_new_n104_));
AOI22X1 AOI22X1_126 ( .A(obct_cs_2_), .B(1'h0), .C(obct_cs_4_), .D(1'h0), .Y(u2__abc_74202_new_n107_));
AOI22X1 AOI22X1_127 ( .A(obct_cs_3_), .B(1'h0), .C(obct_cs_5_), .D(1'h0), .Y(u2__abc_74202_new_n108_));
AOI22X1 AOI22X1_128 ( .A(obct_cs_0_), .B(u2_row_same_0), .C(obct_cs_1_), .D(u2_row_same_1), .Y(u2__abc_74202_new_n110_));
AOI22X1 AOI22X1_129 ( .A(obct_cs_6_), .B(1'h0), .C(obct_cs_7_), .D(1'h0), .Y(u2__abc_74202_new_n111_));
AOI22X1 AOI22X1_13 ( .A(u0__abc_74894_new_n3699_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3779_));
AOI22X1 AOI22X1_130 ( .A(u2_u0__abc_73914_new_n267_), .B(row_adr_9_), .C(u2_u0_b3_last_row_11_), .D(u2_u0__abc_73914_new_n173_), .Y(u2_u0__abc_73914_new_n270_));
AOI22X1 AOI22X1_131 ( .A(u2_u0__abc_73914_new_n152_), .B(u2_u0_b3_last_row_4_), .C(u2_u0__abc_73914_new_n271_), .D(row_adr_11_), .Y(u2_u0__abc_73914_new_n272_));
AOI22X1 AOI22X1_132 ( .A(u2_u0__abc_73914_new_n278_), .B(u2_u0__abc_73914_new_n277_), .C(u2_u0__abc_73914_new_n279_), .D(u2_u0__abc_73914_new_n280_), .Y(u2_u0__abc_73914_new_n281_));
AOI22X1 AOI22X1_133 ( .A(u2_u0__abc_73914_new_n143_), .B(u2_u0_b3_last_row_1_), .C(u2_u0__abc_73914_new_n290_), .D(row_adr_2_), .Y(u2_u0__abc_73914_new_n291_));
AOI22X1 AOI22X1_134 ( .A(u2_u0__abc_73914_new_n307_), .B(u2_u0__abc_73914_new_n306_), .C(u2_u0__abc_73914_new_n308_), .D(u2_u0__abc_73914_new_n309_), .Y(u2_u0__abc_73914_new_n310_));
AOI22X1 AOI22X1_135 ( .A(u2_u0__abc_73914_new_n161_), .B(u2_u0_b1_last_row_7_), .C(row_adr_9_), .D(u2_u0__abc_73914_new_n324_), .Y(u2_u0__abc_73914_new_n325_));
AOI22X1 AOI22X1_136 ( .A(u2_u0__abc_73914_new_n314_), .B(u2_u0__abc_73914_new_n328_), .C(u2_u0__abc_73914_new_n283_), .D(u2_u0__abc_73914_new_n297_), .Y(u2_u0__abc_73914_new_n329_));
AOI22X1 AOI22X1_137 ( .A(u2_u0__abc_73914_new_n176_), .B(u2_u0_b0_last_row_12_), .C(row_adr_3_), .D(u2_u0__abc_73914_new_n334_), .Y(u2_u0__abc_73914_new_n335_));
AOI22X1 AOI22X1_138 ( .A(u2_u0__abc_73914_new_n341_), .B(row_adr_6_), .C(row_adr_12_), .D(u2_u0__abc_73914_new_n342_), .Y(u2_u0__abc_73914_new_n343_));
AOI22X1 AOI22X1_139 ( .A(u2_u0__abc_73914_new_n346_), .B(u2_u0__abc_73914_new_n347_), .C(u2_u0__abc_73914_new_n348_), .D(u2_u0__abc_73914_new_n349_), .Y(u2_u0__abc_73914_new_n350_));
AOI22X1 AOI22X1_14 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3781_));
AOI22X1 AOI22X1_140 ( .A(u2_u0__abc_73914_new_n152_), .B(u2_u0_b0_last_row_4_), .C(u2_u0__abc_73914_new_n173_), .D(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_73914_new_n354_));
AOI22X1 AOI22X1_141 ( .A(u2_u0__abc_73914_new_n355_), .B(row_adr_2_), .C(row_adr_4_), .D(u2_u0__abc_73914_new_n356_), .Y(u2_u0__abc_73914_new_n357_));
AOI22X1 AOI22X1_142 ( .A(u2_u0__abc_73914_new_n359_), .B(u2_u0__abc_73914_new_n358_), .C(u2_u0__abc_73914_new_n360_), .D(u2_u0__abc_73914_new_n361_), .Y(u2_u0__abc_73914_new_n362_));
AOI22X1 AOI22X1_143 ( .A(u2_u0__abc_73914_new_n167_), .B(u2_u0_b2_last_row_9_), .C(row_adr_11_), .D(u2_u0__abc_73914_new_n367_), .Y(u2_u0__abc_73914_new_n368_));
AOI22X1 AOI22X1_144 ( .A(u2_u0__abc_73914_new_n173_), .B(u2_u0_b2_last_row_11_), .C(row_adr_4_), .D(u2_u0__abc_73914_new_n369_), .Y(u2_u0__abc_73914_new_n370_));
AOI22X1 AOI22X1_145 ( .A(u2_u0__abc_73914_new_n152_), .B(u2_u0_b2_last_row_4_), .C(row_adr_6_), .D(u2_u0__abc_73914_new_n374_), .Y(u2_u0__abc_73914_new_n388_));
AOI22X1 AOI22X1_146 ( .A(u2_u0__abc_73914_new_n364_), .B(u2_u0__abc_73914_new_n345_), .C(u2_u0__abc_73914_new_n383_), .D(u2_u0__abc_73914_new_n395_), .Y(u2_u0__abc_73914_new_n396_));
AOI22X1 AOI22X1_147 ( .A(u2_u0__abc_73914_new_n138_), .B(u2_u0_bank3_open), .C(u2_u0_bank2_open), .D(u2_u0__abc_73914_new_n237_), .Y(u2_u0__abc_73914_new_n400_));
AOI22X1 AOI22X1_148 ( .A(u2_u1__abc_73914_new_n267_), .B(row_adr_9_), .C(u2_u1_b3_last_row_11_), .D(u2_u1__abc_73914_new_n173_), .Y(u2_u1__abc_73914_new_n270_));
AOI22X1 AOI22X1_149 ( .A(u2_u1__abc_73914_new_n152_), .B(u2_u1_b3_last_row_4_), .C(u2_u1__abc_73914_new_n271_), .D(row_adr_11_), .Y(u2_u1__abc_73914_new_n272_));
AOI22X1 AOI22X1_15 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3782_));
AOI22X1 AOI22X1_150 ( .A(u2_u1__abc_73914_new_n278_), .B(u2_u1__abc_73914_new_n277_), .C(u2_u1__abc_73914_new_n279_), .D(u2_u1__abc_73914_new_n280_), .Y(u2_u1__abc_73914_new_n281_));
AOI22X1 AOI22X1_151 ( .A(u2_u1__abc_73914_new_n143_), .B(u2_u1_b3_last_row_1_), .C(u2_u1__abc_73914_new_n290_), .D(row_adr_2_), .Y(u2_u1__abc_73914_new_n291_));
AOI22X1 AOI22X1_152 ( .A(u2_u1__abc_73914_new_n307_), .B(u2_u1__abc_73914_new_n306_), .C(u2_u1__abc_73914_new_n308_), .D(u2_u1__abc_73914_new_n309_), .Y(u2_u1__abc_73914_new_n310_));
AOI22X1 AOI22X1_153 ( .A(u2_u1__abc_73914_new_n161_), .B(u2_u1_b1_last_row_7_), .C(row_adr_9_), .D(u2_u1__abc_73914_new_n324_), .Y(u2_u1__abc_73914_new_n325_));
AOI22X1 AOI22X1_154 ( .A(u2_u1__abc_73914_new_n314_), .B(u2_u1__abc_73914_new_n328_), .C(u2_u1__abc_73914_new_n283_), .D(u2_u1__abc_73914_new_n297_), .Y(u2_u1__abc_73914_new_n329_));
AOI22X1 AOI22X1_155 ( .A(u2_u1__abc_73914_new_n176_), .B(u2_u1_b0_last_row_12_), .C(row_adr_3_), .D(u2_u1__abc_73914_new_n334_), .Y(u2_u1__abc_73914_new_n335_));
AOI22X1 AOI22X1_156 ( .A(u2_u1__abc_73914_new_n341_), .B(row_adr_6_), .C(row_adr_12_), .D(u2_u1__abc_73914_new_n342_), .Y(u2_u1__abc_73914_new_n343_));
AOI22X1 AOI22X1_157 ( .A(u2_u1__abc_73914_new_n346_), .B(u2_u1__abc_73914_new_n347_), .C(u2_u1__abc_73914_new_n348_), .D(u2_u1__abc_73914_new_n349_), .Y(u2_u1__abc_73914_new_n350_));
AOI22X1 AOI22X1_158 ( .A(u2_u1__abc_73914_new_n152_), .B(u2_u1_b0_last_row_4_), .C(u2_u1__abc_73914_new_n173_), .D(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_73914_new_n354_));
AOI22X1 AOI22X1_159 ( .A(u2_u1__abc_73914_new_n355_), .B(row_adr_2_), .C(row_adr_4_), .D(u2_u1__abc_73914_new_n356_), .Y(u2_u1__abc_73914_new_n357_));
AOI22X1 AOI22X1_16 ( .A(u0__abc_74894_new_n3749_), .B(u0_csc_mask_2_), .C(\poc_o[2] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3791_));
AOI22X1 AOI22X1_160 ( .A(u2_u1__abc_73914_new_n359_), .B(u2_u1__abc_73914_new_n358_), .C(u2_u1__abc_73914_new_n360_), .D(u2_u1__abc_73914_new_n361_), .Y(u2_u1__abc_73914_new_n362_));
AOI22X1 AOI22X1_161 ( .A(u2_u1__abc_73914_new_n167_), .B(u2_u1_b2_last_row_9_), .C(row_adr_11_), .D(u2_u1__abc_73914_new_n367_), .Y(u2_u1__abc_73914_new_n368_));
AOI22X1 AOI22X1_162 ( .A(u2_u1__abc_73914_new_n173_), .B(u2_u1_b2_last_row_11_), .C(row_adr_4_), .D(u2_u1__abc_73914_new_n369_), .Y(u2_u1__abc_73914_new_n370_));
AOI22X1 AOI22X1_163 ( .A(u2_u1__abc_73914_new_n152_), .B(u2_u1_b2_last_row_4_), .C(row_adr_6_), .D(u2_u1__abc_73914_new_n374_), .Y(u2_u1__abc_73914_new_n388_));
AOI22X1 AOI22X1_164 ( .A(u2_u1__abc_73914_new_n364_), .B(u2_u1__abc_73914_new_n345_), .C(u2_u1__abc_73914_new_n383_), .D(u2_u1__abc_73914_new_n395_), .Y(u2_u1__abc_73914_new_n396_));
AOI22X1 AOI22X1_165 ( .A(u2_u1__abc_73914_new_n138_), .B(u2_u1_bank3_open), .C(u2_u1_bank2_open), .D(u2_u1__abc_73914_new_n237_), .Y(u2_u1__abc_73914_new_n400_));
AOI22X1 AOI22X1_166 ( .A(csc_5_), .B(mc_data_ir_16_), .C(mc_data_ir_0_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n563_));
AOI22X1 AOI22X1_167 ( .A(u3__abc_73372_new_n562_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n564_), .D(u3__abc_73372_new_n563_), .Y(mem_dout_16_));
AOI22X1 AOI22X1_168 ( .A(csc_5_), .B(mc_data_ir_17_), .C(mc_data_ir_1_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n567_));
AOI22X1 AOI22X1_169 ( .A(u3__abc_73372_new_n566_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n568_), .D(u3__abc_73372_new_n567_), .Y(mem_dout_17_));
AOI22X1 AOI22X1_17 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_2_), .C(u0_tms0_2_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3793_));
AOI22X1 AOI22X1_170 ( .A(csc_5_), .B(mc_data_ir_18_), .C(mc_data_ir_2_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n571_));
AOI22X1 AOI22X1_171 ( .A(u3__abc_73372_new_n570_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n572_), .D(u3__abc_73372_new_n571_), .Y(mem_dout_18_));
AOI22X1 AOI22X1_172 ( .A(csc_5_), .B(mc_data_ir_19_), .C(mc_data_ir_3_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n575_));
AOI22X1 AOI22X1_173 ( .A(u3__abc_73372_new_n574_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n576_), .D(u3__abc_73372_new_n575_), .Y(mem_dout_19_));
AOI22X1 AOI22X1_174 ( .A(csc_5_), .B(mc_data_ir_20_), .C(mc_data_ir_4_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n579_));
AOI22X1 AOI22X1_175 ( .A(u3__abc_73372_new_n578_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n580_), .D(u3__abc_73372_new_n579_), .Y(mem_dout_20_));
AOI22X1 AOI22X1_176 ( .A(csc_5_), .B(mc_data_ir_21_), .C(mc_data_ir_5_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n583_));
AOI22X1 AOI22X1_177 ( .A(u3__abc_73372_new_n582_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n584_), .D(u3__abc_73372_new_n583_), .Y(mem_dout_21_));
AOI22X1 AOI22X1_178 ( .A(csc_5_), .B(mc_data_ir_22_), .C(mc_data_ir_6_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n587_));
AOI22X1 AOI22X1_179 ( .A(u3__abc_73372_new_n586_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n588_), .D(u3__abc_73372_new_n587_), .Y(mem_dout_22_));
AOI22X1 AOI22X1_18 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_3_), .C(u0_tms0_3_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3801_));
AOI22X1 AOI22X1_180 ( .A(csc_5_), .B(mc_data_ir_23_), .C(mc_data_ir_7_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n591_));
AOI22X1 AOI22X1_181 ( .A(u3__abc_73372_new_n590_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n592_), .D(u3__abc_73372_new_n591_), .Y(mem_dout_23_));
AOI22X1 AOI22X1_182 ( .A(csc_5_), .B(mc_data_ir_24_), .C(mc_data_ir_8_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n595_));
AOI22X1 AOI22X1_183 ( .A(u3__abc_73372_new_n594_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n596_), .D(u3__abc_73372_new_n595_), .Y(mem_dout_24_));
AOI22X1 AOI22X1_184 ( .A(csc_5_), .B(mc_data_ir_25_), .C(mc_data_ir_9_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n599_));
AOI22X1 AOI22X1_185 ( .A(u3__abc_73372_new_n598_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n600_), .D(u3__abc_73372_new_n599_), .Y(mem_dout_25_));
AOI22X1 AOI22X1_186 ( .A(csc_5_), .B(mc_data_ir_26_), .C(mc_data_ir_10_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n603_));
AOI22X1 AOI22X1_187 ( .A(u3__abc_73372_new_n602_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n604_), .D(u3__abc_73372_new_n603_), .Y(mem_dout_26_));
AOI22X1 AOI22X1_188 ( .A(csc_5_), .B(mc_data_ir_27_), .C(mc_data_ir_11_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n607_));
AOI22X1 AOI22X1_189 ( .A(u3__abc_73372_new_n606_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n608_), .D(u3__abc_73372_new_n607_), .Y(mem_dout_27_));
AOI22X1 AOI22X1_19 ( .A(u0__abc_74894_new_n3749_), .B(u0_csc_mask_3_), .C(u0_tms1_3_), .D(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n3803_));
AOI22X1 AOI22X1_190 ( .A(csc_5_), .B(mc_data_ir_28_), .C(mc_data_ir_12_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n611_));
AOI22X1 AOI22X1_191 ( .A(u3__abc_73372_new_n610_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n612_), .D(u3__abc_73372_new_n611_), .Y(mem_dout_28_));
AOI22X1 AOI22X1_192 ( .A(csc_5_), .B(mc_data_ir_29_), .C(mc_data_ir_13_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n615_));
AOI22X1 AOI22X1_193 ( .A(u3__abc_73372_new_n614_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n616_), .D(u3__abc_73372_new_n615_), .Y(mem_dout_29_));
AOI22X1 AOI22X1_194 ( .A(csc_5_), .B(mc_data_ir_30_), .C(mc_data_ir_14_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n619_));
AOI22X1 AOI22X1_195 ( .A(u3__abc_73372_new_n618_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n620_), .D(u3__abc_73372_new_n619_), .Y(mem_dout_30_));
AOI22X1 AOI22X1_196 ( .A(csc_5_), .B(mc_data_ir_31_), .C(mc_data_ir_15_), .D(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n623_));
AOI22X1 AOI22X1_197 ( .A(u3__abc_73372_new_n622_), .B(u3__abc_73372_new_n275_), .C(u3__abc_73372_new_n624_), .D(u3__abc_73372_new_n623_), .Y(mem_dout_31_));
AOI22X1 AOI22X1_198 ( .A(u3__abc_73372_new_n647_), .B(u3__abc_73372_new_n649_), .C(u3__abc_73372_new_n674_), .D(u3__abc_73372_new_n677_), .Y(u3__abc_73372_new_n678_));
AOI22X1 AOI22X1_199 ( .A(u3__abc_73372_new_n695_), .B(u3__abc_73372_new_n699_), .C(u3__abc_73372_new_n724_), .D(u3__abc_73372_new_n727_), .Y(u3__abc_73372_new_n728_));
AOI22X1 AOI22X1_2 ( .A(u0__abc_74894_new_n3713_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3714_));
AOI22X1 AOI22X1_20 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n3808_));
AOI22X1 AOI22X1_200 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_0_), .C(u3_u0_r2_0_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n748_));
AOI22X1 AOI22X1_201 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_1_), .C(u3_u0_r2_1_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n752_));
AOI22X1 AOI22X1_202 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_2_), .C(u3_u0_r2_2_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n756_));
AOI22X1 AOI22X1_203 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_3_), .C(u3_u0_r2_3_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n760_));
AOI22X1 AOI22X1_204 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_4_), .C(u3_u0_r2_4_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n764_));
AOI22X1 AOI22X1_205 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_5_), .C(u3_u0_r2_5_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n768_));
AOI22X1 AOI22X1_206 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_6_), .C(u3_u0_r2_6_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n772_));
AOI22X1 AOI22X1_207 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_7_), .C(u3_u0_r2_7_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n776_));
AOI22X1 AOI22X1_208 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_8_), .C(u3_u0_r2_8_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n780_));
AOI22X1 AOI22X1_209 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_9_), .C(u3_u0_r2_9_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n784_));
AOI22X1 AOI22X1_21 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n3810_));
AOI22X1 AOI22X1_210 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_10_), .C(u3_u0_r2_10_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n788_));
AOI22X1 AOI22X1_211 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_11_), .C(u3_u0_r2_11_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n792_));
AOI22X1 AOI22X1_212 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_12_), .C(u3_u0_r2_12_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n796_));
AOI22X1 AOI22X1_213 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_13_), .C(u3_u0_r2_13_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n800_));
AOI22X1 AOI22X1_214 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_14_), .C(u3_u0_r2_14_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n804_));
AOI22X1 AOI22X1_215 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_15_), .C(u3_u0_r2_15_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n808_));
AOI22X1 AOI22X1_216 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_16_), .C(u3_u0_r2_16_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n812_));
AOI22X1 AOI22X1_217 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_17_), .C(u3_u0_r2_17_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n816_));
AOI22X1 AOI22X1_218 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_18_), .C(u3_u0_r2_18_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n820_));
AOI22X1 AOI22X1_219 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_19_), .C(u3_u0_r2_19_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n824_));
AOI22X1 AOI22X1_22 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(u0_csc1_3_), .D(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n3817_));
AOI22X1 AOI22X1_220 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_20_), .C(u3_u0_r2_20_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n828_));
AOI22X1 AOI22X1_221 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_21_), .C(u3_u0_r2_21_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n832_));
AOI22X1 AOI22X1_222 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_22_), .C(u3_u0_r2_22_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n836_));
AOI22X1 AOI22X1_223 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_23_), .C(u3_u0_r2_23_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n840_));
AOI22X1 AOI22X1_224 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_24_), .C(u3_u0_r2_24_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n844_));
AOI22X1 AOI22X1_225 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_25_), .C(u3_u0_r2_25_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n848_));
AOI22X1 AOI22X1_226 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_26_), .C(u3_u0_r2_26_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n852_));
AOI22X1 AOI22X1_227 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_27_), .C(u3_u0_r2_27_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n856_));
AOI22X1 AOI22X1_228 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_28_), .C(u3_u0_r2_28_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n860_));
AOI22X1 AOI22X1_229 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_29_), .C(u3_u0_r2_29_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n864_));
AOI22X1 AOI22X1_23 ( .A(u0__abc_74894_new_n3701_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3818_));
AOI22X1 AOI22X1_230 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_30_), .C(u3_u0_r2_30_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n868_));
AOI22X1 AOI22X1_231 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_31_), .C(u3_u0_r2_31_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n872_));
AOI22X1 AOI22X1_232 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_32_), .C(u3_u0_r2_32_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n876_));
AOI22X1 AOI22X1_233 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_33_), .C(u3_u0_r2_33_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n880_));
AOI22X1 AOI22X1_234 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_34_), .C(u3_u0_r2_34_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n884_));
AOI22X1 AOI22X1_235 ( .A(u3_u0__abc_74260_new_n744_), .B(u3_u0_r1_35_), .C(u3_u0_r2_35_), .D(u3_u0__abc_74260_new_n747_), .Y(u3_u0__abc_74260_new_n888_));
AOI22X1 AOI22X1_236 ( .A(u4__abc_74770_new_n71_), .B(u4__abc_74770_new_n72_), .C(u4__abc_74770_new_n73_), .D(u4__abc_74770_new_n74_), .Y(u4__abc_74770_new_n75_));
AOI22X1 AOI22X1_237 ( .A(u4__abc_74770_new_n76_), .B(u4__abc_74770_new_n77_), .C(u4__abc_74770_new_n78_), .D(u4__abc_74770_new_n79_), .Y(u4__abc_74770_new_n80_));
AOI22X1 AOI22X1_238 ( .A(u4__abc_74770_new_n84_), .B(u4__abc_74770_new_n85_), .C(u4__abc_74770_new_n86_), .D(u4__abc_74770_new_n87_), .Y(u4__abc_74770_new_n88_));
AOI22X1 AOI22X1_239 ( .A(u4__abc_74770_new_n135_), .B(u4__abc_74770_new_n137_), .C(u4__abc_74770_new_n132_), .D(u4__0rfr_early_0_0_), .Y(u4__0ps_cnt_7_0__0_));
AOI22X1 AOI22X1_24 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3824_));
AOI22X1 AOI22X1_240 ( .A(u4__abc_74770_new_n144_), .B(u4__abc_74770_new_n145_), .C(u4__abc_74770_new_n132_), .D(u4__0rfr_early_0_0_), .Y(u4__0ps_cnt_7_0__2_));
AOI22X1 AOI22X1_241 ( .A(u4__abc_74770_new_n162_), .B(u4__abc_74770_new_n163_), .C(u4__abc_74770_new_n132_), .D(u4__0rfr_early_0_0_), .Y(u4__0ps_cnt_7_0__6_));
AOI22X1 AOI22X1_242 ( .A(u5__abc_78290_new_n844_), .B(u5__abc_78290_new_n455_), .C(u5__abc_78290_new_n838_), .D(u5__abc_78290_new_n839_), .Y(u5__abc_78290_new_n845_));
AOI22X1 AOI22X1_243 ( .A(u5__abc_78290_new_n1257_), .B(u5__abc_78290_new_n1613_), .C(u5__abc_78290_new_n1273_), .D(u5__abc_78290_new_n1611_), .Y(u5__abc_78290_new_n1614_));
AOI22X1 AOI22X1_244 ( .A(u5__abc_78290_new_n1262_), .B(u5__abc_78290_new_n1610_), .C(u5__abc_78290_new_n1621_), .D(u5__abc_78290_new_n1619_), .Y(u5__abc_78290_new_n1622_));
AOI22X1 AOI22X1_245 ( .A(u5__abc_78290_new_n1662_), .B(u5__abc_78290_new_n1659_), .C(1'h0), .D(u5__abc_78290_new_n1654_), .Y(u5__abc_78290_new_n1663_));
AOI22X1 AOI22X1_246 ( .A(u5__abc_78290_new_n1187_), .B(u5__abc_78290_new_n1316_), .C(u5__abc_78290_new_n1706_), .D(u5__abc_78290_new_n1699_), .Y(u5__abc_78290_new_n1707_));
AOI22X1 AOI22X1_247 ( .A(u5__abc_78290_new_n2223_), .B(u5__abc_78290_new_n2228_), .C(u5__abc_78290_new_n2227_), .D(u5__abc_78290_new_n2213_), .Y(u5__0timer_7_0__0_));
AOI22X1 AOI22X1_248 ( .A(u5__abc_78290_new_n2223_), .B(u5__abc_78290_new_n2230_), .C(u5__abc_78290_new_n2261_), .D(u5__abc_78290_new_n2258_), .Y(u5__0timer_7_0__1_));
AOI22X1 AOI22X1_249 ( .A(u5__abc_78290_new_n2281_), .B(u5__abc_78290_new_n2288_), .C(u5__abc_78290_new_n1187_), .D(u5__abc_78290_new_n2290_), .Y(u5__abc_78290_new_n2291_));
AOI22X1 AOI22X1_25 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3826_));
AOI22X1 AOI22X1_250 ( .A(u5__abc_78290_new_n2274_), .B(u5__abc_78290_new_n2164_), .C(u5__abc_78290_new_n2299_), .D(u5__abc_78290_new_n2298_), .Y(u5__abc_78290_new_n2300_));
AOI22X1 AOI22X1_251 ( .A(u5__abc_78290_new_n2223_), .B(u5__abc_78290_new_n2306_), .C(u5__abc_78290_new_n2305_), .D(u5__abc_78290_new_n2302_), .Y(u5__0timer_7_0__2_));
AOI22X1 AOI22X1_252 ( .A(u5__abc_78290_new_n2033_), .B(u5__abc_78290_new_n2310_), .C(u5__abc_78290_new_n2319_), .D(u5__abc_78290_new_n2320_), .Y(u5__abc_78290_new_n2321_));
AOI22X1 AOI22X1_253 ( .A(u5__abc_78290_new_n2145_), .B(u5__abc_78290_new_n2223_), .C(u5__abc_78290_new_n2327_), .D(u5__abc_78290_new_n2325_), .Y(u5__0timer_7_0__3_));
AOI22X1 AOI22X1_254 ( .A(u5__abc_78290_new_n1990_), .B(u5__abc_78290_new_n2417_), .C(u5__abc_78290_new_n2421_), .D(u5__abc_78290_new_n2208_), .Y(u5__abc_78290_new_n2422_));
AOI22X1 AOI22X1_255 ( .A(u5__abc_78290_new_n2225_), .B(u5__abc_78290_new_n2437_), .C(u5__abc_78290_new_n2451_), .D(u5__abc_78290_new_n2454_), .Y(u5__abc_78290_new_n2455_));
AOI22X1 AOI22X1_256 ( .A(u5__abc_78290_new_n2464_), .B(u5__abc_78290_new_n2367_), .C(u5__abc_78290_new_n2481_), .D(u5__abc_78290_new_n2477_), .Y(u5__0timer2_8_0__2_));
AOI22X1 AOI22X1_257 ( .A(u5__abc_78290_new_n2303_), .B(u5__abc_78290_new_n2437_), .C(u5__abc_78290_new_n2486_), .D(u5__abc_78290_new_n2490_), .Y(u5__abc_78290_new_n2491_));
AOI22X1 AOI22X1_258 ( .A(u5__abc_78290_new_n1472_), .B(u5__abc_78290_new_n2385_), .C(u5__abc_78290_new_n2507_), .D(u5__abc_78290_new_n2505_), .Y(u5__abc_78290_new_n2508_));
AOI22X1 AOI22X1_259 ( .A(u5__abc_78290_new_n2405_), .B(u5__abc_78290_new_n2520_), .C(u5__abc_78290_new_n2393_), .D(u5__abc_78290_new_n2406_), .Y(u5__abc_78290_new_n2521_));
AOI22X1 AOI22X1_26 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3827_));
AOI22X1 AOI22X1_260 ( .A(u5__abc_78290_new_n2652_), .B(u5__abc_78290_new_n2654_), .C(u5_state_4_), .D(u5__abc_78290_new_n2592_), .Y(u5__abc_78290_new_n2655_));
AOI22X1 AOI22X1_261 ( .A(u5__abc_78290_new_n2670_), .B(u5__abc_78290_new_n2674_), .C(u5__abc_78290_new_n2671_), .D(u5__abc_78290_new_n2675_), .Y(u5__abc_78290_new_n2676_));
AOI22X1 AOI22X1_262 ( .A(u5__abc_78290_new_n1456_), .B(u5__abc_78290_new_n2682_), .C(u5__abc_78290_new_n2684_), .D(u5__abc_78290_new_n1619_), .Y(u5__abc_78290_new_n2685_));
AOI22X1 AOI22X1_263 ( .A(u5__abc_78290_new_n2687_), .B(u5_state_8_), .C(row_same), .D(u5__abc_78290_new_n2652_), .Y(u5__abc_78290_new_n2688_));
AOI22X1 AOI22X1_264 ( .A(u5__abc_78290_new_n1375_), .B(u5__abc_78290_new_n1551_), .C(u5_cmd_asserted), .D(u5__abc_78290_new_n1268_), .Y(u5__abc_78290_new_n2710_));
AOI22X1 AOI22X1_265 ( .A(u5__abc_78290_new_n1551_), .B(u5__abc_78290_new_n2718_), .C(u5__abc_78290_new_n2717_), .D(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2719_));
AOI22X1 AOI22X1_266 ( .A(u5__abc_78290_new_n2629_), .B(u5__abc_78290_new_n2723_), .C(u5__abc_78290_new_n2722_), .D(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2724_));
AOI22X1 AOI22X1_267 ( .A(u5__abc_78290_new_n2697_), .B(u5__abc_78290_new_n2743_), .C(u5__abc_78290_new_n763_), .D(u5__abc_78290_new_n2742_), .Y(u5__abc_78290_new_n2744_));
AOI22X1 AOI22X1_268 ( .A(u5__abc_78290_new_n2069_), .B(u5__abc_78290_new_n2746_), .C(u5__abc_78290_new_n2744_), .D(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2747_));
AOI22X1 AOI22X1_269 ( .A(u5__abc_78290_new_n1554_), .B(u5__abc_78290_new_n2779_), .C(u5__abc_78290_new_n2776_), .D(u5__abc_78290_new_n2777_), .Y(u5__abc_78290_new_n2780_));
AOI22X1 AOI22X1_27 ( .A(u0__abc_74894_new_n3713_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3830_));
AOI22X1 AOI22X1_270 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1221_), .C(u5__abc_78290_new_n2805_), .D(u5__abc_78290_new_n1982_), .Y(u5__abc_78290_new_n2806_));
AOI22X1 AOI22X1_271 ( .A(u5__abc_78290_new_n1200_), .B(u5__abc_78290_new_n2810_), .C(u5__abc_78290_new_n2809_), .D(u5__abc_78290_new_n1982_), .Y(u5__abc_78290_new_n2811_));
AOI22X1 AOI22X1_272 ( .A(u5__abc_78290_new_n500_), .B(u5__abc_78290_new_n1375_), .C(u5__abc_78290_new_n594_), .D(u5__abc_78290_new_n505_), .Y(u5__abc_78290_new_n2816_));
AOI22X1 AOI22X1_273 ( .A(u5__abc_78290_new_n1197_), .B(u5__abc_78290_new_n2826_), .C(u5__abc_78290_new_n2827_), .D(u5__abc_78290_new_n2618_), .Y(u5__abc_78290_new_n2828_));
AOI22X1 AOI22X1_274 ( .A(u5__abc_78290_new_n1361_), .B(u5__abc_78290_new_n2886_), .C(u5__abc_78290_new_n2887_), .D(u5__abc_78290_new_n1380_), .Y(u5__abc_78290_new_n2888_));
AOI22X1 AOI22X1_275 ( .A(u5__abc_78290_new_n2440_), .B(u5__abc_78290_new_n2893_), .C(u5_state_44_), .D(u5__abc_78290_new_n2659_), .Y(u5__abc_78290_new_n2894_));
AOI22X1 AOI22X1_276 ( .A(u5__abc_78290_new_n2578_), .B(u5__abc_78290_new_n2905_), .C(u5_state_47_), .D(u5__abc_78290_new_n2592_), .Y(u5__abc_78290_new_n2906_));
AOI22X1 AOI22X1_277 ( .A(u5__abc_78290_new_n632_), .B(u5__abc_78290_new_n2912_), .C(u5__abc_78290_new_n1441_), .D(u5__abc_78290_new_n2584_), .Y(u5_next_state_49_));
AOI22X1 AOI22X1_278 ( .A(u5__abc_78290_new_n1139_), .B(u5__abc_78290_new_n1142_), .C(u5__abc_78290_new_n2565_), .D(u5__abc_78290_new_n2914_), .Y(u5__abc_78290_new_n2915_));
AOI22X1 AOI22X1_279 ( .A(u5__abc_78290_new_n619_), .B(u5__abc_78290_new_n2917_), .C(u5__abc_78290_new_n1495_), .D(u5__abc_78290_new_n2584_), .Y(u5_next_state_51_));
AOI22X1 AOI22X1_28 ( .A(u0__abc_74894_new_n3749_), .B(u0_csc_mask_4_), .C(\poc_o[4] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3834_));
AOI22X1 AOI22X1_280 ( .A(u5__abc_78290_new_n2218_), .B(u5__abc_78290_new_n2927_), .C(u5__abc_78290_new_n2565_), .D(u5__abc_78290_new_n2926_), .Y(u5__abc_78290_new_n2928_));
AOI22X1 AOI22X1_281 ( .A(u5__abc_78290_new_n2697_), .B(u5__abc_78290_new_n2935_), .C(u5__abc_78290_new_n976_), .D(u5__abc_78290_new_n2742_), .Y(u5__abc_78290_new_n2936_));
AOI22X1 AOI22X1_282 ( .A(u3_wb_read_go), .B(u5__abc_78290_new_n2937_), .C(u5__abc_78290_new_n2936_), .D(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2938_));
AOI22X1 AOI22X1_283 ( .A(u5__abc_78290_new_n2949_), .B(u5__abc_78290_new_n2960_), .C(u5__abc_78290_new_n1325_), .D(u5__abc_78290_new_n1517_), .Y(u5__abc_78290_new_n2961_));
AOI22X1 AOI22X1_284 ( .A(u5__abc_78290_new_n2949_), .B(u5__abc_78290_new_n2964_), .C(u5_wb_wait), .D(u5__abc_78290_new_n1517_), .Y(u5__abc_78290_new_n2965_));
AOI22X1 AOI22X1_285 ( .A(u5__abc_78290_new_n1616_), .B(u5__abc_78290_new_n2974_), .C(u5__abc_78290_new_n2973_), .D(u5__abc_78290_new_n2976_), .Y(u5__abc_78290_new_n2977_));
AOI22X1 AOI22X1_286 ( .A(u5__abc_78290_new_n1065_), .B(u5__abc_78290_new_n2979_), .C(u5__abc_78290_new_n1615_), .D(u5__abc_78290_new_n2584_), .Y(u5_next_state_62_));
AOI22X1 AOI22X1_287 ( .A(u5__abc_78290_new_n2975_), .B(u5__abc_78290_new_n2197_), .C(u5_state_65_), .D(u5__abc_78290_new_n2659_), .Y(u5__abc_78290_new_n2991_));
AOI22X1 AOI22X1_288 ( .A(u5__abc_78290_new_n433_), .B(u5__abc_78290_new_n440_), .C(u5_wb_wait), .D(u5__abc_78290_new_n3133_), .Y(u5__abc_78290_new_n3134_));
AOI22X1 AOI22X1_29 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_4_), .C(u0_tms0_4_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3836_));
AOI22X1 AOI22X1_3 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n3721_));
AOI22X1 AOI22X1_30 ( .A(u0__abc_74894_new_n3802_), .B(u0_tms1_5_), .C(u0_csc0_5_), .D(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n3851_));
AOI22X1 AOI22X1_31 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n3853_));
AOI22X1 AOI22X1_32 ( .A(u0_csc1_5_), .B(u0__abc_74894_new_n3816_), .C(\poc_o[5] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3858_));
AOI22X1 AOI22X1_33 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n3859_));
AOI22X1 AOI22X1_34 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3865_));
AOI22X1 AOI22X1_35 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3867_));
AOI22X1 AOI22X1_36 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3868_));
AOI22X1 AOI22X1_37 ( .A(u0__abc_74894_new_n3713_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3871_));
AOI22X1 AOI22X1_38 ( .A(u0__abc_74894_new_n3749_), .B(u0_csc_mask_6_), .C(\poc_o[6] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3875_));
AOI22X1 AOI22X1_39 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_6_), .C(u0_tms0_6_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3877_));
AOI22X1 AOI22X1_4 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_0_), .C(u0_tms0_0_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3738_));
AOI22X1 AOI22X1_40 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3881_));
AOI22X1 AOI22X1_41 ( .A(u0__abc_74894_new_n3699_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3882_));
AOI22X1 AOI22X1_42 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3894_));
AOI22X1 AOI22X1_43 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3902_));
AOI22X1 AOI22X1_44 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3904_));
AOI22X1 AOI22X1_45 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3905_));
AOI22X1 AOI22X1_46 ( .A(u0__abc_74894_new_n3713_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3908_));
AOI22X1 AOI22X1_47 ( .A(u0__abc_74894_new_n3749_), .B(u0_csc_mask_8_), .C(\poc_o[8] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3912_));
AOI22X1 AOI22X1_48 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_9_), .C(u0_tms0_9_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3921_));
AOI22X1 AOI22X1_49 ( .A(u0__abc_74894_new_n3751_), .B(\poc_o[9] ), .C(u0_tms1_9_), .D(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n3922_));
AOI22X1 AOI22X1_5 ( .A(u0__abc_74894_new_n3749_), .B(u0_csc_mask_0_), .C(\poc_o[0] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3752_));
AOI22X1 AOI22X1_50 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n3927_));
AOI22X1 AOI22X1_51 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n3929_));
AOI22X1 AOI22X1_52 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(u0_csc1_9_), .D(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n3934_));
AOI22X1 AOI22X1_53 ( .A(u0__abc_74894_new_n3701_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3935_));
AOI22X1 AOI22X1_54 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3941_));
AOI22X1 AOI22X1_55 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3943_));
AOI22X1 AOI22X1_56 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3944_));
AOI22X1 AOI22X1_57 ( .A(u0__abc_74894_new_n3713_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3947_));
AOI22X1 AOI22X1_58 ( .A(u0__abc_74894_new_n3749_), .B(u0_csc_mask_10_), .C(\poc_o[10] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3951_));
AOI22X1 AOI22X1_59 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_10_), .C(u0_tms0_10_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3953_));
AOI22X1 AOI22X1_6 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3756_));
AOI22X1 AOI22X1_60 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3960_));
AOI22X1 AOI22X1_61 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3964_));
AOI22X1 AOI22X1_62 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_11_), .C(u0_tms0_11_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3967_));
AOI22X1 AOI22X1_63 ( .A(u0_csc1_11_), .B(u0__abc_74894_new_n3816_), .C(u0_tms1_11_), .D(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n3968_));
AOI22X1 AOI22X1_64 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n3972_));
AOI22X1 AOI22X1_65 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3979_));
AOI22X1 AOI22X1_66 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3983_));
AOI22X1 AOI22X1_67 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_12_), .C(u0_tms0_12_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3986_));
AOI22X1 AOI22X1_68 ( .A(u0_csc1_12_), .B(u0__abc_74894_new_n3816_), .C(u0_tms1_12_), .D(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n3987_));
AOI22X1 AOI22X1_69 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n3991_));
AOI22X1 AOI22X1_7 ( .A(u0__abc_74894_new_n3699_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3757_));
AOI22X1 AOI22X1_70 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4009_));
AOI22X1 AOI22X1_71 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4031_));
AOI22X1 AOI22X1_72 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(\poc_o[16] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4063_));
AOI22X1 AOI22X1_73 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4071_));
AOI22X1 AOI22X1_74 ( .A(u0__abc_74894_new_n3745_), .B(1'h0), .C(u0_tms1_16_), .D(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4075_));
AOI22X1 AOI22X1_75 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4139_));
AOI22X1 AOI22X1_76 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4150_));
AOI22X1 AOI22X1_77 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4154_));
AOI22X1 AOI22X1_78 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_20_), .C(u0_tms0_20_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4157_));
AOI22X1 AOI22X1_79 ( .A(u0_csc1_20_), .B(u0__abc_74894_new_n3816_), .C(u0_tms1_20_), .D(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4158_));
AOI22X1 AOI22X1_8 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3759_));
AOI22X1 AOI22X1_80 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4162_));
AOI22X1 AOI22X1_81 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4181_));
AOI22X1 AOI22X1_82 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4192_));
AOI22X1 AOI22X1_83 ( .A(u0__abc_74894_new_n3741_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4196_));
AOI22X1 AOI22X1_84 ( .A(u0__abc_74894_new_n3734_), .B(u0_csc0_22_), .C(u0_tms0_22_), .D(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4199_));
AOI22X1 AOI22X1_85 ( .A(u0_csc1_22_), .B(u0__abc_74894_new_n3816_), .C(u0_tms1_22_), .D(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4200_));
AOI22X1 AOI22X1_86 ( .A(u0__abc_74894_new_n3717_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4204_));
AOI22X1 AOI22X1_87 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(\poc_o[23] ), .D(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4210_));
AOI22X1 AOI22X1_88 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4218_));
AOI22X1 AOI22X1_89 ( .A(u0__abc_74894_new_n3745_), .B(1'h0), .C(u0_tms1_23_), .D(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4222_));
AOI22X1 AOI22X1_9 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .C(1'h0), .D(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3760_));
AOI22X1 AOI22X1_90 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .C(1'h0), .D(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4274_));
AOI22X1 AOI22X1_91 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4363_));
AOI22X1 AOI22X1_92 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4364_));
AOI22X1 AOI22X1_93 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4387_));
AOI22X1 AOI22X1_94 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4388_));
AOI22X1 AOI22X1_95 ( .A(u0__abc_74894_new_n3693_), .B(1'h0), .C(1'h0), .D(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4411_));
AOI22X1 AOI22X1_96 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .C(1'h0), .D(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4412_));
AOI22X1 AOI22X1_97 ( .A(u1__abc_72801_new_n278_), .B(u1__abc_72801_new_n279_), .C(u1__abc_72801_new_n280_), .D(u1__abc_72801_new_n281_), .Y(u1__abc_72801_new_n282_));
AOI22X1 AOI22X1_98 ( .A(\wb_addr_i[10] ), .B(page_size_8_), .C(\wb_addr_i[11] ), .D(page_size_9_), .Y(u1__abc_72801_new_n284_));
AOI22X1 AOI22X1_99 ( .A(u1__abc_72801_new_n280_), .B(u1__abc_72801_new_n265_), .C(u1__abc_72801_new_n262_), .D(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n293_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_i), .D(mem_ack), .Q(mem_ack_r));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_i), .D(u0__0poc_31_0__6_), .Q(\poc_o[6] ));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__26_), .Q(u0_csc0_26_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__27_), .Q(u0_csc0_27_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__28_), .Q(u0_csc0_28_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__29_), .Q(u0_csc0_29_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__30_), .Q(u0_csc0_30_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__31_), .Q(u0_csc0_31_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_i), .D(\wb_addr_i[2] ), .Q(u0_u0_addr_r_2_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_i), .D(\wb_addr_i[3] ), .Q(u0_u0_addr_r_3_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_i), .D(\wb_addr_i[4] ), .Q(u0_u0_addr_r_4_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_i), .D(\wb_addr_i[5] ), .Q(u0_u0_addr_r_5_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_i), .D(u0__0poc_31_0__7_), .Q(\poc_o[7] ));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_i), .D(\wb_addr_i[6] ), .Q(u0_u0_addr_r_6_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__0_), .Q(u0_tms1_0_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__1_), .Q(u0_tms1_1_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__2_), .Q(u0_tms1_2_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__3_), .Q(u0_tms1_3_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__4_), .Q(u0_tms1_4_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__5_), .Q(u0_tms1_5_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__6_), .Q(u0_tms1_6_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__7_), .Q(u0_tms1_7_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__8_), .Q(u0_tms1_8_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_i), .D(u0__0poc_31_0__8_), .Q(\poc_o[8] ));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__9_), .Q(u0_tms1_9_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__10_), .Q(u0_tms1_10_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__11_), .Q(u0_tms1_11_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__12_), .Q(u0_tms1_12_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__13_), .Q(u0_tms1_13_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__14_), .Q(u0_tms1_14_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__15_), .Q(u0_tms1_15_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__16_), .Q(u0_tms1_16_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__17_), .Q(u0_tms1_17_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__18_), .Q(u0_tms1_18_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_i), .D(u0__0poc_31_0__9_), .Q(\poc_o[9] ));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__19_), .Q(u0_tms1_19_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__20_), .Q(u0_tms1_20_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__21_), .Q(u0_tms1_21_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__22_), .Q(u0_tms1_22_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__23_), .Q(u0_tms1_23_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__24_), .Q(u0_tms1_24_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__25_), .Q(u0_tms1_25_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__26_), .Q(u0_tms1_26_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__27_), .Q(u0_tms1_27_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__28_), .Q(u0_tms1_28_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_i), .D(u0__0poc_31_0__10_), .Q(\poc_o[10] ));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__29_), .Q(u0_tms1_29_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__30_), .Q(u0_tms1_30_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_i), .D(u0_u1__0tms_31_0__31_), .Q(u0_tms1_31_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__0_), .Q(u0_csc1_0_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__1_), .Q(u0_csc1_1_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__2_), .Q(u0_csc1_2_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__3_), .Q(u0_csc1_3_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__4_), .Q(u0_csc1_4_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__5_), .Q(u0_csc1_5_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__6_), .Q(u0_csc1_6_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_i), .D(u0__0poc_31_0__11_), .Q(\poc_o[11] ));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__7_), .Q(u0_csc1_7_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__8_), .Q(u0_csc1_8_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__9_), .Q(u0_csc1_9_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__10_), .Q(u0_csc1_10_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__11_), .Q(u0_csc1_11_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__12_), .Q(u0_csc1_12_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__13_), .Q(u0_csc1_13_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__14_), .Q(u0_csc1_14_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__15_), .Q(u0_csc1_15_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__16_), .Q(u0_csc1_16_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_i), .D(u0__0poc_31_0__12_), .Q(\poc_o[12] ));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__17_), .Q(u0_csc1_17_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__18_), .Q(u0_csc1_18_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__19_), .Q(u0_csc1_19_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__20_), .Q(u0_csc1_20_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__21_), .Q(u0_csc1_21_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__22_), .Q(u0_csc1_22_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__23_), .Q(u0_csc1_23_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__24_), .Q(u0_csc1_24_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__25_), .Q(u0_csc1_25_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__26_), .Q(u0_csc1_26_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_i), .D(u0__0poc_31_0__13_), .Q(\poc_o[13] ));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__27_), .Q(u0_csc1_27_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__28_), .Q(u0_csc1_28_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__29_), .Q(u0_csc1_29_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__30_), .Q(u0_csc1_30_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_i), .D(u0_u1__0csc_31_0__31_), .Q(u0_csc1_31_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_i), .D(\wb_addr_i[2] ), .Q(u0_u1_addr_r_2_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_i), .D(\wb_addr_i[3] ), .Q(u0_u1_addr_r_3_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_i), .D(\wb_addr_i[4] ), .Q(u0_u1_addr_r_4_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_i), .D(\wb_addr_i[5] ), .Q(u0_u1_addr_r_5_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_i), .D(\wb_addr_i[6] ), .Q(u0_u1_addr_r_6_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_i), .D(u0__0poc_31_0__14_), .Q(\poc_o[14] ));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_i), .D(u1__0bank_adr_1_0__0_), .Q(bank_adr_0_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_i), .D(u1__0bank_adr_1_0__1_), .Q(bank_adr_1_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_i), .D(u1__0row_adr_12_0__0_), .Q(row_adr_0_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_i), .D(u1__0row_adr_12_0__1_), .Q(row_adr_1_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_i), .D(u1__0row_adr_12_0__2_), .Q(row_adr_2_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_i), .D(u1__0row_adr_12_0__3_), .Q(row_adr_3_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_i), .D(u1__0row_adr_12_0__4_), .Q(row_adr_4_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_i), .D(u1__0row_adr_12_0__5_), .Q(row_adr_5_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_i), .D(u1__0row_adr_12_0__6_), .Q(row_adr_6_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_i), .D(u1__0row_adr_12_0__7_), .Q(row_adr_7_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_i), .D(u0__0poc_31_0__15_), .Q(\poc_o[15] ));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_i), .D(u1__0row_adr_12_0__8_), .Q(row_adr_8_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_i), .D(u1__0row_adr_12_0__9_), .Q(row_adr_9_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_i), .D(u1__0row_adr_12_0__10_), .Q(row_adr_10_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_i), .D(u1__0row_adr_12_0__11_), .Q(row_adr_11_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_i), .D(u1__0row_adr_12_0__12_), .Q(row_adr_12_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_i), .D(u1__0col_adr_9_0__0_), .Q(u1_col_adr_0_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_i), .D(u1__0col_adr_9_0__1_), .Q(u1_col_adr_1_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_i), .D(u1__0col_adr_9_0__2_), .Q(u1_col_adr_2_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_i), .D(u1__0col_adr_9_0__3_), .Q(u1_col_adr_3_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_i), .D(u1__0col_adr_9_0__4_), .Q(u1_col_adr_4_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_i), .D(lmr_ack), .Q(u0_lmr_ack_r));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_i), .D(u0__0poc_31_0__16_), .Q(\poc_o[16] ));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_i), .D(u1__0col_adr_9_0__5_), .Q(u1_col_adr_5_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_i), .D(u1__0col_adr_9_0__6_), .Q(u1_col_adr_6_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_i), .D(u1__0col_adr_9_0__7_), .Q(u1_col_adr_7_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_i), .D(u1__0col_adr_9_0__8_), .Q(u1_col_adr_8_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_i), .D(u1__0col_adr_9_0__9_), .Q(u1_col_adr_9_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__0_), .Q(u1_acs_addr_0_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__1_), .Q(u1_acs_addr_1_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__2_), .Q(u1_acs_addr_2_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__3_), .Q(u1_acs_addr_3_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__4_), .Q(u1_acs_addr_4_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_i), .D(u0__0poc_31_0__17_), .Q(\poc_o[17] ));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__5_), .Q(u1_acs_addr_5_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__6_), .Q(u1_acs_addr_6_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__7_), .Q(u1_acs_addr_7_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__8_), .Q(u1_acs_addr_8_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__9_), .Q(u1_acs_addr_9_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__10_), .Q(u1_acs_addr_10_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__11_), .Q(u1_acs_addr_11_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__12_), .Q(u1_acs_addr_12_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__13_), .Q(u1_acs_addr_13_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__14_), .Q(u1_acs_addr_14_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_i), .D(u0__0poc_31_0__18_), .Q(\poc_o[18] ));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__15_), .Q(u1_acs_addr_15_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__16_), .Q(u1_acs_addr_16_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__17_), .Q(u1_acs_addr_17_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__18_), .Q(u1_acs_addr_18_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__19_), .Q(u1_acs_addr_19_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__20_), .Q(u1_acs_addr_20_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__21_), .Q(u1_acs_addr_21_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__22_), .Q(u1_acs_addr_22_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_i), .D(u1__0acs_addr_23_0__23_), .Q(u1_acs_addr_23_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__0_), .Q(u1_sram_addr_0_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_i), .D(u0__0poc_31_0__19_), .Q(\poc_o[19] ));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__1_), .Q(u1_sram_addr_1_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__2_), .Q(u1_sram_addr_2_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__3_), .Q(u1_sram_addr_3_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__4_), .Q(u1_sram_addr_4_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__5_), .Q(u1_sram_addr_5_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__6_), .Q(u1_sram_addr_6_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__7_), .Q(u1_sram_addr_7_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__8_), .Q(u1_sram_addr_8_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__9_), .Q(u1_sram_addr_9_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__10_), .Q(u1_sram_addr_10_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_i), .D(u0__0poc_31_0__20_), .Q(\poc_o[20] ));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__11_), .Q(u1_sram_addr_11_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__12_), .Q(u1_sram_addr_12_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__13_), .Q(u1_sram_addr_13_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__14_), .Q(u1_sram_addr_14_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__15_), .Q(u1_sram_addr_15_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__16_), .Q(u1_sram_addr_16_));
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__17_), .Q(u1_sram_addr_17_));
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__18_), .Q(u1_sram_addr_18_));
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__19_), .Q(u1_sram_addr_19_));
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__20_), .Q(u1_sram_addr_20_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_i), .D(u0__0poc_31_0__21_), .Q(\poc_o[21] ));
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__21_), .Q(u1_sram_addr_21_));
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__22_), .Q(u1_sram_addr_22_));
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_i), .D(u1__0sram_addr_23_0__23_), .Q(u1_sram_addr_23_));
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__0_), .Q(u1_acs_addr_pl1_0_));
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__1_), .Q(u1_acs_addr_pl1_1_));
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__2_), .Q(u1_acs_addr_pl1_2_));
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__3_), .Q(u1_acs_addr_pl1_3_));
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__4_), .Q(u1_acs_addr_pl1_4_));
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__5_), .Q(u1_acs_addr_pl1_5_));
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__6_), .Q(u1_acs_addr_pl1_6_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_i), .D(u0__0poc_31_0__22_), .Q(\poc_o[22] ));
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__7_), .Q(u1_acs_addr_pl1_7_));
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__8_), .Q(u1_acs_addr_pl1_8_));
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__9_), .Q(u1_acs_addr_pl1_9_));
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__10_), .Q(u1_acs_addr_pl1_10_));
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__11_), .Q(u1_acs_addr_pl1_11_));
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_i), .D(u1_u0__0out_r_12_0__12_), .Q(u1_u0_inc_next));
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_i), .D(u2__0row_same_0_0_), .Q(row_same));
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_i), .D(u2__0bank_open_0_0_), .Q(bank_open));
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__0_), .Q(u2_u0_b3_last_row_0_));
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__1_), .Q(u2_u0_b3_last_row_1_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_i), .D(u0__0poc_31_0__23_), .Q(\poc_o[23] ));
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__2_), .Q(u2_u0_b3_last_row_2_));
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__3_), .Q(u2_u0_b3_last_row_3_));
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__4_), .Q(u2_u0_b3_last_row_4_));
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__5_), .Q(u2_u0_b3_last_row_5_));
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__6_), .Q(u2_u0_b3_last_row_6_));
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__7_), .Q(u2_u0_b3_last_row_7_));
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__8_), .Q(u2_u0_b3_last_row_8_));
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__9_), .Q(u2_u0_b3_last_row_9_));
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__10_), .Q(u2_u0_b3_last_row_10_));
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__11_), .Q(u2_u0_b3_last_row_11_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_i), .D(u0__0poc_31_0__24_), .Q(\poc_o[24] ));
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_i), .D(u2_u0__0b3_last_row_12_0__12_), .Q(u2_u0_b3_last_row_12_));
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__0_), .Q(u2_u0_b2_last_row_0_));
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__1_), .Q(u2_u0_b2_last_row_1_));
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__2_), .Q(u2_u0_b2_last_row_2_));
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__3_), .Q(u2_u0_b2_last_row_3_));
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__4_), .Q(u2_u0_b2_last_row_4_));
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__5_), .Q(u2_u0_b2_last_row_5_));
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__6_), .Q(u2_u0_b2_last_row_6_));
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__7_), .Q(u2_u0_b2_last_row_7_));
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__8_), .Q(u2_u0_b2_last_row_8_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_i), .D(u0__0poc_31_0__25_), .Q(\poc_o[25] ));
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__9_), .Q(u2_u0_b2_last_row_9_));
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__10_), .Q(u2_u0_b2_last_row_10_));
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__11_), .Q(u2_u0_b2_last_row_11_));
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_i), .D(u2_u0__0b2_last_row_12_0__12_), .Q(u2_u0_b2_last_row_12_));
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__0_), .Q(u2_u0_b1_last_row_0_));
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__1_), .Q(u2_u0_b1_last_row_1_));
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__2_), .Q(u2_u0_b1_last_row_2_));
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__3_), .Q(u2_u0_b1_last_row_3_));
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__4_), .Q(u2_u0_b1_last_row_4_));
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__5_), .Q(u2_u0_b1_last_row_5_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_i), .D(init_ack), .Q(u0_init_ack_r));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_i), .D(u0__0poc_31_0__26_), .Q(\poc_o[26] ));
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__6_), .Q(u2_u0_b1_last_row_6_));
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__7_), .Q(u2_u0_b1_last_row_7_));
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__8_), .Q(u2_u0_b1_last_row_8_));
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__9_), .Q(u2_u0_b1_last_row_9_));
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__10_), .Q(u2_u0_b1_last_row_10_));
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__11_), .Q(u2_u0_b1_last_row_11_));
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_i), .D(u2_u0__0b1_last_row_12_0__12_), .Q(u2_u0_b1_last_row_12_));
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__0_), .Q(u2_u0_b0_last_row_0_));
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__1_), .Q(u2_u0_b0_last_row_1_));
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__2_), .Q(u2_u0_b0_last_row_2_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_i), .D(u0__0poc_31_0__27_), .Q(\poc_o[27] ));
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__3_), .Q(u2_u0_b0_last_row_3_));
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__4_), .Q(u2_u0_b0_last_row_4_));
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__5_), .Q(u2_u0_b0_last_row_5_));
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__6_), .Q(u2_u0_b0_last_row_6_));
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__7_), .Q(u2_u0_b0_last_row_7_));
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__8_), .Q(u2_u0_b0_last_row_8_));
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__9_), .Q(u2_u0_b0_last_row_9_));
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__10_), .Q(u2_u0_b0_last_row_10_));
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__11_), .Q(u2_u0_b0_last_row_11_));
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_i), .D(u2_u0__0b0_last_row_12_0__12_), .Q(u2_u0_b0_last_row_12_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_i), .D(u0__0poc_31_0__28_), .Q(\poc_o[28] ));
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__0_), .Q(u2_u1_b3_last_row_0_));
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__1_), .Q(u2_u1_b3_last_row_1_));
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__2_), .Q(u2_u1_b3_last_row_2_));
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__3_), .Q(u2_u1_b3_last_row_3_));
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__4_), .Q(u2_u1_b3_last_row_4_));
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__5_), .Q(u2_u1_b3_last_row_5_));
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__6_), .Q(u2_u1_b3_last_row_6_));
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__7_), .Q(u2_u1_b3_last_row_7_));
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__8_), .Q(u2_u1_b3_last_row_8_));
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__9_), .Q(u2_u1_b3_last_row_9_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_i), .D(u0__0poc_31_0__29_), .Q(\poc_o[29] ));
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__10_), .Q(u2_u1_b3_last_row_10_));
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__11_), .Q(u2_u1_b3_last_row_11_));
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_i), .D(u2_u1__0b3_last_row_12_0__12_), .Q(u2_u1_b3_last_row_12_));
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__0_), .Q(u2_u1_b2_last_row_0_));
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__1_), .Q(u2_u1_b2_last_row_1_));
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__2_), .Q(u2_u1_b2_last_row_2_));
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__3_), .Q(u2_u1_b2_last_row_3_));
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__4_), .Q(u2_u1_b2_last_row_4_));
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__5_), .Q(u2_u1_b2_last_row_5_));
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__6_), .Q(u2_u1_b2_last_row_6_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_i), .D(u0__0poc_31_0__30_), .Q(\poc_o[30] ));
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__7_), .Q(u2_u1_b2_last_row_7_));
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__8_), .Q(u2_u1_b2_last_row_8_));
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__9_), .Q(u2_u1_b2_last_row_9_));
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__10_), .Q(u2_u1_b2_last_row_10_));
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__11_), .Q(u2_u1_b2_last_row_11_));
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_i), .D(u2_u1__0b2_last_row_12_0__12_), .Q(u2_u1_b2_last_row_12_));
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__0_), .Q(u2_u1_b1_last_row_0_));
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__1_), .Q(u2_u1_b1_last_row_1_));
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__2_), .Q(u2_u1_b1_last_row_2_));
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__3_), .Q(u2_u1_b1_last_row_3_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_i), .D(u0__0poc_31_0__31_), .Q(\poc_o[31] ));
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__4_), .Q(u2_u1_b1_last_row_4_));
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__5_), .Q(u2_u1_b1_last_row_5_));
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__6_), .Q(u2_u1_b1_last_row_6_));
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__7_), .Q(u2_u1_b1_last_row_7_));
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__8_), .Q(u2_u1_b1_last_row_8_));
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__9_), .Q(u2_u1_b1_last_row_9_));
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__10_), .Q(u2_u1_b1_last_row_10_));
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__11_), .Q(u2_u1_b1_last_row_11_));
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_i), .D(u2_u1__0b1_last_row_12_0__12_), .Q(u2_u1_b1_last_row_12_));
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__0_), .Q(u2_u1_b0_last_row_0_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_i), .D(mc_sts_ir), .Q(u0_csr_0_));
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__1_), .Q(u2_u1_b0_last_row_1_));
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__2_), .Q(u2_u1_b0_last_row_2_));
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__3_), .Q(u2_u1_b0_last_row_3_));
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__4_), .Q(u2_u1_b0_last_row_4_));
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__5_), .Q(u2_u1_b0_last_row_5_));
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__6_), .Q(u2_u1_b0_last_row_6_));
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__7_), .Q(u2_u1_b0_last_row_7_));
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__8_), .Q(u2_u1_b0_last_row_8_));
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__9_), .Q(u2_u1_b0_last_row_9_));
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__10_), .Q(u2_u1_b0_last_row_10_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_i), .D(\wb_addr_i[2] ), .Q(u0_wb_addr_r_2_));
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__11_), .Q(u2_u1_b0_last_row_11_));
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_i), .D(u2_u1__0b0_last_row_12_0__12_), .Q(u2_u1_b0_last_row_12_));
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_i), .D(u3__0mc_dp_o_3_0__0_), .Q(mc_dp_od_0_));
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_i), .D(u3__0mc_dp_o_3_0__1_), .Q(mc_dp_od_1_));
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_i), .D(u3__0mc_dp_o_3_0__2_), .Q(mc_dp_od_2_));
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_i), .D(u3__0mc_dp_o_3_0__3_), .Q(mc_dp_od_3_));
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_i), .D(u3__0byte2_7_0__0_), .Q(u3_byte2_0_));
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_i), .D(u3__0byte2_7_0__1_), .Q(u3_byte2_1_));
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_i), .D(u3__0byte2_7_0__2_), .Q(u3_byte2_2_));
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_i), .D(u3__0byte2_7_0__3_), .Q(u3_byte2_3_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_i), .D(\wb_addr_i[3] ), .Q(u0_wb_addr_r_3_));
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_i), .D(u3__0byte2_7_0__4_), .Q(u3_byte2_4_));
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_i), .D(u3__0byte2_7_0__5_), .Q(u3_byte2_5_));
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_i), .D(u3__0byte2_7_0__6_), .Q(u3_byte2_6_));
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_i), .D(u3__0byte2_7_0__7_), .Q(u3_byte2_7_));
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_i), .D(u3__0byte1_7_0__0_), .Q(u3_byte1_0_));
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_i), .D(u3__0byte1_7_0__1_), .Q(u3_byte1_1_));
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_i), .D(u3__0byte1_7_0__2_), .Q(u3_byte1_2_));
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_i), .D(u3__0byte1_7_0__3_), .Q(u3_byte1_3_));
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_i), .D(u3__0byte1_7_0__4_), .Q(u3_byte1_4_));
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_i), .D(u3__0byte1_7_0__5_), .Q(u3_byte1_5_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_i), .D(\wb_addr_i[4] ), .Q(u0_wb_addr_r_4_));
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_i), .D(u3__0byte1_7_0__6_), .Q(u3_byte1_6_));
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_i), .D(u3__0byte1_7_0__7_), .Q(u3_byte1_7_));
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_i), .D(u3__0byte0_7_0__0_), .Q(u3_byte0_0_));
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_i), .D(u3__0byte0_7_0__1_), .Q(u3_byte0_1_));
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_i), .D(u3__0byte0_7_0__2_), .Q(u3_byte0_2_));
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_i), .D(u3__0byte0_7_0__3_), .Q(u3_byte0_3_));
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_i), .D(u3__0byte0_7_0__4_), .Q(u3_byte0_4_));
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_i), .D(u3__0byte0_7_0__5_), .Q(u3_byte0_5_));
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_i), .D(u3__0byte0_7_0__6_), .Q(u3_byte0_6_));
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_i), .D(u3__0byte0_7_0__7_), .Q(u3_byte0_7_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_i), .D(u0__0poc_31_0__0_), .Q(\poc_o[0] ));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_i), .D(\wb_addr_i[5] ), .Q(u0_wb_addr_r_5_));
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__0_), .Q(mc_data_od_0_));
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__1_), .Q(mc_data_od_1_));
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__2_), .Q(mc_data_od_2_));
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__3_), .Q(mc_data_od_3_));
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__4_), .Q(mc_data_od_4_));
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__5_), .Q(mc_data_od_5_));
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__6_), .Q(mc_data_od_6_));
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__7_), .Q(mc_data_od_7_));
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__8_), .Q(mc_data_od_8_));
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__9_), .Q(mc_data_od_9_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_i), .D(\wb_addr_i[6] ), .Q(u0_wb_addr_r_6_));
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__10_), .Q(mc_data_od_10_));
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__11_), .Q(mc_data_od_11_));
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__12_), .Q(mc_data_od_12_));
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__13_), .Q(mc_data_od_13_));
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__14_), .Q(mc_data_od_14_));
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__15_), .Q(mc_data_od_15_));
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__16_), .Q(mc_data_od_16_));
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__17_), .Q(mc_data_od_17_));
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__18_), .Q(mc_data_od_18_));
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__19_), .Q(mc_data_od_19_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__0_), .Q(u0_tms0_0_));
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__20_), .Q(mc_data_od_20_));
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__21_), .Q(mc_data_od_21_));
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__22_), .Q(mc_data_od_22_));
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__23_), .Q(mc_data_od_23_));
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__24_), .Q(mc_data_od_24_));
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__25_), .Q(mc_data_od_25_));
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__26_), .Q(mc_data_od_26_));
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__27_), .Q(mc_data_od_27_));
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__28_), .Q(mc_data_od_28_));
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__29_), .Q(mc_data_od_29_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__1_), .Q(u0_tms0_1_));
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__30_), .Q(mc_data_od_30_));
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_i), .D(u3__0mc_data_o_31_0__31_), .Q(mc_data_od_31_));
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__0_), .Q(u3_u0_r3_0_));
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__1_), .Q(u3_u0_r3_1_));
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__2_), .Q(u3_u0_r3_2_));
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__3_), .Q(u3_u0_r3_3_));
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__4_), .Q(u3_u0_r3_4_));
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__5_), .Q(u3_u0_r3_5_));
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__6_), .Q(u3_u0_r3_6_));
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__7_), .Q(u3_u0_r3_7_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__2_), .Q(u0_tms0_2_));
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__8_), .Q(u3_u0_r3_8_));
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__9_), .Q(u3_u0_r3_9_));
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__10_), .Q(u3_u0_r3_10_));
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__11_), .Q(u3_u0_r3_11_));
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__12_), .Q(u3_u0_r3_12_));
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__13_), .Q(u3_u0_r3_13_));
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__14_), .Q(u3_u0_r3_14_));
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__15_), .Q(u3_u0_r3_15_));
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__16_), .Q(u3_u0_r3_16_));
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__17_), .Q(u3_u0_r3_17_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__3_), .Q(u0_tms0_3_));
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__18_), .Q(u3_u0_r3_18_));
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__19_), .Q(u3_u0_r3_19_));
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__20_), .Q(u3_u0_r3_20_));
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__21_), .Q(u3_u0_r3_21_));
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__22_), .Q(u3_u0_r3_22_));
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__23_), .Q(u3_u0_r3_23_));
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__24_), .Q(u3_u0_r3_24_));
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__25_), .Q(u3_u0_r3_25_));
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__26_), .Q(u3_u0_r3_26_));
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__27_), .Q(u3_u0_r3_27_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__4_), .Q(u0_tms0_4_));
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__28_), .Q(u3_u0_r3_28_));
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__29_), .Q(u3_u0_r3_29_));
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__30_), .Q(u3_u0_r3_30_));
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__31_), .Q(u3_u0_r3_31_));
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__32_), .Q(u3_u0_r3_32_));
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__33_), .Q(u3_u0_r3_33_));
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__34_), .Q(u3_u0_r3_34_));
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_i), .D(u3_u0__0r3_35_0__35_), .Q(u3_u0_r3_35_));
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__0_), .Q(u3_u0_r2_0_));
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__1_), .Q(u3_u0_r2_1_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__5_), .Q(u0_tms0_5_));
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__2_), .Q(u3_u0_r2_2_));
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__3_), .Q(u3_u0_r2_3_));
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__4_), .Q(u3_u0_r2_4_));
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__5_), .Q(u3_u0_r2_5_));
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__6_), .Q(u3_u0_r2_6_));
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__7_), .Q(u3_u0_r2_7_));
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__8_), .Q(u3_u0_r2_8_));
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__9_), .Q(u3_u0_r2_9_));
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__10_), .Q(u3_u0_r2_10_));
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__11_), .Q(u3_u0_r2_11_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__6_), .Q(u0_tms0_6_));
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__12_), .Q(u3_u0_r2_12_));
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__13_), .Q(u3_u0_r2_13_));
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__14_), .Q(u3_u0_r2_14_));
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__15_), .Q(u3_u0_r2_15_));
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__16_), .Q(u3_u0_r2_16_));
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__17_), .Q(u3_u0_r2_17_));
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__18_), .Q(u3_u0_r2_18_));
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__19_), .Q(u3_u0_r2_19_));
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__20_), .Q(u3_u0_r2_20_));
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__21_), .Q(u3_u0_r2_21_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__7_), .Q(u0_tms0_7_));
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__22_), .Q(u3_u0_r2_22_));
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__23_), .Q(u3_u0_r2_23_));
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__24_), .Q(u3_u0_r2_24_));
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__25_), .Q(u3_u0_r2_25_));
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__26_), .Q(u3_u0_r2_26_));
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__27_), .Q(u3_u0_r2_27_));
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__28_), .Q(u3_u0_r2_28_));
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__29_), .Q(u3_u0_r2_29_));
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__30_), .Q(u3_u0_r2_30_));
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__31_), .Q(u3_u0_r2_31_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_i), .D(u0__0poc_31_0__1_), .Q(\poc_o[1] ));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__8_), .Q(u0_tms0_8_));
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__32_), .Q(u3_u0_r2_32_));
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__33_), .Q(u3_u0_r2_33_));
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__34_), .Q(u3_u0_r2_34_));
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_i), .D(u3_u0__0r2_35_0__35_), .Q(u3_u0_r2_35_));
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__0_), .Q(u3_u0_r1_0_));
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__1_), .Q(u3_u0_r1_1_));
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__2_), .Q(u3_u0_r1_2_));
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__3_), .Q(u3_u0_r1_3_));
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__4_), .Q(u3_u0_r1_4_));
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__5_), .Q(u3_u0_r1_5_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__9_), .Q(u0_tms0_9_));
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__6_), .Q(u3_u0_r1_6_));
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__7_), .Q(u3_u0_r1_7_));
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__8_), .Q(u3_u0_r1_8_));
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__9_), .Q(u3_u0_r1_9_));
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__10_), .Q(u3_u0_r1_10_));
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__11_), .Q(u3_u0_r1_11_));
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__12_), .Q(u3_u0_r1_12_));
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__13_), .Q(u3_u0_r1_13_));
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__14_), .Q(u3_u0_r1_14_));
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__15_), .Q(u3_u0_r1_15_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__10_), .Q(u0_tms0_10_));
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__16_), .Q(u3_u0_r1_16_));
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__17_), .Q(u3_u0_r1_17_));
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__18_), .Q(u3_u0_r1_18_));
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__19_), .Q(u3_u0_r1_19_));
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__20_), .Q(u3_u0_r1_20_));
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__21_), .Q(u3_u0_r1_21_));
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__22_), .Q(u3_u0_r1_22_));
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__23_), .Q(u3_u0_r1_23_));
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__24_), .Q(u3_u0_r1_24_));
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__25_), .Q(u3_u0_r1_25_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__11_), .Q(u0_tms0_11_));
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__26_), .Q(u3_u0_r1_26_));
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__27_), .Q(u3_u0_r1_27_));
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__28_), .Q(u3_u0_r1_28_));
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__29_), .Q(u3_u0_r1_29_));
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__30_), .Q(u3_u0_r1_30_));
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__31_), .Q(u3_u0_r1_31_));
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__32_), .Q(u3_u0_r1_32_));
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__33_), .Q(u3_u0_r1_33_));
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__34_), .Q(u3_u0_r1_34_));
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_i), .D(u3_u0__0r1_35_0__35_), .Q(u3_u0_r1_35_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__12_), .Q(u0_tms0_12_));
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__0_), .Q(u3_u0_r0_0_));
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__1_), .Q(u3_u0_r0_1_));
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__2_), .Q(u3_u0_r0_2_));
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__3_), .Q(u3_u0_r0_3_));
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__4_), .Q(u3_u0_r0_4_));
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__5_), .Q(u3_u0_r0_5_));
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__6_), .Q(u3_u0_r0_6_));
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__7_), .Q(u3_u0_r0_7_));
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__8_), .Q(u3_u0_r0_8_));
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__9_), .Q(u3_u0_r0_9_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__13_), .Q(u0_tms0_13_));
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__10_), .Q(u3_u0_r0_10_));
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__11_), .Q(u3_u0_r0_11_));
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__12_), .Q(u3_u0_r0_12_));
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__13_), .Q(u3_u0_r0_13_));
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__14_), .Q(u3_u0_r0_14_));
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__15_), .Q(u3_u0_r0_15_));
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__16_), .Q(u3_u0_r0_16_));
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__17_), .Q(u3_u0_r0_17_));
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__18_), .Q(u3_u0_r0_18_));
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__19_), .Q(u3_u0_r0_19_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__14_), .Q(u0_tms0_14_));
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__20_), .Q(u3_u0_r0_20_));
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__21_), .Q(u3_u0_r0_21_));
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__22_), .Q(u3_u0_r0_22_));
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__23_), .Q(u3_u0_r0_23_));
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__24_), .Q(u3_u0_r0_24_));
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__25_), .Q(u3_u0_r0_25_));
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__26_), .Q(u3_u0_r0_26_));
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__27_), .Q(u3_u0_r0_27_));
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__28_), .Q(u3_u0_r0_28_));
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__29_), .Q(u3_u0_r0_29_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__15_), .Q(u0_tms0_15_));
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__30_), .Q(u3_u0_r0_30_));
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__31_), .Q(u3_u0_r0_31_));
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__32_), .Q(u3_u0_r0_32_));
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__33_), .Q(u3_u0_r0_33_));
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__34_), .Q(u3_u0_r0_34_));
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_i), .D(u3_u0__0r0_35_0__35_), .Q(u3_u0_r0_35_));
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_i), .D(u4__0rfr_clr_0_0_), .Q(u4_rfr_clr));
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_i), .D(u1_wb_write_go), .Q(u5_wb_write_go_r));
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_i), .D(cmd_a10), .Q(u5_cmd_a10_r));
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_i), .D(u5__0burst_act_rd_0_0_), .Q(u5_burst_act_rd));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__16_), .Q(u0_tms0_16_));
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__0_), .Q(u5_burst_cnt_0_));
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__1_), .Q(u5_burst_cnt_1_));
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__2_), .Q(u5_burst_cnt_2_));
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__3_), .Q(u5_burst_cnt_3_));
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__4_), .Q(u5_burst_cnt_4_));
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__5_), .Q(u5_burst_cnt_5_));
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__6_), .Q(u5_burst_cnt_6_));
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__7_), .Q(u5_burst_cnt_7_));
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__8_), .Q(u5_burst_cnt_8_));
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__9_), .Q(u5_burst_cnt_9_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__17_), .Q(u0_tms0_17_));
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_i), .D(u5__0burst_cnt_10_0__10_), .Q(u5_burst_cnt_10_));
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_i), .D(u5__0ir_cnt_done_0_0_), .Q(u5_ir_cnt_done));
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_i), .D(u5__0ir_cnt_3_0__0_), .Q(u5_ir_cnt_0_));
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_i), .D(u5__0ir_cnt_3_0__1_), .Q(u5_ir_cnt_1_));
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_i), .D(u5__0ir_cnt_3_0__2_), .Q(u5_ir_cnt_2_));
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_i), .D(u5__0ir_cnt_3_0__3_), .Q(u5_ir_cnt_3_));
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_i), .D(u5__0timer2_8_0__0_), .Q(u5_timer2_0_));
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_i), .D(u5__0timer2_8_0__1_), .Q(u5_timer2_1_));
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_i), .D(u5__0timer2_8_0__2_), .Q(u5_timer2_2_));
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_i), .D(u5__0timer2_8_0__3_), .Q(u5_timer2_3_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_i), .D(u0__0poc_31_0__2_), .Q(\poc_o[2] ));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__18_), .Q(u0_tms0_18_));
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_i), .D(u5__0timer2_8_0__4_), .Q(u5_timer2_4_));
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_i), .D(u5__0timer2_8_0__5_), .Q(u5_timer2_5_));
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_i), .D(u5__0timer2_8_0__6_), .Q(u5_timer2_6_));
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_i), .D(u5__0timer2_8_0__7_), .Q(u5_timer2_7_));
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_i), .D(u5__0timer2_8_0__8_), .Q(u5_timer2_8_));
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_i), .D(u5_cnt_next), .Q(u5_cnt));
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_i), .D(u5_wb_wait_r2), .Q(u5_wb_wait_r));
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_i), .D(u5_wb_wait), .Q(u5_wb_wait_r2));
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_i), .D(u5_cke_o_r2), .Q(u5_cke_o_del));
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_i), .D(u5_cke_o_r1), .Q(u5_cke_o_r2));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__19_), .Q(u0_tms0_19_));
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_i), .D(mc_cke_pad_o_), .Q(u5_cke_o_r1));
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_i), .D(u5__0cke__0_0_), .Q(mc_cke_pad_o_));
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_i), .D(u5_cke_d), .Q(u5_cke_r));
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_i), .D(u5_pack_le2_d), .Q(pack_le2));
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_i), .D(u5_pack_le1_d), .Q(pack_le1));
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_i), .D(u5_pack_le0_d), .Q(pack_le0));
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_i), .D(cs_le_d), .Q(cs_le));
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_i), .D(cs_le), .Q(u5_cs_le_r1));
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_i), .D(u5_cs_le_r1), .Q(u5_cs_le_r));
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_i), .D(u5_lmr_ack_d), .Q(lmr_ack));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__20_), .Q(u0_tms0_20_));
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__0_), .Q(\wb_data_o[0] ));
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__1_), .Q(\wb_data_o[1] ));
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__2_), .Q(\wb_data_o[2] ));
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__3_), .Q(\wb_data_o[3] ));
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__4_), .Q(\wb_data_o[4] ));
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__5_), .Q(\wb_data_o[5] ));
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__6_), .Q(\wb_data_o[6] ));
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__7_), .Q(\wb_data_o[7] ));
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__8_), .Q(\wb_data_o[8] ));
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__9_), .Q(\wb_data_o[9] ));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__21_), .Q(u0_tms0_21_));
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__10_), .Q(\wb_data_o[10] ));
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__11_), .Q(\wb_data_o[11] ));
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__12_), .Q(\wb_data_o[12] ));
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__13_), .Q(\wb_data_o[13] ));
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__14_), .Q(\wb_data_o[14] ));
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__15_), .Q(\wb_data_o[15] ));
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__16_), .Q(\wb_data_o[16] ));
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__17_), .Q(\wb_data_o[17] ));
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__18_), .Q(\wb_data_o[18] ));
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__19_), .Q(\wb_data_o[19] ));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__22_), .Q(u0_tms0_22_));
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__20_), .Q(\wb_data_o[20] ));
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__21_), .Q(\wb_data_o[21] ));
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__22_), .Q(\wb_data_o[22] ));
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__23_), .Q(\wb_data_o[23] ));
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__24_), .Q(\wb_data_o[24] ));
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__25_), .Q(\wb_data_o[25] ));
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__26_), .Q(\wb_data_o[26] ));
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__27_), .Q(\wb_data_o[27] ));
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__28_), .Q(\wb_data_o[28] ));
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__29_), .Q(\wb_data_o[29] ));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__23_), .Q(u0_tms0_23_));
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__30_), .Q(\wb_data_o[30] ));
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_i), .D(u6__0wb_data_o_31_0__31_), .Q(\wb_data_o[31] ));
DFFPOSX1 DFFPOSX1_652 ( .CLK(mc_clk_i), .D(u7__0mc_adv__0_0_), .Q(mc_adv_pad_o_));
DFFPOSX1 DFFPOSX1_653 ( .CLK(mc_clk_i), .D(u7__0mc_adsc__0_0_), .Q(mc_adsc_pad_o_));
DFFPOSX1 DFFPOSX1_654 ( .CLK(mc_clk_i), .D(ras_), .Q(mc_ras_pad_o_));
DFFPOSX1 DFFPOSX1_655 ( .CLK(mc_clk_i), .D(cas_), .Q(mc_cas_pad_o_));
DFFPOSX1 DFFPOSX1_656 ( .CLK(mc_clk_i), .D(u5_we_), .Q(mc_we_pad_o_));
DFFPOSX1 DFFPOSX1_657 ( .CLK(mc_clk_i), .D(u7__0mc_dqm_3_0__0_), .Q(\mc_dqm_pad_o[0] ));
DFFPOSX1 DFFPOSX1_658 ( .CLK(mc_clk_i), .D(u7__0mc_dqm_3_0__1_), .Q(\mc_dqm_pad_o[1] ));
DFFPOSX1 DFFPOSX1_659 ( .CLK(mc_clk_i), .D(u7__0mc_dqm_3_0__2_), .Q(\mc_dqm_pad_o[2] ));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__24_), .Q(u0_tms0_24_));
DFFPOSX1 DFFPOSX1_660 ( .CLK(mc_clk_i), .D(u7__0mc_dqm_3_0__3_), .Q(\mc_dqm_pad_o[3] ));
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_i), .D(u7_mc_dqm_r_0_), .Q(u7_mc_dqm_r2_0_));
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_i), .D(u7_mc_dqm_r_1_), .Q(u7_mc_dqm_r2_1_));
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_i), .D(u7_mc_dqm_r_2_), .Q(u7_mc_dqm_r2_2_));
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_i), .D(u7_mc_dqm_r_3_), .Q(u7_mc_dqm_r2_3_));
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_i), .D(u7__0mc_dqm_r_3_0__0_), .Q(u7_mc_dqm_r_0_));
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_i), .D(u7__0mc_dqm_r_3_0__1_), .Q(u7_mc_dqm_r_1_));
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_i), .D(u7__0mc_dqm_r_3_0__2_), .Q(u7_mc_dqm_r_2_));
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_i), .D(u7__0mc_dqm_r_3_0__3_), .Q(u7_mc_dqm_r_3_));
DFFPOSX1 DFFPOSX1_669 ( .CLK(mc_clk_i), .D(mc_addr_d_0_), .Q(\mc_addr_pad_o[0] ));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__25_), .Q(u0_tms0_25_));
DFFPOSX1 DFFPOSX1_670 ( .CLK(mc_clk_i), .D(mc_addr_d_1_), .Q(\mc_addr_pad_o[1] ));
DFFPOSX1 DFFPOSX1_671 ( .CLK(mc_clk_i), .D(mc_addr_d_2_), .Q(\mc_addr_pad_o[2] ));
DFFPOSX1 DFFPOSX1_672 ( .CLK(mc_clk_i), .D(mc_addr_d_3_), .Q(\mc_addr_pad_o[3] ));
DFFPOSX1 DFFPOSX1_673 ( .CLK(mc_clk_i), .D(mc_addr_d_4_), .Q(\mc_addr_pad_o[4] ));
DFFPOSX1 DFFPOSX1_674 ( .CLK(mc_clk_i), .D(mc_addr_d_5_), .Q(\mc_addr_pad_o[5] ));
DFFPOSX1 DFFPOSX1_675 ( .CLK(mc_clk_i), .D(mc_addr_d_6_), .Q(\mc_addr_pad_o[6] ));
DFFPOSX1 DFFPOSX1_676 ( .CLK(mc_clk_i), .D(mc_addr_d_7_), .Q(\mc_addr_pad_o[7] ));
DFFPOSX1 DFFPOSX1_677 ( .CLK(mc_clk_i), .D(mc_addr_d_8_), .Q(\mc_addr_pad_o[8] ));
DFFPOSX1 DFFPOSX1_678 ( .CLK(mc_clk_i), .D(mc_addr_d_9_), .Q(\mc_addr_pad_o[9] ));
DFFPOSX1 DFFPOSX1_679 ( .CLK(mc_clk_i), .D(mc_addr_d_10_), .Q(\mc_addr_pad_o[10] ));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__26_), .Q(u0_tms0_26_));
DFFPOSX1 DFFPOSX1_680 ( .CLK(mc_clk_i), .D(mc_addr_d_11_), .Q(\mc_addr_pad_o[11] ));
DFFPOSX1 DFFPOSX1_681 ( .CLK(mc_clk_i), .D(mc_addr_d_12_), .Q(\mc_addr_pad_o[12] ));
DFFPOSX1 DFFPOSX1_682 ( .CLK(mc_clk_i), .D(mc_addr_d_13_), .Q(\mc_addr_pad_o[13] ));
DFFPOSX1 DFFPOSX1_683 ( .CLK(mc_clk_i), .D(mc_addr_d_14_), .Q(\mc_addr_pad_o[14] ));
DFFPOSX1 DFFPOSX1_684 ( .CLK(mc_clk_i), .D(mc_addr_d_15_), .Q(\mc_addr_pad_o[15] ));
DFFPOSX1 DFFPOSX1_685 ( .CLK(mc_clk_i), .D(mc_addr_d_16_), .Q(\mc_addr_pad_o[16] ));
DFFPOSX1 DFFPOSX1_686 ( .CLK(mc_clk_i), .D(mc_addr_d_17_), .Q(\mc_addr_pad_o[17] ));
DFFPOSX1 DFFPOSX1_687 ( .CLK(mc_clk_i), .D(mc_addr_d_18_), .Q(\mc_addr_pad_o[18] ));
DFFPOSX1 DFFPOSX1_688 ( .CLK(mc_clk_i), .D(mc_addr_d_19_), .Q(\mc_addr_pad_o[19] ));
DFFPOSX1 DFFPOSX1_689 ( .CLK(mc_clk_i), .D(mc_addr_d_20_), .Q(\mc_addr_pad_o[20] ));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__27_), .Q(u0_tms0_27_));
DFFPOSX1 DFFPOSX1_690 ( .CLK(mc_clk_i), .D(mc_addr_d_21_), .Q(\mc_addr_pad_o[21] ));
DFFPOSX1 DFFPOSX1_691 ( .CLK(mc_clk_i), .D(mc_addr_d_22_), .Q(\mc_addr_pad_o[22] ));
DFFPOSX1 DFFPOSX1_692 ( .CLK(mc_clk_i), .D(mc_addr_d_23_), .Q(\mc_addr_pad_o[23] ));
DFFPOSX1 DFFPOSX1_693 ( .CLK(mc_clk_i), .D(mc_dp_od_0_), .Q(\mc_dp_pad_o[0] ));
DFFPOSX1 DFFPOSX1_694 ( .CLK(mc_clk_i), .D(mc_dp_od_1_), .Q(\mc_dp_pad_o[1] ));
DFFPOSX1 DFFPOSX1_695 ( .CLK(mc_clk_i), .D(mc_dp_od_2_), .Q(\mc_dp_pad_o[2] ));
DFFPOSX1 DFFPOSX1_696 ( .CLK(mc_clk_i), .D(mc_dp_od_3_), .Q(\mc_dp_pad_o[3] ));
DFFPOSX1 DFFPOSX1_697 ( .CLK(mc_clk_i), .D(mc_data_od_0_), .Q(\mc_data_pad_o[0] ));
DFFPOSX1 DFFPOSX1_698 ( .CLK(mc_clk_i), .D(mc_data_od_1_), .Q(\mc_data_pad_o[1] ));
DFFPOSX1 DFFPOSX1_699 ( .CLK(mc_clk_i), .D(mc_data_od_2_), .Q(\mc_data_pad_o[2] ));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_i), .D(u0__0poc_31_0__3_), .Q(\poc_o[3] ));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__28_), .Q(u0_tms0_28_));
DFFPOSX1 DFFPOSX1_700 ( .CLK(mc_clk_i), .D(mc_data_od_3_), .Q(\mc_data_pad_o[3] ));
DFFPOSX1 DFFPOSX1_701 ( .CLK(mc_clk_i), .D(mc_data_od_4_), .Q(\mc_data_pad_o[4] ));
DFFPOSX1 DFFPOSX1_702 ( .CLK(mc_clk_i), .D(mc_data_od_5_), .Q(\mc_data_pad_o[5] ));
DFFPOSX1 DFFPOSX1_703 ( .CLK(mc_clk_i), .D(mc_data_od_6_), .Q(\mc_data_pad_o[6] ));
DFFPOSX1 DFFPOSX1_704 ( .CLK(mc_clk_i), .D(mc_data_od_7_), .Q(\mc_data_pad_o[7] ));
DFFPOSX1 DFFPOSX1_705 ( .CLK(mc_clk_i), .D(mc_data_od_8_), .Q(\mc_data_pad_o[8] ));
DFFPOSX1 DFFPOSX1_706 ( .CLK(mc_clk_i), .D(mc_data_od_9_), .Q(\mc_data_pad_o[9] ));
DFFPOSX1 DFFPOSX1_707 ( .CLK(mc_clk_i), .D(mc_data_od_10_), .Q(\mc_data_pad_o[10] ));
DFFPOSX1 DFFPOSX1_708 ( .CLK(mc_clk_i), .D(mc_data_od_11_), .Q(\mc_data_pad_o[11] ));
DFFPOSX1 DFFPOSX1_709 ( .CLK(mc_clk_i), .D(mc_data_od_12_), .Q(\mc_data_pad_o[12] ));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__29_), .Q(u0_tms0_29_));
DFFPOSX1 DFFPOSX1_710 ( .CLK(mc_clk_i), .D(mc_data_od_13_), .Q(\mc_data_pad_o[13] ));
DFFPOSX1 DFFPOSX1_711 ( .CLK(mc_clk_i), .D(mc_data_od_14_), .Q(\mc_data_pad_o[14] ));
DFFPOSX1 DFFPOSX1_712 ( .CLK(mc_clk_i), .D(mc_data_od_15_), .Q(\mc_data_pad_o[15] ));
DFFPOSX1 DFFPOSX1_713 ( .CLK(mc_clk_i), .D(mc_data_od_16_), .Q(\mc_data_pad_o[16] ));
DFFPOSX1 DFFPOSX1_714 ( .CLK(mc_clk_i), .D(mc_data_od_17_), .Q(\mc_data_pad_o[17] ));
DFFPOSX1 DFFPOSX1_715 ( .CLK(mc_clk_i), .D(mc_data_od_18_), .Q(\mc_data_pad_o[18] ));
DFFPOSX1 DFFPOSX1_716 ( .CLK(mc_clk_i), .D(mc_data_od_19_), .Q(\mc_data_pad_o[19] ));
DFFPOSX1 DFFPOSX1_717 ( .CLK(mc_clk_i), .D(mc_data_od_20_), .Q(\mc_data_pad_o[20] ));
DFFPOSX1 DFFPOSX1_718 ( .CLK(mc_clk_i), .D(mc_data_od_21_), .Q(\mc_data_pad_o[21] ));
DFFPOSX1 DFFPOSX1_719 ( .CLK(mc_clk_i), .D(mc_data_od_22_), .Q(\mc_data_pad_o[22] ));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__30_), .Q(u0_tms0_30_));
DFFPOSX1 DFFPOSX1_720 ( .CLK(mc_clk_i), .D(mc_data_od_23_), .Q(\mc_data_pad_o[23] ));
DFFPOSX1 DFFPOSX1_721 ( .CLK(mc_clk_i), .D(mc_data_od_24_), .Q(\mc_data_pad_o[24] ));
DFFPOSX1 DFFPOSX1_722 ( .CLK(mc_clk_i), .D(mc_data_od_25_), .Q(\mc_data_pad_o[25] ));
DFFPOSX1 DFFPOSX1_723 ( .CLK(mc_clk_i), .D(mc_data_od_26_), .Q(\mc_data_pad_o[26] ));
DFFPOSX1 DFFPOSX1_724 ( .CLK(mc_clk_i), .D(mc_data_od_27_), .Q(\mc_data_pad_o[27] ));
DFFPOSX1 DFFPOSX1_725 ( .CLK(mc_clk_i), .D(mc_data_od_28_), .Q(\mc_data_pad_o[28] ));
DFFPOSX1 DFFPOSX1_726 ( .CLK(mc_clk_i), .D(mc_data_od_29_), .Q(\mc_data_pad_o[29] ));
DFFPOSX1 DFFPOSX1_727 ( .CLK(mc_clk_i), .D(mc_data_od_30_), .Q(\mc_data_pad_o[30] ));
DFFPOSX1 DFFPOSX1_728 ( .CLK(mc_clk_i), .D(mc_data_od_31_), .Q(\mc_data_pad_o[31] ));
DFFPOSX1 DFFPOSX1_729 ( .CLK(mc_clk_i), .D(mc_bg_d), .Q(mc_bg_pad_o));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_i), .D(u0_u0__0tms_31_0__31_), .Q(u0_tms0_31_));
DFFPOSX1 DFFPOSX1_730 ( .CLK(mc_clk_i), .D(mc_ack_pad_i), .Q(mc_ack_r));
DFFPOSX1 DFFPOSX1_731 ( .CLK(mc_clk_i), .D(mc_br_pad_i), .Q(mc_br_r));
DFFPOSX1 DFFPOSX1_732 ( .CLK(mc_clk_i), .D(u7__0mc_rp_0_0_), .Q(mc_rp_pad_o_));
DFFPOSX1 DFFPOSX1_733 ( .CLK(mc_clk_i), .D(mc_c_oe_d), .Q(mc_coe_pad_coe_o));
DFFPOSX1 DFFPOSX1_734 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[0] ), .Q(mc_data_ir_0_));
DFFPOSX1 DFFPOSX1_735 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[1] ), .Q(mc_data_ir_1_));
DFFPOSX1 DFFPOSX1_736 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[2] ), .Q(mc_data_ir_2_));
DFFPOSX1 DFFPOSX1_737 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[3] ), .Q(mc_data_ir_3_));
DFFPOSX1 DFFPOSX1_738 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[4] ), .Q(mc_data_ir_4_));
DFFPOSX1 DFFPOSX1_739 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[5] ), .Q(mc_data_ir_5_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__0_), .Q(u0_csc0_0_));
DFFPOSX1 DFFPOSX1_740 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[6] ), .Q(mc_data_ir_6_));
DFFPOSX1 DFFPOSX1_741 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[7] ), .Q(mc_data_ir_7_));
DFFPOSX1 DFFPOSX1_742 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[8] ), .Q(mc_data_ir_8_));
DFFPOSX1 DFFPOSX1_743 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[9] ), .Q(mc_data_ir_9_));
DFFPOSX1 DFFPOSX1_744 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[10] ), .Q(mc_data_ir_10_));
DFFPOSX1 DFFPOSX1_745 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[11] ), .Q(mc_data_ir_11_));
DFFPOSX1 DFFPOSX1_746 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[12] ), .Q(mc_data_ir_12_));
DFFPOSX1 DFFPOSX1_747 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[13] ), .Q(mc_data_ir_13_));
DFFPOSX1 DFFPOSX1_748 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[14] ), .Q(mc_data_ir_14_));
DFFPOSX1 DFFPOSX1_749 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[15] ), .Q(mc_data_ir_15_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__1_), .Q(u0_csc0_1_));
DFFPOSX1 DFFPOSX1_750 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[16] ), .Q(mc_data_ir_16_));
DFFPOSX1 DFFPOSX1_751 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[17] ), .Q(mc_data_ir_17_));
DFFPOSX1 DFFPOSX1_752 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[18] ), .Q(mc_data_ir_18_));
DFFPOSX1 DFFPOSX1_753 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[19] ), .Q(mc_data_ir_19_));
DFFPOSX1 DFFPOSX1_754 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[20] ), .Q(mc_data_ir_20_));
DFFPOSX1 DFFPOSX1_755 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[21] ), .Q(mc_data_ir_21_));
DFFPOSX1 DFFPOSX1_756 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[22] ), .Q(mc_data_ir_22_));
DFFPOSX1 DFFPOSX1_757 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[23] ), .Q(mc_data_ir_23_));
DFFPOSX1 DFFPOSX1_758 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[24] ), .Q(mc_data_ir_24_));
DFFPOSX1 DFFPOSX1_759 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[25] ), .Q(mc_data_ir_25_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__2_), .Q(u0_csc0_2_));
DFFPOSX1 DFFPOSX1_760 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[26] ), .Q(mc_data_ir_26_));
DFFPOSX1 DFFPOSX1_761 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[27] ), .Q(mc_data_ir_27_));
DFFPOSX1 DFFPOSX1_762 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[28] ), .Q(mc_data_ir_28_));
DFFPOSX1 DFFPOSX1_763 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[29] ), .Q(mc_data_ir_29_));
DFFPOSX1 DFFPOSX1_764 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[30] ), .Q(mc_data_ir_30_));
DFFPOSX1 DFFPOSX1_765 ( .CLK(mc_clk_i), .D(\mc_data_pad_i[31] ), .Q(mc_data_ir_31_));
DFFPOSX1 DFFPOSX1_766 ( .CLK(mc_clk_i), .D(\mc_dp_pad_i[0] ), .Q(mc_data_ir_32_));
DFFPOSX1 DFFPOSX1_767 ( .CLK(mc_clk_i), .D(\mc_dp_pad_i[1] ), .Q(mc_data_ir_33_));
DFFPOSX1 DFFPOSX1_768 ( .CLK(mc_clk_i), .D(\mc_dp_pad_i[2] ), .Q(mc_data_ir_34_));
DFFPOSX1 DFFPOSX1_769 ( .CLK(mc_clk_i), .D(\mc_dp_pad_i[3] ), .Q(mc_data_ir_35_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__3_), .Q(u0_csc0_3_));
DFFPOSX1 DFFPOSX1_770 ( .CLK(mc_clk_i), .D(mc_sts_pad_i), .Q(mc_sts_ir));
DFFPOSX1 DFFPOSX1_771 ( .CLK(mc_clk_i), .D(suspended_o), .Q(mc_zz_pad_o));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__4_), .Q(u0_csc0_4_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__5_), .Q(u0_csc0_5_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_i), .D(u0__0poc_31_0__4_), .Q(\poc_o[4] ));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__6_), .Q(u0_csc0_6_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__7_), .Q(u0_csc0_7_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__8_), .Q(u0_csc0_8_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__9_), .Q(u0_csc0_9_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__10_), .Q(u0_csc0_10_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__11_), .Q(u0_csc0_11_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__12_), .Q(u0_csc0_12_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__13_), .Q(u0_csc0_13_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__14_), .Q(u0_csc0_14_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__15_), .Q(u0_csc0_15_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_i), .D(u0__0poc_31_0__5_), .Q(\poc_o[5] ));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__16_), .Q(u0_csc0_16_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__17_), .Q(u0_csc0_17_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__18_), .Q(u0_csc0_18_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__19_), .Q(u0_csc0_19_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__20_), .Q(u0_csc0_20_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__21_), .Q(u0_csc0_21_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__22_), .Q(u0_csc0_22_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__23_), .Q(u0_csc0_23_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__24_), .Q(u0_csc0_24_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_i), .D(u0_u0__0csc_31_0__25_), .Q(u0_csc0_25_));
DFFSR DFFSR_1 ( .CLK(clk_i), .D(u0__0lmr_req_0_0_), .Q(lmr_req), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_10 ( .CLK(clk_i), .D(u0__0spec_req_cs_7_0__6_), .Q(spec_req_cs_6_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_100 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__2_), .Q(u0_csc_mask_2_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_101 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__3_), .Q(u0_csc_mask_3_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_102 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__4_), .Q(u0_csc_mask_4_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_103 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__5_), .Q(u0_csc_mask_5_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_104 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__6_), .Q(u0_csc_mask_6_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_105 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__7_), .Q(u0_csc_mask_7_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_106 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__8_), .Q(u0_csc_mask_8_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_107 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__9_), .Q(u0_csc_mask_9_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_108 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__10_), .Q(u0_csc_mask_10_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_109 ( .CLK(clk_i), .D(u0__0csr_r_10_1__0_), .Q(mc_vpen_pad_o), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_11 ( .CLK(clk_i), .D(u0__0spec_req_cs_7_0__7_), .Q(spec_req_cs_7_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_110 ( .CLK(clk_i), .D(u0__0csr_r_10_1__1_), .Q(fs), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_111 ( .CLK(clk_i), .D(u0__0csr_r_10_1__2_), .Q(u0_csr_3_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_112 ( .CLK(clk_i), .D(u0__0csr_r_10_1__3_), .Q(u0_csr_4_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_113 ( .CLK(clk_i), .D(u0__0csr_r_10_1__4_), .Q(u0_csr_5_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_114 ( .CLK(clk_i), .D(u0__0csr_r_10_1__5_), .Q(u0_csr_6_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_115 ( .CLK(clk_i), .D(u0__0csr_r_10_1__6_), .Q(u0_csr_7_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_116 ( .CLK(clk_i), .D(u0__0csr_r_10_1__7_), .Q(ref_int_0_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_117 ( .CLK(clk_i), .D(u0__0csr_r_10_1__8_), .Q(ref_int_1_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_118 ( .CLK(clk_i), .D(u0__0csr_r_10_1__9_), .Q(ref_int_2_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_119 ( .CLK(clk_i), .D(u0__0csr_r2_7_0__0_), .Q(rfr_ps_val_0_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_12 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__0_), .Q(sp_tms_0_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_120 ( .CLK(clk_i), .D(u0__0csr_r2_7_0__1_), .Q(rfr_ps_val_1_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_121 ( .CLK(clk_i), .D(u0__0csr_r2_7_0__2_), .Q(rfr_ps_val_2_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_122 ( .CLK(clk_i), .D(u0__0csr_r2_7_0__3_), .Q(rfr_ps_val_3_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_123 ( .CLK(clk_i), .D(u0__0csr_r2_7_0__4_), .Q(rfr_ps_val_4_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_124 ( .CLK(clk_i), .D(u0__0csr_r2_7_0__5_), .Q(rfr_ps_val_5_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_125 ( .CLK(clk_i), .D(u0__0csr_r2_7_0__6_), .Q(rfr_ps_val_6_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_126 ( .CLK(clk_i), .D(u0__0csr_r2_7_0__7_), .Q(rfr_ps_val_7_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_127 ( .CLK(clk_i), .D(u0__0rf_we_0_0_), .Q(u0_rf_we), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_128 ( .CLK(clk_i), .D(u0_u0__0inited_0_0_), .Q(u0_u0_inited), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_129 ( .CLK(clk_i), .D(u0_u0__0init_req_0_0_), .Q(u0_init_req0), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_13 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__1_), .Q(sp_tms_1_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_130 ( .CLK(clk_i), .D(u0_u0__0init_req_we_0_0_), .Q(u0_u0_init_req_we), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_131 ( .CLK(clk_i), .D(u0_u0__0lmr_req_0_0_), .Q(u0_lmr_req0), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_132 ( .CLK(clk_i), .D(u0_u0__0lmr_req_we_0_0_), .Q(u0_u0_lmr_req_we), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_133 ( .CLK(clk_i), .D(1'h0), .Q(u0_u0_rst_r2), .R(1'h1), .S(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494));
DFFSR DFFSR_134 ( .CLK(clk_i), .D(u0_u1__0inited_0_0_), .Q(u0_u1_inited), .R(u0_u1__abc_72470_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_135 ( .CLK(clk_i), .D(u0_u1__0init_req_0_0_), .Q(u0_init_req1), .R(u0_u1__abc_72470_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_136 ( .CLK(clk_i), .D(u0_u1__0init_req_we_0_0_), .Q(u0_u1_init_req_we), .R(u0_u1__abc_72470_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_137 ( .CLK(clk_i), .D(u0_u1__0lmr_req_0_0_), .Q(u0_lmr_req1), .R(u0_u1__abc_72470_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_138 ( .CLK(clk_i), .D(u0_u1__0lmr_req_we_0_0_), .Q(u0_u1_lmr_req_we), .R(u0_u1__abc_72470_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_139 ( .CLK(clk_i), .D(1'h0), .Q(u0_u1_rst_r2), .R(1'h1), .S(u0_u1__abc_72470_auto_rtlil_cc_1942_NotGate_71506));
DFFSR DFFSR_14 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__2_), .Q(sp_tms_2_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_140 ( .CLK(clk_i), .D(u2_u0__0bank3_open_0_0_), .Q(u2_u0_bank3_open), .R(u2_u0__abc_73914_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_141 ( .CLK(clk_i), .D(u2_u0__0bank2_open_0_0_), .Q(u2_u0_bank2_open), .R(u2_u0__abc_73914_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_142 ( .CLK(clk_i), .D(u2_u0__0bank1_open_0_0_), .Q(u2_u0_bank1_open), .R(u2_u0__abc_73914_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_143 ( .CLK(clk_i), .D(u2_u0__0bank0_open_0_0_), .Q(u2_u0_bank0_open), .R(u2_u0__abc_73914_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_144 ( .CLK(clk_i), .D(u2_u1__0bank3_open_0_0_), .Q(u2_u1_bank3_open), .R(u2_u1__abc_73914_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_145 ( .CLK(clk_i), .D(u2_u1__0bank2_open_0_0_), .Q(u2_u1_bank2_open), .R(u2_u1__abc_73914_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_146 ( .CLK(clk_i), .D(u2_u1__0bank1_open_0_0_), .Q(u2_u1_bank1_open), .R(u2_u1__abc_73914_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_147 ( .CLK(clk_i), .D(u2_u1__0bank0_open_0_0_), .Q(u2_u1_bank0_open), .R(u2_u1__abc_73914_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_148 ( .CLK(clk_i), .D(u3_u0__0wr_adr_3_0__0_), .Q(u3_u0_wr_adr_0_), .R(1'h1), .S(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546));
DFFSR DFFSR_149 ( .CLK(clk_i), .D(u3_u0__0wr_adr_3_0__1_), .Q(u3_u0_wr_adr_1_), .R(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_15 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__3_), .Q(sp_tms_3_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_150 ( .CLK(clk_i), .D(u3_u0__0wr_adr_3_0__2_), .Q(u3_u0_wr_adr_2_), .R(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_151 ( .CLK(clk_i), .D(u3_u0__0wr_adr_3_0__3_), .Q(u3_u0_wr_adr_3_), .R(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_152 ( .CLK(clk_i), .D(u3_u0__0rd_adr_3_0__0_), .Q(u3_u0_rd_adr_0_), .R(1'h1), .S(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546));
DFFSR DFFSR_153 ( .CLK(clk_i), .D(u3_u0__0rd_adr_3_0__1_), .Q(u3_u0_rd_adr_1_), .R(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_154 ( .CLK(clk_i), .D(u3_u0__0rd_adr_3_0__2_), .Q(u3_u0_rd_adr_2_), .R(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_155 ( .CLK(clk_i), .D(u3_u0__0rd_adr_3_0__3_), .Q(u3_u0_rd_adr_3_), .R(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_156 ( .CLK(clk_i), .D(u4__0rfr_req_0_0_), .Q(rfr_req), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_157 ( .CLK(clk_i), .D(u4__0rfr_cnt_7_0__0_), .Q(u4_rfr_cnt_0_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_158 ( .CLK(clk_i), .D(u4__0rfr_cnt_7_0__1_), .Q(u4_rfr_cnt_1_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_159 ( .CLK(clk_i), .D(u4__0rfr_cnt_7_0__2_), .Q(u4_rfr_cnt_2_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_16 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__4_), .Q(sp_tms_4_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_160 ( .CLK(clk_i), .D(u4__0rfr_cnt_7_0__3_), .Q(u4_rfr_cnt_3_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_161 ( .CLK(clk_i), .D(u4__0rfr_cnt_7_0__4_), .Q(u4_rfr_cnt_4_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_162 ( .CLK(clk_i), .D(u4__0rfr_cnt_7_0__5_), .Q(u4_rfr_cnt_5_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_163 ( .CLK(clk_i), .D(u4__0rfr_cnt_7_0__6_), .Q(u4_rfr_cnt_6_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_164 ( .CLK(clk_i), .D(u4__0rfr_cnt_7_0__7_), .Q(u4_rfr_cnt_7_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_165 ( .CLK(clk_i), .D(u4_ps_cnt_clr), .Q(u4_rfr_ce), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_166 ( .CLK(clk_i), .D(u4__0rfr_early_0_0_), .Q(u4_rfr_early), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_167 ( .CLK(clk_i), .D(u4__0ps_cnt_7_0__0_), .Q(u4_ps_cnt_0_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_168 ( .CLK(clk_i), .D(u4__0ps_cnt_7_0__1_), .Q(u4_ps_cnt_1_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_169 ( .CLK(clk_i), .D(u4__0ps_cnt_7_0__2_), .Q(u4_ps_cnt_2_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_17 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__5_), .Q(sp_tms_5_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_170 ( .CLK(clk_i), .D(u4__0ps_cnt_7_0__3_), .Q(u4_ps_cnt_3_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_171 ( .CLK(clk_i), .D(u4__0ps_cnt_7_0__4_), .Q(u4_ps_cnt_4_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_172 ( .CLK(clk_i), .D(u4__0ps_cnt_7_0__5_), .Q(u4_ps_cnt_5_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_173 ( .CLK(clk_i), .D(u4__0ps_cnt_7_0__6_), .Q(u4_ps_cnt_6_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_174 ( .CLK(clk_i), .D(u4__0ps_cnt_7_0__7_), .Q(u4_ps_cnt_7_), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_175 ( .CLK(clk_i), .D(u4__0rfr_en_0_0_), .Q(u4_rfr_en), .R(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562), .S(1'h1));
DFFSR DFFSR_176 ( .CLK(clk_i), .D(u5_next_state_0_), .Q(u5_state_0_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_177 ( .CLK(clk_i), .D(u5_next_state_1_), .Q(u5_state_1_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_178 ( .CLK(clk_i), .D(u5_next_state_2_), .Q(u5_state_2_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_179 ( .CLK(clk_i), .D(u5_next_state_3_), .Q(u5_state_3_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_18 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__6_), .Q(sp_tms_6_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_180 ( .CLK(clk_i), .D(u5_next_state_4_), .Q(u5_state_4_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_181 ( .CLK(clk_i), .D(u5_next_state_5_), .Q(u5_state_5_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_182 ( .CLK(clk_i), .D(u5_next_state_6_), .Q(u5_state_6_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_183 ( .CLK(clk_i), .D(u5_next_state_7_), .Q(u5_state_7_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_184 ( .CLK(clk_i), .D(u5_next_state_8_), .Q(u5_state_8_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_185 ( .CLK(clk_i), .D(u5_next_state_9_), .Q(u5_state_9_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_186 ( .CLK(clk_i), .D(u5_next_state_10_), .Q(u5_state_10_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_187 ( .CLK(clk_i), .D(u5_next_state_11_), .Q(u5_state_11_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_188 ( .CLK(clk_i), .D(u5_next_state_12_), .Q(u5_state_12_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_189 ( .CLK(clk_i), .D(u5_next_state_13_), .Q(u5_state_13_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_19 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__7_), .Q(sp_tms_7_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_190 ( .CLK(clk_i), .D(u5_next_state_14_), .Q(u5_state_14_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_191 ( .CLK(clk_i), .D(u5_next_state_15_), .Q(u5_state_15_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_192 ( .CLK(clk_i), .D(u5_next_state_16_), .Q(u5_state_16_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_193 ( .CLK(clk_i), .D(u5_next_state_17_), .Q(u5_state_17_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_194 ( .CLK(clk_i), .D(u5_next_state_18_), .Q(u5_state_18_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_195 ( .CLK(clk_i), .D(u5_next_state_19_), .Q(u5_state_19_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_196 ( .CLK(clk_i), .D(u5_next_state_20_), .Q(u5_state_20_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_197 ( .CLK(clk_i), .D(u5_next_state_21_), .Q(u5_state_21_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_198 ( .CLK(clk_i), .D(u5_next_state_22_), .Q(u5_state_22_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_199 ( .CLK(clk_i), .D(u5_next_state_23_), .Q(u5_state_23_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_2 ( .CLK(clk_i), .D(u0__0init_req_0_0_), .Q(init_req), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_20 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__8_), .Q(sp_tms_8_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_200 ( .CLK(clk_i), .D(u5_next_state_24_), .Q(u5_state_24_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_201 ( .CLK(clk_i), .D(u5_next_state_25_), .Q(u5_state_25_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_202 ( .CLK(clk_i), .D(u5_next_state_26_), .Q(u5_state_26_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_203 ( .CLK(clk_i), .D(u5_next_state_27_), .Q(u5_state_27_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_204 ( .CLK(clk_i), .D(u5_next_state_28_), .Q(u5_state_28_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_205 ( .CLK(clk_i), .D(u5_next_state_29_), .Q(u5_state_29_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_206 ( .CLK(clk_i), .D(u5_next_state_30_), .Q(u5_state_30_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_207 ( .CLK(clk_i), .D(u5_next_state_31_), .Q(u5_state_31_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_208 ( .CLK(clk_i), .D(u5_next_state_32_), .Q(u5_state_32_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_209 ( .CLK(clk_i), .D(u5_next_state_33_), .Q(u5_state_33_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_21 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__9_), .Q(sp_tms_9_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_210 ( .CLK(clk_i), .D(u5_next_state_34_), .Q(u5_state_34_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_211 ( .CLK(clk_i), .D(u5_next_state_35_), .Q(u5_state_35_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_212 ( .CLK(clk_i), .D(u5_next_state_36_), .Q(u5_state_36_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_213 ( .CLK(clk_i), .D(u5_next_state_37_), .Q(u5_state_37_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_214 ( .CLK(clk_i), .D(u5_next_state_38_), .Q(u5_state_38_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_215 ( .CLK(clk_i), .D(u5_next_state_39_), .Q(u5_state_39_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_216 ( .CLK(clk_i), .D(u5_next_state_40_), .Q(u5_state_40_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_217 ( .CLK(clk_i), .D(u5_next_state_41_), .Q(u5_state_41_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_218 ( .CLK(clk_i), .D(u5_next_state_42_), .Q(u5_state_42_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_219 ( .CLK(clk_i), .D(u5_next_state_43_), .Q(u5_state_43_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_22 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__10_), .Q(sp_tms_10_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_220 ( .CLK(clk_i), .D(u5_next_state_44_), .Q(u5_state_44_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_221 ( .CLK(clk_i), .D(u5_next_state_45_), .Q(u5_state_45_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_222 ( .CLK(clk_i), .D(u5_next_state_46_), .Q(u5_state_46_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_223 ( .CLK(clk_i), .D(u5_next_state_47_), .Q(u5_state_47_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_224 ( .CLK(clk_i), .D(u5_next_state_48_), .Q(u5_state_48_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_225 ( .CLK(clk_i), .D(u5_next_state_49_), .Q(u5_state_49_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_226 ( .CLK(clk_i), .D(u5_next_state_50_), .Q(u5_state_50_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_227 ( .CLK(clk_i), .D(u5_next_state_51_), .Q(u5_state_51_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_228 ( .CLK(clk_i), .D(u5_next_state_52_), .Q(u5_state_52_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_229 ( .CLK(clk_i), .D(u5_next_state_53_), .Q(u5_state_53_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_23 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__11_), .Q(sp_tms_11_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_230 ( .CLK(clk_i), .D(u5_next_state_54_), .Q(u5_state_54_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_231 ( .CLK(clk_i), .D(u5_next_state_55_), .Q(u5_state_55_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_232 ( .CLK(clk_i), .D(u5_next_state_56_), .Q(u5_state_56_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_233 ( .CLK(clk_i), .D(u5_next_state_57_), .Q(u5_state_57_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_234 ( .CLK(clk_i), .D(u5_next_state_58_), .Q(u5_state_58_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_235 ( .CLK(clk_i), .D(u5_next_state_59_), .Q(u5_state_59_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_236 ( .CLK(clk_i), .D(u5_next_state_60_), .Q(u5_state_60_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_237 ( .CLK(clk_i), .D(u5_next_state_61_), .Q(u5_state_61_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_238 ( .CLK(clk_i), .D(u5_next_state_62_), .Q(u5_state_62_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_239 ( .CLK(clk_i), .D(u5_next_state_63_), .Q(u5_state_63_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_24 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__12_), .Q(sp_tms_12_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_240 ( .CLK(clk_i), .D(u5_next_state_64_), .Q(u5_state_64_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_241 ( .CLK(clk_i), .D(u5_next_state_65_), .Q(u5_state_65_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_242 ( .CLK(clk_i), .D(u5__0wb_stb_first_0_0_), .Q(u5_wb_stb_first), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_243 ( .CLK(clk_i), .D(dv), .Q(u5_dv_r), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_244 ( .CLK(clk_i), .D(u5__0ap_en_0_0_), .Q(u5_ap_en), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_245 ( .CLK(clk_i), .D(u5_timer_is_zero), .Q(u5_tmr_done), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_246 ( .CLK(clk_i), .D(u5__0timer_7_0__0_), .Q(u5_timer_0_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_247 ( .CLK(clk_i), .D(u5__0timer_7_0__1_), .Q(u5_timer_1_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_248 ( .CLK(clk_i), .D(u5__0timer_7_0__2_), .Q(u5_timer_2_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_249 ( .CLK(clk_i), .D(u5__0timer_7_0__3_), .Q(u5_timer_3_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_25 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__13_), .Q(sp_tms_13_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_250 ( .CLK(clk_i), .D(u5__0timer_7_0__4_), .Q(u5_timer_4_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_251 ( .CLK(clk_i), .D(u5__0timer_7_0__5_), .Q(u5_timer_5_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_252 ( .CLK(clk_i), .D(u5__0timer_7_0__6_), .Q(u5_timer_6_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_253 ( .CLK(clk_i), .D(u5__0timer_7_0__7_), .Q(u5_timer_7_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_254 ( .CLK(clk_i), .D(u5__0tmr2_done_0_0_), .Q(u5_tmr2_done), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_255 ( .CLK(clk_i), .D(u5__0susp_sel_r_0_0_), .Q(susp_sel), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_256 ( .CLK(clk_i), .D(u5_rfr_ack_d), .Q(rfr_ack), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_257 ( .CLK(clk_i), .D(u5_suspended_d), .Q(suspended_o), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_258 ( .CLK(clk_i), .D(resume_req_i), .Q(u5_resume_req_r), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_259 ( .CLK(clk_i), .D(susp_req_i), .Q(u5_susp_req_r), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_26 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__14_), .Q(sp_tms_14_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_260 ( .CLK(clk_i), .D(u5__0ack_cnt_3_0__0_), .Q(u5_ack_cnt_0_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_261 ( .CLK(clk_i), .D(u5__0ack_cnt_3_0__1_), .Q(u5_ack_cnt_1_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_262 ( .CLK(clk_i), .D(u5__0ack_cnt_3_0__2_), .Q(u5_ack_cnt_2_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_263 ( .CLK(clk_i), .D(u5__0ack_cnt_3_0__3_), .Q(u5_ack_cnt_3_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_264 ( .CLK(clk_i), .D(u5__0no_wb_cycle_0_0_), .Q(u5_no_wb_cycle), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_265 ( .CLK(clk_i), .D(u5__0wb_cycle_0_0_), .Q(u5_wb_cycle), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_266 ( .CLK(clk_i), .D(u5__0wr_cycle_0_0_), .Q(u1_wr_cycle), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_267 ( .CLK(clk_i), .D(u5__0lookup_ready2_0_0_), .Q(u5_lookup_ready2), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_268 ( .CLK(clk_i), .D(u5__0lookup_ready1_0_0_), .Q(u5_lookup_ready1), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_269 ( .CLK(clk_i), .D(u5__0data_oe_0_0_), .Q(data_oe), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_27 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__15_), .Q(sp_tms_15_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_270 ( .CLK(clk_i), .D(u5_data_oe_r), .Q(u5_data_oe_r2), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_271 ( .CLK(clk_i), .D(u5_data_oe_d), .Q(u5_data_oe_r), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_272 ( .CLK(clk_i), .D(u5__0oe__0_0_), .Q(oe_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_273 ( .CLK(clk_i), .D(u5__0cmd_asserted2_0_0_), .Q(u5_cmd_asserted2), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_274 ( .CLK(clk_i), .D(u5__0cmd_asserted_0_0_), .Q(u5_cmd_asserted), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_275 ( .CLK(clk_i), .D(u5_cmd_r_0_), .Q(u5_cmd_del_0_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_276 ( .CLK(clk_i), .D(u5_cmd_r_1_), .Q(u5_cmd_del_1_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_277 ( .CLK(clk_i), .D(u5_cmd_r_2_), .Q(u5_cmd_del_2_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_278 ( .CLK(clk_i), .D(u5_cmd_r_3_), .Q(u5_cmd_del_3_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_279 ( .CLK(clk_i), .D(u5_cmd_0_), .Q(u5_cmd_r_0_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_28 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__16_), .Q(sp_tms_16_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_280 ( .CLK(clk_i), .D(u5_cmd_1_), .Q(u5_cmd_r_1_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_281 ( .CLK(clk_i), .D(u5_cmd_2_), .Q(u5_cmd_r_2_), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_282 ( .CLK(clk_i), .D(u5_cmd_3_), .Q(u5_cmd_r_3_), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_283 ( .CLK(clk_i), .D(mem_ack), .Q(u5_mem_ack_r), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_284 ( .CLK(clk_i), .D(u5__0mc_adv_r_0_0_), .Q(u5_mc_adv_r), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_285 ( .CLK(clk_i), .D(u5__0mc_adv_r1_0_0_), .Q(u5_mc_adv_r1), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_286 ( .CLK(clk_i), .D(u5__0mc_le_0_0_), .Q(u5_mc_le), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_72182), .S(1'h1));
DFFSR DFFSR_287 ( .CLK(clk_i), .D(u5_mc_c_oe_d), .Q(mc_c_oe_d), .R(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962), .S(1'h1));
DFFSR DFFSR_288 ( .CLK(clk_i), .D(1'h0), .Q(u5_rsts), .R(1'h1), .S(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
DFFSR DFFSR_289 ( .CLK(clk_i), .D(u6__0wb_err_0_0_), .Q(wb_err_o), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_29 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__17_), .Q(sp_tms_17_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_290 ( .CLK(clk_i), .D(u6__0wb_ack_o_0_0_), .Q(wb_ack_o), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_291 ( .CLK(clk_i), .D(u6__0wr_hold_0_0_), .Q(u1_wr_hold), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_292 ( .CLK(clk_i), .D(u6__0wb_first_r_0_0_), .Q(u6_wb_first_r), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_293 ( .CLK(clk_i), .D(u6__0write_go_r_0_0_), .Q(u6_write_go_r), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_294 ( .CLK(clk_i), .D(u6__0write_go_r1_0_0_), .Q(u6_write_go_r1), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_295 ( .CLK(clk_i), .D(u6__0read_go_r_0_0_), .Q(u6_read_go_r), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_296 ( .CLK(clk_i), .D(u6__0read_go_r1_0_0_), .Q(u6_read_go_r1), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_297 ( .CLK(clk_i), .D(u6__0rmw_r_0_0_), .Q(u6_rmw_r), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_298 ( .CLK(clk_i), .D(u6__0rmw_en_0_0_), .Q(u6_rmw_en), .R(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_299 ( .CLK(mc_clk_i), .D(u7__0mc_cs__7_7_), .Q(\mc_cs_pad_o_[7] ), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_3 ( .CLK(clk_i), .D(u0__0sreq_cs_le_0_0_), .Q(u0_sreq_cs_le), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_30 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__18_), .Q(sp_tms_18_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_300 ( .CLK(mc_clk_i), .D(u7__0mc_cs__6_6_), .Q(\mc_cs_pad_o_[6] ), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_301 ( .CLK(mc_clk_i), .D(u7__0mc_cs__5_5_), .Q(\mc_cs_pad_o_[5] ), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_302 ( .CLK(mc_clk_i), .D(u7__0mc_cs__4_4_), .Q(\mc_cs_pad_o_[4] ), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_303 ( .CLK(mc_clk_i), .D(u7__0mc_cs__3_3_), .Q(\mc_cs_pad_o_[3] ), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_304 ( .CLK(mc_clk_i), .D(u7__0mc_cs__2_2_), .Q(\mc_cs_pad_o_[2] ), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_305 ( .CLK(mc_clk_i), .D(u7__0mc_cs__1_1_), .Q(\mc_cs_pad_o_[1] ), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_306 ( .CLK(mc_clk_i), .D(u7__0mc_cs__0_0_), .Q(\mc_cs_pad_o_[0] ), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_307 ( .CLK(mc_clk_i), .D(u7__0mc_oe__0_0_), .Q(mc_oe_pad_o_), .R(1'h1), .S(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_308 ( .CLK(mc_clk_i), .D(u7__0mc_data_oe_0_0_), .Q(mc_doe_pad_doe_o), .R(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518), .S(1'h1));
DFFSR DFFSR_31 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__19_), .Q(sp_tms_19_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_32 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__20_), .Q(sp_tms_20_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_33 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__21_), .Q(sp_tms_21_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_34 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__22_), .Q(sp_tms_22_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_35 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__23_), .Q(sp_tms_23_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_36 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__24_), .Q(sp_tms_24_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_37 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__25_), .Q(sp_tms_25_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_38 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__26_), .Q(sp_tms_26_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_39 ( .CLK(clk_i), .D(u0__0sp_tms_31_0__27_), .Q(sp_tms_27_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_4 ( .CLK(clk_i), .D(u0__0spec_req_cs_7_0__0_), .Q(spec_req_cs_0_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_40 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__1_), .Q(sp_csc_1_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_41 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__2_), .Q(sp_csc_2_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_42 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__3_), .Q(sp_csc_3_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_43 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__4_), .Q(sp_csc_4_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_44 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__5_), .Q(sp_csc_5_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_45 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__6_), .Q(sp_csc_6_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_46 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__7_), .Q(sp_csc_7_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_47 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__9_), .Q(sp_csc_9_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_48 ( .CLK(clk_i), .D(u0__0sp_csc_31_0__10_), .Q(sp_csc_10_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_49 ( .CLK(clk_i), .D(u0__0tms_31_0__0_), .Q(tms_0_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_5 ( .CLK(clk_i), .D(u0__0spec_req_cs_7_0__1_), .Q(spec_req_cs_1_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_50 ( .CLK(clk_i), .D(u0__0tms_31_0__1_), .Q(tms_1_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_51 ( .CLK(clk_i), .D(u0__0tms_31_0__2_), .Q(tms_2_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_52 ( .CLK(clk_i), .D(u0__0tms_31_0__3_), .Q(tms_3_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_53 ( .CLK(clk_i), .D(u0__0tms_31_0__4_), .Q(tms_4_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_54 ( .CLK(clk_i), .D(u0__0tms_31_0__5_), .Q(tms_5_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_55 ( .CLK(clk_i), .D(u0__0tms_31_0__6_), .Q(tms_6_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_56 ( .CLK(clk_i), .D(u0__0tms_31_0__7_), .Q(tms_7_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_57 ( .CLK(clk_i), .D(u0__0tms_31_0__8_), .Q(tms_8_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_58 ( .CLK(clk_i), .D(u0__0tms_31_0__9_), .Q(tms_9_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_59 ( .CLK(clk_i), .D(u0__0tms_31_0__10_), .Q(tms_10_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_6 ( .CLK(clk_i), .D(u0__0spec_req_cs_7_0__2_), .Q(spec_req_cs_2_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_60 ( .CLK(clk_i), .D(u0__0tms_31_0__11_), .Q(tms_11_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_61 ( .CLK(clk_i), .D(u0__0tms_31_0__12_), .Q(tms_12_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_62 ( .CLK(clk_i), .D(u0__0tms_31_0__13_), .Q(tms_13_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_63 ( .CLK(clk_i), .D(u0__0tms_31_0__14_), .Q(tms_14_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_64 ( .CLK(clk_i), .D(u0__0tms_31_0__15_), .Q(tms_15_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_65 ( .CLK(clk_i), .D(u0__0tms_31_0__16_), .Q(tms_16_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_66 ( .CLK(clk_i), .D(u0__0tms_31_0__17_), .Q(tms_17_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_67 ( .CLK(clk_i), .D(u0__0tms_31_0__18_), .Q(tms_18_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_68 ( .CLK(clk_i), .D(u0__0tms_31_0__19_), .Q(tms_19_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_69 ( .CLK(clk_i), .D(u0__0tms_31_0__20_), .Q(tms_20_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_7 ( .CLK(clk_i), .D(u0__0spec_req_cs_7_0__3_), .Q(spec_req_cs_3_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_70 ( .CLK(clk_i), .D(u0__0tms_31_0__21_), .Q(tms_21_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_71 ( .CLK(clk_i), .D(u0__0tms_31_0__22_), .Q(tms_22_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_72 ( .CLK(clk_i), .D(u0__0tms_31_0__23_), .Q(tms_23_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_73 ( .CLK(clk_i), .D(u0__0tms_31_0__24_), .Q(tms_24_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_74 ( .CLK(clk_i), .D(u0__0tms_31_0__25_), .Q(tms_25_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_75 ( .CLK(clk_i), .D(u0__0tms_31_0__26_), .Q(tms_26_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_76 ( .CLK(clk_i), .D(u0__0tms_31_0__27_), .Q(tms_27_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_77 ( .CLK(clk_i), .D(u0__0csc_31_0__1_), .Q(csc_1_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_78 ( .CLK(clk_i), .D(u0__0csc_31_0__2_), .Q(csc_2_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_79 ( .CLK(clk_i), .D(u0__0csc_31_0__3_), .Q(csc_3_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_8 ( .CLK(clk_i), .D(u0__0spec_req_cs_7_0__4_), .Q(spec_req_cs_4_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_80 ( .CLK(clk_i), .D(u0__0csc_31_0__4_), .Q(csc_4_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_81 ( .CLK(clk_i), .D(u0__0csc_31_0__5_), .Q(csc_5_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_82 ( .CLK(clk_i), .D(u0__0csc_31_0__6_), .Q(csc_6_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_83 ( .CLK(clk_i), .D(u0__0csc_31_0__7_), .Q(csc_7_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_84 ( .CLK(clk_i), .D(u0__0csc_31_0__9_), .Q(csc_9_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_85 ( .CLK(clk_i), .D(u0__0csc_31_0__10_), .Q(csc_10_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_86 ( .CLK(clk_i), .D(u0__0csc_31_0__11_), .Q(u3_pen), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_87 ( .CLK(clk_i), .D(u0__0wp_err_0_0_), .Q(u0_wp_err), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_88 ( .CLK(clk_i), .D(u0__0cs_7_0__0_), .Q(cs_0_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_89 ( .CLK(clk_i), .D(u0__0cs_7_0__1_), .Q(cs_1_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_9 ( .CLK(clk_i), .D(u0__0spec_req_cs_7_0__5_), .Q(spec_req_cs_5_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_90 ( .CLK(clk_i), .D(u0__0cs_7_0__2_), .Q(cs_2_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_91 ( .CLK(clk_i), .D(u0__0cs_7_0__3_), .Q(cs_3_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_92 ( .CLK(clk_i), .D(u0__0cs_7_0__4_), .Q(cs_4_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_93 ( .CLK(clk_i), .D(u0__0cs_7_0__5_), .Q(cs_5_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_94 ( .CLK(clk_i), .D(u0__0cs_7_0__6_), .Q(cs_6_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_95 ( .CLK(clk_i), .D(u0__0cs_7_0__7_), .Q(cs_7_), .R(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602), .S(1'h1));
DFFSR DFFSR_96 ( .CLK(clk_i), .D(u0_rst_r2), .Q(u0_rst_r3), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_97 ( .CLK(clk_i), .D(1'h0), .Q(u0_rst_r2), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_98 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__0_), .Q(u0_csc_mask_0_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
DFFSR DFFSR_99 ( .CLK(clk_i), .D(u0__0csc_mask_r_10_0__1_), .Q(u0_csc_mask_1_), .R(1'h1), .S(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
INVX1 INVX1_1 ( .A(_abc_81086_new_n236_), .Y(lmr_sel));
INVX1 INVX1_10 ( .A(tms_8_), .Y(_abc_81086_new_n295_));
INVX1 INVX1_100 ( .A(u0_tms0_9_), .Y(u0__abc_74894_new_n1352_));
INVX1 INVX1_1000 ( .A(u5__abc_78290_new_n2588_), .Y(u5__abc_78290_new_n2589_));
INVX1 INVX1_1001 ( .A(u5__abc_78290_new_n1061_), .Y(u5__abc_78290_new_n2590_));
INVX1 INVX1_1002 ( .A(u5__abc_78290_new_n2591_), .Y(u5__abc_78290_new_n2592_));
INVX1 INVX1_1003 ( .A(u5_kro), .Y(u5__abc_78290_new_n2598_));
INVX1 INVX1_1004 ( .A(u5__abc_78290_new_n2599_), .Y(u5__abc_78290_new_n2600_));
INVX1 INVX1_1005 ( .A(u5__abc_78290_new_n1609_), .Y(u5__abc_78290_new_n2605_));
INVX1 INVX1_1006 ( .A(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2613_));
INVX1 INVX1_1007 ( .A(u5__abc_78290_new_n1363_), .Y(u5__abc_78290_new_n2620_));
INVX1 INVX1_1008 ( .A(u5__abc_78290_new_n2624_), .Y(u5__abc_78290_new_n2625_));
INVX1 INVX1_1009 ( .A(u5__abc_78290_new_n2627_), .Y(u5__abc_78290_new_n2628_));
INVX1 INVX1_101 ( .A(1'h0), .Y(u0__abc_74894_new_n1357_));
INVX1 INVX1_1010 ( .A(u5__abc_78290_new_n2639_), .Y(u5__abc_78290_new_n2640_));
INVX1 INVX1_1011 ( .A(u5__abc_78290_new_n1514_), .Y(u5__abc_78290_new_n2653_));
INVX1 INVX1_1012 ( .A(u5__abc_78290_new_n2584_), .Y(u5__abc_78290_new_n2659_));
INVX1 INVX1_1013 ( .A(u5__abc_78290_new_n2582_), .Y(u5__abc_78290_new_n2663_));
INVX1 INVX1_1014 ( .A(u5__abc_78290_new_n1023_), .Y(u5__abc_78290_new_n2670_));
INVX1 INVX1_1015 ( .A(rfr_ack), .Y(u5__abc_78290_new_n2672_));
INVX1 INVX1_1016 ( .A(u5__abc_78290_new_n2666_), .Y(u5__abc_78290_new_n2687_));
INVX1 INVX1_1017 ( .A(u5__abc_78290_new_n2740_), .Y(u5__abc_78290_new_n2741_));
INVX1 INVX1_1018 ( .A(u5__abc_78290_new_n2732_), .Y(u5__abc_78290_new_n2745_));
INVX1 INVX1_1019 ( .A(u5__abc_78290_new_n1533_), .Y(u5__abc_78290_new_n2773_));
INVX1 INVX1_102 ( .A(1'h0), .Y(u0__abc_74894_new_n1359_));
INVX1 INVX1_1020 ( .A(u5__abc_78290_new_n2673_), .Y(u5__abc_78290_new_n2778_));
INVX1 INVX1_1021 ( .A(u5__abc_78290_new_n2577_), .Y(u5__abc_78290_new_n2783_));
INVX1 INVX1_1022 ( .A(u5__abc_78290_new_n2593_), .Y(u5__abc_78290_new_n2788_));
INVX1 INVX1_1023 ( .A(u5__abc_78290_new_n2795_), .Y(u5__abc_78290_new_n2796_));
INVX1 INVX1_1024 ( .A(u5__abc_78290_new_n1436_), .Y(u5__abc_78290_new_n2835_));
INVX1 INVX1_1025 ( .A(u5__abc_78290_new_n2863_), .Y(u5__abc_78290_new_n2864_));
INVX1 INVX1_1026 ( .A(u5__abc_78290_new_n1386_), .Y(u5__abc_78290_new_n2877_));
INVX1 INVX1_1027 ( .A(u5__abc_78290_new_n1174_), .Y(u5__abc_78290_new_n2886_));
INVX1 INVX1_1028 ( .A(u5__abc_78290_new_n1380_), .Y(u5__abc_78290_new_n2890_));
INVX1 INVX1_1029 ( .A(csc_s_4_), .Y(u5__abc_78290_new_n2896_));
INVX1 INVX1_103 ( .A(u0_tms1_10_), .Y(u0__abc_74894_new_n1370_));
INVX1 INVX1_1030 ( .A(u5__abc_78290_new_n1495_), .Y(u5__abc_78290_new_n2914_));
INVX1 INVX1_1031 ( .A(u5__abc_78290_new_n1093_), .Y(u5__abc_78290_new_n2926_));
INVX1 INVX1_1032 ( .A(u5__abc_78290_new_n2947_), .Y(u5__abc_78290_new_n2948_));
INVX1 INVX1_1033 ( .A(u5__abc_78290_new_n1104_), .Y(u5__abc_78290_new_n2949_));
INVX1 INVX1_1034 ( .A(u5__abc_78290_new_n2950_), .Y(u5__abc_78290_new_n2963_));
INVX1 INVX1_1035 ( .A(u5__abc_78290_new_n2196_), .Y(u5__abc_78290_new_n2973_));
INVX1 INVX1_1036 ( .A(mc_ack_r), .Y(u5__abc_78290_new_n2975_));
INVX1 INVX1_1037 ( .A(u5__abc_78290_new_n2981_), .Y(u5__abc_78290_new_n2987_));
INVX1 INVX1_1038 ( .A(u5__abc_78290_new_n2208_), .Y(u5__abc_78290_new_n2994_));
INVX1 INVX1_1039 ( .A(u5__abc_78290_new_n1384_), .Y(u5__abc_78290_new_n2995_));
INVX1 INVX1_104 ( .A(u0_tms0_10_), .Y(u0__abc_74894_new_n1372_));
INVX1 INVX1_1040 ( .A(u5__abc_78290_new_n487_), .Y(u5__abc_78290_new_n3005_));
INVX1 INVX1_1041 ( .A(u5__abc_78290_new_n2330_), .Y(u5__abc_78290_new_n3008_));
INVX1 INVX1_1042 ( .A(u5__abc_78290_new_n1209_), .Y(u5__abc_78290_new_n3016_));
INVX1 INVX1_1043 ( .A(u5__abc_78290_new_n1058_), .Y(u5__abc_78290_new_n3038_));
INVX1 INVX1_1044 ( .A(u5__abc_78290_new_n2678_), .Y(u5__abc_78290_new_n3050_));
INVX1 INVX1_1045 ( .A(u5__abc_78290_new_n1438_), .Y(u5__abc_78290_new_n3060_));
INVX1 INVX1_1046 ( .A(u5__abc_78290_new_n1642_), .Y(u5__abc_78290_new_n3072_));
INVX1 INVX1_1047 ( .A(u5__abc_78290_new_n1555_), .Y(u5__abc_78290_new_n3075_));
INVX1 INVX1_1048 ( .A(u5__abc_78290_new_n3096_), .Y(u5__abc_78290_new_n3097_));
INVX1 INVX1_1049 ( .A(u5__abc_78290_new_n3141_), .Y(u5__0lookup_ready1_0_0_));
INVX1 INVX1_105 ( .A(1'h0), .Y(u0__abc_74894_new_n1377_));
INVX1 INVX1_1050 ( .A(u5__abc_78290_new_n3143_), .Y(u5__0lookup_ready2_0_0_));
INVX1 INVX1_1051 ( .A(u5_rsts), .Y(u5__abc_78290_auto_rtlil_cc_1942_NotGate_72182));
INVX1 INVX1_1052 ( .A(rst_i), .Y(u5__abc_78290_auto_rtlil_cc_1942_NotGate_71962));
INVX1 INVX1_1053 ( .A(\wb_addr_i[29] ), .Y(u6__abc_81318_new_n133_));
INVX1 INVX1_1054 ( .A(wb_cyc_i), .Y(u6__abc_81318_new_n136_));
INVX1 INVX1_1055 ( .A(wb_stb_i), .Y(u6__abc_81318_new_n137_));
INVX1 INVX1_1056 ( .A(wb_ack_o), .Y(u6__abc_81318_new_n143_));
INVX1 INVX1_1057 ( .A(mem_dout_0_), .Y(u6__abc_81318_new_n146_));
INVX1 INVX1_1058 ( .A(mem_dout_1_), .Y(u6__abc_81318_new_n149_));
INVX1 INVX1_1059 ( .A(mem_dout_2_), .Y(u6__abc_81318_new_n152_));
INVX1 INVX1_106 ( .A(1'h0), .Y(u0__abc_74894_new_n1379_));
INVX1 INVX1_1060 ( .A(mem_dout_3_), .Y(u6__abc_81318_new_n155_));
INVX1 INVX1_1061 ( .A(mem_dout_4_), .Y(u6__abc_81318_new_n158_));
INVX1 INVX1_1062 ( .A(mem_dout_5_), .Y(u6__abc_81318_new_n161_));
INVX1 INVX1_1063 ( .A(mem_dout_6_), .Y(u6__abc_81318_new_n164_));
INVX1 INVX1_1064 ( .A(mem_dout_7_), .Y(u6__abc_81318_new_n167_));
INVX1 INVX1_1065 ( .A(mem_dout_8_), .Y(u6__abc_81318_new_n170_));
INVX1 INVX1_1066 ( .A(mem_dout_9_), .Y(u6__abc_81318_new_n173_));
INVX1 INVX1_1067 ( .A(mem_dout_10_), .Y(u6__abc_81318_new_n176_));
INVX1 INVX1_1068 ( .A(mem_dout_11_), .Y(u6__abc_81318_new_n179_));
INVX1 INVX1_1069 ( .A(mem_dout_12_), .Y(u6__abc_81318_new_n182_));
INVX1 INVX1_107 ( .A(u0_tms1_11_), .Y(u0__abc_74894_new_n1390_));
INVX1 INVX1_1070 ( .A(mem_dout_13_), .Y(u6__abc_81318_new_n185_));
INVX1 INVX1_1071 ( .A(mem_dout_14_), .Y(u6__abc_81318_new_n188_));
INVX1 INVX1_1072 ( .A(mem_dout_15_), .Y(u6__abc_81318_new_n191_));
INVX1 INVX1_1073 ( .A(mem_dout_16_), .Y(u6__abc_81318_new_n194_));
INVX1 INVX1_1074 ( .A(mem_dout_17_), .Y(u6__abc_81318_new_n197_));
INVX1 INVX1_1075 ( .A(mem_dout_18_), .Y(u6__abc_81318_new_n200_));
INVX1 INVX1_1076 ( .A(mem_dout_19_), .Y(u6__abc_81318_new_n203_));
INVX1 INVX1_1077 ( .A(mem_dout_20_), .Y(u6__abc_81318_new_n206_));
INVX1 INVX1_1078 ( .A(mem_dout_21_), .Y(u6__abc_81318_new_n209_));
INVX1 INVX1_1079 ( .A(mem_dout_22_), .Y(u6__abc_81318_new_n212_));
INVX1 INVX1_108 ( .A(u0_tms0_11_), .Y(u0__abc_74894_new_n1392_));
INVX1 INVX1_1080 ( .A(mem_dout_23_), .Y(u6__abc_81318_new_n215_));
INVX1 INVX1_1081 ( .A(mem_dout_24_), .Y(u6__abc_81318_new_n218_));
INVX1 INVX1_1082 ( .A(mem_dout_25_), .Y(u6__abc_81318_new_n221_));
INVX1 INVX1_1083 ( .A(mem_dout_26_), .Y(u6__abc_81318_new_n224_));
INVX1 INVX1_1084 ( .A(mem_dout_27_), .Y(u6__abc_81318_new_n227_));
INVX1 INVX1_1085 ( .A(mem_dout_28_), .Y(u6__abc_81318_new_n230_));
INVX1 INVX1_1086 ( .A(mem_dout_29_), .Y(u6__abc_81318_new_n233_));
INVX1 INVX1_1087 ( .A(mem_dout_30_), .Y(u6__abc_81318_new_n236_));
INVX1 INVX1_1088 ( .A(mem_dout_31_), .Y(u6__abc_81318_new_n239_));
INVX1 INVX1_1089 ( .A(u1_wr_hold), .Y(u6__abc_81318_new_n242_));
INVX1 INVX1_109 ( .A(1'h0), .Y(u0__abc_74894_new_n1397_));
INVX1 INVX1_1090 ( .A(u6_read_go_r), .Y(u6__abc_81318_new_n247_));
INVX1 INVX1_1091 ( .A(wb_we_i), .Y(u6__abc_81318_new_n248_));
INVX1 INVX1_1092 ( .A(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n249_));
INVX1 INVX1_1093 ( .A(u6_rmw_r), .Y(u6__abc_81318_new_n251_));
INVX1 INVX1_1094 ( .A(u6__abc_81318_new_n243_), .Y(u6__abc_81318_new_n252_));
INVX1 INVX1_1095 ( .A(u6_rmw_en), .Y(u6__abc_81318_new_n253_));
INVX1 INVX1_1096 ( .A(u6__abc_81318_new_n258_), .Y(u6__0read_go_r_0_0_));
INVX1 INVX1_1097 ( .A(u6__abc_81318_new_n260_), .Y(u3_wb_read_go));
INVX1 INVX1_1098 ( .A(u6_write_go_r), .Y(u6__abc_81318_new_n262_));
INVX1 INVX1_1099 ( .A(u6__abc_81318_new_n267_), .Y(u1_wb_write_go));
INVX1 INVX1_11 ( .A(tms_9_), .Y(_abc_81086_new_n298_));
INVX1 INVX1_110 ( .A(1'h0), .Y(u0__abc_74894_new_n1399_));
INVX1 INVX1_1100 ( .A(wb_err_o), .Y(u6__abc_81318_new_n270_));
INVX1 INVX1_1101 ( .A(rst_i), .Y(u6__abc_81318_auto_rtlil_cc_1942_NotGate_72188));
INVX1 INVX1_1102 ( .A(susp_sel), .Y(u7__abc_73829_new_n75_));
INVX1 INVX1_1103 ( .A(data_oe), .Y(u7__abc_73829_new_n76_));
INVX1 INVX1_1104 ( .A(u5_wb_cycle), .Y(u7__abc_73829_new_n78_));
INVX1 INVX1_1105 ( .A(\wb_sel_i[0] ), .Y(u7__abc_73829_new_n87_));
INVX1 INVX1_1106 ( .A(\wb_sel_i[1] ), .Y(u7__abc_73829_new_n91_));
INVX1 INVX1_1107 ( .A(\wb_sel_i[2] ), .Y(u7__abc_73829_new_n94_));
INVX1 INVX1_1108 ( .A(\wb_sel_i[3] ), .Y(u7__abc_73829_new_n97_));
INVX1 INVX1_1109 ( .A(lmr_sel), .Y(u7__abc_73829_new_n101_));
INVX1 INVX1_111 ( .A(u0_tms1_12_), .Y(u0__abc_74894_new_n1410_));
INVX1 INVX1_1110 ( .A(cs_need_rfr_0_), .Y(u7__abc_73829_new_n105_));
INVX1 INVX1_1111 ( .A(cs_en), .Y(u7__abc_73829_new_n106_));
INVX1 INVX1_1112 ( .A(cs_need_rfr_1_), .Y(u7__abc_73829_new_n113_));
INVX1 INVX1_1113 ( .A(cs_need_rfr_2_), .Y(u7__abc_73829_new_n119_));
INVX1 INVX1_1114 ( .A(cs_need_rfr_3_), .Y(u7__abc_73829_new_n125_));
INVX1 INVX1_1115 ( .A(cs_need_rfr_4_), .Y(u7__abc_73829_new_n131_));
INVX1 INVX1_1116 ( .A(cs_need_rfr_5_), .Y(u7__abc_73829_new_n137_));
INVX1 INVX1_1117 ( .A(cs_need_rfr_6_), .Y(u7__abc_73829_new_n143_));
INVX1 INVX1_1118 ( .A(cs_need_rfr_7_), .Y(u7__abc_73829_new_n149_));
INVX1 INVX1_1119 ( .A(mc_adsc_d), .Y(u7__0mc_adsc__0_0_));
INVX1 INVX1_112 ( .A(u0_tms0_12_), .Y(u0__abc_74894_new_n1412_));
INVX1 INVX1_1120 ( .A(mc_adv_d), .Y(u7__0mc_adv__0_0_));
INVX1 INVX1_1121 ( .A(rst_i), .Y(u7__abc_73829_auto_rtlil_cc_1942_NotGate_71518));
INVX1 INVX1_113 ( .A(1'h0), .Y(u0__abc_74894_new_n1417_));
INVX1 INVX1_114 ( .A(1'h0), .Y(u0__abc_74894_new_n1419_));
INVX1 INVX1_115 ( .A(u0_tms1_13_), .Y(u0__abc_74894_new_n1430_));
INVX1 INVX1_116 ( .A(u0_tms0_13_), .Y(u0__abc_74894_new_n1432_));
INVX1 INVX1_117 ( .A(1'h0), .Y(u0__abc_74894_new_n1437_));
INVX1 INVX1_118 ( .A(1'h0), .Y(u0__abc_74894_new_n1439_));
INVX1 INVX1_119 ( .A(u0_tms1_14_), .Y(u0__abc_74894_new_n1450_));
INVX1 INVX1_12 ( .A(tms_10_), .Y(_abc_81086_new_n301_));
INVX1 INVX1_120 ( .A(u0_tms0_14_), .Y(u0__abc_74894_new_n1452_));
INVX1 INVX1_121 ( .A(1'h0), .Y(u0__abc_74894_new_n1457_));
INVX1 INVX1_122 ( .A(1'h0), .Y(u0__abc_74894_new_n1459_));
INVX1 INVX1_123 ( .A(u0_tms1_15_), .Y(u0__abc_74894_new_n1470_));
INVX1 INVX1_124 ( .A(u0_tms0_15_), .Y(u0__abc_74894_new_n1472_));
INVX1 INVX1_125 ( .A(1'h0), .Y(u0__abc_74894_new_n1477_));
INVX1 INVX1_126 ( .A(1'h0), .Y(u0__abc_74894_new_n1479_));
INVX1 INVX1_127 ( .A(u0_tms1_16_), .Y(u0__abc_74894_new_n1490_));
INVX1 INVX1_128 ( .A(u0_tms0_16_), .Y(u0__abc_74894_new_n1492_));
INVX1 INVX1_129 ( .A(1'h0), .Y(u0__abc_74894_new_n1497_));
INVX1 INVX1_13 ( .A(tms_11_), .Y(_abc_81086_new_n304_));
INVX1 INVX1_130 ( .A(1'h0), .Y(u0__abc_74894_new_n1499_));
INVX1 INVX1_131 ( .A(u0_tms1_17_), .Y(u0__abc_74894_new_n1510_));
INVX1 INVX1_132 ( .A(u0_tms0_17_), .Y(u0__abc_74894_new_n1512_));
INVX1 INVX1_133 ( .A(1'h0), .Y(u0__abc_74894_new_n1517_));
INVX1 INVX1_134 ( .A(1'h0), .Y(u0__abc_74894_new_n1519_));
INVX1 INVX1_135 ( .A(u0_tms1_18_), .Y(u0__abc_74894_new_n1530_));
INVX1 INVX1_136 ( .A(u0_tms0_18_), .Y(u0__abc_74894_new_n1532_));
INVX1 INVX1_137 ( .A(1'h0), .Y(u0__abc_74894_new_n1537_));
INVX1 INVX1_138 ( .A(1'h0), .Y(u0__abc_74894_new_n1539_));
INVX1 INVX1_139 ( .A(u0_tms1_19_), .Y(u0__abc_74894_new_n1550_));
INVX1 INVX1_14 ( .A(tms_12_), .Y(_abc_81086_new_n307_));
INVX1 INVX1_140 ( .A(u0_tms0_19_), .Y(u0__abc_74894_new_n1552_));
INVX1 INVX1_141 ( .A(1'h0), .Y(u0__abc_74894_new_n1557_));
INVX1 INVX1_142 ( .A(1'h0), .Y(u0__abc_74894_new_n1559_));
INVX1 INVX1_143 ( .A(u0_tms1_20_), .Y(u0__abc_74894_new_n1570_));
INVX1 INVX1_144 ( .A(u0_tms0_20_), .Y(u0__abc_74894_new_n1572_));
INVX1 INVX1_145 ( .A(1'h0), .Y(u0__abc_74894_new_n1577_));
INVX1 INVX1_146 ( .A(1'h0), .Y(u0__abc_74894_new_n1579_));
INVX1 INVX1_147 ( .A(u0_tms1_21_), .Y(u0__abc_74894_new_n1590_));
INVX1 INVX1_148 ( .A(u0_tms0_21_), .Y(u0__abc_74894_new_n1592_));
INVX1 INVX1_149 ( .A(1'h0), .Y(u0__abc_74894_new_n1597_));
INVX1 INVX1_15 ( .A(tms_13_), .Y(_abc_81086_new_n310_));
INVX1 INVX1_150 ( .A(1'h0), .Y(u0__abc_74894_new_n1599_));
INVX1 INVX1_151 ( .A(u0_tms1_22_), .Y(u0__abc_74894_new_n1610_));
INVX1 INVX1_152 ( .A(u0_tms0_22_), .Y(u0__abc_74894_new_n1612_));
INVX1 INVX1_153 ( .A(1'h0), .Y(u0__abc_74894_new_n1617_));
INVX1 INVX1_154 ( .A(1'h0), .Y(u0__abc_74894_new_n1619_));
INVX1 INVX1_155 ( .A(u0_tms1_23_), .Y(u0__abc_74894_new_n1630_));
INVX1 INVX1_156 ( .A(u0_tms0_23_), .Y(u0__abc_74894_new_n1632_));
INVX1 INVX1_157 ( .A(1'h0), .Y(u0__abc_74894_new_n1637_));
INVX1 INVX1_158 ( .A(1'h0), .Y(u0__abc_74894_new_n1639_));
INVX1 INVX1_159 ( .A(u0_tms1_24_), .Y(u0__abc_74894_new_n1650_));
INVX1 INVX1_16 ( .A(tms_14_), .Y(_abc_81086_new_n313_));
INVX1 INVX1_160 ( .A(u0_tms0_24_), .Y(u0__abc_74894_new_n1652_));
INVX1 INVX1_161 ( .A(1'h0), .Y(u0__abc_74894_new_n1657_));
INVX1 INVX1_162 ( .A(1'h0), .Y(u0__abc_74894_new_n1659_));
INVX1 INVX1_163 ( .A(u0_tms1_25_), .Y(u0__abc_74894_new_n1670_));
INVX1 INVX1_164 ( .A(u0_tms0_25_), .Y(u0__abc_74894_new_n1672_));
INVX1 INVX1_165 ( .A(1'h0), .Y(u0__abc_74894_new_n1677_));
INVX1 INVX1_166 ( .A(1'h0), .Y(u0__abc_74894_new_n1679_));
INVX1 INVX1_167 ( .A(u0_tms1_26_), .Y(u0__abc_74894_new_n1690_));
INVX1 INVX1_168 ( .A(u0_tms0_26_), .Y(u0__abc_74894_new_n1692_));
INVX1 INVX1_169 ( .A(1'h0), .Y(u0__abc_74894_new_n1697_));
INVX1 INVX1_17 ( .A(tms_15_), .Y(_abc_81086_new_n316_));
INVX1 INVX1_170 ( .A(1'h0), .Y(u0__abc_74894_new_n1699_));
INVX1 INVX1_171 ( .A(u0_tms1_27_), .Y(u0__abc_74894_new_n1710_));
INVX1 INVX1_172 ( .A(u0_tms0_27_), .Y(u0__abc_74894_new_n1712_));
INVX1 INVX1_173 ( .A(1'h0), .Y(u0__abc_74894_new_n1717_));
INVX1 INVX1_174 ( .A(1'h0), .Y(u0__abc_74894_new_n1737_));
INVX1 INVX1_175 ( .A(1'h0), .Y(u0__abc_74894_new_n1757_));
INVX1 INVX1_176 ( .A(u0_csc1_0_), .Y(u0__abc_74894_new_n1811_));
INVX1 INVX1_177 ( .A(1'h0), .Y(u0__abc_74894_new_n1818_));
INVX1 INVX1_178 ( .A(1'h0), .Y(u0__abc_74894_new_n1820_));
INVX1 INVX1_179 ( .A(u0_csc1_1_), .Y(u0__abc_74894_new_n1831_));
INVX1 INVX1_18 ( .A(tms_16_), .Y(_abc_81086_new_n319_));
INVX1 INVX1_180 ( .A(u0_csc0_1_), .Y(u0__abc_74894_new_n1833_));
INVX1 INVX1_181 ( .A(1'h0), .Y(u0__abc_74894_new_n1838_));
INVX1 INVX1_182 ( .A(1'h0), .Y(u0__abc_74894_new_n1840_));
INVX1 INVX1_183 ( .A(u0_csc1_2_), .Y(u0__abc_74894_new_n1851_));
INVX1 INVX1_184 ( .A(u0_csc0_2_), .Y(u0__abc_74894_new_n1853_));
INVX1 INVX1_185 ( .A(1'h0), .Y(u0__abc_74894_new_n1858_));
INVX1 INVX1_186 ( .A(1'h0), .Y(u0__abc_74894_new_n1860_));
INVX1 INVX1_187 ( .A(u0_csc1_3_), .Y(u0__abc_74894_new_n1871_));
INVX1 INVX1_188 ( .A(u0_csc0_3_), .Y(u0__abc_74894_new_n1873_));
INVX1 INVX1_189 ( .A(1'h0), .Y(u0__abc_74894_new_n1878_));
INVX1 INVX1_19 ( .A(tms_17_), .Y(_abc_81086_new_n322_));
INVX1 INVX1_190 ( .A(1'h0), .Y(u0__abc_74894_new_n1880_));
INVX1 INVX1_191 ( .A(u0_csc1_4_), .Y(u0__abc_74894_new_n1891_));
INVX1 INVX1_192 ( .A(u0_csc0_4_), .Y(u0__abc_74894_new_n1893_));
INVX1 INVX1_193 ( .A(1'h0), .Y(u0__abc_74894_new_n1898_));
INVX1 INVX1_194 ( .A(1'h0), .Y(u0__abc_74894_new_n1900_));
INVX1 INVX1_195 ( .A(u0_csc1_5_), .Y(u0__abc_74894_new_n1911_));
INVX1 INVX1_196 ( .A(u0_csc0_5_), .Y(u0__abc_74894_new_n1913_));
INVX1 INVX1_197 ( .A(1'h0), .Y(u0__abc_74894_new_n1918_));
INVX1 INVX1_198 ( .A(1'h0), .Y(u0__abc_74894_new_n1920_));
INVX1 INVX1_199 ( .A(u0_csc1_6_), .Y(u0__abc_74894_new_n1931_));
INVX1 INVX1_2 ( .A(tms_0_), .Y(_abc_81086_new_n271_));
INVX1 INVX1_20 ( .A(tms_18_), .Y(_abc_81086_new_n325_));
INVX1 INVX1_200 ( .A(u0_csc0_6_), .Y(u0__abc_74894_new_n1933_));
INVX1 INVX1_201 ( .A(1'h0), .Y(u0__abc_74894_new_n1938_));
INVX1 INVX1_202 ( .A(1'h0), .Y(u0__abc_74894_new_n1940_));
INVX1 INVX1_203 ( .A(u0_csc1_7_), .Y(u0__abc_74894_new_n1951_));
INVX1 INVX1_204 ( .A(u0_csc0_7_), .Y(u0__abc_74894_new_n1953_));
INVX1 INVX1_205 ( .A(1'h0), .Y(u0__abc_74894_new_n1958_));
INVX1 INVX1_206 ( .A(u0_csc0_8_), .Y(u0__abc_74894_new_n1973_));
INVX1 INVX1_207 ( .A(1'h0), .Y(u0__abc_74894_new_n1978_));
INVX1 INVX1_208 ( .A(1'h0), .Y(u0__abc_74894_new_n1980_));
INVX1 INVX1_209 ( .A(u0_csc1_9_), .Y(u0__abc_74894_new_n1991_));
INVX1 INVX1_21 ( .A(tms_19_), .Y(_abc_81086_new_n328_));
INVX1 INVX1_210 ( .A(u0_csc0_9_), .Y(u0__abc_74894_new_n1993_));
INVX1 INVX1_211 ( .A(1'h0), .Y(u0__abc_74894_new_n1998_));
INVX1 INVX1_212 ( .A(1'h0), .Y(u0__abc_74894_new_n2000_));
INVX1 INVX1_213 ( .A(u0_csc1_10_), .Y(u0__abc_74894_new_n2011_));
INVX1 INVX1_214 ( .A(u0_csc0_10_), .Y(u0__abc_74894_new_n2013_));
INVX1 INVX1_215 ( .A(1'h0), .Y(u0__abc_74894_new_n2018_));
INVX1 INVX1_216 ( .A(1'h0), .Y(u0__abc_74894_new_n2020_));
INVX1 INVX1_217 ( .A(u0_csc1_11_), .Y(u0__abc_74894_new_n2031_));
INVX1 INVX1_218 ( .A(1'h0), .Y(u0__abc_74894_new_n2058_));
INVX1 INVX1_219 ( .A(u0_csc0_13_), .Y(u0__abc_74894_new_n2073_));
INVX1 INVX1_22 ( .A(tms_20_), .Y(_abc_81086_new_n331_));
INVX1 INVX1_220 ( .A(1'h0), .Y(u0__abc_74894_new_n2078_));
INVX1 INVX1_221 ( .A(u0_csc1_15_), .Y(u0__abc_74894_new_n2111_));
INVX1 INVX1_222 ( .A(u0_csc0_16_), .Y(u0__abc_74894_new_n2133_));
INVX1 INVX1_223 ( .A(u0_csc1_17_), .Y(u0__abc_74894_new_n2151_));
INVX1 INVX1_224 ( .A(u0_csc1_18_), .Y(u0__abc_74894_new_n2171_));
INVX1 INVX1_225 ( .A(1'h0), .Y(u0__abc_74894_new_n2178_));
INVX1 INVX1_226 ( .A(u0_csc0_19_), .Y(u0__abc_74894_new_n2193_));
INVX1 INVX1_227 ( .A(1'h0), .Y(u0__abc_74894_new_n2218_));
INVX1 INVX1_228 ( .A(u0_csc0_23_), .Y(u0__abc_74894_new_n2273_));
INVX1 INVX1_229 ( .A(1'h0), .Y(u0__abc_74894_new_n2438_));
INVX1 INVX1_23 ( .A(tms_21_), .Y(_abc_81086_new_n334_));
INVX1 INVX1_230 ( .A(1'h0), .Y(u0__abc_74894_new_n2440_));
INVX1 INVX1_231 ( .A(1'h0), .Y(u0__abc_74894_new_n2441_));
INVX1 INVX1_232 ( .A(1'h0), .Y(u0__abc_74894_new_n2443_));
INVX1 INVX1_233 ( .A(1'h0), .Y(u0__abc_74894_new_n2444_));
INVX1 INVX1_234 ( .A(u0_cs1), .Y(u0__abc_74894_new_n2454_));
INVX1 INVX1_235 ( .A(u0_cs0), .Y(u0__abc_74894_new_n2455_));
INVX1 INVX1_236 ( .A(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n2970_));
INVX1 INVX1_237 ( .A(u0__abc_74894_new_n3469_), .Y(u0__abc_74894_new_n3470_));
INVX1 INVX1_238 ( .A(cs_7_), .Y(u0__abc_74894_new_n3493_));
INVX1 INVX1_239 ( .A(\poc_o[0] ), .Y(u0__abc_74894_new_n3496_));
INVX1 INVX1_24 ( .A(tms_22_), .Y(_abc_81086_new_n337_));
INVX1 INVX1_240 ( .A(\poc_o[1] ), .Y(u0__abc_74894_new_n3499_));
INVX1 INVX1_241 ( .A(\poc_o[2] ), .Y(u0__abc_74894_new_n3502_));
INVX1 INVX1_242 ( .A(\poc_o[3] ), .Y(u0__abc_74894_new_n3505_));
INVX1 INVX1_243 ( .A(\poc_o[4] ), .Y(u0__abc_74894_new_n3508_));
INVX1 INVX1_244 ( .A(\poc_o[5] ), .Y(u0__abc_74894_new_n3511_));
INVX1 INVX1_245 ( .A(\poc_o[6] ), .Y(u0__abc_74894_new_n3514_));
INVX1 INVX1_246 ( .A(\poc_o[7] ), .Y(u0__abc_74894_new_n3517_));
INVX1 INVX1_247 ( .A(\poc_o[8] ), .Y(u0__abc_74894_new_n3520_));
INVX1 INVX1_248 ( .A(\poc_o[9] ), .Y(u0__abc_74894_new_n3523_));
INVX1 INVX1_249 ( .A(\poc_o[10] ), .Y(u0__abc_74894_new_n3526_));
INVX1 INVX1_25 ( .A(tms_23_), .Y(_abc_81086_new_n340_));
INVX1 INVX1_250 ( .A(\poc_o[11] ), .Y(u0__abc_74894_new_n3529_));
INVX1 INVX1_251 ( .A(\poc_o[12] ), .Y(u0__abc_74894_new_n3532_));
INVX1 INVX1_252 ( .A(\poc_o[13] ), .Y(u0__abc_74894_new_n3535_));
INVX1 INVX1_253 ( .A(\poc_o[14] ), .Y(u0__abc_74894_new_n3538_));
INVX1 INVX1_254 ( .A(\poc_o[15] ), .Y(u0__abc_74894_new_n3541_));
INVX1 INVX1_255 ( .A(\poc_o[16] ), .Y(u0__abc_74894_new_n3544_));
INVX1 INVX1_256 ( .A(\poc_o[17] ), .Y(u0__abc_74894_new_n3547_));
INVX1 INVX1_257 ( .A(\poc_o[18] ), .Y(u0__abc_74894_new_n3550_));
INVX1 INVX1_258 ( .A(\poc_o[19] ), .Y(u0__abc_74894_new_n3553_));
INVX1 INVX1_259 ( .A(\poc_o[20] ), .Y(u0__abc_74894_new_n3556_));
INVX1 INVX1_26 ( .A(tms_24_), .Y(_abc_81086_new_n343_));
INVX1 INVX1_260 ( .A(\poc_o[21] ), .Y(u0__abc_74894_new_n3559_));
INVX1 INVX1_261 ( .A(\poc_o[22] ), .Y(u0__abc_74894_new_n3562_));
INVX1 INVX1_262 ( .A(\poc_o[23] ), .Y(u0__abc_74894_new_n3565_));
INVX1 INVX1_263 ( .A(\poc_o[24] ), .Y(u0__abc_74894_new_n3568_));
INVX1 INVX1_264 ( .A(\poc_o[25] ), .Y(u0__abc_74894_new_n3571_));
INVX1 INVX1_265 ( .A(\poc_o[26] ), .Y(u0__abc_74894_new_n3574_));
INVX1 INVX1_266 ( .A(\poc_o[27] ), .Y(u0__abc_74894_new_n3577_));
INVX1 INVX1_267 ( .A(\poc_o[28] ), .Y(u0__abc_74894_new_n3580_));
INVX1 INVX1_268 ( .A(\poc_o[29] ), .Y(u0__abc_74894_new_n3583_));
INVX1 INVX1_269 ( .A(\poc_o[30] ), .Y(u0__abc_74894_new_n3586_));
INVX1 INVX1_27 ( .A(tms_25_), .Y(_abc_81086_new_n346_));
INVX1 INVX1_270 ( .A(\poc_o[31] ), .Y(u0__abc_74894_new_n3589_));
INVX1 INVX1_271 ( .A(u0_csc_mask_0_), .Y(u0__abc_74894_new_n3592_));
INVX1 INVX1_272 ( .A(u0_wb_addr_r_6_), .Y(u0__abc_74894_new_n3593_));
INVX1 INVX1_273 ( .A(u0_wb_addr_r_2_), .Y(u0__abc_74894_new_n3596_));
INVX1 INVX1_274 ( .A(u0_csc_mask_1_), .Y(u0__abc_74894_new_n3601_));
INVX1 INVX1_275 ( .A(u0_csc_mask_2_), .Y(u0__abc_74894_new_n3604_));
INVX1 INVX1_276 ( .A(u0_csc_mask_3_), .Y(u0__abc_74894_new_n3607_));
INVX1 INVX1_277 ( .A(u0_csc_mask_4_), .Y(u0__abc_74894_new_n3610_));
INVX1 INVX1_278 ( .A(u0_csc_mask_5_), .Y(u0__abc_74894_new_n3613_));
INVX1 INVX1_279 ( .A(u0_csc_mask_6_), .Y(u0__abc_74894_new_n3616_));
INVX1 INVX1_28 ( .A(tms_26_), .Y(_abc_81086_new_n349_));
INVX1 INVX1_280 ( .A(u0_csc_mask_7_), .Y(u0__abc_74894_new_n3619_));
INVX1 INVX1_281 ( .A(u0_csc_mask_8_), .Y(u0__abc_74894_new_n3622_));
INVX1 INVX1_282 ( .A(u0_csc_mask_9_), .Y(u0__abc_74894_new_n3625_));
INVX1 INVX1_283 ( .A(u0_csc_mask_10_), .Y(u0__abc_74894_new_n3628_));
INVX1 INVX1_284 ( .A(mc_vpen_pad_o), .Y(u0__abc_74894_new_n3631_));
INVX1 INVX1_285 ( .A(u0_wb_addr_r_3_), .Y(u0__abc_74894_new_n3632_));
INVX1 INVX1_286 ( .A(fs), .Y(u0__abc_74894_new_n3637_));
INVX1 INVX1_287 ( .A(u0_csr_3_), .Y(u0__abc_74894_new_n3640_));
INVX1 INVX1_288 ( .A(u0_csr_4_), .Y(u0__abc_74894_new_n3643_));
INVX1 INVX1_289 ( .A(u0_csr_5_), .Y(u0__abc_74894_new_n3646_));
INVX1 INVX1_29 ( .A(tms_27_), .Y(_abc_81086_new_n352_));
INVX1 INVX1_290 ( .A(u0_csr_6_), .Y(u0__abc_74894_new_n3649_));
INVX1 INVX1_291 ( .A(u0_csr_7_), .Y(u0__abc_74894_new_n3652_));
INVX1 INVX1_292 ( .A(ref_int_0_), .Y(u0__abc_74894_new_n3655_));
INVX1 INVX1_293 ( .A(ref_int_1_), .Y(u0__abc_74894_new_n3658_));
INVX1 INVX1_294 ( .A(ref_int_2_), .Y(u0__abc_74894_new_n3661_));
INVX1 INVX1_295 ( .A(rfr_ps_val_0_), .Y(u0__abc_74894_new_n3664_));
INVX1 INVX1_296 ( .A(rfr_ps_val_1_), .Y(u0__abc_74894_new_n3667_));
INVX1 INVX1_297 ( .A(rfr_ps_val_2_), .Y(u0__abc_74894_new_n3670_));
INVX1 INVX1_298 ( .A(rfr_ps_val_3_), .Y(u0__abc_74894_new_n3673_));
INVX1 INVX1_299 ( .A(rfr_ps_val_4_), .Y(u0__abc_74894_new_n3676_));
INVX1 INVX1_3 ( .A(tms_1_), .Y(_abc_81086_new_n274_));
INVX1 INVX1_30 ( .A(csc_1_), .Y(_abc_81086_new_n370_));
INVX1 INVX1_300 ( .A(rfr_ps_val_5_), .Y(u0__abc_74894_new_n3679_));
INVX1 INVX1_301 ( .A(rfr_ps_val_6_), .Y(u0__abc_74894_new_n3682_));
INVX1 INVX1_302 ( .A(rfr_ps_val_7_), .Y(u0__abc_74894_new_n3685_));
INVX1 INVX1_303 ( .A(\wb_addr_i[3] ), .Y(u0__abc_74894_new_n3690_));
INVX1 INVX1_304 ( .A(\wb_addr_i[2] ), .Y(u0__abc_74894_new_n3691_));
INVX1 INVX1_305 ( .A(\wb_addr_i[5] ), .Y(u0__abc_74894_new_n3704_));
INVX1 INVX1_306 ( .A(u0__abc_74894_new_n3707_), .Y(u0__abc_74894_new_n3708_));
INVX1 INVX1_307 ( .A(u0__abc_74894_new_n3716_), .Y(u0__abc_74894_new_n3717_));
INVX1 INVX1_308 ( .A(u0__abc_74894_new_n3719_), .Y(u0__abc_74894_new_n3720_));
INVX1 INVX1_309 ( .A(\wb_addr_i[6] ), .Y(u0__abc_74894_new_n3724_));
INVX1 INVX1_31 ( .A(csc_2_), .Y(_abc_81086_new_n373_));
INVX1 INVX1_310 ( .A(u0__abc_74894_new_n3698_), .Y(u0__abc_74894_new_n3725_));
INVX1 INVX1_311 ( .A(u0__abc_74894_new_n3692_), .Y(u0__abc_74894_new_n3726_));
INVX1 INVX1_312 ( .A(u0__abc_74894_new_n3733_), .Y(u0__abc_74894_new_n3734_));
INVX1 INVX1_313 ( .A(u0__abc_74894_new_n3695_), .Y(u0__abc_74894_new_n3735_));
INVX1 INVX1_314 ( .A(u0__abc_74894_new_n3736_), .Y(u0__abc_74894_new_n3737_));
INVX1 INVX1_315 ( .A(u0__abc_74894_new_n3750_), .Y(u0__abc_74894_new_n3751_));
INVX1 INVX1_316 ( .A(1'h0), .Y(u0__abc_74894_new_n3764_));
INVX1 INVX1_317 ( .A(1'h0), .Y(u0__abc_74894_new_n3785_));
INVX1 INVX1_318 ( .A(1'h0), .Y(u0__abc_74894_new_n3797_));
INVX1 INVX1_319 ( .A(u0__abc_74894_new_n3693_), .Y(u0__abc_74894_new_n3798_));
INVX1 INVX1_32 ( .A(csc_3_), .Y(_abc_81086_new_n376_));
INVX1 INVX1_320 ( .A(u0__abc_74894_new_n3748_), .Y(u0__abc_74894_new_n3802_));
INVX1 INVX1_321 ( .A(1'h0), .Y(u0__abc_74894_new_n3840_));
INVX1 INVX1_322 ( .A(1'h0), .Y(u0__abc_74894_new_n3918_));
INVX1 INVX1_323 ( .A(1'h0), .Y(u0__abc_74894_new_n4001_));
INVX1 INVX1_324 ( .A(1'h0), .Y(u0__abc_74894_new_n4023_));
INVX1 INVX1_325 ( .A(1'h0), .Y(u0__abc_74894_new_n4052_));
INVX1 INVX1_326 ( .A(1'h0), .Y(u0__abc_74894_new_n4094_));
INVX1 INVX1_327 ( .A(1'h0), .Y(u0__abc_74894_new_n4116_));
INVX1 INVX1_328 ( .A(1'h0), .Y(u0__abc_74894_new_n4131_));
INVX1 INVX1_329 ( .A(1'h0), .Y(u0__abc_74894_new_n4173_));
INVX1 INVX1_33 ( .A(csc_4_), .Y(_abc_81086_new_n379_));
INVX1 INVX1_330 ( .A(1'h0), .Y(u0__abc_74894_new_n4272_));
INVX1 INVX1_331 ( .A(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4273_));
INVX1 INVX1_332 ( .A(1'h0), .Y(u0__abc_74894_new_n4328_));
INVX1 INVX1_333 ( .A(lmr_ack), .Y(u0__abc_74894_new_n4461_));
INVX1 INVX1_334 ( .A(init_ack), .Y(u0__abc_74894_new_n4463_));
INVX1 INVX1_335 ( .A(rst_i), .Y(u0__abc_74894_auto_rtlil_cc_1942_NotGate_71602));
INVX1 INVX1_336 ( .A(u0_u0_lmr_req_we), .Y(u0_u0__abc_72207_new_n205_));
INVX1 INVX1_337 ( .A(u0_csc0_3_), .Y(u0_u0__abc_72207_new_n206_));
INVX1 INVX1_338 ( .A(u0_lmr_ack0), .Y(u0_u0__abc_72207_new_n211_));
INVX1 INVX1_339 ( .A(u0_u0_addr_r_3_), .Y(u0_u0__abc_72207_new_n214_));
INVX1 INVX1_34 ( .A(csc_5_), .Y(_abc_81086_new_n382_));
INVX1 INVX1_340 ( .A(u0_u0_addr_r_6_), .Y(u0_u0__abc_72207_new_n216_));
INVX1 INVX1_341 ( .A(u0_u0_addr_r_5_), .Y(u0_u0__abc_72207_new_n217_));
INVX1 INVX1_342 ( .A(u0_u0__abc_72207_new_n220_), .Y(u0_u0__0lmr_req_we_0_0_));
INVX1 INVX1_343 ( .A(u0_u0_addr_r_2_), .Y(u0_u0__abc_72207_new_n318_));
INVX1 INVX1_344 ( .A(u0_rf_we), .Y(u0_u0__abc_72207_new_n320_));
INVX1 INVX1_345 ( .A(u0_u0__abc_72207_new_n322_), .Y(u0_u0__0init_req_we_0_0_));
INVX1 INVX1_346 ( .A(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n324_));
INVX1 INVX1_347 ( .A(u0_csc0_0_), .Y(u0_u0__abc_72207_new_n325_));
INVX1 INVX1_348 ( .A(\wb_data_i[0] ), .Y(u0_u0__abc_72207_new_n327_));
INVX1 INVX1_349 ( .A(u0_csc0_4_), .Y(u0_u0__abc_72207_new_n343_));
INVX1 INVX1_35 ( .A(csc_6_), .Y(_abc_81086_new_n385_));
INVX1 INVX1_350 ( .A(\wb_data_i[4] ), .Y(u0_u0__abc_72207_new_n345_));
INVX1 INVX1_351 ( .A(u0_csc0_5_), .Y(u0_u0__abc_72207_new_n350_));
INVX1 INVX1_352 ( .A(\wb_data_i[5] ), .Y(u0_u0__abc_72207_new_n352_));
INVX1 INVX1_353 ( .A(u0_csc0_6_), .Y(u0_u0__abc_72207_new_n356_));
INVX1 INVX1_354 ( .A(u0_csc0_7_), .Y(u0_u0__abc_72207_new_n359_));
INVX1 INVX1_355 ( .A(u0_csc0_8_), .Y(u0_u0__abc_72207_new_n362_));
INVX1 INVX1_356 ( .A(u0_csc0_9_), .Y(u0_u0__abc_72207_new_n365_));
INVX1 INVX1_357 ( .A(u0_csc0_10_), .Y(u0_u0__abc_72207_new_n368_));
INVX1 INVX1_358 ( .A(u0_csc0_11_), .Y(u0_u0__abc_72207_new_n371_));
INVX1 INVX1_359 ( .A(u0_csc0_12_), .Y(u0_u0__abc_72207_new_n374_));
INVX1 INVX1_36 ( .A(csc_7_), .Y(_abc_81086_new_n388_));
INVX1 INVX1_360 ( .A(u0_csc0_13_), .Y(u0_u0__abc_72207_new_n377_));
INVX1 INVX1_361 ( .A(u0_csc0_14_), .Y(u0_u0__abc_72207_new_n380_));
INVX1 INVX1_362 ( .A(u0_csc0_15_), .Y(u0_u0__abc_72207_new_n383_));
INVX1 INVX1_363 ( .A(u0_csc0_16_), .Y(u0_u0__abc_72207_new_n386_));
INVX1 INVX1_364 ( .A(u0_csc0_17_), .Y(u0_u0__abc_72207_new_n389_));
INVX1 INVX1_365 ( .A(u0_csc0_18_), .Y(u0_u0__abc_72207_new_n392_));
INVX1 INVX1_366 ( .A(u0_csc0_19_), .Y(u0_u0__abc_72207_new_n395_));
INVX1 INVX1_367 ( .A(u0_csc0_20_), .Y(u0_u0__abc_72207_new_n398_));
INVX1 INVX1_368 ( .A(u0_csc0_21_), .Y(u0_u0__abc_72207_new_n401_));
INVX1 INVX1_369 ( .A(u0_csc0_22_), .Y(u0_u0__abc_72207_new_n404_));
INVX1 INVX1_37 ( .A(csc_9_), .Y(_abc_81086_new_n394_));
INVX1 INVX1_370 ( .A(u0_csc0_23_), .Y(u0_u0__abc_72207_new_n407_));
INVX1 INVX1_371 ( .A(u0_csc0_24_), .Y(u0_u0__abc_72207_new_n410_));
INVX1 INVX1_372 ( .A(u0_csc0_25_), .Y(u0_u0__abc_72207_new_n413_));
INVX1 INVX1_373 ( .A(u0_csc0_26_), .Y(u0_u0__abc_72207_new_n416_));
INVX1 INVX1_374 ( .A(u0_csc0_27_), .Y(u0_u0__abc_72207_new_n419_));
INVX1 INVX1_375 ( .A(u0_csc0_28_), .Y(u0_u0__abc_72207_new_n422_));
INVX1 INVX1_376 ( .A(u0_csc0_29_), .Y(u0_u0__abc_72207_new_n425_));
INVX1 INVX1_377 ( .A(u0_csc0_30_), .Y(u0_u0__abc_72207_new_n428_));
INVX1 INVX1_378 ( .A(u0_csc0_31_), .Y(u0_u0__abc_72207_new_n431_));
INVX1 INVX1_379 ( .A(u0_u0__abc_72207_new_n439_), .Y(u0_u0__abc_72207_new_n440_));
INVX1 INVX1_38 ( .A(csc_10_), .Y(_abc_81086_new_n397_));
INVX1 INVX1_380 ( .A(u0_init_req0), .Y(u0_u0__abc_72207_new_n462_));
INVX1 INVX1_381 ( .A(rst_i), .Y(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494));
INVX1 INVX1_382 ( .A(u0_u1_lmr_req_we), .Y(u0_u1__abc_72470_new_n201_));
INVX1 INVX1_383 ( .A(u0_csc1_3_), .Y(u0_u1__abc_72470_new_n202_));
INVX1 INVX1_384 ( .A(u0_lmr_ack1), .Y(u0_u1__abc_72470_new_n207_));
INVX1 INVX1_385 ( .A(u0_u1_addr_r_2_), .Y(u0_u1__abc_72470_new_n210_));
INVX1 INVX1_386 ( .A(u0_u1_addr_r_5_), .Y(u0_u1__abc_72470_new_n211_));
INVX1 INVX1_387 ( .A(u0_u1_addr_r_6_), .Y(u0_u1__abc_72470_new_n213_));
INVX1 INVX1_388 ( .A(u0_u1__abc_72470_new_n416_), .Y(u0_u1__abc_72470_new_n417_));
INVX1 INVX1_389 ( .A(u0_init_req1), .Y(u0_u1__abc_72470_new_n438_));
INVX1 INVX1_39 ( .A(\wb_addr_i[31] ), .Y(_abc_81086_new_n463_));
INVX1 INVX1_390 ( .A(u0_u1_inited), .Y(u0_u1__abc_72470_new_n439_));
INVX1 INVX1_391 ( .A(rst_i), .Y(u0_u1__abc_72470_auto_rtlil_cc_1942_NotGate_71506));
INVX1 INVX1_392 ( .A(csc_s_5_), .Y(u1__abc_72801_new_n260_));
INVX1 INVX1_393 ( .A(csc_s_7_), .Y(u1__abc_72801_new_n262_));
INVX1 INVX1_394 ( .A(csc_s_6_), .Y(u1__abc_72801_new_n265_));
INVX1 INVX1_395 ( .A(csc_s_4_), .Y(u1__abc_72801_new_n269_));
INVX1 INVX1_396 ( .A(page_size_8_), .Y(u1__abc_72801_new_n273_));
INVX1 INVX1_397 ( .A(u1__abc_72801_new_n274_), .Y(page_size_10_));
INVX1 INVX1_398 ( .A(bank_adr_0_), .Y(u1__abc_72801_new_n276_));
INVX1 INVX1_399 ( .A(\wb_addr_i[12] ), .Y(u1__abc_72801_new_n277_));
INVX1 INVX1_4 ( .A(tms_2_), .Y(_abc_81086_new_n277_));
INVX1 INVX1_40 ( .A(spec_req_cs_0_), .Y(u0__abc_74894_new_n1100_));
INVX1 INVX1_400 ( .A(\wb_addr_i[25] ), .Y(u1__abc_72801_new_n287_));
INVX1 INVX1_401 ( .A(\wb_addr_i[21] ), .Y(u1__abc_72801_new_n300_));
INVX1 INVX1_402 ( .A(bank_adr_1_), .Y(u1__abc_72801_new_n307_));
INVX1 INVX1_403 ( .A(\wb_addr_i[13] ), .Y(u1__abc_72801_new_n308_));
INVX1 INVX1_404 ( .A(\wb_addr_i[26] ), .Y(u1__abc_72801_new_n312_));
INVX1 INVX1_405 ( .A(cs_le), .Y(u1__abc_72801_new_n322_));
INVX1 INVX1_406 ( .A(\wb_addr_i[14] ), .Y(u1__abc_72801_new_n324_));
INVX1 INVX1_407 ( .A(u1_bas), .Y(u1__abc_72801_new_n328_));
INVX1 INVX1_408 ( .A(\wb_addr_i[15] ), .Y(u1__abc_72801_new_n332_));
INVX1 INVX1_409 ( .A(row_adr_2_), .Y(u1__abc_72801_new_n346_));
INVX1 INVX1_41 ( .A(init_req), .Y(u0__abc_74894_new_n1101_));
INVX1 INVX1_410 ( .A(\wb_addr_i[19] ), .Y(u1__abc_72801_new_n399_));
INVX1 INVX1_411 ( .A(\wb_addr_i[20] ), .Y(u1__abc_72801_new_n408_));
INVX1 INVX1_412 ( .A(row_adr_9_), .Y(u1__abc_72801_new_n417_));
INVX1 INVX1_413 ( .A(\wb_addr_i[22] ), .Y(u1__abc_72801_new_n422_));
INVX1 INVX1_414 ( .A(\wb_addr_i[23] ), .Y(u1__abc_72801_new_n423_));
INVX1 INVX1_415 ( .A(\wb_addr_i[24] ), .Y(u1__abc_72801_new_n432_));
INVX1 INVX1_416 ( .A(row_adr_11_), .Y(u1__abc_72801_new_n441_));
INVX1 INVX1_417 ( .A(\wb_addr_i[2] ), .Y(u1__abc_72801_new_n460_));
INVX1 INVX1_418 ( .A(\wb_addr_i[3] ), .Y(u1__abc_72801_new_n464_));
INVX1 INVX1_419 ( .A(\wb_addr_i[4] ), .Y(u1__abc_72801_new_n467_));
INVX1 INVX1_42 ( .A(u0_lmr_req0), .Y(u0__abc_74894_new_n1102_));
INVX1 INVX1_420 ( .A(\wb_addr_i[5] ), .Y(u1__abc_72801_new_n470_));
INVX1 INVX1_421 ( .A(\wb_addr_i[6] ), .Y(u1__abc_72801_new_n473_));
INVX1 INVX1_422 ( .A(\wb_addr_i[7] ), .Y(u1__abc_72801_new_n476_));
INVX1 INVX1_423 ( .A(\wb_addr_i[8] ), .Y(u1__abc_72801_new_n479_));
INVX1 INVX1_424 ( .A(\wb_addr_i[9] ), .Y(u1__abc_72801_new_n482_));
INVX1 INVX1_425 ( .A(u1__abc_72801_new_n491_), .Y(u1__abc_72801_new_n498_));
INVX1 INVX1_426 ( .A(\wb_addr_i[10] ), .Y(u1__abc_72801_new_n537_));
INVX1 INVX1_427 ( .A(\wb_addr_i[11] ), .Y(u1__abc_72801_new_n543_));
INVX1 INVX1_428 ( .A(\wb_addr_i[16] ), .Y(u1__abc_72801_new_n580_));
INVX1 INVX1_429 ( .A(u1_sram_addr_14_), .Y(u1__abc_72801_new_n648_));
INVX1 INVX1_43 ( .A(spec_req_cs_1_), .Y(u0__abc_74894_new_n1106_));
INVX1 INVX1_430 ( .A(u1_sram_addr_15_), .Y(u1__abc_72801_new_n651_));
INVX1 INVX1_431 ( .A(u1_sram_addr_16_), .Y(u1__abc_72801_new_n654_));
INVX1 INVX1_432 ( .A(u1__abc_72801_new_n672_), .Y(u1__abc_72801_new_n673_));
INVX1 INVX1_433 ( .A(u1__abc_72801_new_n675_), .Y(u1__abc_72801_new_n676_));
INVX1 INVX1_434 ( .A(lmr_sel), .Y(u1__abc_72801_new_n682_));
INVX1 INVX1_435 ( .A(u1__abc_72801_new_n683_), .Y(u1__abc_72801_new_n684_));
INVX1 INVX1_436 ( .A(row_sel), .Y(u1__abc_72801_new_n767_));
INVX1 INVX1_437 ( .A(row_adr_12_), .Y(u1__abc_72801_new_n775_));
INVX1 INVX1_438 ( .A(u1_acs_addr_4_), .Y(u1_u0__abc_72719_new_n56_));
INVX1 INVX1_439 ( .A(u1_u0__abc_72719_new_n61_), .Y(u1_u0__abc_72719_new_n62_));
INVX1 INVX1_44 ( .A(u0_lmr_req1), .Y(u0__abc_74894_new_n1108_));
INVX1 INVX1_440 ( .A(u1_acs_addr_6_), .Y(u1_u0__abc_72719_new_n65_));
INVX1 INVX1_441 ( .A(u1_acs_addr_7_), .Y(u1_u0__abc_72719_new_n66_));
INVX1 INVX1_442 ( .A(u1_acs_addr_8_), .Y(u1_u0__abc_72719_new_n74_));
INVX1 INVX1_443 ( .A(u1_acs_addr_9_), .Y(u1_u0__abc_72719_new_n75_));
INVX1 INVX1_444 ( .A(u1_acs_addr_10_), .Y(u1_u0__abc_72719_new_n81_));
INVX1 INVX1_445 ( .A(u1_acs_addr_11_), .Y(u1_u0__abc_72719_new_n82_));
INVX1 INVX1_446 ( .A(u1_acs_addr_0_), .Y(u1_u0__0out_r_12_0__0_));
INVX1 INVX1_447 ( .A(u1_acs_addr_14_), .Y(u1_u0__abc_72719_new_n93_));
INVX1 INVX1_448 ( .A(u1_acs_addr_15_), .Y(u1_u0__abc_72719_new_n94_));
INVX1 INVX1_449 ( .A(u1_acs_addr_20_), .Y(u1_u0__abc_72719_new_n112_));
INVX1 INVX1_45 ( .A(spec_req_cs_2_), .Y(u0__abc_74894_new_n1112_));
INVX1 INVX1_450 ( .A(u1_u0__abc_72719_new_n119_), .Y(u1_u0__abc_72719_new_n120_));
INVX1 INVX1_451 ( .A(u1_acs_addr_22_), .Y(u1_u0__abc_72719_new_n123_));
INVX1 INVX1_452 ( .A(u1_acs_addr_23_), .Y(u1_u0__abc_72719_new_n125_));
INVX1 INVX1_453 ( .A(u1_u0__abc_72719_new_n85_), .Y(u1_u0__0out_r_12_0__12_));
INVX1 INVX1_454 ( .A(bank_set), .Y(u2__abc_74202_new_n64_));
INVX1 INVX1_455 ( .A(obct_cs_0_), .Y(u2__abc_74202_new_n65_));
INVX1 INVX1_456 ( .A(obct_cs_1_), .Y(u2__abc_74202_new_n67_));
INVX1 INVX1_457 ( .A(bank_clr), .Y(u2__abc_74202_new_n81_));
INVX1 INVX1_458 ( .A(bank_clr_all), .Y(u2__abc_74202_new_n90_));
INVX1 INVX1_459 ( .A(rfr_ack), .Y(u2__abc_74202_new_n91_));
INVX1 INVX1_46 ( .A(1'h0), .Y(u0__abc_74894_new_n1113_));
INVX1 INVX1_460 ( .A(row_adr_0_), .Y(u2_u0__abc_73914_new_n136_));
INVX1 INVX1_461 ( .A(u2_u0__abc_73914_new_n137_), .Y(u2_u0__abc_73914_new_n138_));
INVX1 INVX1_462 ( .A(u2_bank_set_0), .Y(u2_u0__abc_73914_new_n140_));
INVX1 INVX1_463 ( .A(row_adr_1_), .Y(u2_u0__abc_73914_new_n143_));
INVX1 INVX1_464 ( .A(row_adr_2_), .Y(u2_u0__abc_73914_new_n146_));
INVX1 INVX1_465 ( .A(row_adr_3_), .Y(u2_u0__abc_73914_new_n149_));
INVX1 INVX1_466 ( .A(row_adr_4_), .Y(u2_u0__abc_73914_new_n152_));
INVX1 INVX1_467 ( .A(row_adr_5_), .Y(u2_u0__abc_73914_new_n155_));
INVX1 INVX1_468 ( .A(row_adr_6_), .Y(u2_u0__abc_73914_new_n158_));
INVX1 INVX1_469 ( .A(row_adr_7_), .Y(u2_u0__abc_73914_new_n161_));
INVX1 INVX1_47 ( .A(u0__abc_74894_new_n1107_), .Y(u0__abc_74894_new_n1116_));
INVX1 INVX1_470 ( .A(row_adr_8_), .Y(u2_u0__abc_73914_new_n164_));
INVX1 INVX1_471 ( .A(row_adr_9_), .Y(u2_u0__abc_73914_new_n167_));
INVX1 INVX1_472 ( .A(row_adr_10_), .Y(u2_u0__abc_73914_new_n170_));
INVX1 INVX1_473 ( .A(row_adr_11_), .Y(u2_u0__abc_73914_new_n173_));
INVX1 INVX1_474 ( .A(row_adr_12_), .Y(u2_u0__abc_73914_new_n176_));
INVX1 INVX1_475 ( .A(u2_u0__abc_73914_new_n180_), .Y(u2_u0__abc_73914_new_n181_));
INVX1 INVX1_476 ( .A(bank_adr_1_), .Y(u2_u0__abc_73914_new_n208_));
INVX1 INVX1_477 ( .A(u2_u0__abc_73914_new_n237_), .Y(u2_u0__abc_73914_new_n239_));
INVX1 INVX1_478 ( .A(u2_u0_b3_last_row_8_), .Y(u2_u0__abc_73914_new_n266_));
INVX1 INVX1_479 ( .A(u2_u0_b3_last_row_9_), .Y(u2_u0__abc_73914_new_n267_));
INVX1 INVX1_48 ( .A(spec_req_cs_3_), .Y(u0__abc_74894_new_n1119_));
INVX1 INVX1_480 ( .A(u2_u0_b3_last_row_11_), .Y(u2_u0__abc_73914_new_n271_));
INVX1 INVX1_481 ( .A(u2_u0_b3_last_row_1_), .Y(u2_u0__abc_73914_new_n275_));
INVX1 INVX1_482 ( .A(u2_u0_b3_last_row_2_), .Y(u2_u0__abc_73914_new_n290_));
INVX1 INVX1_483 ( .A(u2_u0_b3_last_row_6_), .Y(u2_u0__abc_73914_new_n293_));
INVX1 INVX1_484 ( .A(u2_u0_b1_last_row_3_), .Y(u2_u0__abc_73914_new_n302_));
INVX1 INVX1_485 ( .A(u2_u0_b1_last_row_9_), .Y(u2_u0__abc_73914_new_n324_));
INVX1 INVX1_486 ( .A(u2_u0_b0_last_row_3_), .Y(u2_u0__abc_73914_new_n334_));
INVX1 INVX1_487 ( .A(u2_u0_b0_last_row_6_), .Y(u2_u0__abc_73914_new_n341_));
INVX1 INVX1_488 ( .A(u2_u0_b0_last_row_12_), .Y(u2_u0__abc_73914_new_n342_));
INVX1 INVX1_489 ( .A(u2_u0_b0_last_row_2_), .Y(u2_u0__abc_73914_new_n355_));
INVX1 INVX1_49 ( .A(1'h0), .Y(u0__abc_74894_new_n1120_));
INVX1 INVX1_490 ( .A(u2_u0_b0_last_row_4_), .Y(u2_u0__abc_73914_new_n356_));
INVX1 INVX1_491 ( .A(u2_u0_b2_last_row_11_), .Y(u2_u0__abc_73914_new_n367_));
INVX1 INVX1_492 ( .A(u2_u0_b2_last_row_4_), .Y(u2_u0__abc_73914_new_n369_));
INVX1 INVX1_493 ( .A(u2_u0_b2_last_row_6_), .Y(u2_u0__abc_73914_new_n374_));
INVX1 INVX1_494 ( .A(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_73914_new_n379_));
INVX1 INVX1_495 ( .A(u2_u0_bank0_open), .Y(u2_u0__abc_73914_new_n398_));
INVX1 INVX1_496 ( .A(u2_u0_bank1_open), .Y(u2_u0__abc_73914_new_n399_));
INVX1 INVX1_497 ( .A(u2_u0__abc_73914_new_n401_), .Y(u2_u0__abc_73914_new_n402_));
INVX1 INVX1_498 ( .A(u2_bank_clr_0), .Y(u2_u0__abc_73914_new_n404_));
INVX1 INVX1_499 ( .A(u2_u0_bank2_open), .Y(u2_u0__abc_73914_new_n405_));
INVX1 INVX1_5 ( .A(tms_3_), .Y(_abc_81086_new_n280_));
INVX1 INVX1_50 ( .A(spec_req_cs_4_), .Y(u0__abc_74894_new_n1125_));
INVX1 INVX1_500 ( .A(u2_u0_bank3_open), .Y(u2_u0__abc_73914_new_n409_));
INVX1 INVX1_501 ( .A(rst_i), .Y(u2_u0__abc_73914_auto_rtlil_cc_1942_NotGate_71538));
INVX1 INVX1_502 ( .A(row_adr_0_), .Y(u2_u1__abc_73914_new_n136_));
INVX1 INVX1_503 ( .A(u2_u1__abc_73914_new_n137_), .Y(u2_u1__abc_73914_new_n138_));
INVX1 INVX1_504 ( .A(u2_bank_set_1), .Y(u2_u1__abc_73914_new_n140_));
INVX1 INVX1_505 ( .A(row_adr_1_), .Y(u2_u1__abc_73914_new_n143_));
INVX1 INVX1_506 ( .A(row_adr_2_), .Y(u2_u1__abc_73914_new_n146_));
INVX1 INVX1_507 ( .A(row_adr_3_), .Y(u2_u1__abc_73914_new_n149_));
INVX1 INVX1_508 ( .A(row_adr_4_), .Y(u2_u1__abc_73914_new_n152_));
INVX1 INVX1_509 ( .A(row_adr_5_), .Y(u2_u1__abc_73914_new_n155_));
INVX1 INVX1_51 ( .A(1'h0), .Y(u0__abc_74894_new_n1126_));
INVX1 INVX1_510 ( .A(row_adr_6_), .Y(u2_u1__abc_73914_new_n158_));
INVX1 INVX1_511 ( .A(row_adr_7_), .Y(u2_u1__abc_73914_new_n161_));
INVX1 INVX1_512 ( .A(row_adr_8_), .Y(u2_u1__abc_73914_new_n164_));
INVX1 INVX1_513 ( .A(row_adr_9_), .Y(u2_u1__abc_73914_new_n167_));
INVX1 INVX1_514 ( .A(row_adr_10_), .Y(u2_u1__abc_73914_new_n170_));
INVX1 INVX1_515 ( .A(row_adr_11_), .Y(u2_u1__abc_73914_new_n173_));
INVX1 INVX1_516 ( .A(row_adr_12_), .Y(u2_u1__abc_73914_new_n176_));
INVX1 INVX1_517 ( .A(u2_u1__abc_73914_new_n180_), .Y(u2_u1__abc_73914_new_n181_));
INVX1 INVX1_518 ( .A(bank_adr_1_), .Y(u2_u1__abc_73914_new_n208_));
INVX1 INVX1_519 ( .A(u2_u1__abc_73914_new_n237_), .Y(u2_u1__abc_73914_new_n239_));
INVX1 INVX1_52 ( .A(u0__abc_74894_new_n1128_), .Y(u0__abc_74894_new_n1129_));
INVX1 INVX1_520 ( .A(u2_u1_b3_last_row_8_), .Y(u2_u1__abc_73914_new_n266_));
INVX1 INVX1_521 ( .A(u2_u1_b3_last_row_9_), .Y(u2_u1__abc_73914_new_n267_));
INVX1 INVX1_522 ( .A(u2_u1_b3_last_row_11_), .Y(u2_u1__abc_73914_new_n271_));
INVX1 INVX1_523 ( .A(u2_u1_b3_last_row_1_), .Y(u2_u1__abc_73914_new_n275_));
INVX1 INVX1_524 ( .A(u2_u1_b3_last_row_2_), .Y(u2_u1__abc_73914_new_n290_));
INVX1 INVX1_525 ( .A(u2_u1_b3_last_row_6_), .Y(u2_u1__abc_73914_new_n293_));
INVX1 INVX1_526 ( .A(u2_u1_b1_last_row_3_), .Y(u2_u1__abc_73914_new_n302_));
INVX1 INVX1_527 ( .A(u2_u1_b1_last_row_9_), .Y(u2_u1__abc_73914_new_n324_));
INVX1 INVX1_528 ( .A(u2_u1_b0_last_row_3_), .Y(u2_u1__abc_73914_new_n334_));
INVX1 INVX1_529 ( .A(u2_u1_b0_last_row_6_), .Y(u2_u1__abc_73914_new_n341_));
INVX1 INVX1_53 ( .A(u0__abc_74894_new_n1122_), .Y(u0__abc_74894_new_n1130_));
INVX1 INVX1_530 ( .A(u2_u1_b0_last_row_12_), .Y(u2_u1__abc_73914_new_n342_));
INVX1 INVX1_531 ( .A(u2_u1_b0_last_row_2_), .Y(u2_u1__abc_73914_new_n355_));
INVX1 INVX1_532 ( .A(u2_u1_b0_last_row_4_), .Y(u2_u1__abc_73914_new_n356_));
INVX1 INVX1_533 ( .A(u2_u1_b2_last_row_11_), .Y(u2_u1__abc_73914_new_n367_));
INVX1 INVX1_534 ( .A(u2_u1_b2_last_row_4_), .Y(u2_u1__abc_73914_new_n369_));
INVX1 INVX1_535 ( .A(u2_u1_b2_last_row_6_), .Y(u2_u1__abc_73914_new_n374_));
INVX1 INVX1_536 ( .A(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_73914_new_n379_));
INVX1 INVX1_537 ( .A(u2_u1_bank0_open), .Y(u2_u1__abc_73914_new_n398_));
INVX1 INVX1_538 ( .A(u2_u1_bank1_open), .Y(u2_u1__abc_73914_new_n399_));
INVX1 INVX1_539 ( .A(u2_u1__abc_73914_new_n401_), .Y(u2_u1__abc_73914_new_n402_));
INVX1 INVX1_54 ( .A(spec_req_cs_5_), .Y(u0__abc_74894_new_n1134_));
INVX1 INVX1_540 ( .A(u2_bank_clr_1), .Y(u2_u1__abc_73914_new_n404_));
INVX1 INVX1_541 ( .A(u2_u1_bank2_open), .Y(u2_u1__abc_73914_new_n405_));
INVX1 INVX1_542 ( .A(u2_u1_bank3_open), .Y(u2_u1__abc_73914_new_n409_));
INVX1 INVX1_543 ( .A(rst_i), .Y(u2_u1__abc_73914_auto_rtlil_cc_1942_NotGate_71538));
INVX1 INVX1_544 ( .A(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n278_));
INVX1 INVX1_545 ( .A(mc_data_ir_0_), .Y(u3__abc_73372_new_n315_));
INVX1 INVX1_546 ( .A(mc_data_ir_1_), .Y(u3__abc_73372_new_n318_));
INVX1 INVX1_547 ( .A(mc_data_ir_2_), .Y(u3__abc_73372_new_n321_));
INVX1 INVX1_548 ( .A(mc_data_ir_3_), .Y(u3__abc_73372_new_n324_));
INVX1 INVX1_549 ( .A(mc_data_ir_4_), .Y(u3__abc_73372_new_n327_));
INVX1 INVX1_55 ( .A(1'h0), .Y(u0__abc_74894_new_n1135_));
INVX1 INVX1_550 ( .A(mc_data_ir_5_), .Y(u3__abc_73372_new_n330_));
INVX1 INVX1_551 ( .A(mc_data_ir_6_), .Y(u3__abc_73372_new_n333_));
INVX1 INVX1_552 ( .A(mc_data_ir_7_), .Y(u3__abc_73372_new_n336_));
INVX1 INVX1_553 ( .A(pack_le1), .Y(u3__abc_73372_new_n341_));
INVX1 INVX1_554 ( .A(u3__abc_73372_new_n339_), .Y(u3__abc_73372_new_n342_));
INVX1 INVX1_555 ( .A(mc_data_ir_8_), .Y(u3__abc_73372_new_n343_));
INVX1 INVX1_556 ( .A(csc_4_), .Y(u3__abc_73372_new_n344_));
INVX1 INVX1_557 ( .A(mc_data_ir_9_), .Y(u3__abc_73372_new_n351_));
INVX1 INVX1_558 ( .A(mc_data_ir_10_), .Y(u3__abc_73372_new_n356_));
INVX1 INVX1_559 ( .A(mc_data_ir_11_), .Y(u3__abc_73372_new_n361_));
INVX1 INVX1_56 ( .A(spec_req_cs_6_), .Y(u0__abc_74894_new_n1140_));
INVX1 INVX1_560 ( .A(mc_data_ir_12_), .Y(u3__abc_73372_new_n366_));
INVX1 INVX1_561 ( .A(mc_data_ir_13_), .Y(u3__abc_73372_new_n371_));
INVX1 INVX1_562 ( .A(mc_data_ir_14_), .Y(u3__abc_73372_new_n376_));
INVX1 INVX1_563 ( .A(mc_data_ir_15_), .Y(u3__abc_73372_new_n381_));
INVX1 INVX1_564 ( .A(mc_data_od_0_), .Y(u3__abc_73372_new_n402_));
INVX1 INVX1_565 ( .A(mc_data_od_1_), .Y(u3__abc_73372_new_n405_));
INVX1 INVX1_566 ( .A(mc_data_od_2_), .Y(u3__abc_73372_new_n408_));
INVX1 INVX1_567 ( .A(mc_data_od_3_), .Y(u3__abc_73372_new_n411_));
INVX1 INVX1_568 ( .A(mc_data_od_4_), .Y(u3__abc_73372_new_n414_));
INVX1 INVX1_569 ( .A(mc_data_od_5_), .Y(u3__abc_73372_new_n417_));
INVX1 INVX1_57 ( .A(1'h0), .Y(u0__abc_74894_new_n1141_));
INVX1 INVX1_570 ( .A(mc_data_od_6_), .Y(u3__abc_73372_new_n420_));
INVX1 INVX1_571 ( .A(mc_data_od_7_), .Y(u3__abc_73372_new_n423_));
INVX1 INVX1_572 ( .A(mc_data_od_8_), .Y(u3__abc_73372_new_n426_));
INVX1 INVX1_573 ( .A(mc_data_od_9_), .Y(u3__abc_73372_new_n429_));
INVX1 INVX1_574 ( .A(mc_data_od_10_), .Y(u3__abc_73372_new_n432_));
INVX1 INVX1_575 ( .A(mc_data_od_11_), .Y(u3__abc_73372_new_n435_));
INVX1 INVX1_576 ( .A(mc_data_od_12_), .Y(u3__abc_73372_new_n438_));
INVX1 INVX1_577 ( .A(mc_data_od_13_), .Y(u3__abc_73372_new_n441_));
INVX1 INVX1_578 ( .A(mc_data_od_14_), .Y(u3__abc_73372_new_n444_));
INVX1 INVX1_579 ( .A(mc_data_od_15_), .Y(u3__abc_73372_new_n447_));
INVX1 INVX1_58 ( .A(spec_req_cs_7_), .Y(u0__abc_74894_new_n1147_));
INVX1 INVX1_580 ( .A(mc_data_od_16_), .Y(u3__abc_73372_new_n450_));
INVX1 INVX1_581 ( .A(mc_data_od_17_), .Y(u3__abc_73372_new_n453_));
INVX1 INVX1_582 ( .A(mc_data_od_18_), .Y(u3__abc_73372_new_n456_));
INVX1 INVX1_583 ( .A(mc_data_od_19_), .Y(u3__abc_73372_new_n459_));
INVX1 INVX1_584 ( .A(mc_data_od_20_), .Y(u3__abc_73372_new_n462_));
INVX1 INVX1_585 ( .A(mc_data_od_21_), .Y(u3__abc_73372_new_n465_));
INVX1 INVX1_586 ( .A(mc_data_od_22_), .Y(u3__abc_73372_new_n468_));
INVX1 INVX1_587 ( .A(mc_data_od_23_), .Y(u3__abc_73372_new_n471_));
INVX1 INVX1_588 ( .A(mc_data_od_24_), .Y(u3__abc_73372_new_n474_));
INVX1 INVX1_589 ( .A(mc_data_od_25_), .Y(u3__abc_73372_new_n477_));
INVX1 INVX1_59 ( .A(u0__abc_74894_new_n1143_), .Y(u0__abc_74894_new_n1148_));
INVX1 INVX1_590 ( .A(mc_data_od_26_), .Y(u3__abc_73372_new_n480_));
INVX1 INVX1_591 ( .A(mc_data_od_27_), .Y(u3__abc_73372_new_n483_));
INVX1 INVX1_592 ( .A(mc_data_od_28_), .Y(u3__abc_73372_new_n486_));
INVX1 INVX1_593 ( .A(mc_data_od_29_), .Y(u3__abc_73372_new_n489_));
INVX1 INVX1_594 ( .A(mc_data_od_30_), .Y(u3__abc_73372_new_n492_));
INVX1 INVX1_595 ( .A(mc_data_od_31_), .Y(u3__abc_73372_new_n495_));
INVX1 INVX1_596 ( .A(u3_rd_fifo_out_16_), .Y(u3__abc_73372_new_n562_));
INVX1 INVX1_597 ( .A(u3_rd_fifo_out_17_), .Y(u3__abc_73372_new_n566_));
INVX1 INVX1_598 ( .A(u3_rd_fifo_out_18_), .Y(u3__abc_73372_new_n570_));
INVX1 INVX1_599 ( .A(u3_rd_fifo_out_19_), .Y(u3__abc_73372_new_n574_));
INVX1 INVX1_6 ( .A(tms_4_), .Y(_abc_81086_new_n283_));
INVX1 INVX1_60 ( .A(1'h0), .Y(u0__abc_74894_new_n1149_));
INVX1 INVX1_600 ( .A(u3_rd_fifo_out_20_), .Y(u3__abc_73372_new_n578_));
INVX1 INVX1_601 ( .A(u3_rd_fifo_out_21_), .Y(u3__abc_73372_new_n582_));
INVX1 INVX1_602 ( .A(u3_rd_fifo_out_22_), .Y(u3__abc_73372_new_n586_));
INVX1 INVX1_603 ( .A(u3_rd_fifo_out_23_), .Y(u3__abc_73372_new_n590_));
INVX1 INVX1_604 ( .A(u3_rd_fifo_out_24_), .Y(u3__abc_73372_new_n594_));
INVX1 INVX1_605 ( .A(u3_rd_fifo_out_25_), .Y(u3__abc_73372_new_n598_));
INVX1 INVX1_606 ( .A(u3_rd_fifo_out_26_), .Y(u3__abc_73372_new_n602_));
INVX1 INVX1_607 ( .A(u3_rd_fifo_out_27_), .Y(u3__abc_73372_new_n606_));
INVX1 INVX1_608 ( .A(u3_rd_fifo_out_28_), .Y(u3__abc_73372_new_n610_));
INVX1 INVX1_609 ( .A(u3_rd_fifo_out_29_), .Y(u3__abc_73372_new_n614_));
INVX1 INVX1_61 ( .A(1'h0), .Y(u0__abc_74894_new_n1157_));
INVX1 INVX1_610 ( .A(u3_rd_fifo_out_30_), .Y(u3__abc_73372_new_n618_));
INVX1 INVX1_611 ( .A(u3_rd_fifo_out_31_), .Y(u3__abc_73372_new_n622_));
INVX1 INVX1_612 ( .A(wb_stb_i), .Y(u3__abc_73372_new_n626_));
INVX1 INVX1_613 ( .A(wb_we_i), .Y(u3__abc_73372_new_n627_));
INVX1 INVX1_614 ( .A(u3_rd_fifo_out_33_), .Y(u3__abc_73372_new_n634_));
INVX1 INVX1_615 ( .A(\wb_sel_i[1] ), .Y(u3__abc_73372_new_n648_));
INVX1 INVX1_616 ( .A(u3__abc_73372_new_n650_), .Y(u3__abc_73372_new_n651_));
INVX1 INVX1_617 ( .A(u3_rd_fifo_out_34_), .Y(u3__abc_73372_new_n652_));
INVX1 INVX1_618 ( .A(u3__abc_73372_new_n680_), .Y(u3__abc_73372_new_n681_));
INVX1 INVX1_619 ( .A(u3_rd_fifo_out_32_), .Y(u3__abc_73372_new_n684_));
INVX1 INVX1_62 ( .A(1'h0), .Y(u0__abc_74894_new_n1159_));
INVX1 INVX1_620 ( .A(\wb_sel_i[0] ), .Y(u3__abc_73372_new_n696_));
INVX1 INVX1_621 ( .A(u3__abc_73372_new_n700_), .Y(u3__abc_73372_new_n701_));
INVX1 INVX1_622 ( .A(u3_rd_fifo_out_35_), .Y(u3__abc_73372_new_n702_));
INVX1 INVX1_623 ( .A(mc_data_ir_0_), .Y(u3_u0__abc_74260_new_n382_));
INVX1 INVX1_624 ( .A(mc_data_ir_1_), .Y(u3_u0__abc_74260_new_n386_));
INVX1 INVX1_625 ( .A(mc_data_ir_2_), .Y(u3_u0__abc_74260_new_n389_));
INVX1 INVX1_626 ( .A(mc_data_ir_3_), .Y(u3_u0__abc_74260_new_n392_));
INVX1 INVX1_627 ( .A(mc_data_ir_4_), .Y(u3_u0__abc_74260_new_n395_));
INVX1 INVX1_628 ( .A(mc_data_ir_5_), .Y(u3_u0__abc_74260_new_n398_));
INVX1 INVX1_629 ( .A(mc_data_ir_6_), .Y(u3_u0__abc_74260_new_n401_));
INVX1 INVX1_63 ( .A(u0_tms1_0_), .Y(u0__abc_74894_new_n1170_));
INVX1 INVX1_630 ( .A(mc_data_ir_7_), .Y(u3_u0__abc_74260_new_n404_));
INVX1 INVX1_631 ( .A(mc_data_ir_8_), .Y(u3_u0__abc_74260_new_n407_));
INVX1 INVX1_632 ( .A(mc_data_ir_9_), .Y(u3_u0__abc_74260_new_n410_));
INVX1 INVX1_633 ( .A(mc_data_ir_10_), .Y(u3_u0__abc_74260_new_n413_));
INVX1 INVX1_634 ( .A(mc_data_ir_11_), .Y(u3_u0__abc_74260_new_n416_));
INVX1 INVX1_635 ( .A(mc_data_ir_12_), .Y(u3_u0__abc_74260_new_n419_));
INVX1 INVX1_636 ( .A(mc_data_ir_13_), .Y(u3_u0__abc_74260_new_n422_));
INVX1 INVX1_637 ( .A(mc_data_ir_14_), .Y(u3_u0__abc_74260_new_n425_));
INVX1 INVX1_638 ( .A(mc_data_ir_15_), .Y(u3_u0__abc_74260_new_n428_));
INVX1 INVX1_639 ( .A(mc_data_ir_16_), .Y(u3_u0__abc_74260_new_n431_));
INVX1 INVX1_64 ( .A(u0_tms0_0_), .Y(u0__abc_74894_new_n1172_));
INVX1 INVX1_640 ( .A(mc_data_ir_17_), .Y(u3_u0__abc_74260_new_n434_));
INVX1 INVX1_641 ( .A(mc_data_ir_18_), .Y(u3_u0__abc_74260_new_n437_));
INVX1 INVX1_642 ( .A(mc_data_ir_19_), .Y(u3_u0__abc_74260_new_n440_));
INVX1 INVX1_643 ( .A(mc_data_ir_20_), .Y(u3_u0__abc_74260_new_n443_));
INVX1 INVX1_644 ( .A(mc_data_ir_21_), .Y(u3_u0__abc_74260_new_n446_));
INVX1 INVX1_645 ( .A(mc_data_ir_22_), .Y(u3_u0__abc_74260_new_n449_));
INVX1 INVX1_646 ( .A(mc_data_ir_23_), .Y(u3_u0__abc_74260_new_n452_));
INVX1 INVX1_647 ( .A(mc_data_ir_24_), .Y(u3_u0__abc_74260_new_n455_));
INVX1 INVX1_648 ( .A(mc_data_ir_25_), .Y(u3_u0__abc_74260_new_n458_));
INVX1 INVX1_649 ( .A(mc_data_ir_26_), .Y(u3_u0__abc_74260_new_n461_));
INVX1 INVX1_65 ( .A(1'h0), .Y(u0__abc_74894_new_n1177_));
INVX1 INVX1_650 ( .A(mc_data_ir_27_), .Y(u3_u0__abc_74260_new_n464_));
INVX1 INVX1_651 ( .A(mc_data_ir_28_), .Y(u3_u0__abc_74260_new_n467_));
INVX1 INVX1_652 ( .A(mc_data_ir_29_), .Y(u3_u0__abc_74260_new_n470_));
INVX1 INVX1_653 ( .A(mc_data_ir_30_), .Y(u3_u0__abc_74260_new_n473_));
INVX1 INVX1_654 ( .A(mc_data_ir_31_), .Y(u3_u0__abc_74260_new_n476_));
INVX1 INVX1_655 ( .A(mc_data_ir_32_), .Y(u3_u0__abc_74260_new_n479_));
INVX1 INVX1_656 ( .A(mc_data_ir_33_), .Y(u3_u0__abc_74260_new_n482_));
INVX1 INVX1_657 ( .A(mc_data_ir_34_), .Y(u3_u0__abc_74260_new_n485_));
INVX1 INVX1_658 ( .A(mc_data_ir_35_), .Y(u3_u0__abc_74260_new_n488_));
INVX1 INVX1_659 ( .A(u3_u0_rd_adr_0_), .Y(u3_u0__abc_74260_new_n637_));
INVX1 INVX1_66 ( .A(1'h0), .Y(u0__abc_74894_new_n1179_));
INVX1 INVX1_660 ( .A(u3_re), .Y(u3_u0__abc_74260_new_n640_));
INVX1 INVX1_661 ( .A(u3_u0_rd_adr_1_), .Y(u3_u0__abc_74260_new_n641_));
INVX1 INVX1_662 ( .A(u3_rd_fifo_clr), .Y(u3_u0__abc_74260_new_n642_));
INVX1 INVX1_663 ( .A(u3_u0_rd_adr_2_), .Y(u3_u0__abc_74260_new_n645_));
INVX1 INVX1_664 ( .A(u3_u0_rd_adr_3_), .Y(u3_u0__abc_74260_new_n648_));
INVX1 INVX1_665 ( .A(u3_u0_wr_adr_0_), .Y(u3_u0__abc_74260_new_n651_));
INVX1 INVX1_666 ( .A(dv), .Y(u3_u0__abc_74260_new_n654_));
INVX1 INVX1_667 ( .A(rst_i), .Y(u3_u0__abc_74260_auto_rtlil_cc_1942_NotGate_71546));
INVX1 INVX1_668 ( .A(rfr_ack), .Y(u4__abc_74770_new_n94_));
INVX1 INVX1_669 ( .A(u4__abc_74770_new_n97_), .Y(u4__abc_74770_new_n98_));
INVX1 INVX1_67 ( .A(u0_tms1_1_), .Y(u0__abc_74894_new_n1190_));
INVX1 INVX1_670 ( .A(u4_rfr_ce), .Y(u4__abc_74770_new_n101_));
INVX1 INVX1_671 ( .A(u4_rfr_cnt_3_), .Y(u4__abc_74770_new_n106_));
INVX1 INVX1_672 ( .A(u4_rfr_cnt_6_), .Y(u4__abc_74770_new_n117_));
INVX1 INVX1_673 ( .A(u4_rfr_cnt_7_), .Y(u4__abc_74770_new_n122_));
INVX1 INVX1_674 ( .A(u4__abc_74770_new_n123_), .Y(u4__abc_74770_new_n124_));
INVX1 INVX1_675 ( .A(u4_rfr_en), .Y(u4__abc_74770_new_n134_));
INVX1 INVX1_676 ( .A(u4_ps_cnt_0_), .Y(u4__abc_74770_new_n136_));
INVX1 INVX1_677 ( .A(u4_ps_cnt_1_), .Y(u4__abc_74770_new_n140_));
INVX1 INVX1_678 ( .A(u4_ps_cnt_2_), .Y(u4__abc_74770_new_n147_));
INVX1 INVX1_679 ( .A(u4__abc_74770_new_n154_), .Y(u4__abc_74770_new_n155_));
INVX1 INVX1_68 ( .A(u0_tms0_1_), .Y(u0__abc_74894_new_n1192_));
INVX1 INVX1_680 ( .A(u4_ps_cnt_5_), .Y(u4__abc_74770_new_n157_));
INVX1 INVX1_681 ( .A(u4_ps_cnt_7_), .Y(u4__abc_74770_new_n167_));
INVX1 INVX1_682 ( .A(u4_rfr_early), .Y(u4__abc_74770_new_n172_));
INVX1 INVX1_683 ( .A(ref_int_2_), .Y(u4__abc_74770_new_n173_));
INVX1 INVX1_684 ( .A(ref_int_0_), .Y(u4__abc_74770_new_n174_));
INVX1 INVX1_685 ( .A(ref_int_1_), .Y(u4__abc_74770_new_n177_));
INVX1 INVX1_686 ( .A(rst_i), .Y(u4__abc_74770_auto_rtlil_cc_1942_NotGate_71562));
INVX1 INVX1_687 ( .A(u5_burst_cnt_2_), .Y(u5__abc_78290_new_n366_));
INVX1 INVX1_688 ( .A(u5_burst_cnt_10_), .Y(u5__abc_78290_new_n373_));
INVX1 INVX1_689 ( .A(u5_state_31_), .Y(u5__abc_78290_new_n437_));
INVX1 INVX1_69 ( .A(1'h0), .Y(u0__abc_74894_new_n1197_));
INVX1 INVX1_690 ( .A(u5__abc_78290_new_n403_), .Y(u5__abc_78290_new_n466_));
INVX1 INVX1_691 ( .A(u5_state_33_), .Y(u5__abc_78290_new_n467_));
INVX1 INVX1_692 ( .A(u5_state_30_), .Y(u5__abc_78290_new_n481_));
INVX1 INVX1_693 ( .A(u5_wb_cycle), .Y(u5__abc_78290_new_n486_));
INVX1 INVX1_694 ( .A(u5_state_65_), .Y(u5__abc_78290_new_n489_));
INVX1 INVX1_695 ( .A(u5_state_64_), .Y(u5__abc_78290_new_n490_));
INVX1 INVX1_696 ( .A(u5_state_11_), .Y(u5__abc_78290_new_n492_));
INVX1 INVX1_697 ( .A(u5_state_24_), .Y(u5__abc_78290_new_n500_));
INVX1 INVX1_698 ( .A(u5_state_27_), .Y(u5__abc_78290_new_n506_));
INVX1 INVX1_699 ( .A(u5_state_35_), .Y(u5__abc_78290_new_n513_));
INVX1 INVX1_7 ( .A(tms_5_), .Y(_abc_81086_new_n286_));
INVX1 INVX1_70 ( .A(1'h0), .Y(u0__abc_74894_new_n1199_));
INVX1 INVX1_700 ( .A(u5_state_34_), .Y(u5__abc_78290_new_n515_));
INVX1 INVX1_701 ( .A(u5__abc_78290_new_n519_), .Y(u5__abc_78290_new_n520_));
INVX1 INVX1_702 ( .A(u5_state_29_), .Y(u5__abc_78290_new_n522_));
INVX1 INVX1_703 ( .A(u5_state_28_), .Y(u5__abc_78290_new_n523_));
INVX1 INVX1_704 ( .A(u5_state_32_), .Y(u5__abc_78290_new_n530_));
INVX1 INVX1_705 ( .A(u5__abc_78290_new_n542_), .Y(u5__abc_78290_new_n543_));
INVX1 INVX1_706 ( .A(u5_state_26_), .Y(u5__abc_78290_new_n548_));
INVX1 INVX1_707 ( .A(u5_state_18_), .Y(u5__abc_78290_new_n558_));
INVX1 INVX1_708 ( .A(u5__abc_78290_new_n424_), .Y(u5__abc_78290_new_n563_));
INVX1 INVX1_709 ( .A(u5_state_16_), .Y(u5__abc_78290_new_n564_));
INVX1 INVX1_71 ( .A(u0_tms1_2_), .Y(u0__abc_74894_new_n1210_));
INVX1 INVX1_710 ( .A(u5_state_17_), .Y(u5__abc_78290_new_n571_));
INVX1 INVX1_711 ( .A(u5__abc_78290_new_n577_), .Y(u5__abc_78290_new_n578_));
INVX1 INVX1_712 ( .A(u5__abc_78290_new_n434_), .Y(u5__abc_78290_new_n581_));
INVX1 INVX1_713 ( .A(u5_state_25_), .Y(u5__abc_78290_new_n582_));
INVX1 INVX1_714 ( .A(u5_state_23_), .Y(u5__abc_78290_new_n590_));
INVX1 INVX1_715 ( .A(u5_state_22_), .Y(u5__abc_78290_new_n596_));
INVX1 INVX1_716 ( .A(u5__abc_78290_new_n601_), .Y(u5__abc_78290_new_n602_));
INVX1 INVX1_717 ( .A(u5_state_20_), .Y(u5__abc_78290_new_n603_));
INVX1 INVX1_718 ( .A(u5_state_50_), .Y(u5__abc_78290_new_n614_));
INVX1 INVX1_719 ( .A(u5_state_51_), .Y(u5__abc_78290_new_n619_));
INVX1 INVX1_72 ( .A(u0_tms0_2_), .Y(u0__abc_74894_new_n1212_));
INVX1 INVX1_720 ( .A(u5__abc_78290_new_n624_), .Y(u5__abc_78290_new_n625_));
INVX1 INVX1_721 ( .A(u5_state_4_), .Y(u5__abc_78290_new_n627_));
INVX1 INVX1_722 ( .A(u5_state_49_), .Y(u5__abc_78290_new_n632_));
INVX1 INVX1_723 ( .A(u5_state_48_), .Y(u5__abc_78290_new_n634_));
INVX1 INVX1_724 ( .A(u5_state_41_), .Y(u5__abc_78290_new_n643_));
INVX1 INVX1_725 ( .A(u5_state_40_), .Y(u5__abc_78290_new_n644_));
INVX1 INVX1_726 ( .A(u5_state_46_), .Y(u5__abc_78290_new_n655_));
INVX1 INVX1_727 ( .A(u5_state_38_), .Y(u5__abc_78290_new_n662_));
INVX1 INVX1_728 ( .A(u5__abc_78290_new_n666_), .Y(u5__abc_78290_new_n667_));
INVX1 INVX1_729 ( .A(u5__abc_78290_new_n661_), .Y(u5__abc_78290_new_n670_));
INVX1 INVX1_73 ( .A(1'h0), .Y(u0__abc_74894_new_n1217_));
INVX1 INVX1_730 ( .A(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n671_));
INVX1 INVX1_731 ( .A(u5__abc_78290_new_n397_), .Y(u5__abc_78290_new_n672_));
INVX1 INVX1_732 ( .A(u5_state_36_), .Y(u5__abc_78290_new_n677_));
INVX1 INVX1_733 ( .A(u5_state_47_), .Y(u5__abc_78290_new_n686_));
INVX1 INVX1_734 ( .A(u5__abc_78290_new_n687_), .Y(u5__abc_78290_new_n688_));
INVX1 INVX1_735 ( .A(u5_state_44_), .Y(u5__abc_78290_new_n692_));
INVX1 INVX1_736 ( .A(u5_state_39_), .Y(u5__abc_78290_new_n698_));
INVX1 INVX1_737 ( .A(u5_state_45_), .Y(u5__abc_78290_new_n703_));
INVX1 INVX1_738 ( .A(u5_state_42_), .Y(u5__abc_78290_new_n711_));
INVX1 INVX1_739 ( .A(u5_state_9_), .Y(u5__abc_78290_new_n726_));
INVX1 INVX1_74 ( .A(1'h0), .Y(u0__abc_74894_new_n1219_));
INVX1 INVX1_740 ( .A(u5__abc_78290_new_n731_), .Y(u5__abc_78290_new_n732_));
INVX1 INVX1_741 ( .A(u5_state_6_), .Y(u5__abc_78290_new_n733_));
INVX1 INVX1_742 ( .A(u5_state_8_), .Y(u5__abc_78290_new_n741_));
INVX1 INVX1_743 ( .A(u5_state_12_), .Y(u5__abc_78290_new_n747_));
INVX1 INVX1_744 ( .A(u5_state_10_), .Y(u5__abc_78290_new_n757_));
INVX1 INVX1_745 ( .A(u5_state_15_), .Y(u5__abc_78290_new_n763_));
INVX1 INVX1_746 ( .A(u5__abc_78290_new_n764_), .Y(u5__abc_78290_new_n765_));
INVX1 INVX1_747 ( .A(u5_state_5_), .Y(u5__abc_78290_new_n771_));
INVX1 INVX1_748 ( .A(u5_state_7_), .Y(u5__abc_78290_new_n777_));
INVX1 INVX1_749 ( .A(u5__abc_78290_new_n778_), .Y(u5__abc_78290_new_n779_));
INVX1 INVX1_75 ( .A(u0_tms1_3_), .Y(u0__abc_74894_new_n1230_));
INVX1 INVX1_750 ( .A(u5_state_0_), .Y(u5__abc_78290_new_n787_));
INVX1 INVX1_751 ( .A(u5_state_1_), .Y(u5__abc_78290_new_n793_));
INVX1 INVX1_752 ( .A(u5_state_13_), .Y(u5__abc_78290_new_n823_));
INVX1 INVX1_753 ( .A(u5_state_14_), .Y(u5__abc_78290_new_n829_));
INVX1 INVX1_754 ( .A(u5_state_63_), .Y(u5__abc_78290_new_n840_));
INVX1 INVX1_755 ( .A(u5_state_60_), .Y(u5__abc_78290_new_n846_));
INVX1 INVX1_756 ( .A(u5__abc_78290_new_n847_), .Y(u5__abc_78290_new_n848_));
INVX1 INVX1_757 ( .A(u5__abc_78290_new_n378_), .Y(u5__abc_78290_new_n849_));
INVX1 INVX1_758 ( .A(u5_state_61_), .Y(u5__abc_78290_new_n854_));
INVX1 INVX1_759 ( .A(u5__abc_78290_new_n855_), .Y(u5__abc_78290_new_n856_));
INVX1 INVX1_76 ( .A(u0_tms0_3_), .Y(u0__abc_74894_new_n1232_));
INVX1 INVX1_760 ( .A(u5_state_2_), .Y(u5__abc_78290_new_n862_));
INVX1 INVX1_761 ( .A(u5__abc_78290_new_n420_), .Y(u5__abc_78290_new_n864_));
INVX1 INVX1_762 ( .A(u5_state_3_), .Y(u5__abc_78290_new_n869_));
INVX1 INVX1_763 ( .A(u5_mc_adv_r), .Y(u5__abc_78290_new_n887_));
INVX1 INVX1_764 ( .A(u5__abc_78290_new_n894_), .Y(u5__abc_78290_new_n895_));
INVX1 INVX1_765 ( .A(u5_state_37_), .Y(u5__abc_78290_new_n898_));
INVX1 INVX1_766 ( .A(u5_state_59_), .Y(u5__abc_78290_new_n902_));
INVX1 INVX1_767 ( .A(u5_state_58_), .Y(u5__abc_78290_new_n904_));
INVX1 INVX1_768 ( .A(u5_state_57_), .Y(u5__abc_78290_new_n909_));
INVX1 INVX1_769 ( .A(u5_state_56_), .Y(u5__abc_78290_new_n911_));
INVX1 INVX1_77 ( .A(1'h0), .Y(u0__abc_74894_new_n1237_));
INVX1 INVX1_770 ( .A(u5_state_54_), .Y(u5__abc_78290_new_n929_));
INVX1 INVX1_771 ( .A(u5__abc_78290_new_n930_), .Y(u5__abc_78290_new_n931_));
INVX1 INVX1_772 ( .A(u5__abc_78290_new_n386_), .Y(u5__abc_78290_new_n932_));
INVX1 INVX1_773 ( .A(u5_state_53_), .Y(u5__abc_78290_new_n938_));
INVX1 INVX1_774 ( .A(u5__abc_78290_new_n939_), .Y(u5__abc_78290_new_n940_));
INVX1 INVX1_775 ( .A(u5__abc_78290_new_n385_), .Y(u5__abc_78290_new_n941_));
INVX1 INVX1_776 ( .A(u5_state_52_), .Y(u5__abc_78290_new_n946_));
INVX1 INVX1_777 ( .A(u5__abc_78290_new_n947_), .Y(u5__abc_78290_new_n948_));
INVX1 INVX1_778 ( .A(u5_mc_le), .Y(u5__0mc_le_0_0_));
INVX1 INVX1_779 ( .A(u5_timer_6_), .Y(u5__abc_78290_new_n961_));
INVX1 INVX1_78 ( .A(1'h0), .Y(u0__abc_74894_new_n1239_));
INVX1 INVX1_780 ( .A(u5_timer_0_), .Y(u5__abc_78290_new_n962_));
INVX1 INVX1_781 ( .A(u5_ir_cnt_0_), .Y(u5__abc_78290_new_n969_));
INVX1 INVX1_782 ( .A(rfr_req), .Y(u5__abc_78290_new_n974_));
INVX1 INVX1_783 ( .A(u5_state_55_), .Y(u5__abc_78290_new_n976_));
INVX1 INVX1_784 ( .A(u5__abc_78290_new_n977_), .Y(u5__abc_78290_new_n978_));
INVX1 INVX1_785 ( .A(u5__abc_78290_new_n560_), .Y(u5__abc_78290_new_n1013_));
INVX1 INVX1_786 ( .A(u5__abc_78290_new_n379_), .Y(u5__abc_78290_new_n1064_));
INVX1 INVX1_787 ( .A(u5_state_62_), .Y(u5__abc_78290_new_n1065_));
INVX1 INVX1_788 ( .A(u5__abc_78290_new_n1116_), .Y(u5__abc_78290_new_n1117_));
INVX1 INVX1_789 ( .A(u5__abc_78290_new_n622_), .Y(u5__abc_78290_new_n1134_));
INVX1 INVX1_79 ( .A(u0_tms1_4_), .Y(u0__abc_74894_new_n1250_));
INVX1 INVX1_790 ( .A(u5__abc_78290_new_n1135_), .Y(u5__abc_78290_new_n1136_));
INVX1 INVX1_791 ( .A(u5__abc_78290_new_n1147_), .Y(u5__abc_78290_new_n1148_));
INVX1 INVX1_792 ( .A(u5__abc_78290_new_n1156_), .Y(u5__abc_78290_new_n1157_));
INVX1 INVX1_793 ( .A(u5__abc_78290_new_n1186_), .Y(u5__abc_78290_new_n1187_));
INVX1 INVX1_794 ( .A(u5__abc_78290_new_n1190_), .Y(u5__abc_78290_new_n1191_));
INVX1 INVX1_795 ( .A(u5__abc_78290_new_n1196_), .Y(u5__abc_78290_new_n1197_));
INVX1 INVX1_796 ( .A(u5__abc_78290_new_n1199_), .Y(u5__abc_78290_new_n1200_));
INVX1 INVX1_797 ( .A(u5__abc_78290_new_n1211_), .Y(u5__abc_78290_new_n1212_));
INVX1 INVX1_798 ( .A(u5__abc_78290_new_n1224_), .Y(u5__abc_78290_new_n1225_));
INVX1 INVX1_799 ( .A(u5__abc_78290_new_n1267_), .Y(u5__abc_78290_new_n1268_));
INVX1 INVX1_8 ( .A(tms_6_), .Y(_abc_81086_new_n289_));
INVX1 INVX1_80 ( .A(u0_tms0_4_), .Y(u0__abc_74894_new_n1252_));
INVX1 INVX1_800 ( .A(u5__abc_78290_new_n1300_), .Y(u5__abc_78290_new_n1301_));
INVX1 INVX1_801 ( .A(u5__abc_78290_new_n1302_), .Y(u5__abc_78290_new_n1303_));
INVX1 INVX1_802 ( .A(u5__abc_78290_new_n1317_), .Y(u5__abc_78290_new_n1318_));
INVX1 INVX1_803 ( .A(csc_s_1_), .Y(u5__abc_78290_new_n1319_));
INVX1 INVX1_804 ( .A(csc_s_2_), .Y(u5__abc_78290_new_n1320_));
INVX1 INVX1_805 ( .A(u5__abc_78290_new_n1321_), .Y(u5__abc_78290_new_n1322_));
INVX1 INVX1_806 ( .A(u1_wb_write_go), .Y(u5__abc_78290_new_n1324_));
INVX1 INVX1_807 ( .A(u5__abc_78290_new_n1333_), .Y(u5__abc_78290_new_n1334_));
INVX1 INVX1_808 ( .A(u5_lookup_ready2), .Y(u5__abc_78290_new_n1336_));
INVX1 INVX1_809 ( .A(lmr_req), .Y(u5__abc_78290_new_n1337_));
INVX1 INVX1_81 ( .A(1'h0), .Y(u0__abc_74894_new_n1257_));
INVX1 INVX1_810 ( .A(u5_susp_req_r), .Y(u5__abc_78290_new_n1338_));
INVX1 INVX1_811 ( .A(u5__abc_78290_new_n1339_), .Y(u5__abc_78290_new_n1340_));
INVX1 INVX1_812 ( .A(u5__abc_78290_new_n1341_), .Y(u5__abc_78290_new_n1342_));
INVX1 INVX1_813 ( .A(u5__abc_78290_new_n1345_), .Y(u5__abc_78290_new_n1346_));
INVX1 INVX1_814 ( .A(u5__abc_78290_new_n1216_), .Y(u5__abc_78290_new_n1348_));
INVX1 INVX1_815 ( .A(u5__abc_78290_new_n1084_), .Y(u5__abc_78290_new_n1349_));
INVX1 INVX1_816 ( .A(u5__abc_78290_new_n1351_), .Y(u5__abc_78290_new_n1352_));
INVX1 INVX1_817 ( .A(u5__abc_78290_new_n1356_), .Y(u5__abc_78290_new_n1357_));
INVX1 INVX1_818 ( .A(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1361_));
INVX1 INVX1_819 ( .A(u5__abc_78290_new_n574_), .Y(u5__abc_78290_new_n1374_));
INVX1 INVX1_82 ( .A(1'h0), .Y(u0__abc_74894_new_n1259_));
INVX1 INVX1_820 ( .A(u5_tmr_done), .Y(u5__abc_78290_new_n1375_));
INVX1 INVX1_821 ( .A(u5__abc_78290_new_n1052_), .Y(u5__abc_78290_new_n1391_));
INVX1 INVX1_822 ( .A(u5__abc_78290_new_n1120_), .Y(u5__abc_78290_new_n1392_));
INVX1 INVX1_823 ( .A(u5__abc_78290_new_n1394_), .Y(u5__abc_78290_new_n1395_));
INVX1 INVX1_824 ( .A(u5__abc_78290_new_n1085_), .Y(u5__abc_78290_new_n1399_));
INVX1 INVX1_825 ( .A(u5__abc_78290_new_n1401_), .Y(u5__abc_78290_new_n1402_));
INVX1 INVX1_826 ( .A(u5__abc_78290_new_n1404_), .Y(u5__abc_78290_new_n1405_));
INVX1 INVX1_827 ( .A(u5__abc_78290_new_n1273_), .Y(u5__abc_78290_new_n1408_));
INVX1 INVX1_828 ( .A(tms_s_9_), .Y(u5__abc_78290_new_n1409_));
INVX1 INVX1_829 ( .A(u5__abc_78290_new_n1410_), .Y(u5__abc_78290_new_n1411_));
INVX1 INVX1_83 ( .A(u0_tms1_5_), .Y(u0__abc_74894_new_n1270_));
INVX1 INVX1_830 ( .A(u5_wb_wait), .Y(u5__abc_78290_new_n1414_));
INVX1 INVX1_831 ( .A(u5_cke_r), .Y(u5__abc_78290_new_n1416_));
INVX1 INVX1_832 ( .A(u5__abc_78290_new_n1418_), .Y(u5__abc_78290_new_n1419_));
INVX1 INVX1_833 ( .A(u5_cmd_del_0_), .Y(u5__abc_78290_new_n1428_));
INVX1 INVX1_834 ( .A(u1_wr_cycle), .Y(u5__abc_78290_new_n1429_));
INVX1 INVX1_835 ( .A(u5__abc_78290_new_n1316_), .Y(u5__abc_78290_new_n1432_));
INVX1 INVX1_836 ( .A(u5__abc_78290_new_n877_), .Y(u5__abc_78290_new_n1433_));
INVX1 INVX1_837 ( .A(u5__abc_78290_new_n579_), .Y(u5__abc_78290_new_n1437_));
INVX1 INVX1_838 ( .A(u5__abc_78290_new_n1407_), .Y(u5__abc_78290_new_n1446_));
INVX1 INVX1_839 ( .A(u5_cmd_del_1_), .Y(u5__abc_78290_new_n1451_));
INVX1 INVX1_84 ( .A(u0_tms0_5_), .Y(u0__abc_74894_new_n1272_));
INVX1 INVX1_840 ( .A(u5_wb_wait_r), .Y(u5__abc_78290_new_n1455_));
INVX1 INVX1_841 ( .A(u5__abc_78290_new_n1456_), .Y(u5__abc_78290_new_n1457_));
INVX1 INVX1_842 ( .A(u5__abc_78290_new_n1257_), .Y(u5__abc_78290_new_n1458_));
INVX1 INVX1_843 ( .A(u5__abc_78290_new_n1459_), .Y(u5__abc_78290_new_n1460_));
INVX1 INVX1_844 ( .A(u5_cmd_del_2_), .Y(u5__abc_78290_new_n1465_));
INVX1 INVX1_845 ( .A(tms_s_18_), .Y(u5__abc_78290_new_n1473_));
INVX1 INVX1_846 ( .A(u5__abc_78290_new_n1019_), .Y(u5__abc_78290_new_n1478_));
INVX1 INVX1_847 ( .A(u5__abc_78290_new_n1323_), .Y(u5__abc_78290_new_n1486_));
INVX1 INVX1_848 ( .A(u5__abc_78290_new_n1479_), .Y(u5__abc_78290_new_n1488_));
INVX1 INVX1_849 ( .A(u5__abc_78290_new_n1376_), .Y(u5__abc_78290_new_n1490_));
INVX1 INVX1_85 ( .A(1'h0), .Y(u0__abc_74894_new_n1277_));
INVX1 INVX1_850 ( .A(u5__abc_78290_new_n1496_), .Y(u5__abc_78290_new_n1497_));
INVX1 INVX1_851 ( .A(u5__abc_78290_new_n1413_), .Y(u5__abc_78290_new_n1500_));
INVX1 INVX1_852 ( .A(u5__abc_78290_new_n1508_), .Y(u5_cmd_3_));
INVX1 INVX1_853 ( .A(u5__abc_78290_new_n1325_), .Y(u5__abc_78290_new_n1512_));
INVX1 INVX1_854 ( .A(csc_s_3_), .Y(u5__abc_78290_new_n1513_));
INVX1 INVX1_855 ( .A(u5__abc_78290_new_n1368_), .Y(u5__abc_78290_new_n1517_));
INVX1 INVX1_856 ( .A(u5_data_oe_r2), .Y(u5__abc_78290_new_n1522_));
INVX1 INVX1_857 ( .A(u5__abc_78290_new_n986_), .Y(u5__abc_78290_new_n1525_));
INVX1 INVX1_858 ( .A(u5__abc_78290_new_n1527_), .Y(u5__abc_78290_new_n1528_));
INVX1 INVX1_859 ( .A(u5__abc_78290_new_n472_), .Y(u5__abc_78290_new_n1532_));
INVX1 INVX1_86 ( .A(1'h0), .Y(u0__abc_74894_new_n1279_));
INVX1 INVX1_860 ( .A(u5__abc_78290_new_n1305_), .Y(u5__abc_78290_new_n1543_));
INVX1 INVX1_861 ( .A(u5__abc_78290_new_n1544_), .Y(u5__abc_78290_new_n1545_));
INVX1 INVX1_862 ( .A(u5__abc_78290_new_n1282_), .Y(u5__abc_78290_new_n1551_));
INVX1 INVX1_863 ( .A(u5__abc_78290_new_n1563_), .Y(u5__abc_78290_new_n1564_));
INVX1 INVX1_864 ( .A(u5__abc_78290_new_n1567_), .Y(u5__abc_78290_new_n1568_));
INVX1 INVX1_865 ( .A(u5__abc_78290_new_n1570_), .Y(u5__abc_78290_new_n1571_));
INVX1 INVX1_866 ( .A(u5__abc_78290_new_n1562_), .Y(u5__abc_78290_new_n1577_));
INVX1 INVX1_867 ( .A(u5__abc_78290_new_n1534_), .Y(u5__abc_78290_new_n1579_));
INVX1 INVX1_868 ( .A(u5__abc_78290_new_n1535_), .Y(u5__abc_78290_new_n1581_));
INVX1 INVX1_869 ( .A(u5__abc_78290_new_n1542_), .Y(u5__abc_78290_new_n1582_));
INVX1 INVX1_87 ( .A(u0_tms1_6_), .Y(u0__abc_74894_new_n1290_));
INVX1 INVX1_870 ( .A(u5__abc_78290_new_n1593_), .Y(u5__abc_78290_new_n1594_));
INVX1 INVX1_871 ( .A(u5__abc_78290_new_n1595_), .Y(u5__abc_78290_new_n1596_));
INVX1 INVX1_872 ( .A(wb_we_i), .Y(u5__abc_78290_new_n1598_));
INVX1 INVX1_873 ( .A(wb_stb_i), .Y(u5__abc_78290_new_n1599_));
INVX1 INVX1_874 ( .A(u3_wb_read_go), .Y(u5__abc_78290_new_n1600_));
INVX1 INVX1_875 ( .A(u5__abc_78290_new_n1601_), .Y(u5__abc_78290_new_n1602_));
INVX1 INVX1_876 ( .A(u5__abc_78290_new_n1406_), .Y(u5__abc_78290_new_n1608_));
INVX1 INVX1_877 ( .A(u5__abc_78290_new_n1615_), .Y(u5__abc_78290_new_n1616_));
INVX1 INVX1_878 ( .A(u5__abc_78290_new_n1291_), .Y(u5__abc_78290_new_n1619_));
INVX1 INVX1_879 ( .A(u5_ap_en), .Y(u5__abc_78290_new_n1631_));
INVX1 INVX1_88 ( .A(u0_tms0_6_), .Y(u0__abc_74894_new_n1292_));
INVX1 INVX1_880 ( .A(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n1632_));
INVX1 INVX1_881 ( .A(u5__abc_78290_new_n1637_), .Y(u5__abc_78290_new_n1638_));
INVX1 INVX1_882 ( .A(u5__abc_78290_new_n1105_), .Y(u5__abc_78290_new_n1643_));
INVX1 INVX1_883 ( .A(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1649_));
INVX1 INVX1_884 ( .A(tms_s_1_), .Y(u5__abc_78290_new_n1650_));
INVX1 INVX1_885 ( .A(tms_s_0_), .Y(u5__abc_78290_new_n1651_));
INVX1 INVX1_886 ( .A(tms_s_2_), .Y(u5__abc_78290_new_n1656_));
INVX1 INVX1_887 ( .A(u5__abc_78290_new_n1658_), .Y(u5__abc_78290_new_n1659_));
INVX1 INVX1_888 ( .A(u5__abc_78290_new_n1652_), .Y(u5__abc_78290_new_n1660_));
INVX1 INVX1_889 ( .A(u5__abc_78290_new_n1668_), .Y(u5__abc_78290_new_n1669_));
INVX1 INVX1_89 ( .A(1'h0), .Y(u0__abc_74894_new_n1297_));
INVX1 INVX1_890 ( .A(u5__abc_78290_new_n1653_), .Y(u5__abc_78290_new_n1675_));
INVX1 INVX1_891 ( .A(u5__abc_78290_new_n368_), .Y(u5__abc_78290_new_n1679_));
INVX1 INVX1_892 ( .A(u5_burst_cnt_4_), .Y(u5__abc_78290_new_n1692_));
INVX1 INVX1_893 ( .A(u5__abc_78290_new_n1694_), .Y(u5__abc_78290_new_n1695_));
INVX1 INVX1_894 ( .A(u5__abc_78290_new_n1699_), .Y(u5__abc_78290_new_n1700_));
INVX1 INVX1_895 ( .A(u5_burst_cnt_6_), .Y(u5__abc_78290_new_n1706_));
INVX1 INVX1_896 ( .A(u5__abc_78290_new_n1028_), .Y(u5__abc_78290_new_n1711_));
INVX1 INVX1_897 ( .A(u5__abc_78290_new_n1035_), .Y(u5__abc_78290_new_n1712_));
INVX1 INVX1_898 ( .A(u5__abc_78290_new_n1717_), .Y(u5__abc_78290_new_n1718_));
INVX1 INVX1_899 ( .A(u5__abc_78290_new_n1728_), .Y(u5__abc_78290_new_n1729_));
INVX1 INVX1_9 ( .A(tms_7_), .Y(_abc_81086_new_n292_));
INVX1 INVX1_90 ( .A(1'h0), .Y(u0__abc_74894_new_n1299_));
INVX1 INVX1_900 ( .A(u5__abc_78290_new_n1736_), .Y(u5__abc_78290_new_n1737_));
INVX1 INVX1_901 ( .A(u5__abc_78290_new_n1751_), .Y(u5__abc_78290_new_n1752_));
INVX1 INVX1_902 ( .A(u5__abc_78290_new_n1820_), .Y(u5__abc_78290_new_n1821_));
INVX1 INVX1_903 ( .A(u5__abc_78290_new_n1861_), .Y(u5__abc_78290_new_n1862_));
INVX1 INVX1_904 ( .A(u5_burst_cnt_8_), .Y(u5__abc_78290_new_n1961_));
INVX1 INVX1_905 ( .A(u5__abc_78290_new_n369_), .Y(u5__abc_78290_new_n1967_));
INVX1 INVX1_906 ( .A(u5__abc_78290_new_n1193_), .Y(u5__abc_78290_new_n1982_));
INVX1 INVX1_907 ( .A(u5_cmd_asserted), .Y(u5__abc_78290_new_n1990_));
INVX1 INVX1_908 ( .A(u5__abc_78290_new_n536_), .Y(u5__abc_78290_new_n1991_));
INVX1 INVX1_909 ( .A(u5__abc_78290_new_n1283_), .Y(u5__abc_78290_new_n1996_));
INVX1 INVX1_91 ( .A(u0_tms1_7_), .Y(u0__abc_74894_new_n1310_));
INVX1 INVX1_910 ( .A(u5__abc_78290_new_n2005_), .Y(u5__abc_78290_new_n2006_));
INVX1 INVX1_911 ( .A(u5__abc_78290_new_n2010_), .Y(u5__abc_78290_new_n2011_));
INVX1 INVX1_912 ( .A(u5__abc_78290_new_n2018_), .Y(u5__0ir_cnt_3_0__2_));
INVX1 INVX1_913 ( .A(u5__abc_78290_new_n2021_), .Y(u5__0ir_cnt_3_0__3_));
INVX1 INVX1_914 ( .A(u5__abc_78290_new_n1537_), .Y(u5__abc_78290_new_n2023_));
INVX1 INVX1_915 ( .A(u5__abc_78290_new_n2033_), .Y(u5__abc_78290_new_n2034_));
INVX1 INVX1_916 ( .A(u5__abc_78290_new_n768_), .Y(u5__abc_78290_new_n2068_));
INVX1 INVX1_917 ( .A(u5__abc_78290_new_n752_), .Y(u5__abc_78290_new_n2069_));
INVX1 INVX1_918 ( .A(u5__abc_78290_new_n2084_), .Y(u5__abc_78290_new_n2085_));
INVX1 INVX1_919 ( .A(u5__abc_78290_new_n1759_), .Y(u5__abc_78290_new_n2119_));
INVX1 INVX1_92 ( .A(u0_tms0_7_), .Y(u0__abc_74894_new_n1312_));
INVX1 INVX1_920 ( .A(u5__abc_78290_new_n2124_), .Y(u5__abc_78290_new_n2125_));
INVX1 INVX1_921 ( .A(u5__abc_78290_new_n2133_), .Y(u5__abc_78290_new_n2134_));
INVX1 INVX1_922 ( .A(u5__abc_78290_new_n1003_), .Y(u5__abc_78290_new_n2135_));
INVX1 INVX1_923 ( .A(u5__abc_78290_new_n2140_), .Y(u5__abc_78290_new_n2141_));
INVX1 INVX1_924 ( .A(u5__abc_78290_new_n1482_), .Y(u5__abc_78290_new_n2147_));
INVX1 INVX1_925 ( .A(u5__abc_78290_new_n2155_), .Y(u5__abc_78290_new_n2156_));
INVX1 INVX1_926 ( .A(u5__abc_78290_new_n2167_), .Y(u5__abc_78290_new_n2168_));
INVX1 INVX1_927 ( .A(u5__abc_78290_new_n1989_), .Y(u5__abc_78290_new_n2169_));
INVX1 INVX1_928 ( .A(u5__abc_78290_new_n2172_), .Y(u5__abc_78290_new_n2173_));
INVX1 INVX1_929 ( .A(u5__abc_78290_new_n1565_), .Y(u5__abc_78290_new_n2177_));
INVX1 INVX1_93 ( .A(1'h0), .Y(u0__abc_74894_new_n1317_));
INVX1 INVX1_930 ( .A(u5__abc_78290_new_n1062_), .Y(u5__abc_78290_new_n2182_));
INVX1 INVX1_931 ( .A(u5__abc_78290_new_n2188_), .Y(u5__abc_78290_new_n2189_));
INVX1 INVX1_932 ( .A(u5__abc_78290_new_n2199_), .Y(u5__abc_78290_new_n2200_));
INVX1 INVX1_933 ( .A(u5__abc_78290_new_n2210_), .Y(u5__abc_78290_new_n2211_));
INVX1 INVX1_934 ( .A(u5__abc_78290_new_n1043_), .Y(u5__abc_78290_new_n2216_));
INVX1 INVX1_935 ( .A(u5__abc_78290_new_n1063_), .Y(u5__abc_78290_new_n2217_));
INVX1 INVX1_936 ( .A(u5__abc_78290_new_n1089_), .Y(u5__abc_78290_new_n2218_));
INVX1 INVX1_937 ( .A(u5__abc_78290_new_n2225_), .Y(u5__abc_78290_new_n2226_));
INVX1 INVX1_938 ( .A(u5__abc_78290_new_n2234_), .Y(u5__abc_78290_new_n2235_));
INVX1 INVX1_939 ( .A(u5__abc_78290_new_n2244_), .Y(u5__abc_78290_new_n2245_));
INVX1 INVX1_94 ( .A(1'h0), .Y(u0__abc_74894_new_n1319_));
INVX1 INVX1_940 ( .A(tms_s_16_), .Y(u5__abc_78290_new_n2249_));
INVX1 INVX1_941 ( .A(tms_s_21_), .Y(u5__abc_78290_new_n2250_));
INVX1 INVX1_942 ( .A(u5__abc_78290_new_n1655_), .Y(u5__abc_78290_new_n2256_));
INVX1 INVX1_943 ( .A(u5__abc_78290_new_n2259_), .Y(u5__abc_78290_new_n2260_));
INVX1 INVX1_944 ( .A(u5__abc_78290_new_n2264_), .Y(u5__abc_78290_new_n2265_));
INVX1 INVX1_945 ( .A(u5__abc_78290_new_n2248_), .Y(u5__abc_78290_new_n2266_));
INVX1 INVX1_946 ( .A(u5__abc_78290_new_n2251_), .Y(u5__abc_78290_new_n2267_));
INVX1 INVX1_947 ( .A(u5__abc_78290_new_n2276_), .Y(u5__abc_78290_new_n2277_));
INVX1 INVX1_948 ( .A(u5__abc_78290_new_n1580_), .Y(u5__abc_78290_new_n2278_));
INVX1 INVX1_949 ( .A(u5__abc_78290_new_n1185_), .Y(u5__abc_78290_new_n2282_));
INVX1 INVX1_95 ( .A(u0_tms1_8_), .Y(u0__abc_74894_new_n1330_));
INVX1 INVX1_950 ( .A(u5__abc_78290_new_n1999_), .Y(u5__abc_78290_new_n2283_));
INVX1 INVX1_951 ( .A(u5__abc_78290_new_n1201_), .Y(u5__abc_78290_new_n2285_));
INVX1 INVX1_952 ( .A(u5__abc_78290_new_n2292_), .Y(u5__abc_78290_new_n2293_));
INVX1 INVX1_953 ( .A(u5__abc_78290_new_n2303_), .Y(u5__abc_78290_new_n2304_));
INVX1 INVX1_954 ( .A(u5__abc_78290_new_n2308_), .Y(u5__abc_78290_new_n2310_));
INVX1 INVX1_955 ( .A(u5__abc_78290_new_n965_), .Y(u5__abc_78290_new_n2314_));
INVX1 INVX1_956 ( .A(u5__abc_78290_new_n2206_), .Y(u5__abc_78290_new_n2329_));
INVX1 INVX1_957 ( .A(u5__abc_78290_new_n2339_), .Y(u5__abc_78290_new_n2340_));
INVX1 INVX1_958 ( .A(u5__abc_78290_new_n2341_), .Y(u5__abc_78290_new_n2342_));
INVX1 INVX1_959 ( .A(u5__abc_78290_new_n2224_), .Y(u5__abc_78290_new_n2352_));
INVX1 INVX1_96 ( .A(u0_tms0_8_), .Y(u0__abc_74894_new_n1332_));
INVX1 INVX1_960 ( .A(u5__abc_78290_new_n2231_), .Y(u5__abc_78290_new_n2353_));
INVX1 INVX1_961 ( .A(u5__abc_78290_new_n2379_), .Y(u5__abc_78290_new_n2380_));
INVX1 INVX1_962 ( .A(u5__abc_78290_new_n1184_), .Y(u5__abc_78290_new_n2381_));
INVX1 INVX1_963 ( .A(u5_timer2_0_), .Y(u5__abc_78290_new_n2392_));
INVX1 INVX1_964 ( .A(u5_timer2_8_), .Y(u5__abc_78290_new_n2393_));
INVX1 INVX1_965 ( .A(u5_timer2_5_), .Y(u5__abc_78290_new_n2394_));
INVX1 INVX1_966 ( .A(u5_timer2_4_), .Y(u5__abc_78290_new_n2395_));
INVX1 INVX1_967 ( .A(u5__abc_78290_new_n2396_), .Y(u5__abc_78290_new_n2397_));
INVX1 INVX1_968 ( .A(u5__abc_78290_new_n2398_), .Y(u5__abc_78290_new_n2399_));
INVX1 INVX1_969 ( .A(u5__abc_78290_new_n2401_), .Y(u5__abc_78290_new_n2402_));
INVX1 INVX1_97 ( .A(1'h0), .Y(u0__abc_74894_new_n1337_));
INVX1 INVX1_970 ( .A(u5__abc_78290_new_n2404_), .Y(u5__abc_78290_new_n2405_));
INVX1 INVX1_971 ( .A(u5__abc_78290_new_n2281_), .Y(u5__abc_78290_new_n2408_));
INVX1 INVX1_972 ( .A(u5__abc_78290_new_n1986_), .Y(u5__abc_78290_new_n2409_));
INVX1 INVX1_973 ( .A(u5__abc_78290_new_n1441_), .Y(u5__abc_78290_new_n2417_));
INVX1 INVX1_974 ( .A(u5__abc_78290_new_n2228_), .Y(u5__abc_78290_new_n2424_));
INVX1 INVX1_975 ( .A(u5__abc_78290_new_n2367_), .Y(u5__abc_78290_new_n2425_));
INVX1 INVX1_976 ( .A(u5__abc_78290_new_n2426_), .Y(u5__abc_78290_new_n2427_));
INVX1 INVX1_977 ( .A(u5__abc_78290_new_n2429_), .Y(u5__abc_78290_new_n2430_));
INVX1 INVX1_978 ( .A(u5__abc_78290_new_n2422_), .Y(u5__abc_78290_new_n2458_));
INVX1 INVX1_979 ( .A(u5__abc_78290_new_n2230_), .Y(u5__abc_78290_new_n2461_));
INVX1 INVX1_98 ( .A(1'h0), .Y(u0__abc_74894_new_n1339_));
INVX1 INVX1_980 ( .A(u5__abc_78290_new_n2385_), .Y(u5__abc_78290_new_n2465_));
INVX1 INVX1_981 ( .A(u5__abc_78290_new_n2306_), .Y(u5__abc_78290_new_n2478_));
INVX1 INVX1_982 ( .A(u5__abc_78290_new_n2479_), .Y(u5__abc_78290_new_n2480_));
INVX1 INVX1_983 ( .A(u5__abc_78290_new_n2145_), .Y(u5__abc_78290_new_n2484_));
INVX1 INVX1_984 ( .A(u5__abc_78290_new_n2400_), .Y(u5__abc_78290_new_n2487_));
INVX1 INVX1_985 ( .A(u5__abc_78290_new_n2323_), .Y(u5__abc_78290_new_n2499_));
INVX1 INVX1_986 ( .A(u5__abc_78290_new_n2413_), .Y(u5__abc_78290_new_n2500_));
INVX1 INVX1_987 ( .A(u5__abc_78290_new_n2403_), .Y(u5__abc_78290_new_n2511_));
INVX1 INVX1_988 ( .A(u5__abc_78290_new_n2406_), .Y(u5__abc_78290_new_n2526_));
INVX1 INVX1_989 ( .A(u5__abc_78290_new_n2535_), .Y(u5__abc_78290_new_n2536_));
INVX1 INVX1_99 ( .A(u0_tms1_9_), .Y(u0__abc_74894_new_n1350_));
INVX1 INVX1_990 ( .A(u5_no_wb_cycle), .Y(u5__abc_78290_new_n2538_));
INVX1 INVX1_991 ( .A(u5__abc_78290_new_n2541_), .Y(u5__abc_78290_new_n2542_));
INVX1 INVX1_992 ( .A(u5_ack_cnt_2_), .Y(u5__abc_78290_new_n2548_));
INVX1 INVX1_993 ( .A(u5_mc_adv_r1), .Y(u5__abc_78290_new_n2562_));
INVX1 INVX1_994 ( .A(u5_tmr2_done), .Y(u5__abc_78290_new_n2565_));
INVX1 INVX1_995 ( .A(u5__abc_78290_new_n1109_), .Y(u5__abc_78290_new_n2567_));
INVX1 INVX1_996 ( .A(u5__abc_78290_new_n1335_), .Y(u5__abc_78290_new_n2578_));
INVX1 INVX1_997 ( .A(mc_br_r), .Y(u5__abc_78290_new_n2579_));
INVX1 INVX1_998 ( .A(u5__abc_78290_new_n2580_), .Y(u5__abc_78290_new_n2581_));
INVX1 INVX1_999 ( .A(u5__abc_78290_new_n2586_), .Y(u5__abc_78290_new_n2587_));
MUX2X1 MUX2X1_1 ( .A(u0__abc_74894_new_n1104_), .B(u0__abc_74894_new_n1100_), .S(u0_sreq_cs_le), .Y(u0__0spec_req_cs_7_0__0_));
MUX2X1 MUX2X1_10 ( .A(u1_acs_addr_pl1_7_), .B(u1_acs_addr_7_), .S(next_adr), .Y(u1__abc_72801_new_n530_));
MUX2X1 MUX2X1_11 ( .A(u1_acs_addr_pl1_8_), .B(u1_acs_addr_8_), .S(next_adr), .Y(u1__abc_72801_new_n535_));
MUX2X1 MUX2X1_12 ( .A(u1_acs_addr_pl1_9_), .B(u1_acs_addr_9_), .S(next_adr), .Y(u1__abc_72801_new_n541_));
MUX2X1 MUX2X1_13 ( .A(u1_acs_addr_pl1_10_), .B(u1_acs_addr_10_), .S(next_adr), .Y(u1__abc_72801_new_n548_));
MUX2X1 MUX2X1_14 ( .A(u1_acs_addr_pl1_11_), .B(u1_acs_addr_11_), .S(next_adr), .Y(u1__abc_72801_new_n553_));
MUX2X1 MUX2X1_15 ( .A(u1_acs_addr_pl1_12_), .B(u1_acs_addr_12_), .S(next_adr), .Y(u1__abc_72801_new_n558_));
MUX2X1 MUX2X1_16 ( .A(u1_acs_addr_pl1_13_), .B(u1_acs_addr_13_), .S(next_adr), .Y(u1__abc_72801_new_n563_));
MUX2X1 MUX2X1_17 ( .A(u1_acs_addr_pl1_14_), .B(u1_acs_addr_14_), .S(next_adr), .Y(u1__abc_72801_new_n568_));
MUX2X1 MUX2X1_18 ( .A(u1_acs_addr_pl1_15_), .B(u1_acs_addr_15_), .S(next_adr), .Y(u1__abc_72801_new_n573_));
MUX2X1 MUX2X1_19 ( .A(u1_acs_addr_pl1_16_), .B(u1_acs_addr_16_), .S(next_adr), .Y(u1__abc_72801_new_n579_));
MUX2X1 MUX2X1_2 ( .A(mem_ack_r), .B(wb_stb_i), .S(u1_wr_cycle), .Y(u1__abc_72801_new_n461_));
MUX2X1 MUX2X1_20 ( .A(u1_acs_addr_pl1_17_), .B(u1_acs_addr_17_), .S(next_adr), .Y(u1__abc_72801_new_n585_));
MUX2X1 MUX2X1_21 ( .A(u1_acs_addr_pl1_18_), .B(u1_acs_addr_18_), .S(next_adr), .Y(u1__abc_72801_new_n591_));
MUX2X1 MUX2X1_22 ( .A(u1_acs_addr_pl1_19_), .B(u1_acs_addr_19_), .S(next_adr), .Y(u1__abc_72801_new_n596_));
MUX2X1 MUX2X1_23 ( .A(u1_acs_addr_pl1_20_), .B(u1_acs_addr_20_), .S(next_adr), .Y(u1__abc_72801_new_n601_));
MUX2X1 MUX2X1_24 ( .A(u1__abc_72801_new_n603_), .B(u1__abc_72801_new_n601_), .S(u1__abc_72801_new_n498_), .Y(u1__0acs_addr_23_0__20_));
MUX2X1 MUX2X1_25 ( .A(u1_acs_addr_pl1_21_), .B(u1_acs_addr_21_), .S(next_adr), .Y(u1__abc_72801_new_n605_));
MUX2X1 MUX2X1_26 ( .A(u1_acs_addr_pl1_22_), .B(u1_acs_addr_22_), .S(next_adr), .Y(u1__abc_72801_new_n610_));
MUX2X1 MUX2X1_27 ( .A(u1_acs_addr_pl1_23_), .B(u1_acs_addr_23_), .S(next_adr), .Y(u1__abc_72801_new_n615_));
MUX2X1 MUX2X1_28 ( .A(row_adr_0_), .B(u1_col_adr_0_), .S(row_sel), .Y(u1__abc_72801_new_n685_));
MUX2X1 MUX2X1_29 ( .A(row_adr_1_), .B(u1_col_adr_1_), .S(row_sel), .Y(u1__abc_72801_new_n693_));
MUX2X1 MUX2X1_3 ( .A(u1_acs_addr_pl1_0_), .B(u1_acs_addr_0_), .S(next_adr), .Y(u1__abc_72801_new_n492_));
MUX2X1 MUX2X1_30 ( .A(row_adr_3_), .B(u1_col_adr_3_), .S(row_sel), .Y(u1__abc_72801_new_n710_));
MUX2X1 MUX2X1_31 ( .A(row_adr_4_), .B(u1_col_adr_4_), .S(row_sel), .Y(u1__abc_72801_new_n718_));
MUX2X1 MUX2X1_32 ( .A(row_adr_5_), .B(u1_col_adr_5_), .S(row_sel), .Y(u1__abc_72801_new_n726_));
MUX2X1 MUX2X1_33 ( .A(row_adr_6_), .B(u1_col_adr_6_), .S(row_sel), .Y(u1__abc_72801_new_n734_));
MUX2X1 MUX2X1_34 ( .A(row_adr_7_), .B(u1_col_adr_7_), .S(row_sel), .Y(u1__abc_72801_new_n742_));
MUX2X1 MUX2X1_35 ( .A(row_adr_8_), .B(u1_col_adr_8_), .S(row_sel), .Y(u1__abc_72801_new_n750_));
MUX2X1 MUX2X1_36 ( .A(u1_sram_addr_17_), .B(\wb_addr_i[19] ), .S(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n798_));
MUX2X1 MUX2X1_37 ( .A(u1_sram_addr_18_), .B(\wb_addr_i[20] ), .S(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n801_));
MUX2X1 MUX2X1_38 ( .A(u1_sram_addr_19_), .B(\wb_addr_i[21] ), .S(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n804_));
MUX2X1 MUX2X1_39 ( .A(u1_sram_addr_20_), .B(\wb_addr_i[22] ), .S(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n807_));
MUX2X1 MUX2X1_4 ( .A(u1_acs_addr_pl1_1_), .B(u1_acs_addr_1_), .S(next_adr), .Y(u1__abc_72801_new_n499_));
MUX2X1 MUX2X1_40 ( .A(u1_sram_addr_21_), .B(\wb_addr_i[23] ), .S(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n810_));
MUX2X1 MUX2X1_41 ( .A(u1_sram_addr_22_), .B(\wb_addr_i[24] ), .S(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n813_));
MUX2X1 MUX2X1_42 ( .A(u1_sram_addr_23_), .B(\wb_addr_i[25] ), .S(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n816_));
MUX2X1 MUX2X1_43 ( .A(row_adr_10_), .B(cmd_a10), .S(row_sel), .Y(u1__abc_72801_new_n823_));
MUX2X1 MUX2X1_44 ( .A(u5__abc_78290_new_n1954_), .B(u5_burst_cnt_7_), .S(u5__abc_78290_new_n1673_), .Y(u5__abc_78290_new_n1955_));
MUX2X1 MUX2X1_45 ( .A(u5__abc_78290_new_n1970_), .B(u5_burst_cnt_9_), .S(u5__abc_78290_new_n1673_), .Y(u5__abc_78290_new_n1971_));
MUX2X1 MUX2X1_46 ( .A(u5__abc_78290_new_n2360_), .B(u5__abc_78290_new_n2528_), .S(u5__abc_78290_new_n2450_), .Y(u5__abc_78290_new_n2529_));
MUX2X1 MUX2X1_47 ( .A(u5__abc_78290_new_n1416_), .B(u5_wb_wait), .S(u5_cnt), .Y(u5__abc_78290_new_n3009_));
MUX2X1 MUX2X1_5 ( .A(u1_acs_addr_pl1_2_), .B(u1_acs_addr_2_), .S(next_adr), .Y(u1__abc_72801_new_n505_));
MUX2X1 MUX2X1_6 ( .A(u1_acs_addr_pl1_3_), .B(u1_acs_addr_3_), .S(next_adr), .Y(u1__abc_72801_new_n510_));
MUX2X1 MUX2X1_7 ( .A(u1_acs_addr_pl1_4_), .B(u1_acs_addr_4_), .S(next_adr), .Y(u1__abc_72801_new_n515_));
MUX2X1 MUX2X1_8 ( .A(u1_acs_addr_pl1_5_), .B(u1_acs_addr_5_), .S(next_adr), .Y(u1__abc_72801_new_n520_));
MUX2X1 MUX2X1_9 ( .A(u1_acs_addr_pl1_6_), .B(u1_acs_addr_6_), .S(next_adr), .Y(u1__abc_72801_new_n525_));
NAND2X1 NAND2X1_1 ( .A(wb_stb_i), .B(wb_cyc_i), .Y(_abc_81086_new_n465_));
NAND2X1 NAND2X1_10 ( .A(u0__abc_74894_new_n1115_), .B(u0__abc_74894_new_n1130_), .Y(u0__abc_74894_new_n1131_));
NAND2X1 NAND2X1_100 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1362_));
NAND2X1 NAND2X1_1000 ( .A(u0_u0__abc_72207_new_n270_), .B(u0_u0__abc_72207_new_n271_), .Y(u0_u0__0tms_31_0__16_));
NAND2X1 NAND2X1_1001 ( .A(u0_u0__abc_72207_new_n273_), .B(u0_u0__abc_72207_new_n274_), .Y(u0_u0__0tms_31_0__17_));
NAND2X1 NAND2X1_1002 ( .A(u0_u0__abc_72207_new_n276_), .B(u0_u0__abc_72207_new_n277_), .Y(u0_u0__0tms_31_0__18_));
NAND2X1 NAND2X1_1003 ( .A(u0_u0__abc_72207_new_n279_), .B(u0_u0__abc_72207_new_n280_), .Y(u0_u0__0tms_31_0__19_));
NAND2X1 NAND2X1_1004 ( .A(u0_u0__abc_72207_new_n282_), .B(u0_u0__abc_72207_new_n283_), .Y(u0_u0__0tms_31_0__20_));
NAND2X1 NAND2X1_1005 ( .A(u0_u0__abc_72207_new_n285_), .B(u0_u0__abc_72207_new_n286_), .Y(u0_u0__0tms_31_0__21_));
NAND2X1 NAND2X1_1006 ( .A(u0_u0__abc_72207_new_n288_), .B(u0_u0__abc_72207_new_n289_), .Y(u0_u0__0tms_31_0__22_));
NAND2X1 NAND2X1_1007 ( .A(u0_u0__abc_72207_new_n291_), .B(u0_u0__abc_72207_new_n292_), .Y(u0_u0__0tms_31_0__23_));
NAND2X1 NAND2X1_1008 ( .A(u0_u0__abc_72207_new_n294_), .B(u0_u0__abc_72207_new_n295_), .Y(u0_u0__0tms_31_0__24_));
NAND2X1 NAND2X1_1009 ( .A(u0_u0__abc_72207_new_n297_), .B(u0_u0__abc_72207_new_n298_), .Y(u0_u0__0tms_31_0__25_));
NAND2X1 NAND2X1_101 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1365_));
NAND2X1 NAND2X1_1010 ( .A(u0_u0__abc_72207_new_n300_), .B(u0_u0__abc_72207_new_n301_), .Y(u0_u0__0tms_31_0__26_));
NAND2X1 NAND2X1_1011 ( .A(u0_u0__abc_72207_new_n303_), .B(u0_u0__abc_72207_new_n304_), .Y(u0_u0__0tms_31_0__27_));
NAND2X1 NAND2X1_1012 ( .A(u0_u0__abc_72207_new_n306_), .B(u0_u0__abc_72207_new_n307_), .Y(u0_u0__0tms_31_0__28_));
NAND2X1 NAND2X1_1013 ( .A(u0_u0__abc_72207_new_n309_), .B(u0_u0__abc_72207_new_n310_), .Y(u0_u0__0tms_31_0__29_));
NAND2X1 NAND2X1_1014 ( .A(u0_u0__abc_72207_new_n312_), .B(u0_u0__abc_72207_new_n313_), .Y(u0_u0__0tms_31_0__30_));
NAND2X1 NAND2X1_1015 ( .A(u0_u0__abc_72207_new_n315_), .B(u0_u0__abc_72207_new_n316_), .Y(u0_u0__0tms_31_0__31_));
NAND2X1 NAND2X1_1016 ( .A(u0_u0__abc_72207_new_n325_), .B(u0_u0__abc_72207_new_n322_), .Y(u0_u0__abc_72207_new_n326_));
NAND2X1 NAND2X1_1017 ( .A(u0_u0__abc_72207_new_n330_), .B(u0_u0__abc_72207_new_n329_), .Y(u0_u0__0csc_31_0__0_));
NAND2X1 NAND2X1_1018 ( .A(u0_u0_rst_r2), .B(\poc_o[2] ), .Y(u0_u0__abc_72207_new_n332_));
NAND2X1 NAND2X1_1019 ( .A(u0_u0_rst_r2), .B(\poc_o[3] ), .Y(u0_u0__abc_72207_new_n336_));
NAND2X1 NAND2X1_102 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1368_));
NAND2X1 NAND2X1_1020 ( .A(u0_u0_rst_r2), .B(\poc_o[0] ), .Y(u0_u0__abc_72207_new_n342_));
NAND2X1 NAND2X1_1021 ( .A(u0_u0__abc_72207_new_n343_), .B(u0_u0__abc_72207_new_n322_), .Y(u0_u0__abc_72207_new_n344_));
NAND2X1 NAND2X1_1022 ( .A(u0_u0__abc_72207_new_n342_), .B(u0_u0__abc_72207_new_n347_), .Y(u0_u0__0csc_31_0__4_));
NAND2X1 NAND2X1_1023 ( .A(u0_u0_rst_r2), .B(\poc_o[1] ), .Y(u0_u0__abc_72207_new_n349_));
NAND2X1 NAND2X1_1024 ( .A(u0_u0__abc_72207_new_n350_), .B(u0_u0__abc_72207_new_n322_), .Y(u0_u0__abc_72207_new_n351_));
NAND2X1 NAND2X1_1025 ( .A(u0_u0__abc_72207_new_n349_), .B(u0_u0__abc_72207_new_n354_), .Y(u0_u0__0csc_31_0__5_));
NAND2X1 NAND2X1_1026 ( .A(u0_csc0_8_), .B(wb_we_i), .Y(u0_u0__abc_72207_new_n434_));
NAND2X1 NAND2X1_1027 ( .A(u0_u0_init_req_we), .B(u0_u0__abc_72207_new_n463_), .Y(u0_u0__abc_72207_new_n464_));
NAND2X1 NAND2X1_1028 ( .A(u0_u1__abc_72470_new_n202_), .B(u0_u1__abc_72470_new_n203_), .Y(u0_u1__abc_72470_new_n204_));
NAND2X1 NAND2X1_1029 ( .A(u0_u1_inited), .B(u0_u1__abc_72470_new_n205_), .Y(u0_u1__abc_72470_new_n206_));
NAND2X1 NAND2X1_103 ( .A(u0__abc_74894_new_n1356_), .B(u0__abc_74894_new_n1374_), .Y(u0__0sp_tms_31_0__10_));
NAND2X1 NAND2X1_1030 ( .A(u0_lmr_req1), .B(u0_u1__abc_72470_new_n207_), .Y(u0_u1__abc_72470_new_n208_));
NAND2X1 NAND2X1_1031 ( .A(u0_rf_we), .B(u0_u1__abc_72470_new_n211_), .Y(u0_u1__abc_72470_new_n212_));
NAND2X1 NAND2X1_1032 ( .A(u0_csc1_8_), .B(wb_we_i), .Y(u0_u1__abc_72470_new_n411_));
NAND2X1 NAND2X1_1033 ( .A(csc_s_4_), .B(u1__abc_72801_new_n260_), .Y(u1__abc_72801_new_n261_));
NAND2X1 NAND2X1_1034 ( .A(csc_s_6_), .B(u1__abc_72801_new_n262_), .Y(u1__abc_72801_new_n263_));
NAND2X1 NAND2X1_1035 ( .A(csc_s_7_), .B(u1__abc_72801_new_n265_), .Y(u1__abc_72801_new_n266_));
NAND2X1 NAND2X1_1036 ( .A(csc_s_7_), .B(csc_s_6_), .Y(u1__abc_72801_new_n270_));
NAND2X1 NAND2X1_1037 ( .A(u1__abc_72801_new_n273_), .B(u1__abc_72801_new_n268_), .Y(u1__abc_72801_new_n274_));
NAND2X1 NAND2X1_1038 ( .A(csc_s_5_), .B(u1__abc_72801_new_n269_), .Y(u1__abc_72801_new_n288_));
NAND2X1 NAND2X1_1039 ( .A(u1__abc_72801_new_n278_), .B(u1__abc_72801_new_n281_), .Y(u1__abc_72801_new_n291_));
NAND2X1 NAND2X1_104 ( .A(sp_tms_11_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1376_));
NAND2X1 NAND2X1_1040 ( .A(\wb_addr_i[24] ), .B(u1__abc_72801_new_n297_), .Y(u1__abc_72801_new_n298_));
NAND2X1 NAND2X1_1041 ( .A(u1__abc_72801_new_n279_), .B(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n301_));
NAND2X1 NAND2X1_1042 ( .A(\wb_addr_i[23] ), .B(u1__abc_72801_new_n299_), .Y(u1__abc_72801_new_n315_));
NAND2X1 NAND2X1_1043 ( .A(row_adr_0_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n323_));
NAND2X1 NAND2X1_1044 ( .A(row_adr_1_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n331_));
NAND2X1 NAND2X1_1045 ( .A(u1__abc_72801_new_n278_), .B(u1__abc_72801_new_n335_), .Y(u1__abc_72801_new_n336_));
NAND2X1 NAND2X1_1046 ( .A(row_adr_3_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n359_));
NAND2X1 NAND2X1_1047 ( .A(u1__abc_72801_new_n359_), .B(u1__abc_72801_new_n369_), .Y(u1__0row_adr_12_0__3_));
NAND2X1 NAND2X1_1048 ( .A(row_adr_4_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n371_));
NAND2X1 NAND2X1_1049 ( .A(u1__abc_72801_new_n371_), .B(u1__abc_72801_new_n378_), .Y(u1__0row_adr_12_0__4_));
NAND2X1 NAND2X1_105 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1377_), .Y(u0__abc_74894_new_n1378_));
NAND2X1 NAND2X1_1050 ( .A(row_adr_5_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n380_));
NAND2X1 NAND2X1_1051 ( .A(u1__abc_72801_new_n380_), .B(u1__abc_72801_new_n387_), .Y(u1__0row_adr_12_0__5_));
NAND2X1 NAND2X1_1052 ( .A(row_adr_6_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n389_));
NAND2X1 NAND2X1_1053 ( .A(u1__abc_72801_new_n389_), .B(u1__abc_72801_new_n396_), .Y(u1__0row_adr_12_0__6_));
NAND2X1 NAND2X1_1054 ( .A(row_adr_7_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n398_));
NAND2X1 NAND2X1_1055 ( .A(u1__abc_72801_new_n384_), .B(u1__abc_72801_new_n383_), .Y(u1__abc_72801_new_n401_));
NAND2X1 NAND2X1_1056 ( .A(row_adr_8_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n407_));
NAND2X1 NAND2X1_1057 ( .A(u1__abc_72801_new_n412_), .B(u1__abc_72801_new_n413_), .Y(u1__abc_72801_new_n414_));
NAND2X1 NAND2X1_1058 ( .A(row_adr_10_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n430_));
NAND2X1 NAND2X1_1059 ( .A(\wb_addr_i[22] ), .B(u1__abc_72801_new_n267_), .Y(u1__abc_72801_new_n443_));
NAND2X1 NAND2X1_106 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1379_), .Y(u0__abc_74894_new_n1380_));
NAND2X1 NAND2X1_1060 ( .A(\wb_addr_i[24] ), .B(u1__abc_72801_new_n289_), .Y(u1__abc_72801_new_n453_));
NAND2X1 NAND2X1_1061 ( .A(row_adr_12_), .B(u1__abc_72801_new_n322_), .Y(u1__abc_72801_new_n458_));
NAND2X1 NAND2X1_1062 ( .A(u1_col_adr_0_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n462_));
NAND2X1 NAND2X1_1063 ( .A(u1_col_adr_1_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n465_));
NAND2X1 NAND2X1_1064 ( .A(u1_col_adr_2_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n468_));
NAND2X1 NAND2X1_1065 ( .A(u1_col_adr_3_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n471_));
NAND2X1 NAND2X1_1066 ( .A(u1_col_adr_4_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n474_));
NAND2X1 NAND2X1_1067 ( .A(u1_col_adr_5_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n477_));
NAND2X1 NAND2X1_1068 ( .A(u1_col_adr_6_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n480_));
NAND2X1 NAND2X1_1069 ( .A(u1_col_adr_7_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n483_));
NAND2X1 NAND2X1_107 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1381_));
NAND2X1 NAND2X1_1070 ( .A(\wb_addr_i[10] ), .B(u1__abc_72801_new_n273_), .Y(u1__abc_72801_new_n485_));
NAND2X1 NAND2X1_1071 ( .A(u1_col_adr_8_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n486_));
NAND2X1 NAND2X1_1072 ( .A(\wb_addr_i[11] ), .B(page_size_10_), .Y(u1__abc_72801_new_n488_));
NAND2X1 NAND2X1_1073 ( .A(u1_col_adr_9_), .B(u1__abc_72801_new_n461_), .Y(u1__abc_72801_new_n489_));
NAND2X1 NAND2X1_1074 ( .A(\wb_addr_i[1] ), .B(u1__abc_72801_new_n493_), .Y(u1__abc_72801_new_n501_));
NAND2X1 NAND2X1_1075 ( .A(\wb_addr_i[9] ), .B(u1__abc_72801_new_n493_), .Y(u1__abc_72801_new_n544_));
NAND2X1 NAND2X1_1076 ( .A(u1__abc_72801_new_n261_), .B(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n574_));
NAND2X1 NAND2X1_1077 ( .A(\wb_addr_i[18] ), .B(u1__abc_72801_new_n280_), .Y(u1__abc_72801_new_n587_));
NAND2X1 NAND2X1_1078 ( .A(\wb_addr_i[16] ), .B(wb_stb_i), .Y(u1__abc_72801_new_n649_));
NAND2X1 NAND2X1_1079 ( .A(\wb_addr_i[17] ), .B(wb_stb_i), .Y(u1__abc_72801_new_n652_));
NAND2X1 NAND2X1_108 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1382_));
NAND2X1 NAND2X1_1080 ( .A(\wb_addr_i[18] ), .B(wb_stb_i), .Y(u1__abc_72801_new_n655_));
NAND2X1 NAND2X1_1081 ( .A(csc_s_2_), .B(u1__abc_72801_new_n674_), .Y(u1__abc_72801_new_n675_));
NAND2X1 NAND2X1_1082 ( .A(csc_s_1_), .B(u1_wr_hold), .Y(u1__abc_72801_new_n677_));
NAND2X1 NAND2X1_1083 ( .A(u1_sram_addr_0_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n679_));
NAND2X1 NAND2X1_1084 ( .A(u1_sram_addr_1_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n690_));
NAND2X1 NAND2X1_1085 ( .A(u1_sram_addr_2_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n698_));
NAND2X1 NAND2X1_1086 ( .A(row_sel), .B(u1__abc_72801_new_n346_), .Y(u1__abc_72801_new_n701_));
NAND2X1 NAND2X1_1087 ( .A(u1_sram_addr_3_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n707_));
NAND2X1 NAND2X1_1088 ( .A(u1_sram_addr_4_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n715_));
NAND2X1 NAND2X1_1089 ( .A(u1_sram_addr_5_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n723_));
NAND2X1 NAND2X1_109 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1385_));
NAND2X1 NAND2X1_1090 ( .A(u1_sram_addr_6_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n731_));
NAND2X1 NAND2X1_1091 ( .A(u1_sram_addr_7_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n739_));
NAND2X1 NAND2X1_1092 ( .A(u1_sram_addr_8_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n747_));
NAND2X1 NAND2X1_1093 ( .A(u1_sram_addr_9_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n755_));
NAND2X1 NAND2X1_1094 ( .A(row_sel), .B(u1__abc_72801_new_n417_), .Y(u1__abc_72801_new_n758_));
NAND2X1 NAND2X1_1095 ( .A(u1_sram_addr_11_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n764_));
NAND2X1 NAND2X1_1096 ( .A(u1_sram_addr_12_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n772_));
NAND2X1 NAND2X1_1097 ( .A(u1_sram_addr_13_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n780_));
NAND2X1 NAND2X1_1098 ( .A(u1_sram_addr_14_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n785_));
NAND2X1 NAND2X1_1099 ( .A(u1__abc_72801_new_n651_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n790_));
NAND2X1 NAND2X1_11 ( .A(init_req), .B(1'h0), .Y(u0__abc_74894_new_n1136_));
NAND2X1 NAND2X1_110 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1388_));
NAND2X1 NAND2X1_1100 ( .A(u1__abc_72801_new_n654_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n794_));
NAND2X1 NAND2X1_1101 ( .A(u1_sram_addr_10_), .B(u1__abc_72801_new_n678_), .Y(u1__abc_72801_new_n819_));
NAND2X1 NAND2X1_1102 ( .A(tms_s_10_), .B(u1__abc_72801_new_n683_), .Y(u1__abc_72801_new_n824_));
NAND2X1 NAND2X1_1103 ( .A(u1_acs_addr_0_), .B(u1_acs_addr_1_), .Y(u1_u0__abc_72719_new_n52_));
NAND2X1 NAND2X1_1104 ( .A(u1_acs_addr_2_), .B(u1_acs_addr_3_), .Y(u1_u0__abc_72719_new_n57_));
NAND2X1 NAND2X1_1105 ( .A(u1_acs_addr_4_), .B(u1_acs_addr_5_), .Y(u1_u0__abc_72719_new_n68_));
NAND2X1 NAND2X1_1106 ( .A(u1_acs_addr_6_), .B(u1_acs_addr_7_), .Y(u1_u0__abc_72719_new_n69_));
NAND2X1 NAND2X1_1107 ( .A(u1_u0__abc_72719_new_n58_), .B(u1_u0__abc_72719_new_n70_), .Y(u1_u0__abc_72719_new_n71_));
NAND2X1 NAND2X1_1108 ( .A(u1_u0__abc_72719_new_n77_), .B(u1_u0__abc_72719_new_n83_), .Y(u1_u0__abc_72719_new_n84_));
NAND2X1 NAND2X1_1109 ( .A(u1_acs_addr_14_), .B(u1_acs_addr_15_), .Y(u1_u0__abc_72719_new_n99_));
NAND2X1 NAND2X1_111 ( .A(u0__abc_74894_new_n1376_), .B(u0__abc_74894_new_n1394_), .Y(u0__0sp_tms_31_0__11_));
NAND2X1 NAND2X1_1110 ( .A(u1_acs_addr_16_), .B(u1_acs_addr_17_), .Y(u1_u0__abc_72719_new_n103_));
NAND2X1 NAND2X1_1111 ( .A(u1_acs_addr_18_), .B(u1_acs_addr_19_), .Y(u1_u0__abc_72719_new_n108_));
NAND2X1 NAND2X1_1112 ( .A(u1_u0__abc_72719_new_n113_), .B(u1_u0__abc_72719_new_n114_), .Y(u1_u0__abc_72719_new_n115_));
NAND2X1 NAND2X1_1113 ( .A(u1_acs_addr_20_), .B(u1_acs_addr_21_), .Y(u1_u0__abc_72719_new_n119_));
NAND2X1 NAND2X1_1114 ( .A(u1_u0__abc_72719_new_n124_), .B(u1_u0__abc_72719_new_n127_), .Y(u1_acs_addr_pl1_23_));
NAND2X1 NAND2X1_1115 ( .A(u2__abc_74202_new_n102_), .B(u2__abc_74202_new_n105_), .Y(u2__0bank_open_0_0_));
NAND2X1 NAND2X1_1116 ( .A(u2__abc_74202_new_n109_), .B(u2__abc_74202_new_n112_), .Y(u2__0row_same_0_0_));
NAND2X1 NAND2X1_1117 ( .A(bank_adr_0_), .B(bank_adr_1_), .Y(u2_u0__abc_73914_new_n137_));
NAND2X1 NAND2X1_1118 ( .A(u2_bank_set_0), .B(u2_u0__abc_73914_new_n138_), .Y(u2_u0__abc_73914_new_n139_));
NAND2X1 NAND2X1_1119 ( .A(bank_adr_0_), .B(u2_u0__abc_73914_new_n208_), .Y(u2_u0__abc_73914_new_n209_));
NAND2X1 NAND2X1_112 ( .A(sp_tms_12_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1396_));
NAND2X1 NAND2X1_1120 ( .A(u2_bank_set_0), .B(u2_u0__abc_73914_new_n237_), .Y(u2_u0__abc_73914_new_n238_));
NAND2X1 NAND2X1_1121 ( .A(u2_u0_b3_last_row_7_), .B(row_adr_7_), .Y(u2_u0__abc_73914_new_n277_));
NAND2X1 NAND2X1_1122 ( .A(u2_u0_b3_last_row_5_), .B(row_adr_5_), .Y(u2_u0__abc_73914_new_n279_));
NAND2X1 NAND2X1_1123 ( .A(row_adr_4_), .B(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_73914_new_n300_));
NAND2X1 NAND2X1_1124 ( .A(u2_u0__abc_73914_new_n299_), .B(u2_u0__abc_73914_new_n304_), .Y(u2_u0__abc_73914_new_n305_));
NAND2X1 NAND2X1_1125 ( .A(row_adr_8_), .B(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_73914_new_n306_));
NAND2X1 NAND2X1_1126 ( .A(row_adr_6_), .B(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_73914_new_n308_));
NAND2X1 NAND2X1_1127 ( .A(u2_u0_b1_last_row_1_), .B(u2_u0__abc_73914_new_n143_), .Y(u2_u0__abc_73914_new_n315_));
NAND2X1 NAND2X1_1128 ( .A(row_adr_3_), .B(u2_u0__abc_73914_new_n302_), .Y(u2_u0__abc_73914_new_n316_));
NAND2X1 NAND2X1_1129 ( .A(u2_u0_b1_last_row_9_), .B(u2_u0__abc_73914_new_n167_), .Y(u2_u0__abc_73914_new_n319_));
NAND2X1 NAND2X1_113 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1397_), .Y(u0__abc_74894_new_n1398_));
NAND2X1 NAND2X1_1130 ( .A(u2_u0_b1_last_row_5_), .B(u2_u0__abc_73914_new_n155_), .Y(u2_u0__abc_73914_new_n326_));
NAND2X1 NAND2X1_1131 ( .A(u2_u0_b0_last_row_9_), .B(u2_u0__abc_73914_new_n167_), .Y(u2_u0__abc_73914_new_n330_));
NAND2X1 NAND2X1_1132 ( .A(u2_u0_b0_last_row_3_), .B(u2_u0__abc_73914_new_n149_), .Y(u2_u0__abc_73914_new_n336_));
NAND2X1 NAND2X1_1133 ( .A(u2_u0_b0_last_row_2_), .B(u2_u0__abc_73914_new_n146_), .Y(u2_u0__abc_73914_new_n339_));
NAND2X1 NAND2X1_1134 ( .A(u2_u0_b0_last_row_6_), .B(u2_u0__abc_73914_new_n158_), .Y(u2_u0__abc_73914_new_n340_));
NAND2X1 NAND2X1_1135 ( .A(row_adr_0_), .B(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_73914_new_n347_));
NAND2X1 NAND2X1_1136 ( .A(row_adr_1_), .B(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_73914_new_n349_));
NAND2X1 NAND2X1_1137 ( .A(row_adr_7_), .B(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_73914_new_n358_));
NAND2X1 NAND2X1_1138 ( .A(row_adr_10_), .B(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_73914_new_n360_));
NAND2X1 NAND2X1_1139 ( .A(row_adr_7_), .B(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_73914_new_n372_));
NAND2X1 NAND2X1_114 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1399_), .Y(u0__abc_74894_new_n1400_));
NAND2X1 NAND2X1_1140 ( .A(row_adr_3_), .B(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_73914_new_n377_));
NAND2X1 NAND2X1_1141 ( .A(u2_u0__abc_73914_new_n376_), .B(u2_u0__abc_73914_new_n381_), .Y(u2_u0__abc_73914_new_n382_));
NAND2X1 NAND2X1_1142 ( .A(u2_u0_b2_last_row_1_), .B(u2_u0__abc_73914_new_n143_), .Y(u2_u0__abc_73914_new_n392_));
NAND2X1 NAND2X1_1143 ( .A(u2_u0__abc_73914_new_n396_), .B(u2_u0__abc_73914_new_n329_), .Y(u2_row_same_0));
NAND2X1 NAND2X1_1144 ( .A(bank_adr_0_), .B(bank_adr_1_), .Y(u2_u1__abc_73914_new_n137_));
NAND2X1 NAND2X1_1145 ( .A(u2_bank_set_1), .B(u2_u1__abc_73914_new_n138_), .Y(u2_u1__abc_73914_new_n139_));
NAND2X1 NAND2X1_1146 ( .A(bank_adr_0_), .B(u2_u1__abc_73914_new_n208_), .Y(u2_u1__abc_73914_new_n209_));
NAND2X1 NAND2X1_1147 ( .A(u2_bank_set_1), .B(u2_u1__abc_73914_new_n237_), .Y(u2_u1__abc_73914_new_n238_));
NAND2X1 NAND2X1_1148 ( .A(u2_u1_b3_last_row_7_), .B(row_adr_7_), .Y(u2_u1__abc_73914_new_n277_));
NAND2X1 NAND2X1_1149 ( .A(u2_u1_b3_last_row_5_), .B(row_adr_5_), .Y(u2_u1__abc_73914_new_n279_));
NAND2X1 NAND2X1_115 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1401_));
NAND2X1 NAND2X1_1150 ( .A(row_adr_4_), .B(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_73914_new_n300_));
NAND2X1 NAND2X1_1151 ( .A(u2_u1__abc_73914_new_n299_), .B(u2_u1__abc_73914_new_n304_), .Y(u2_u1__abc_73914_new_n305_));
NAND2X1 NAND2X1_1152 ( .A(row_adr_8_), .B(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_73914_new_n306_));
NAND2X1 NAND2X1_1153 ( .A(row_adr_6_), .B(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_73914_new_n308_));
NAND2X1 NAND2X1_1154 ( .A(u2_u1_b1_last_row_1_), .B(u2_u1__abc_73914_new_n143_), .Y(u2_u1__abc_73914_new_n315_));
NAND2X1 NAND2X1_1155 ( .A(row_adr_3_), .B(u2_u1__abc_73914_new_n302_), .Y(u2_u1__abc_73914_new_n316_));
NAND2X1 NAND2X1_1156 ( .A(u2_u1_b1_last_row_9_), .B(u2_u1__abc_73914_new_n167_), .Y(u2_u1__abc_73914_new_n319_));
NAND2X1 NAND2X1_1157 ( .A(u2_u1_b1_last_row_5_), .B(u2_u1__abc_73914_new_n155_), .Y(u2_u1__abc_73914_new_n326_));
NAND2X1 NAND2X1_1158 ( .A(u2_u1_b0_last_row_9_), .B(u2_u1__abc_73914_new_n167_), .Y(u2_u1__abc_73914_new_n330_));
NAND2X1 NAND2X1_1159 ( .A(u2_u1_b0_last_row_3_), .B(u2_u1__abc_73914_new_n149_), .Y(u2_u1__abc_73914_new_n336_));
NAND2X1 NAND2X1_116 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1402_));
NAND2X1 NAND2X1_1160 ( .A(u2_u1_b0_last_row_2_), .B(u2_u1__abc_73914_new_n146_), .Y(u2_u1__abc_73914_new_n339_));
NAND2X1 NAND2X1_1161 ( .A(u2_u1_b0_last_row_6_), .B(u2_u1__abc_73914_new_n158_), .Y(u2_u1__abc_73914_new_n340_));
NAND2X1 NAND2X1_1162 ( .A(row_adr_0_), .B(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_73914_new_n347_));
NAND2X1 NAND2X1_1163 ( .A(row_adr_1_), .B(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_73914_new_n349_));
NAND2X1 NAND2X1_1164 ( .A(row_adr_7_), .B(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_73914_new_n358_));
NAND2X1 NAND2X1_1165 ( .A(row_adr_10_), .B(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_73914_new_n360_));
NAND2X1 NAND2X1_1166 ( .A(row_adr_7_), .B(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_73914_new_n372_));
NAND2X1 NAND2X1_1167 ( .A(row_adr_3_), .B(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_73914_new_n377_));
NAND2X1 NAND2X1_1168 ( .A(u2_u1__abc_73914_new_n376_), .B(u2_u1__abc_73914_new_n381_), .Y(u2_u1__abc_73914_new_n382_));
NAND2X1 NAND2X1_1169 ( .A(u2_u1_b2_last_row_1_), .B(u2_u1__abc_73914_new_n143_), .Y(u2_u1__abc_73914_new_n392_));
NAND2X1 NAND2X1_117 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1405_));
NAND2X1 NAND2X1_1170 ( .A(u2_u1__abc_73914_new_n396_), .B(u2_u1__abc_73914_new_n329_), .Y(u2_row_same_1));
NAND2X1 NAND2X1_1171 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n276_), .Y(u3__abc_73372_new_n277_));
NAND2X1 NAND2X1_1172 ( .A(mc_dp_od_0_), .B(u3__abc_73372_new_n278_), .Y(u3__abc_73372_new_n286_));
NAND2X1 NAND2X1_1173 ( .A(mc_dp_od_1_), .B(u3__abc_73372_new_n278_), .Y(u3__abc_73372_new_n295_));
NAND2X1 NAND2X1_1174 ( .A(mc_dp_od_2_), .B(u3__abc_73372_new_n278_), .Y(u3__abc_73372_new_n304_));
NAND2X1 NAND2X1_1175 ( .A(mc_dp_od_3_), .B(u3__abc_73372_new_n278_), .Y(u3__abc_73372_new_n313_));
NAND2X1 NAND2X1_1176 ( .A(pack_le1), .B(u3__abc_73372_new_n339_), .Y(u3__abc_73372_new_n340_));
NAND2X1 NAND2X1_1177 ( .A(pack_le0), .B(u3__abc_73372_new_n345_), .Y(u3__abc_73372_new_n346_));
NAND2X1 NAND2X1_1178 ( .A(u3_byte1_0_), .B(u3__abc_73372_new_n346_), .Y(u3__abc_73372_new_n347_));
NAND2X1 NAND2X1_1179 ( .A(u3_byte1_1_), .B(u3__abc_73372_new_n346_), .Y(u3__abc_73372_new_n352_));
NAND2X1 NAND2X1_118 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1408_));
NAND2X1 NAND2X1_1180 ( .A(u3_byte1_2_), .B(u3__abc_73372_new_n346_), .Y(u3__abc_73372_new_n357_));
NAND2X1 NAND2X1_1181 ( .A(u3_byte1_3_), .B(u3__abc_73372_new_n346_), .Y(u3__abc_73372_new_n362_));
NAND2X1 NAND2X1_1182 ( .A(u3_byte1_4_), .B(u3__abc_73372_new_n346_), .Y(u3__abc_73372_new_n367_));
NAND2X1 NAND2X1_1183 ( .A(u3_byte1_5_), .B(u3__abc_73372_new_n346_), .Y(u3__abc_73372_new_n372_));
NAND2X1 NAND2X1_1184 ( .A(u3_byte1_6_), .B(u3__abc_73372_new_n346_), .Y(u3__abc_73372_new_n377_));
NAND2X1 NAND2X1_1185 ( .A(u3_byte1_7_), .B(u3__abc_73372_new_n346_), .Y(u3__abc_73372_new_n382_));
NAND2X1 NAND2X1_1186 ( .A(\wb_data_i[0] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n403_));
NAND2X1 NAND2X1_1187 ( .A(\wb_data_i[1] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n406_));
NAND2X1 NAND2X1_1188 ( .A(\wb_data_i[2] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n409_));
NAND2X1 NAND2X1_1189 ( .A(\wb_data_i[3] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n412_));
NAND2X1 NAND2X1_119 ( .A(u0__abc_74894_new_n1396_), .B(u0__abc_74894_new_n1414_), .Y(u0__0sp_tms_31_0__12_));
NAND2X1 NAND2X1_1190 ( .A(\wb_data_i[4] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n415_));
NAND2X1 NAND2X1_1191 ( .A(\wb_data_i[5] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n418_));
NAND2X1 NAND2X1_1192 ( .A(\wb_data_i[6] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n421_));
NAND2X1 NAND2X1_1193 ( .A(\wb_data_i[7] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n424_));
NAND2X1 NAND2X1_1194 ( .A(\wb_data_i[8] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n427_));
NAND2X1 NAND2X1_1195 ( .A(\wb_data_i[9] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n430_));
NAND2X1 NAND2X1_1196 ( .A(\wb_data_i[10] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n433_));
NAND2X1 NAND2X1_1197 ( .A(\wb_data_i[11] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n436_));
NAND2X1 NAND2X1_1198 ( .A(\wb_data_i[12] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n439_));
NAND2X1 NAND2X1_1199 ( .A(\wb_data_i[13] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n442_));
NAND2X1 NAND2X1_12 ( .A(u0__abc_74894_new_n1137_), .B(u0__abc_74894_new_n1129_), .Y(u0__abc_74894_new_n1138_));
NAND2X1 NAND2X1_120 ( .A(sp_tms_13_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1416_));
NAND2X1 NAND2X1_1200 ( .A(\wb_data_i[14] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n445_));
NAND2X1 NAND2X1_1201 ( .A(\wb_data_i[15] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n448_));
NAND2X1 NAND2X1_1202 ( .A(\wb_data_i[16] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n451_));
NAND2X1 NAND2X1_1203 ( .A(\wb_data_i[17] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n454_));
NAND2X1 NAND2X1_1204 ( .A(\wb_data_i[18] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n457_));
NAND2X1 NAND2X1_1205 ( .A(\wb_data_i[19] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n460_));
NAND2X1 NAND2X1_1206 ( .A(\wb_data_i[20] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n463_));
NAND2X1 NAND2X1_1207 ( .A(\wb_data_i[21] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n466_));
NAND2X1 NAND2X1_1208 ( .A(\wb_data_i[22] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n469_));
NAND2X1 NAND2X1_1209 ( .A(\wb_data_i[23] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n472_));
NAND2X1 NAND2X1_121 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1417_), .Y(u0__abc_74894_new_n1418_));
NAND2X1 NAND2X1_1210 ( .A(\wb_data_i[24] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n475_));
NAND2X1 NAND2X1_1211 ( .A(\wb_data_i[25] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n478_));
NAND2X1 NAND2X1_1212 ( .A(\wb_data_i[26] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n481_));
NAND2X1 NAND2X1_1213 ( .A(\wb_data_i[27] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n484_));
NAND2X1 NAND2X1_1214 ( .A(\wb_data_i[28] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n487_));
NAND2X1 NAND2X1_1215 ( .A(\wb_data_i[29] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n490_));
NAND2X1 NAND2X1_1216 ( .A(\wb_data_i[30] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n493_));
NAND2X1 NAND2X1_1217 ( .A(\wb_data_i[31] ), .B(u3__abc_73372_new_n277_), .Y(u3__abc_73372_new_n496_));
NAND2X1 NAND2X1_1218 ( .A(csc_5_), .B(u3__abc_73372_new_n315_), .Y(u3__abc_73372_new_n498_));
NAND2X1 NAND2X1_1219 ( .A(u3_rd_fifo_out_0_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n500_));
NAND2X1 NAND2X1_122 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1419_), .Y(u0__abc_74894_new_n1420_));
NAND2X1 NAND2X1_1220 ( .A(csc_5_), .B(u3__abc_73372_new_n318_), .Y(u3__abc_73372_new_n502_));
NAND2X1 NAND2X1_1221 ( .A(u3_rd_fifo_out_1_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n504_));
NAND2X1 NAND2X1_1222 ( .A(csc_5_), .B(u3__abc_73372_new_n321_), .Y(u3__abc_73372_new_n506_));
NAND2X1 NAND2X1_1223 ( .A(u3_rd_fifo_out_2_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n508_));
NAND2X1 NAND2X1_1224 ( .A(csc_5_), .B(u3__abc_73372_new_n324_), .Y(u3__abc_73372_new_n510_));
NAND2X1 NAND2X1_1225 ( .A(u3_rd_fifo_out_3_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n512_));
NAND2X1 NAND2X1_1226 ( .A(csc_5_), .B(u3__abc_73372_new_n327_), .Y(u3__abc_73372_new_n514_));
NAND2X1 NAND2X1_1227 ( .A(u3_rd_fifo_out_4_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n516_));
NAND2X1 NAND2X1_1228 ( .A(csc_5_), .B(u3__abc_73372_new_n330_), .Y(u3__abc_73372_new_n518_));
NAND2X1 NAND2X1_1229 ( .A(u3_rd_fifo_out_5_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n520_));
NAND2X1 NAND2X1_123 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1421_));
NAND2X1 NAND2X1_1230 ( .A(csc_5_), .B(u3__abc_73372_new_n333_), .Y(u3__abc_73372_new_n522_));
NAND2X1 NAND2X1_1231 ( .A(u3_rd_fifo_out_6_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n524_));
NAND2X1 NAND2X1_1232 ( .A(csc_5_), .B(u3__abc_73372_new_n336_), .Y(u3__abc_73372_new_n526_));
NAND2X1 NAND2X1_1233 ( .A(u3_rd_fifo_out_7_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n528_));
NAND2X1 NAND2X1_1234 ( .A(csc_5_), .B(u3__abc_73372_new_n343_), .Y(u3__abc_73372_new_n530_));
NAND2X1 NAND2X1_1235 ( .A(u3_rd_fifo_out_8_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n532_));
NAND2X1 NAND2X1_1236 ( .A(csc_5_), .B(u3__abc_73372_new_n351_), .Y(u3__abc_73372_new_n534_));
NAND2X1 NAND2X1_1237 ( .A(u3_rd_fifo_out_9_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n536_));
NAND2X1 NAND2X1_1238 ( .A(csc_5_), .B(u3__abc_73372_new_n356_), .Y(u3__abc_73372_new_n538_));
NAND2X1 NAND2X1_1239 ( .A(u3_rd_fifo_out_10_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n540_));
NAND2X1 NAND2X1_124 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1422_));
NAND2X1 NAND2X1_1240 ( .A(csc_5_), .B(u3__abc_73372_new_n361_), .Y(u3__abc_73372_new_n542_));
NAND2X1 NAND2X1_1241 ( .A(u3_rd_fifo_out_11_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n544_));
NAND2X1 NAND2X1_1242 ( .A(csc_5_), .B(u3__abc_73372_new_n366_), .Y(u3__abc_73372_new_n546_));
NAND2X1 NAND2X1_1243 ( .A(u3_rd_fifo_out_12_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n548_));
NAND2X1 NAND2X1_1244 ( .A(csc_5_), .B(u3__abc_73372_new_n371_), .Y(u3__abc_73372_new_n550_));
NAND2X1 NAND2X1_1245 ( .A(u3_rd_fifo_out_13_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n552_));
NAND2X1 NAND2X1_1246 ( .A(csc_5_), .B(u3__abc_73372_new_n376_), .Y(u3__abc_73372_new_n554_));
NAND2X1 NAND2X1_1247 ( .A(u3_rd_fifo_out_14_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n556_));
NAND2X1 NAND2X1_1248 ( .A(csc_5_), .B(u3__abc_73372_new_n381_), .Y(u3__abc_73372_new_n558_));
NAND2X1 NAND2X1_1249 ( .A(u3_rd_fifo_out_15_), .B(u3__abc_73372_new_n275_), .Y(u3__abc_73372_new_n560_));
NAND2X1 NAND2X1_125 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1425_));
NAND2X1 NAND2X1_1250 ( .A(u3_rd_fifo_out_8_), .B(u3_rd_fifo_out_9_), .Y(u3__abc_73372_new_n632_));
NAND2X1 NAND2X1_1251 ( .A(u3__abc_73372_new_n638_), .B(u3__abc_73372_new_n642_), .Y(u3__abc_73372_new_n643_));
NAND2X1 NAND2X1_1252 ( .A(u3_rd_fifo_out_16_), .B(u3_rd_fifo_out_17_), .Y(u3__abc_73372_new_n654_));
NAND2X1 NAND2X1_1253 ( .A(u3_rd_fifo_out_16_), .B(u3__abc_73372_new_n566_), .Y(u3__abc_73372_new_n656_));
NAND2X1 NAND2X1_1254 ( .A(u3_rd_fifo_out_17_), .B(u3__abc_73372_new_n562_), .Y(u3__abc_73372_new_n657_));
NAND2X1 NAND2X1_1255 ( .A(u3__abc_73372_new_n662_), .B(u3__abc_73372_new_n659_), .Y(u3__abc_73372_new_n663_));
NAND2X1 NAND2X1_1256 ( .A(u3__abc_73372_new_n668_), .B(u3__abc_73372_new_n673_), .Y(u3__abc_73372_new_n675_));
NAND2X1 NAND2X1_1257 ( .A(u3_rd_fifo_out_0_), .B(u3_rd_fifo_out_1_), .Y(u3__abc_73372_new_n682_));
NAND2X1 NAND2X1_1258 ( .A(u3__abc_73372_new_n687_), .B(u3__abc_73372_new_n691_), .Y(u3__abc_73372_new_n697_));
NAND2X1 NAND2X1_1259 ( .A(u3_rd_fifo_out_24_), .B(u3_rd_fifo_out_25_), .Y(u3__abc_73372_new_n704_));
NAND2X1 NAND2X1_126 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1428_));
NAND2X1 NAND2X1_1260 ( .A(u3_rd_fifo_out_24_), .B(u3__abc_73372_new_n598_), .Y(u3__abc_73372_new_n706_));
NAND2X1 NAND2X1_1261 ( .A(u3_rd_fifo_out_25_), .B(u3__abc_73372_new_n594_), .Y(u3__abc_73372_new_n707_));
NAND2X1 NAND2X1_1262 ( .A(u3__abc_73372_new_n712_), .B(u3__abc_73372_new_n709_), .Y(u3__abc_73372_new_n713_));
NAND2X1 NAND2X1_1263 ( .A(u3__abc_73372_new_n718_), .B(u3__abc_73372_new_n723_), .Y(u3__abc_73372_new_n725_));
NAND2X1 NAND2X1_1264 ( .A(u3_u0_wr_adr_1_), .B(dv), .Y(u3_u0__abc_74260_new_n383_));
NAND2X1 NAND2X1_1265 ( .A(u3_u0_r1_0_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n384_));
NAND2X1 NAND2X1_1266 ( .A(u3_u0_r1_1_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n387_));
NAND2X1 NAND2X1_1267 ( .A(u3_u0_r1_2_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n390_));
NAND2X1 NAND2X1_1268 ( .A(u3_u0_r1_3_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n393_));
NAND2X1 NAND2X1_1269 ( .A(u3_u0_r1_4_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n396_));
NAND2X1 NAND2X1_127 ( .A(u0__abc_74894_new_n1416_), .B(u0__abc_74894_new_n1434_), .Y(u0__0sp_tms_31_0__13_));
NAND2X1 NAND2X1_1270 ( .A(u3_u0_r1_5_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n399_));
NAND2X1 NAND2X1_1271 ( .A(u3_u0_r1_6_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n402_));
NAND2X1 NAND2X1_1272 ( .A(u3_u0_r1_7_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n405_));
NAND2X1 NAND2X1_1273 ( .A(u3_u0_r1_8_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n408_));
NAND2X1 NAND2X1_1274 ( .A(u3_u0_r1_9_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n411_));
NAND2X1 NAND2X1_1275 ( .A(u3_u0_r1_10_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n414_));
NAND2X1 NAND2X1_1276 ( .A(u3_u0_r1_11_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n417_));
NAND2X1 NAND2X1_1277 ( .A(u3_u0_r1_12_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n420_));
NAND2X1 NAND2X1_1278 ( .A(u3_u0_r1_13_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n423_));
NAND2X1 NAND2X1_1279 ( .A(u3_u0_r1_14_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n426_));
NAND2X1 NAND2X1_128 ( .A(sp_tms_14_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1436_));
NAND2X1 NAND2X1_1280 ( .A(u3_u0_r1_15_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n429_));
NAND2X1 NAND2X1_1281 ( .A(u3_u0_r1_16_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n432_));
NAND2X1 NAND2X1_1282 ( .A(u3_u0_r1_17_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n435_));
NAND2X1 NAND2X1_1283 ( .A(u3_u0_r1_18_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n438_));
NAND2X1 NAND2X1_1284 ( .A(u3_u0_r1_19_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n441_));
NAND2X1 NAND2X1_1285 ( .A(u3_u0_r1_20_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n444_));
NAND2X1 NAND2X1_1286 ( .A(u3_u0_r1_21_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n447_));
NAND2X1 NAND2X1_1287 ( .A(u3_u0_r1_22_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n450_));
NAND2X1 NAND2X1_1288 ( .A(u3_u0_r1_23_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n453_));
NAND2X1 NAND2X1_1289 ( .A(u3_u0_r1_24_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n456_));
NAND2X1 NAND2X1_129 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1437_), .Y(u0__abc_74894_new_n1438_));
NAND2X1 NAND2X1_1290 ( .A(u3_u0_r1_25_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n459_));
NAND2X1 NAND2X1_1291 ( .A(u3_u0_r1_26_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n462_));
NAND2X1 NAND2X1_1292 ( .A(u3_u0_r1_27_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n465_));
NAND2X1 NAND2X1_1293 ( .A(u3_u0_r1_28_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n468_));
NAND2X1 NAND2X1_1294 ( .A(u3_u0_r1_29_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n471_));
NAND2X1 NAND2X1_1295 ( .A(u3_u0_r1_30_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n474_));
NAND2X1 NAND2X1_1296 ( .A(u3_u0_r1_31_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n477_));
NAND2X1 NAND2X1_1297 ( .A(u3_u0_r1_32_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n480_));
NAND2X1 NAND2X1_1298 ( .A(u3_u0_r1_33_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n483_));
NAND2X1 NAND2X1_1299 ( .A(u3_u0_r1_34_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n486_));
NAND2X1 NAND2X1_13 ( .A(init_req), .B(1'h0), .Y(u0__abc_74894_new_n1142_));
NAND2X1 NAND2X1_130 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1439_), .Y(u0__abc_74894_new_n1440_));
NAND2X1 NAND2X1_1300 ( .A(u3_u0_r1_35_), .B(u3_u0__abc_74260_new_n383_), .Y(u3_u0__abc_74260_new_n489_));
NAND2X1 NAND2X1_1301 ( .A(dv), .B(u3_u0_wr_adr_3_), .Y(u3_u0__abc_74260_new_n491_));
NAND2X1 NAND2X1_1302 ( .A(u3_u0_r3_0_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n492_));
NAND2X1 NAND2X1_1303 ( .A(u3_u0_r3_1_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n494_));
NAND2X1 NAND2X1_1304 ( .A(u3_u0_r3_2_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n496_));
NAND2X1 NAND2X1_1305 ( .A(u3_u0_r3_3_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n498_));
NAND2X1 NAND2X1_1306 ( .A(u3_u0_r3_4_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n500_));
NAND2X1 NAND2X1_1307 ( .A(u3_u0_r3_5_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n502_));
NAND2X1 NAND2X1_1308 ( .A(u3_u0_r3_6_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n504_));
NAND2X1 NAND2X1_1309 ( .A(u3_u0_r3_7_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n506_));
NAND2X1 NAND2X1_131 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1441_));
NAND2X1 NAND2X1_1310 ( .A(u3_u0_r3_8_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n508_));
NAND2X1 NAND2X1_1311 ( .A(u3_u0_r3_9_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n510_));
NAND2X1 NAND2X1_1312 ( .A(u3_u0_r3_10_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n512_));
NAND2X1 NAND2X1_1313 ( .A(u3_u0_r3_11_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n514_));
NAND2X1 NAND2X1_1314 ( .A(u3_u0_r3_12_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n516_));
NAND2X1 NAND2X1_1315 ( .A(u3_u0_r3_13_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n518_));
NAND2X1 NAND2X1_1316 ( .A(u3_u0_r3_14_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n520_));
NAND2X1 NAND2X1_1317 ( .A(u3_u0_r3_15_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n522_));
NAND2X1 NAND2X1_1318 ( .A(u3_u0_r3_16_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n524_));
NAND2X1 NAND2X1_1319 ( .A(u3_u0_r3_17_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n526_));
NAND2X1 NAND2X1_132 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1442_));
NAND2X1 NAND2X1_1320 ( .A(u3_u0_r3_18_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n528_));
NAND2X1 NAND2X1_1321 ( .A(u3_u0_r3_19_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n530_));
NAND2X1 NAND2X1_1322 ( .A(u3_u0_r3_20_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n532_));
NAND2X1 NAND2X1_1323 ( .A(u3_u0_r3_21_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n534_));
NAND2X1 NAND2X1_1324 ( .A(u3_u0_r3_22_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n536_));
NAND2X1 NAND2X1_1325 ( .A(u3_u0_r3_23_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n538_));
NAND2X1 NAND2X1_1326 ( .A(u3_u0_r3_24_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n540_));
NAND2X1 NAND2X1_1327 ( .A(u3_u0_r3_25_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n542_));
NAND2X1 NAND2X1_1328 ( .A(u3_u0_r3_26_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n544_));
NAND2X1 NAND2X1_1329 ( .A(u3_u0_r3_27_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n546_));
NAND2X1 NAND2X1_133 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1445_));
NAND2X1 NAND2X1_1330 ( .A(u3_u0_r3_28_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n548_));
NAND2X1 NAND2X1_1331 ( .A(u3_u0_r3_29_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n550_));
NAND2X1 NAND2X1_1332 ( .A(u3_u0_r3_30_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n552_));
NAND2X1 NAND2X1_1333 ( .A(u3_u0_r3_31_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n554_));
NAND2X1 NAND2X1_1334 ( .A(u3_u0_r3_32_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n556_));
NAND2X1 NAND2X1_1335 ( .A(u3_u0_r3_33_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n558_));
NAND2X1 NAND2X1_1336 ( .A(u3_u0_r3_34_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n560_));
NAND2X1 NAND2X1_1337 ( .A(u3_u0_r3_35_), .B(u3_u0__abc_74260_new_n491_), .Y(u3_u0__abc_74260_new_n562_));
NAND2X1 NAND2X1_1338 ( .A(dv), .B(u3_u0_wr_adr_2_), .Y(u3_u0__abc_74260_new_n564_));
NAND2X1 NAND2X1_1339 ( .A(u3_u0_r2_0_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n565_));
NAND2X1 NAND2X1_134 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1448_));
NAND2X1 NAND2X1_1340 ( .A(u3_u0_r2_1_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n567_));
NAND2X1 NAND2X1_1341 ( .A(u3_u0_r2_2_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n569_));
NAND2X1 NAND2X1_1342 ( .A(u3_u0_r2_3_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n571_));
NAND2X1 NAND2X1_1343 ( .A(u3_u0_r2_4_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n573_));
NAND2X1 NAND2X1_1344 ( .A(u3_u0_r2_5_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n575_));
NAND2X1 NAND2X1_1345 ( .A(u3_u0_r2_6_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n577_));
NAND2X1 NAND2X1_1346 ( .A(u3_u0_r2_7_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n579_));
NAND2X1 NAND2X1_1347 ( .A(u3_u0_r2_8_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n581_));
NAND2X1 NAND2X1_1348 ( .A(u3_u0_r2_9_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n583_));
NAND2X1 NAND2X1_1349 ( .A(u3_u0_r2_10_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n585_));
NAND2X1 NAND2X1_135 ( .A(u0__abc_74894_new_n1436_), .B(u0__abc_74894_new_n1454_), .Y(u0__0sp_tms_31_0__14_));
NAND2X1 NAND2X1_1350 ( .A(u3_u0_r2_11_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n587_));
NAND2X1 NAND2X1_1351 ( .A(u3_u0_r2_12_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n589_));
NAND2X1 NAND2X1_1352 ( .A(u3_u0_r2_13_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n591_));
NAND2X1 NAND2X1_1353 ( .A(u3_u0_r2_14_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n593_));
NAND2X1 NAND2X1_1354 ( .A(u3_u0_r2_15_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n595_));
NAND2X1 NAND2X1_1355 ( .A(u3_u0_r2_16_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n597_));
NAND2X1 NAND2X1_1356 ( .A(u3_u0_r2_17_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n599_));
NAND2X1 NAND2X1_1357 ( .A(u3_u0_r2_18_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n601_));
NAND2X1 NAND2X1_1358 ( .A(u3_u0_r2_19_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n603_));
NAND2X1 NAND2X1_1359 ( .A(u3_u0_r2_20_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n605_));
NAND2X1 NAND2X1_136 ( .A(sp_tms_15_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1456_));
NAND2X1 NAND2X1_1360 ( .A(u3_u0_r2_21_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n607_));
NAND2X1 NAND2X1_1361 ( .A(u3_u0_r2_22_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n609_));
NAND2X1 NAND2X1_1362 ( .A(u3_u0_r2_23_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n611_));
NAND2X1 NAND2X1_1363 ( .A(u3_u0_r2_24_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n613_));
NAND2X1 NAND2X1_1364 ( .A(u3_u0_r2_25_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n615_));
NAND2X1 NAND2X1_1365 ( .A(u3_u0_r2_26_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n617_));
NAND2X1 NAND2X1_1366 ( .A(u3_u0_r2_27_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n619_));
NAND2X1 NAND2X1_1367 ( .A(u3_u0_r2_28_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n621_));
NAND2X1 NAND2X1_1368 ( .A(u3_u0_r2_29_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n623_));
NAND2X1 NAND2X1_1369 ( .A(u3_u0_r2_30_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n625_));
NAND2X1 NAND2X1_137 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1457_), .Y(u0__abc_74894_new_n1458_));
NAND2X1 NAND2X1_1370 ( .A(u3_u0_r2_31_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n627_));
NAND2X1 NAND2X1_1371 ( .A(u3_u0_r2_32_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n629_));
NAND2X1 NAND2X1_1372 ( .A(u3_u0_r2_33_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n631_));
NAND2X1 NAND2X1_1373 ( .A(u3_u0_r2_34_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n633_));
NAND2X1 NAND2X1_1374 ( .A(u3_u0_r2_35_), .B(u3_u0__abc_74260_new_n564_), .Y(u3_u0__abc_74260_new_n635_));
NAND2X1 NAND2X1_1375 ( .A(u3_u0_wr_adr_2_), .B(u3_u0__abc_74260_new_n654_), .Y(u3_u0__abc_74260_new_n658_));
NAND2X1 NAND2X1_1376 ( .A(u3_u0_wr_adr_3_), .B(u3_u0__abc_74260_new_n654_), .Y(u3_u0__abc_74260_new_n660_));
NAND2X1 NAND2X1_1377 ( .A(u3_u0_rd_adr_1_), .B(u3_u0__abc_74260_new_n645_), .Y(u3_u0__abc_74260_new_n735_));
NAND2X1 NAND2X1_1378 ( .A(u3_u0_r3_0_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n743_));
NAND2X1 NAND2X1_1379 ( .A(u3_u0__abc_74260_new_n637_), .B(u3_u0__abc_74260_new_n641_), .Y(u3_u0__abc_74260_new_n745_));
NAND2X1 NAND2X1_138 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1459_), .Y(u0__abc_74894_new_n1460_));
NAND2X1 NAND2X1_1380 ( .A(u3_u0_rd_adr_2_), .B(u3_u0__abc_74260_new_n648_), .Y(u3_u0__abc_74260_new_n746_));
NAND2X1 NAND2X1_1381 ( .A(u3_u0_r3_1_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n751_));
NAND2X1 NAND2X1_1382 ( .A(u3_u0_r3_2_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n755_));
NAND2X1 NAND2X1_1383 ( .A(u3_u0_r3_3_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n759_));
NAND2X1 NAND2X1_1384 ( .A(u3_u0_r3_4_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n763_));
NAND2X1 NAND2X1_1385 ( .A(u3_u0_r3_5_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n767_));
NAND2X1 NAND2X1_1386 ( .A(u3_u0_r3_6_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n771_));
NAND2X1 NAND2X1_1387 ( .A(u3_u0_r3_7_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n775_));
NAND2X1 NAND2X1_1388 ( .A(u3_u0_r3_8_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n779_));
NAND2X1 NAND2X1_1389 ( .A(u3_u0_r3_9_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n783_));
NAND2X1 NAND2X1_139 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1461_));
NAND2X1 NAND2X1_1390 ( .A(u3_u0_r3_10_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n787_));
NAND2X1 NAND2X1_1391 ( .A(u3_u0_r3_11_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n791_));
NAND2X1 NAND2X1_1392 ( .A(u3_u0_r3_12_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n795_));
NAND2X1 NAND2X1_1393 ( .A(u3_u0_r3_13_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n799_));
NAND2X1 NAND2X1_1394 ( .A(u3_u0_r3_14_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n803_));
NAND2X1 NAND2X1_1395 ( .A(u3_u0_r3_15_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n807_));
NAND2X1 NAND2X1_1396 ( .A(u3_u0_r3_16_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n811_));
NAND2X1 NAND2X1_1397 ( .A(u3_u0_r3_17_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n815_));
NAND2X1 NAND2X1_1398 ( .A(u3_u0_r3_18_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n819_));
NAND2X1 NAND2X1_1399 ( .A(u3_u0_r3_19_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n823_));
NAND2X1 NAND2X1_14 ( .A(u0__abc_74894_new_n1143_), .B(u0__abc_74894_new_n1144_), .Y(u0__abc_74894_new_n1145_));
NAND2X1 NAND2X1_140 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1462_));
NAND2X1 NAND2X1_1400 ( .A(u3_u0_r3_20_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n827_));
NAND2X1 NAND2X1_1401 ( .A(u3_u0_r3_21_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n831_));
NAND2X1 NAND2X1_1402 ( .A(u3_u0_r3_22_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n835_));
NAND2X1 NAND2X1_1403 ( .A(u3_u0_r3_23_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n839_));
NAND2X1 NAND2X1_1404 ( .A(u3_u0_r3_24_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n843_));
NAND2X1 NAND2X1_1405 ( .A(u3_u0_r3_25_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n847_));
NAND2X1 NAND2X1_1406 ( .A(u3_u0_r3_26_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n851_));
NAND2X1 NAND2X1_1407 ( .A(u3_u0_r3_27_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n855_));
NAND2X1 NAND2X1_1408 ( .A(u3_u0_r3_28_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n859_));
NAND2X1 NAND2X1_1409 ( .A(u3_u0_r3_29_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n863_));
NAND2X1 NAND2X1_141 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1465_));
NAND2X1 NAND2X1_1410 ( .A(u3_u0_r3_30_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n867_));
NAND2X1 NAND2X1_1411 ( .A(u3_u0_r3_31_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n871_));
NAND2X1 NAND2X1_1412 ( .A(u3_u0_r3_32_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n875_));
NAND2X1 NAND2X1_1413 ( .A(u3_u0_r3_33_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n879_));
NAND2X1 NAND2X1_1414 ( .A(u3_u0_r3_34_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n883_));
NAND2X1 NAND2X1_1415 ( .A(u3_u0_r3_35_), .B(u3_u0__abc_74260_new_n742_), .Y(u3_u0__abc_74260_new_n887_));
NAND2X1 NAND2X1_1416 ( .A(u4_ps_cnt_3_), .B(rfr_ps_val_3_), .Y(u4__abc_74770_new_n72_));
NAND2X1 NAND2X1_1417 ( .A(u4_ps_cnt_2_), .B(rfr_ps_val_2_), .Y(u4__abc_74770_new_n74_));
NAND2X1 NAND2X1_1418 ( .A(u4_ps_cnt_7_), .B(rfr_ps_val_7_), .Y(u4__abc_74770_new_n77_));
NAND2X1 NAND2X1_1419 ( .A(u4_ps_cnt_6_), .B(rfr_ps_val_6_), .Y(u4__abc_74770_new_n79_));
NAND2X1 NAND2X1_142 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1468_));
NAND2X1 NAND2X1_1420 ( .A(u4__abc_74770_new_n75_), .B(u4__abc_74770_new_n80_), .Y(u4__abc_74770_new_n81_));
NAND2X1 NAND2X1_1421 ( .A(u4_ps_cnt_0_), .B(rfr_ps_val_0_), .Y(u4__abc_74770_new_n85_));
NAND2X1 NAND2X1_1422 ( .A(u4_ps_cnt_1_), .B(rfr_ps_val_1_), .Y(u4__abc_74770_new_n86_));
NAND2X1 NAND2X1_1423 ( .A(u4_rfr_cnt_1_), .B(u4__abc_74770_new_n93_), .Y(u4__abc_74770_new_n97_));
NAND2X1 NAND2X1_1424 ( .A(u4_rfr_cnt_3_), .B(u4_rfr_cnt_4_), .Y(u4__abc_74770_new_n111_));
NAND2X1 NAND2X1_1425 ( .A(u4_rfr_cnt_5_), .B(u4__abc_74770_new_n112_), .Y(u4__abc_74770_new_n118_));
NAND2X1 NAND2X1_1426 ( .A(u4_rfr_cnt_5_), .B(u4_rfr_cnt_6_), .Y(u4__abc_74770_new_n123_));
NAND2X1 NAND2X1_1427 ( .A(u4_ps_cnt_0_), .B(u4__abc_74770_new_n134_), .Y(u4__abc_74770_new_n135_));
NAND2X1 NAND2X1_1428 ( .A(u4_rfr_en), .B(u4__abc_74770_new_n136_), .Y(u4__abc_74770_new_n137_));
NAND2X1 NAND2X1_1429 ( .A(u4__abc_74770_new_n139_), .B(u4__abc_74770_new_n141_), .Y(u4__abc_74770_new_n142_));
NAND2X1 NAND2X1_143 ( .A(u0__abc_74894_new_n1456_), .B(u0__abc_74894_new_n1474_), .Y(u0__0sp_tms_31_0__15_));
NAND2X1 NAND2X1_1430 ( .A(u4_ps_cnt_2_), .B(u4__abc_74770_new_n139_), .Y(u4__abc_74770_new_n145_));
NAND2X1 NAND2X1_1431 ( .A(u4_ps_cnt_3_), .B(u4__abc_74770_new_n148_), .Y(u4__abc_74770_new_n151_));
NAND2X1 NAND2X1_1432 ( .A(u4__abc_74770_new_n155_), .B(u4__abc_74770_new_n148_), .Y(u4__abc_74770_new_n156_));
NAND2X1 NAND2X1_1433 ( .A(u4__abc_74770_new_n157_), .B(u4__abc_74770_new_n158_), .Y(u4__abc_74770_new_n159_));
NAND2X1 NAND2X1_1434 ( .A(u4__abc_74770_new_n156_), .B(u4__abc_74770_new_n159_), .Y(u4__abc_74770_new_n160_));
NAND2X1 NAND2X1_1435 ( .A(u4__abc_74770_new_n167_), .B(u4__abc_74770_new_n168_), .Y(u4__abc_74770_new_n169_));
NAND2X1 NAND2X1_1436 ( .A(u4__abc_74770_new_n166_), .B(u4__abc_74770_new_n169_), .Y(u4__abc_74770_new_n170_));
NAND2X1 NAND2X1_1437 ( .A(u4_rfr_cnt_0_), .B(u4__abc_74770_new_n177_), .Y(u4__abc_74770_new_n178_));
NAND2X1 NAND2X1_1438 ( .A(u4__abc_74770_new_n173_), .B(u4__abc_74770_new_n179_), .Y(u4__abc_74770_new_n180_));
NAND2X1 NAND2X1_1439 ( .A(u5__abc_78290_new_n366_), .B(u5__abc_78290_new_n367_), .Y(u5__abc_78290_new_n368_));
NAND2X1 NAND2X1_144 ( .A(sp_tms_16_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1476_));
NAND2X1 NAND2X1_1440 ( .A(u5__abc_78290_new_n370_), .B(u5__abc_78290_new_n371_), .Y(u5__abc_78290_new_n372_));
NAND2X1 NAND2X1_1441 ( .A(u5__abc_78290_new_n373_), .B(u5__abc_78290_new_n374_), .Y(u5__abc_78290_new_n375_));
NAND2X1 NAND2X1_1442 ( .A(u5__abc_78290_new_n369_), .B(u5__abc_78290_new_n376_), .Y(u5__0burst_act_rd_0_0_));
NAND2X1 NAND2X1_1443 ( .A(u5__abc_78290_new_n380_), .B(u5__abc_78290_new_n383_), .Y(u5__abc_78290_new_n384_));
NAND2X1 NAND2X1_1444 ( .A(u5__abc_78290_new_n387_), .B(u5__abc_78290_new_n390_), .Y(u5__abc_78290_new_n391_));
NAND2X1 NAND2X1_1445 ( .A(u5__abc_78290_new_n395_), .B(u5__abc_78290_new_n398_), .Y(u5__abc_78290_new_n399_));
NAND2X1 NAND2X1_1446 ( .A(u5__abc_78290_new_n402_), .B(u5__abc_78290_new_n405_), .Y(u5__abc_78290_new_n406_));
NAND2X1 NAND2X1_1447 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n408_));
NAND2X1 NAND2X1_1448 ( .A(u5__abc_78290_new_n411_), .B(u5__abc_78290_new_n414_), .Y(u5__abc_78290_new_n415_));
NAND2X1 NAND2X1_1449 ( .A(u5__abc_78290_new_n418_), .B(u5__abc_78290_new_n421_), .Y(u5__abc_78290_new_n422_));
NAND2X1 NAND2X1_145 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1477_), .Y(u0__abc_74894_new_n1478_));
NAND2X1 NAND2X1_1450 ( .A(u5__abc_78290_new_n424_), .B(u5__abc_78290_new_n425_), .Y(u5__abc_78290_new_n426_));
NAND2X1 NAND2X1_1451 ( .A(u5__abc_78290_new_n431_), .B(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n432_));
NAND2X1 NAND2X1_1452 ( .A(u5__abc_78290_new_n434_), .B(u5__abc_78290_new_n435_), .Y(u5__abc_78290_new_n436_));
NAND2X1 NAND2X1_1453 ( .A(u5__abc_78290_new_n440_), .B(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n441_));
NAND2X1 NAND2X1_1454 ( .A(u5__abc_78290_new_n409_), .B(u5__abc_78290_new_n410_), .Y(u5__abc_78290_new_n442_));
NAND2X1 NAND2X1_1455 ( .A(u5__abc_78290_new_n412_), .B(u5__abc_78290_new_n413_), .Y(u5__abc_78290_new_n443_));
NAND2X1 NAND2X1_1456 ( .A(u5__abc_78290_new_n416_), .B(u5__abc_78290_new_n417_), .Y(u5__abc_78290_new_n445_));
NAND2X1 NAND2X1_1457 ( .A(u5__abc_78290_new_n419_), .B(u5__abc_78290_new_n420_), .Y(u5__abc_78290_new_n446_));
NAND2X1 NAND2X1_1458 ( .A(u5__abc_78290_new_n444_), .B(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n448_));
NAND2X1 NAND2X1_1459 ( .A(u5__abc_78290_new_n427_), .B(u5__abc_78290_new_n429_), .Y(u5__abc_78290_new_n449_));
NAND2X1 NAND2X1_146 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1479_), .Y(u0__abc_74894_new_n1480_));
NAND2X1 NAND2X1_1460 ( .A(u5__abc_78290_new_n438_), .B(u5__abc_78290_new_n451_), .Y(u5__abc_78290_new_n452_));
NAND2X1 NAND2X1_1461 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n453_), .Y(u5__abc_78290_new_n454_));
NAND2X1 NAND2X1_1462 ( .A(u5__abc_78290_new_n378_), .B(u5__abc_78290_new_n379_), .Y(u5__abc_78290_new_n456_));
NAND2X1 NAND2X1_1463 ( .A(u5__abc_78290_new_n381_), .B(u5__abc_78290_new_n382_), .Y(u5__abc_78290_new_n457_));
NAND2X1 NAND2X1_1464 ( .A(u5__abc_78290_new_n385_), .B(u5__abc_78290_new_n386_), .Y(u5__abc_78290_new_n459_));
NAND2X1 NAND2X1_1465 ( .A(u5__abc_78290_new_n388_), .B(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n460_));
NAND2X1 NAND2X1_1466 ( .A(u5__abc_78290_new_n458_), .B(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n462_));
NAND2X1 NAND2X1_1467 ( .A(u5__abc_78290_new_n393_), .B(u5__abc_78290_new_n394_), .Y(u5__abc_78290_new_n463_));
NAND2X1 NAND2X1_1468 ( .A(u5__abc_78290_new_n396_), .B(u5__abc_78290_new_n397_), .Y(u5__abc_78290_new_n464_));
NAND2X1 NAND2X1_1469 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n471_), .Y(u5__abc_78290_new_n472_));
NAND2X1 NAND2X1_147 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1481_));
NAND2X1 NAND2X1_1470 ( .A(u5__abc_78290_new_n400_), .B(u5__abc_78290_new_n401_), .Y(u5__abc_78290_new_n474_));
NAND2X1 NAND2X1_1471 ( .A(u5__abc_78290_new_n403_), .B(u5__abc_78290_new_n404_), .Y(u5__abc_78290_new_n475_));
NAND2X1 NAND2X1_1472 ( .A(u5__abc_78290_new_n465_), .B(u5__abc_78290_new_n476_), .Y(u5__abc_78290_new_n477_));
NAND2X1 NAND2X1_1473 ( .A(u5__abc_78290_new_n489_), .B(u5__abc_78290_new_n490_), .Y(u5__abc_78290_new_n491_));
NAND2X1 NAND2X1_1474 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n496_), .Y(u5__abc_78290_new_n497_));
NAND2X1 NAND2X1_1475 ( .A(u5_state_25_), .B(u5__abc_78290_new_n500_), .Y(u5__abc_78290_new_n501_));
NAND2X1 NAND2X1_1476 ( .A(u5_state_26_), .B(u5__abc_78290_new_n506_), .Y(u5__abc_78290_new_n507_));
NAND2X1 NAND2X1_1477 ( .A(u5__abc_78290_new_n505_), .B(u5__abc_78290_new_n511_), .Y(u5__abc_78290_new_n512_));
NAND2X1 NAND2X1_1478 ( .A(u5__abc_78290_new_n515_), .B(u5__abc_78290_new_n404_), .Y(u5__abc_78290_new_n516_));
NAND2X1 NAND2X1_1479 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n520_), .Y(u5__abc_78290_new_n521_));
NAND2X1 NAND2X1_148 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1482_));
NAND2X1 NAND2X1_1480 ( .A(u5__abc_78290_new_n522_), .B(u5__abc_78290_new_n523_), .Y(u5__abc_78290_new_n524_));
NAND2X1 NAND2X1_1481 ( .A(u5__abc_78290_new_n467_), .B(u5__abc_78290_new_n403_), .Y(u5__abc_78290_new_n532_));
NAND2X1 NAND2X1_1482 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n535_), .Y(u5__abc_78290_new_n536_));
NAND2X1 NAND2X1_1483 ( .A(u5__abc_78290_new_n522_), .B(u5__abc_78290_new_n451_), .Y(u5__abc_78290_new_n537_));
NAND2X1 NAND2X1_1484 ( .A(u5__abc_78290_new_n538_), .B(u5__abc_78290_new_n431_), .Y(u5__abc_78290_new_n539_));
NAND2X1 NAND2X1_1485 ( .A(u5__abc_78290_new_n548_), .B(u5__abc_78290_new_n435_), .Y(u5__abc_78290_new_n549_));
NAND2X1 NAND2X1_1486 ( .A(u5__abc_78290_new_n473_), .B(u5__abc_78290_new_n499_), .Y(u5__abc_78290_new_n557_));
NAND2X1 NAND2X1_1487 ( .A(u5__abc_78290_new_n560_), .B(u5__abc_78290_new_n480_), .Y(u5__abc_78290_new_n561_));
NAND2X1 NAND2X1_1488 ( .A(u5_state_17_), .B(u5__abc_78290_new_n564_), .Y(u5__abc_78290_new_n565_));
NAND2X1 NAND2X1_1489 ( .A(u5__abc_78290_new_n479_), .B(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n570_));
NAND2X1 NAND2X1_149 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1485_));
NAND2X1 NAND2X1_1490 ( .A(u5__abc_78290_new_n425_), .B(u5__abc_78290_new_n575_), .Y(u5__abc_78290_new_n576_));
NAND2X1 NAND2X1_1491 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n584_), .Y(u5__abc_78290_new_n585_));
NAND2X1 NAND2X1_1492 ( .A(u5__abc_78290_new_n594_), .B(u5__abc_78290_new_n587_), .Y(u5__abc_78290_new_n595_));
NAND2X1 NAND2X1_1493 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n429_), .Y(u5__abc_78290_new_n601_));
NAND2X1 NAND2X1_1494 ( .A(u5__abc_78290_new_n600_), .B(u5__abc_78290_new_n607_), .Y(u5__abc_78290_new_n608_));
NAND2X1 NAND2X1_1495 ( .A(u5_state_51_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n613_));
NAND2X1 NAND2X1_1496 ( .A(u5__abc_78290_new_n614_), .B(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n615_));
NAND2X1 NAND2X1_1497 ( .A(u5_state_50_), .B(u5__abc_78290_new_n619_), .Y(u5__abc_78290_new_n620_));
NAND2X1 NAND2X1_1498 ( .A(u5__abc_78290_new_n634_), .B(u5__abc_78290_new_n388_), .Y(u5__abc_78290_new_n635_));
NAND2X1 NAND2X1_1499 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n638_), .Y(u5__abc_78290_new_n639_));
NAND2X1 NAND2X1_15 ( .A(init_req), .B(1'h0), .Y(u0__abc_74894_new_n1150_));
NAND2X1 NAND2X1_150 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1488_));
NAND2X1 NAND2X1_1500 ( .A(u5__abc_78290_new_n632_), .B(u5__abc_78290_new_n388_), .Y(u5__abc_78290_new_n650_));
NAND2X1 NAND2X1_1501 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n653_), .Y(u5__abc_78290_new_n654_));
NAND2X1 NAND2X1_1502 ( .A(u5__abc_78290_new_n655_), .B(u5__abc_78290_new_n398_), .Y(u5__abc_78290_new_n656_));
NAND2X1 NAND2X1_1503 ( .A(u5__abc_78290_new_n654_), .B(u5__abc_78290_new_n659_), .Y(u5__abc_78290_new_n660_));
NAND2X1 NAND2X1_1504 ( .A(u5__abc_78290_new_n662_), .B(u5__abc_78290_new_n405_), .Y(u5__abc_78290_new_n663_));
NAND2X1 NAND2X1_1505 ( .A(u5__abc_78290_new_n675_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n676_));
NAND2X1 NAND2X1_1506 ( .A(u5__abc_78290_new_n677_), .B(u5__abc_78290_new_n405_), .Y(u5__abc_78290_new_n678_));
NAND2X1 NAND2X1_1507 ( .A(u5__abc_78290_new_n680_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n681_));
NAND2X1 NAND2X1_1508 ( .A(u5__abc_78290_new_n588_), .B(u5__abc_78290_new_n562_), .Y(u5__abc_78290_new_n683_));
NAND2X1 NAND2X1_1509 ( .A(u5__abc_78290_new_n423_), .B(u5__abc_78290_new_n684_), .Y(u5__abc_78290_new_n685_));
NAND2X1 NAND2X1_151 ( .A(u0__abc_74894_new_n1476_), .B(u0__abc_74894_new_n1494_), .Y(u0__0sp_tms_31_0__16_));
NAND2X1 NAND2X1_1510 ( .A(u5__abc_78290_new_n686_), .B(u5__abc_78290_new_n398_), .Y(u5__abc_78290_new_n687_));
NAND2X1 NAND2X1_1511 ( .A(u5__abc_78290_new_n692_), .B(u5__abc_78290_new_n398_), .Y(u5__abc_78290_new_n693_));
NAND2X1 NAND2X1_1512 ( .A(u5__abc_78290_new_n695_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n696_));
NAND2X1 NAND2X1_1513 ( .A(u5__abc_78290_new_n698_), .B(u5__abc_78290_new_n405_), .Y(u5__abc_78290_new_n699_));
NAND2X1 NAND2X1_1514 ( .A(u5__abc_78290_new_n703_), .B(u5__abc_78290_new_n398_), .Y(u5__abc_78290_new_n704_));
NAND2X1 NAND2X1_1515 ( .A(u5__abc_78290_new_n706_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n707_));
NAND2X1 NAND2X1_1516 ( .A(u5_state_43_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n710_));
NAND2X1 NAND2X1_1517 ( .A(u5__abc_78290_new_n713_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n714_));
NAND2X1 NAND2X1_1518 ( .A(u5__abc_78290_new_n721_), .B(u5__abc_78290_new_n709_), .Y(u5__abc_78290_new_n722_));
NAND2X1 NAND2X1_1519 ( .A(u5_state_13_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n746_));
NAND2X1 NAND2X1_152 ( .A(sp_tms_17_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1496_));
NAND2X1 NAND2X1_1520 ( .A(u5__abc_78290_new_n747_), .B(u5__abc_78290_new_n414_), .Y(u5__abc_78290_new_n748_));
NAND2X1 NAND2X1_1521 ( .A(u5__abc_78290_new_n492_), .B(u5__abc_78290_new_n413_), .Y(u5__abc_78290_new_n754_));
NAND2X1 NAND2X1_1522 ( .A(u5__abc_78290_new_n761_), .B(u5__abc_78290_new_n684_), .Y(u5__abc_78290_new_n762_));
NAND2X1 NAND2X1_1523 ( .A(u5__abc_78290_new_n763_), .B(u5__abc_78290_new_n414_), .Y(u5__abc_78290_new_n764_));
NAND2X1 NAND2X1_1524 ( .A(u5__abc_78290_new_n416_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n770_));
NAND2X1 NAND2X1_1525 ( .A(u5__abc_78290_new_n777_), .B(u5__abc_78290_new_n421_), .Y(u5__abc_78290_new_n778_));
NAND2X1 NAND2X1_1526 ( .A(u5__abc_78290_new_n784_), .B(u5__abc_78290_new_n769_), .Y(u5__abc_78290_new_n785_));
NAND2X1 NAND2X1_1527 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n791_), .Y(u5__abc_78290_new_n792_));
NAND2X1 NAND2X1_1528 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n797_), .Y(u5__abc_78290_new_n798_));
NAND2X1 NAND2X1_1529 ( .A(u5__abc_78290_new_n792_), .B(u5__abc_78290_new_n798_), .Y(u5__abc_78290_new_n799_));
NAND2X1 NAND2X1_153 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1497_), .Y(u0__abc_74894_new_n1498_));
NAND2X1 NAND2X1_1530 ( .A(u5_state_34_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n805_));
NAND2X1 NAND2X1_1531 ( .A(u5__abc_78290_new_n530_), .B(u5__abc_78290_new_n403_), .Y(u5__abc_78290_new_n812_));
NAND2X1 NAND2X1_1532 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n815_), .Y(u5__abc_78290_new_n816_));
NAND2X1 NAND2X1_1533 ( .A(u5_state_21_), .B(u5__abc_78290_new_n603_), .Y(u5__abc_78290_new_n817_));
NAND2X1 NAND2X1_1534 ( .A(u5__abc_78290_new_n818_), .B(u5__abc_78290_new_n453_), .Y(u5__abc_78290_new_n819_));
NAND2X1 NAND2X1_1535 ( .A(u5_state_61_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n850_));
NAND2X1 NAND2X1_1536 ( .A(u5_state_60_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n857_));
NAND2X1 NAND2X1_1537 ( .A(u5__abc_78290_new_n418_), .B(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n872_));
NAND2X1 NAND2X1_1538 ( .A(u5_state_63_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n878_));
NAND2X1 NAND2X1_1539 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n881_), .Y(u5__abc_78290_new_n882_));
NAND2X1 NAND2X1_154 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1499_), .Y(u0__abc_74894_new_n1500_));
NAND2X1 NAND2X1_1540 ( .A(u5__abc_78290_new_n877_), .B(u5__abc_78290_new_n882_), .Y(u5__abc_78290_new_n883_));
NAND2X1 NAND2X1_1541 ( .A(u5__abc_78290_new_n898_), .B(u5__abc_78290_new_n405_), .Y(u5__abc_78290_new_n899_));
NAND2X1 NAND2X1_1542 ( .A(u5__abc_78290_new_n904_), .B(u5__abc_78290_new_n382_), .Y(u5__abc_78290_new_n905_));
NAND2X1 NAND2X1_1543 ( .A(u5__abc_78290_new_n911_), .B(u5__abc_78290_new_n381_), .Y(u5__abc_78290_new_n912_));
NAND2X1 NAND2X1_1544 ( .A(u5__abc_78290_new_n902_), .B(u5__abc_78290_new_n382_), .Y(u5__abc_78290_new_n918_));
NAND2X1 NAND2X1_1545 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n921_), .Y(u5__abc_78290_new_n922_));
NAND2X1 NAND2X1_1546 ( .A(u5__abc_78290_new_n909_), .B(u5__abc_78290_new_n381_), .Y(u5__abc_78290_new_n925_));
NAND2X1 NAND2X1_1547 ( .A(u5_state_55_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n933_));
NAND2X1 NAND2X1_1548 ( .A(u5_state_52_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n942_));
NAND2X1 NAND2X1_1549 ( .A(u5_state_53_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n949_));
NAND2X1 NAND2X1_155 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1501_));
NAND2X1 NAND2X1_1550 ( .A(u5__abc_78290_new_n937_), .B(u5__abc_78290_new_n953_), .Y(u5__abc_78290_new_n954_));
NAND2X1 NAND2X1_1551 ( .A(u5__abc_78290_new_n962_), .B(u5__abc_78290_new_n963_), .Y(u5__abc_78290_new_n964_));
NAND2X1 NAND2X1_1552 ( .A(u5__abc_78290_new_n969_), .B(u5__abc_78290_new_n970_), .Y(u5__abc_78290_new_n971_));
NAND2X1 NAND2X1_1553 ( .A(u5_state_54_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n979_));
NAND2X1 NAND2X1_1554 ( .A(u5__abc_78290_new_n983_), .B(u5__abc_78290_new_n975_), .Y(u5__abc_78290_new_n984_));
NAND2X1 NAND2X1_1555 ( .A(u5__abc_78290_new_n1000_), .B(u5__abc_78290_new_n999_), .Y(u5__abc_78290_new_n1001_));
NAND2X1 NAND2X1_1556 ( .A(u5__abc_78290_new_n547_), .B(u5__abc_78290_new_n569_), .Y(u5__abc_78290_new_n1009_));
NAND2X1 NAND2X1_1557 ( .A(u5__abc_78290_new_n997_), .B(u5__abc_78290_new_n1018_), .Y(u5__abc_78290_new_n1019_));
NAND2X1 NAND2X1_1558 ( .A(u5__abc_78290_new_n1027_), .B(u5__abc_78290_new_n1023_), .Y(u5__abc_78290_new_n1028_));
NAND2X1 NAND2X1_1559 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1030_), .Y(u5__abc_78290_new_n1031_));
NAND2X1 NAND2X1_156 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1502_));
NAND2X1 NAND2X1_1560 ( .A(u5__abc_78290_new_n1034_), .B(u5__abc_78290_new_n1031_), .Y(u5__abc_78290_new_n1035_));
NAND2X1 NAND2X1_1561 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1038_));
NAND2X1 NAND2X1_1562 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1046_), .Y(u5__abc_78290_new_n1047_));
NAND2X1 NAND2X1_1563 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1049_), .Y(u5__abc_78290_new_n1050_));
NAND2X1 NAND2X1_1564 ( .A(u5__abc_78290_new_n684_), .B(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n1053_));
NAND2X1 NAND2X1_1565 ( .A(u5__abc_78290_new_n420_), .B(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1054_));
NAND2X1 NAND2X1_1566 ( .A(u5__abc_78290_new_n1052_), .B(u5__abc_78290_new_n1062_), .Y(u5__abc_78290_new_n1063_));
NAND2X1 NAND2X1_1567 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n1069_), .Y(u5__abc_78290_new_n1070_));
NAND2X1 NAND2X1_1568 ( .A(u5__abc_78290_new_n1070_), .B(u5__abc_78290_new_n877_), .Y(u5__abc_78290_new_n1071_));
NAND2X1 NAND2X1_1569 ( .A(u5__abc_78290_new_n380_), .B(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1073_));
NAND2X1 NAND2X1_157 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1505_));
NAND2X1 NAND2X1_1570 ( .A(u5__abc_78290_new_n1077_), .B(u5__abc_78290_new_n1074_), .Y(u5__abc_78290_new_n1078_));
NAND2X1 NAND2X1_1571 ( .A(u5__abc_78290_new_n1083_), .B(u5__abc_78290_new_n1078_), .Y(u5__abc_78290_new_n1084_));
NAND2X1 NAND2X1_1572 ( .A(u5__abc_78290_new_n1088_), .B(u5__abc_78290_new_n1085_), .Y(u5__abc_78290_new_n1089_));
NAND2X1 NAND2X1_1573 ( .A(u5__abc_78290_new_n1092_), .B(u5__abc_78290_new_n1085_), .Y(u5__abc_78290_new_n1093_));
NAND2X1 NAND2X1_1574 ( .A(u5__abc_78290_new_n1089_), .B(u5__abc_78290_new_n1093_), .Y(u5__abc_78290_new_n1094_));
NAND2X1 NAND2X1_1575 ( .A(u5__abc_78290_new_n1096_), .B(u5__abc_78290_new_n1098_), .Y(u5__abc_78290_new_n1099_));
NAND2X1 NAND2X1_1576 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n1103_), .Y(u5__abc_78290_new_n1104_));
NAND2X1 NAND2X1_1577 ( .A(u5__abc_78290_new_n1108_), .B(u5__abc_78290_new_n1074_), .Y(u5__abc_78290_new_n1109_));
NAND2X1 NAND2X1_1578 ( .A(u5__abc_78290_new_n1112_), .B(u5__abc_78290_new_n1085_), .Y(u5__abc_78290_new_n1113_));
NAND2X1 NAND2X1_1579 ( .A(u5__abc_78290_new_n1113_), .B(u5__abc_78290_new_n1109_), .Y(u5__abc_78290_new_n1114_));
NAND2X1 NAND2X1_158 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1508_));
NAND2X1 NAND2X1_1580 ( .A(u5__abc_78290_new_n1115_), .B(u5__abc_78290_new_n1095_), .Y(u5__abc_78290_new_n1116_));
NAND2X1 NAND2X1_1581 ( .A(u5__abc_78290_new_n1119_), .B(u5__abc_78290_new_n661_), .Y(u5__abc_78290_new_n1120_));
NAND2X1 NAND2X1_1582 ( .A(u5__abc_78290_new_n1122_), .B(u5__abc_78290_new_n661_), .Y(u5__abc_78290_new_n1123_));
NAND2X1 NAND2X1_1583 ( .A(u5__abc_78290_new_n1126_), .B(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n1127_));
NAND2X1 NAND2X1_1584 ( .A(u5__abc_78290_new_n1130_), .B(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n1131_));
NAND2X1 NAND2X1_1585 ( .A(u5__abc_78290_new_n387_), .B(u5__abc_78290_new_n616_), .Y(u5__abc_78290_new_n1135_));
NAND2X1 NAND2X1_1586 ( .A(u5__abc_78290_new_n387_), .B(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1138_));
NAND2X1 NAND2X1_1587 ( .A(u5__abc_78290_new_n1137_), .B(u5__abc_78290_new_n1146_), .Y(u5__abc_78290_new_n1147_));
NAND2X1 NAND2X1_1588 ( .A(u5__abc_78290_new_n1148_), .B(u5__abc_78290_new_n1133_), .Y(u5__abc_78290_new_n1149_));
NAND2X1 NAND2X1_1589 ( .A(u5__abc_78290_new_n1151_), .B(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n1152_));
NAND2X1 NAND2X1_159 ( .A(u0__abc_74894_new_n1496_), .B(u0__abc_74894_new_n1514_), .Y(u0__0sp_tms_31_0__17_));
NAND2X1 NAND2X1_1590 ( .A(u5__abc_78290_new_n1154_), .B(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n1155_));
NAND2X1 NAND2X1_1591 ( .A(u5__abc_78290_new_n1159_), .B(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n1160_));
NAND2X1 NAND2X1_1592 ( .A(u5__abc_78290_new_n1163_), .B(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n1164_));
NAND2X1 NAND2X1_1593 ( .A(u5__abc_78290_new_n397_), .B(u5__abc_78290_new_n1168_), .Y(u5__abc_78290_new_n1169_));
NAND2X1 NAND2X1_1594 ( .A(u5__abc_78290_new_n1170_), .B(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n1171_));
NAND2X1 NAND2X1_1595 ( .A(u5__abc_78290_new_n1173_), .B(u5__abc_78290_new_n642_), .Y(u5__abc_78290_new_n1174_));
NAND2X1 NAND2X1_1596 ( .A(u5__abc_78290_new_n1177_), .B(u5__abc_78290_new_n661_), .Y(u5__abc_78290_new_n1178_));
NAND2X1 NAND2X1_1597 ( .A(u5__abc_78290_new_n1180_), .B(u5__abc_78290_new_n661_), .Y(u5__abc_78290_new_n1181_));
NAND2X1 NAND2X1_1598 ( .A(u5__abc_78290_new_n1183_), .B(u5__abc_78290_new_n1167_), .Y(u5__abc_78290_new_n1184_));
NAND2X1 NAND2X1_1599 ( .A(u5__abc_78290_new_n1192_), .B(u5__abc_78290_new_n1188_), .Y(u5__abc_78290_new_n1193_));
NAND2X1 NAND2X1_16 ( .A(sp_tms_0_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1156_));
NAND2X1 NAND2X1_160 ( .A(sp_tms_18_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1516_));
NAND2X1 NAND2X1_1600 ( .A(u5__abc_78290_new_n1195_), .B(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n1196_));
NAND2X1 NAND2X1_1601 ( .A(u5__abc_78290_new_n1198_), .B(u5__abc_78290_new_n1188_), .Y(u5__abc_78290_new_n1199_));
NAND2X1 NAND2X1_1602 ( .A(u5__abc_78290_new_n1203_), .B(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n1204_));
NAND2X1 NAND2X1_1603 ( .A(u5__abc_78290_new_n499_), .B(u5__abc_78290_new_n584_), .Y(u5__abc_78290_new_n1205_));
NAND2X1 NAND2X1_1604 ( .A(u5__abc_78290_new_n1206_), .B(u5__abc_78290_new_n1188_), .Y(u5__abc_78290_new_n1207_));
NAND2X1 NAND2X1_1605 ( .A(u5__abc_78290_new_n1193_), .B(u5__abc_78290_new_n1209_), .Y(u5__abc_78290_new_n1210_));
NAND2X1 NAND2X1_1606 ( .A(u5__abc_78290_new_n472_), .B(u5__abc_78290_new_n1215_), .Y(u5__abc_78290_new_n1216_));
NAND2X1 NAND2X1_1607 ( .A(u5__abc_78290_new_n1218_), .B(u5__abc_78290_new_n661_), .Y(u5__abc_78290_new_n1219_));
NAND2X1 NAND2X1_1608 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1221_), .Y(u5__abc_78290_new_n1222_));
NAND2X1 NAND2X1_1609 ( .A(u5__abc_78290_new_n409_), .B(u5__abc_78290_new_n414_), .Y(u5__abc_78290_new_n1224_));
NAND2X1 NAND2X1_161 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1517_), .Y(u0__abc_74894_new_n1518_));
NAND2X1 NAND2X1_1610 ( .A(u5_state_12_), .B(u5__abc_78290_new_n823_), .Y(u5__abc_78290_new_n1226_));
NAND2X1 NAND2X1_1611 ( .A(u5__abc_78290_new_n447_), .B(u5__abc_78290_new_n1232_), .Y(u5__abc_78290_new_n1233_));
NAND2X1 NAND2X1_1612 ( .A(u5__abc_78290_new_n1237_), .B(u5__abc_78290_new_n661_), .Y(u5__abc_78290_new_n1238_));
NAND2X1 NAND2X1_1613 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n1247_), .Y(u5__abc_78290_new_n1248_));
NAND2X1 NAND2X1_1614 ( .A(u5__abc_78290_new_n1250_), .B(u5__abc_78290_new_n1240_), .Y(u5__abc_78290_new_n1251_));
NAND2X1 NAND2X1_1615 ( .A(u5_state_13_), .B(u5__abc_78290_new_n747_), .Y(u5__abc_78290_new_n1254_));
NAND2X1 NAND2X1_1616 ( .A(u5__abc_78290_new_n411_), .B(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n1258_));
NAND2X1 NAND2X1_1617 ( .A(u5__abc_78290_new_n447_), .B(u5__abc_78290_new_n1271_), .Y(u5__abc_78290_new_n1272_));
NAND2X1 NAND2X1_1618 ( .A(u5__abc_78290_new_n1263_), .B(u5__abc_78290_new_n1274_), .Y(u5__abc_78290_new_n1275_));
NAND2X1 NAND2X1_1619 ( .A(u5__abc_78290_new_n1281_), .B(u5__abc_78290_new_n1278_), .Y(u5__abc_78290_new_n1282_));
NAND2X1 NAND2X1_162 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1519_), .Y(u0__abc_74894_new_n1520_));
NAND2X1 NAND2X1_1620 ( .A(u5__abc_78290_new_n417_), .B(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n1284_));
NAND2X1 NAND2X1_1621 ( .A(u5__abc_78290_new_n1290_), .B(u5__abc_78290_new_n1278_), .Y(u5__abc_78290_new_n1291_));
NAND2X1 NAND2X1_1622 ( .A(u5__abc_78290_new_n1296_), .B(u5__abc_78290_new_n1278_), .Y(u5__abc_78290_new_n1297_));
NAND2X1 NAND2X1_1623 ( .A(u5__abc_78290_new_n444_), .B(u5__abc_78290_new_n1298_), .Y(u5__abc_78290_new_n1299_));
NAND2X1 NAND2X1_1624 ( .A(u5__abc_78290_new_n545_), .B(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n1302_));
NAND2X1 NAND2X1_1625 ( .A(u5__abc_78290_new_n419_), .B(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n1307_));
NAND2X1 NAND2X1_1626 ( .A(u5__abc_78290_new_n1253_), .B(u5__abc_78290_new_n1314_), .Y(u5__abc_78290_new_n1315_));
NAND2X1 NAND2X1_1627 ( .A(u5__abc_78290_new_n1187_), .B(u5__abc_78290_new_n1316_), .Y(u5__abc_78290_new_n1317_));
NAND2X1 NAND2X1_1628 ( .A(u5__abc_78290_new_n1325_), .B(u5__abc_78290_new_n1323_), .Y(u5__abc_78290_new_n1326_));
NAND2X1 NAND2X1_1629 ( .A(u5__abc_78290_new_n1334_), .B(u5__abc_78290_new_n1332_), .Y(u5__abc_78290_new_n1335_));
NAND2X1 NAND2X1_163 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1521_));
NAND2X1 NAND2X1_1630 ( .A(u5__abc_78290_new_n1343_), .B(u5__abc_78290_new_n1342_), .Y(u5__abc_78290_new_n1344_));
NAND2X1 NAND2X1_1631 ( .A(u5__abc_78290_new_n1350_), .B(u5__abc_78290_new_n1349_), .Y(u5__abc_78290_new_n1351_));
NAND2X1 NAND2X1_1632 ( .A(u5__abc_78290_new_n1361_), .B(u5__abc_78290_new_n1362_), .Y(u5__abc_78290_new_n1363_));
NAND2X1 NAND2X1_1633 ( .A(u5__abc_78290_new_n1382_), .B(u5__abc_78290_new_n1384_), .Y(u5__abc_78290_new_n1385_));
NAND2X1 NAND2X1_1634 ( .A(u5__abc_78290_new_n1392_), .B(u5__abc_78290_new_n1361_), .Y(u5__abc_78290_new_n1393_));
NAND2X1 NAND2X1_1635 ( .A(u5__abc_78290_new_n1397_), .B(u5__abc_78290_new_n1390_), .Y(u5__abc_78290_new_n1398_));
NAND2X1 NAND2X1_1636 ( .A(u5__abc_78290_new_n1142_), .B(u5__abc_78290_new_n1139_), .Y(u5__abc_78290_new_n1400_));
NAND2X1 NAND2X1_1637 ( .A(u5__abc_78290_new_n1411_), .B(u5__0burst_act_rd_0_0_), .Y(u5__abc_78290_new_n1412_));
NAND2X1 NAND2X1_1638 ( .A(u5__abc_78290_new_n1207_), .B(u5__abc_78290_new_n1306_), .Y(u5__abc_78290_new_n1423_));
NAND2X1 NAND2X1_1639 ( .A(u5__abc_78290_new_n1424_), .B(u5__abc_78290_new_n1421_), .Y(u5__abc_78290_new_n1425_));
NAND2X1 NAND2X1_164 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1522_));
NAND2X1 NAND2X1_1640 ( .A(u5__abc_78290_new_n1429_), .B(u5_cmd_0_), .Y(u5__abc_78290_new_n1430_));
NAND2X1 NAND2X1_1641 ( .A(u5__abc_78290_new_n1242_), .B(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n1436_));
NAND2X1 NAND2X1_1642 ( .A(u5__abc_78290_new_n1145_), .B(u5__abc_78290_new_n1139_), .Y(u5__abc_78290_new_n1441_));
NAND2X1 NAND2X1_1643 ( .A(u5__abc_78290_new_n1070_), .B(u5__abc_78290_new_n1104_), .Y(u5__abc_78290_new_n1443_));
NAND2X1 NAND2X1_1644 ( .A(u5__abc_78290_new_n1473_), .B(u5__abc_78290_new_n1474_), .Y(u5__abc_78290_new_n1475_));
NAND2X1 NAND2X1_1645 ( .A(u5__abc_78290_new_n1345_), .B(u5__abc_78290_new_n1478_), .Y(u5__abc_78290_new_n1479_));
NAND2X1 NAND2X1_1646 ( .A(csc_s_1_), .B(u5__abc_78290_new_n1320_), .Y(u5__abc_78290_new_n1480_));
NAND2X1 NAND2X1_1647 ( .A(u5__abc_78290_new_n1320_), .B(u5__abc_78290_new_n1484_), .Y(u5__abc_78290_new_n1485_));
NAND2X1 NAND2X1_1648 ( .A(u5__abc_78290_new_n1487_), .B(u5__abc_78290_new_n1488_), .Y(u5__abc_78290_new_n1489_));
NAND2X1 NAND2X1_1649 ( .A(u5__abc_78290_new_n1189_), .B(u5__abc_78290_new_n1188_), .Y(u5__abc_78290_new_n1491_));
NAND2X1 NAND2X1_165 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1525_));
NAND2X1 NAND2X1_1650 ( .A(u5__abc_78290_new_n1134_), .B(u5__abc_78290_new_n1085_), .Y(u5__abc_78290_new_n1495_));
NAND2X1 NAND2X1_1651 ( .A(u1_wr_cycle), .B(u5_cmd_del_3_), .Y(u5__abc_78290_new_n1510_));
NAND2X1 NAND2X1_1652 ( .A(u5__abc_78290_new_n1429_), .B(u5_data_oe_d), .Y(u5__abc_78290_new_n1523_));
NAND2X1 NAND2X1_1653 ( .A(u5__abc_78290_new_n1215_), .B(u5__abc_78290_new_n1533_), .Y(u5__abc_78290_new_n1534_));
NAND2X1 NAND2X1_1654 ( .A(u5__abc_78290_new_n1204_), .B(u5__abc_78290_new_n1363_), .Y(u5__abc_78290_new_n1535_));
NAND2X1 NAND2X1_1655 ( .A(u5__abc_78290_new_n1207_), .B(u5__abc_78290_new_n1196_), .Y(u5__abc_78290_new_n1536_));
NAND2X1 NAND2X1_1656 ( .A(u5__abc_78290_new_n1558_), .B(u5__abc_78290_new_n1561_), .Y(u5__abc_78290_new_n1562_));
NAND2X1 NAND2X1_1657 ( .A(u5__abc_78290_new_n1550_), .B(u5__abc_78290_new_n1565_), .Y(u5__abc_78290_new_n1566_));
NAND2X1 NAND2X1_1658 ( .A(u5__abc_78290_new_n472_), .B(u5__abc_78290_new_n1579_), .Y(u5__abc_78290_new_n1580_));
NAND2X1 NAND2X1_1659 ( .A(u5__abc_78290_new_n1581_), .B(u5__abc_78290_new_n1582_), .Y(u5__abc_78290_new_n1583_));
NAND2X1 NAND2X1_166 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1528_));
NAND2X1 NAND2X1_1660 ( .A(u5__abc_78290_new_n1325_), .B(u5__abc_78290_new_n1481_), .Y(u5__abc_78290_new_n1606_));
NAND2X1 NAND2X1_1661 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n1610_), .Y(u5__abc_78290_new_n1612_));
NAND2X1 NAND2X1_1662 ( .A(u5__abc_78290_new_n1048_), .B(u5__abc_78290_new_n1045_), .Y(u5__abc_78290_new_n1615_));
NAND2X1 NAND2X1_1663 ( .A(u5__abc_78290_new_n1039_), .B(u5__abc_78290_new_n1359_), .Y(u5__abc_78290_new_n1618_));
NAND2X1 NAND2X1_1664 ( .A(u1_wb_write_go), .B(u5_tmr_done), .Y(u5__abc_78290_new_n1620_));
NAND2X1 NAND2X1_1665 ( .A(u5__abc_78290_new_n1072_), .B(u5__abc_78290_new_n1641_), .Y(u5__abc_78290_new_n1642_));
NAND2X1 NAND2X1_1666 ( .A(u5__abc_78290_new_n1390_), .B(u5__abc_78290_new_n1645_), .Y(u5__abc_78290_new_n1646_));
NAND2X1 NAND2X1_1667 ( .A(u5__abc_78290_new_n1647_), .B(u5__abc_78290_new_n1567_), .Y(u5__abc_78290_new_n1648_));
NAND2X1 NAND2X1_1668 ( .A(u5__abc_78290_new_n1650_), .B(u5__abc_78290_new_n1632_), .Y(u5__abc_78290_new_n1655_));
NAND2X1 NAND2X1_1669 ( .A(tms_s_0_), .B(u5__abc_78290_new_n1656_), .Y(u5__abc_78290_new_n1657_));
NAND2X1 NAND2X1_167 ( .A(u0__abc_74894_new_n1516_), .B(u0__abc_74894_new_n1534_), .Y(u0__0sp_tms_31_0__18_));
NAND2X1 NAND2X1_1670 ( .A(u5__abc_78290_new_n1429_), .B(dv), .Y(u5__abc_78290_new_n1664_));
NAND2X1 NAND2X1_1671 ( .A(u5_burst_cnt_0_), .B(u5__abc_78290_new_n1666_), .Y(u5__abc_78290_new_n1668_));
NAND2X1 NAND2X1_1672 ( .A(u5__abc_78290_new_n1664_), .B(u5__abc_78290_new_n1665_), .Y(u5__abc_78290_new_n1673_));
NAND2X1 NAND2X1_1673 ( .A(u5__abc_78290_new_n1656_), .B(u5__abc_78290_new_n1632_), .Y(u5__abc_78290_new_n1687_));
NAND2X1 NAND2X1_1674 ( .A(1'h0), .B(u5__abc_78290_new_n1675_), .Y(u5__abc_78290_new_n1688_));
NAND2X1 NAND2X1_1675 ( .A(u5__abc_78290_new_n465_), .B(u5__abc_78290_new_n1714_), .Y(u5__abc_78290_new_n1715_));
NAND2X1 NAND2X1_1676 ( .A(u5__abc_78290_new_n1250_), .B(u5__abc_78290_new_n1723_), .Y(u5__abc_78290_new_n1724_));
NAND2X1 NAND2X1_1677 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n1203_), .Y(u5__abc_78290_new_n1726_));
NAND2X1 NAND2X1_1678 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1727_), .Y(u5__abc_78290_new_n1728_));
NAND2X1 NAND2X1_1679 ( .A(u5__abc_78290_new_n1732_), .B(u5__abc_78290_new_n1742_), .Y(u5__abc_78290_new_n1743_));
NAND2X1 NAND2X1_168 ( .A(sp_tms_19_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1536_));
NAND2X1 NAND2X1_1680 ( .A(u5__abc_78290_new_n427_), .B(u5__abc_78290_new_n597_), .Y(u5__abc_78290_new_n1744_));
NAND2X1 NAND2X1_1681 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1750_), .Y(u5__abc_78290_new_n1751_));
NAND2X1 NAND2X1_1682 ( .A(u5__abc_78290_new_n1760_), .B(u5__abc_78290_new_n1753_), .Y(u5__abc_78290_new_n1761_));
NAND2X1 NAND2X1_1683 ( .A(u5__abc_78290_new_n1765_), .B(u5__abc_78290_new_n1767_), .Y(u5__abc_78290_new_n1768_));
NAND2X1 NAND2X1_1684 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1768_), .Y(u5__abc_78290_new_n1769_));
NAND2X1 NAND2X1_1685 ( .A(u5__abc_78290_new_n1775_), .B(u5__abc_78290_new_n1771_), .Y(u5__abc_78290_new_n1776_));
NAND2X1 NAND2X1_1686 ( .A(u5__abc_78290_new_n447_), .B(u5__abc_78290_new_n1778_), .Y(u5__abc_78290_new_n1779_));
NAND2X1 NAND2X1_1687 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1780_), .Y(u5__abc_78290_new_n1781_));
NAND2X1 NAND2X1_1688 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1784_), .Y(u5__abc_78290_new_n1785_));
NAND2X1 NAND2X1_1689 ( .A(u5__abc_78290_new_n1781_), .B(u5__abc_78290_new_n1785_), .Y(u5__abc_78290_new_n1786_));
NAND2X1 NAND2X1_169 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1537_), .Y(u0__abc_74894_new_n1538_));
NAND2X1 NAND2X1_1690 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1799_), .Y(u5__abc_78290_new_n1800_));
NAND2X1 NAND2X1_1691 ( .A(u5__abc_78290_new_n1800_), .B(u5__abc_78290_new_n497_), .Y(u5__abc_78290_new_n1801_));
NAND2X1 NAND2X1_1692 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1801_), .Y(u5__abc_78290_new_n1802_));
NAND2X1 NAND2X1_1693 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1805_), .Y(u5__abc_78290_new_n1806_));
NAND2X1 NAND2X1_1694 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1809_), .Y(u5__abc_78290_new_n1810_));
NAND2X1 NAND2X1_1695 ( .A(u5__abc_78290_new_n1806_), .B(u5__abc_78290_new_n1810_), .Y(u5__abc_78290_new_n1811_));
NAND2X1 NAND2X1_1696 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1811_), .Y(u5__abc_78290_new_n1812_));
NAND2X1 NAND2X1_1697 ( .A(u5__abc_78290_new_n447_), .B(u5__abc_78290_new_n1814_), .Y(u5__abc_78290_new_n1815_));
NAND2X1 NAND2X1_1698 ( .A(u5__abc_78290_new_n478_), .B(u5__abc_78290_new_n1827_), .Y(u5__abc_78290_new_n1828_));
NAND2X1 NAND2X1_1699 ( .A(u5__abc_78290_new_n458_), .B(u5__abc_78290_new_n1835_), .Y(u5__abc_78290_new_n1836_));
NAND2X1 NAND2X1_17 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1157_), .Y(u0__abc_74894_new_n1158_));
NAND2X1 NAND2X1_170 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1539_), .Y(u0__abc_74894_new_n1540_));
NAND2X1 NAND2X1_1700 ( .A(u5__abc_78290_new_n388_), .B(u5__abc_78290_new_n1143_), .Y(u5__abc_78290_new_n1848_));
NAND2X1 NAND2X1_1701 ( .A(u5__abc_78290_new_n1843_), .B(u5__abc_78290_new_n1852_), .Y(u5__abc_78290_new_n1853_));
NAND2X1 NAND2X1_1702 ( .A(u5__abc_78290_new_n476_), .B(u5__abc_78290_new_n1130_), .Y(u5__abc_78290_new_n1854_));
NAND2X1 NAND2X1_1703 ( .A(u5__abc_78290_new_n465_), .B(u5__abc_78290_new_n1122_), .Y(u5__abc_78290_new_n1863_));
NAND2X1 NAND2X1_1704 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1869_), .Y(u5__abc_78290_new_n1870_));
NAND2X1 NAND2X1_1705 ( .A(u5__abc_78290_new_n476_), .B(u5__abc_78290_new_n1154_), .Y(u5__abc_78290_new_n1873_));
NAND2X1 NAND2X1_1706 ( .A(u5__abc_78290_new_n1876_), .B(u5__abc_78290_new_n1870_), .Y(u5__abc_78290_new_n1877_));
NAND2X1 NAND2X1_1707 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1880_), .Y(u5__abc_78290_new_n1881_));
NAND2X1 NAND2X1_1708 ( .A(u5__abc_78290_new_n465_), .B(u5__abc_78290_new_n1180_), .Y(u5__abc_78290_new_n1884_));
NAND2X1 NAND2X1_1709 ( .A(u5__abc_78290_new_n1881_), .B(u5__abc_78290_new_n1887_), .Y(u5__abc_78290_new_n1888_));
NAND2X1 NAND2X1_171 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1541_));
NAND2X1 NAND2X1_1710 ( .A(u5__abc_78290_new_n378_), .B(u5__abc_78290_new_n1049_), .Y(u5__abc_78290_new_n1897_));
NAND2X1 NAND2X1_1711 ( .A(u5__abc_78290_new_n378_), .B(u5__abc_78290_new_n1046_), .Y(u5__abc_78290_new_n1900_));
NAND2X1 NAND2X1_1712 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1903_), .Y(u5__abc_78290_new_n1904_));
NAND2X1 NAND2X1_1713 ( .A(u5__abc_78290_new_n420_), .B(u5__abc_78290_new_n1059_), .Y(u5__abc_78290_new_n1905_));
NAND2X1 NAND2X1_1714 ( .A(u5__abc_78290_new_n385_), .B(u5__abc_78290_new_n1090_), .Y(u5__abc_78290_new_n1916_));
NAND2X1 NAND2X1_1715 ( .A(u5__abc_78290_new_n385_), .B(u5__abc_78290_new_n1086_), .Y(u5__abc_78290_new_n1919_));
NAND2X1 NAND2X1_1716 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1922_), .Y(u5__abc_78290_new_n1923_));
NAND2X1 NAND2X1_1717 ( .A(u5__abc_78290_new_n381_), .B(u5__abc_78290_new_n1075_), .Y(u5__abc_78290_new_n1934_));
NAND2X1 NAND2X1_1718 ( .A(u5__abc_78290_new_n386_), .B(u5__abc_78290_new_n1080_), .Y(u5__abc_78290_new_n1939_));
NAND2X1 NAND2X1_1719 ( .A(u5__abc_78290_new_n369_), .B(u5__abc_78290_new_n1673_), .Y(u5__abc_78290_new_n1959_));
NAND2X1 NAND2X1_172 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1542_));
NAND2X1 NAND2X1_1720 ( .A(u5__abc_78290_new_n1961_), .B(u5__abc_78290_new_n1968_), .Y(u5__abc_78290_new_n1969_));
NAND2X1 NAND2X1_1721 ( .A(u5__abc_78290_new_n374_), .B(u5__abc_78290_new_n1968_), .Y(u5__abc_78290_new_n1975_));
NAND2X1 NAND2X1_1722 ( .A(u5__abc_78290_new_n373_), .B(u5__abc_78290_new_n1666_), .Y(u5__abc_78290_new_n1977_));
NAND2X1 NAND2X1_1723 ( .A(u5__abc_78290_new_n1190_), .B(u5__abc_78290_new_n1986_), .Y(u5__abc_78290_new_n1987_));
NAND2X1 NAND2X1_1724 ( .A(u5__abc_78290_new_n1196_), .B(u5__abc_78290_new_n1581_), .Y(u5__abc_78290_new_n1989_));
NAND2X1 NAND2X1_1725 ( .A(u5__abc_78290_new_n1199_), .B(u5__abc_78290_new_n1992_), .Y(u5__abc_78290_new_n1993_));
NAND2X1 NAND2X1_1726 ( .A(u5__abc_78290_new_n1240_), .B(u5__abc_78290_new_n1996_), .Y(u5__abc_78290_new_n1997_));
NAND2X1 NAND2X1_1727 ( .A(u5__abc_78290_new_n969_), .B(u5__abc_78290_new_n2002_), .Y(u5__abc_78290_new_n2003_));
NAND2X1 NAND2X1_1728 ( .A(u5__abc_78290_new_n1538_), .B(u5__abc_78290_new_n1187_), .Y(u5__abc_78290_new_n2005_));
NAND2X1 NAND2X1_1729 ( .A(u5__abc_78290_new_n2009_), .B(u5__abc_78290_new_n2006_), .Y(u5__abc_78290_new_n2010_));
NAND2X1 NAND2X1_173 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1545_));
NAND2X1 NAND2X1_1730 ( .A(u5__abc_78290_new_n2010_), .B(u5__abc_78290_new_n2020_), .Y(u5__abc_78290_new_n2021_));
NAND2X1 NAND2X1_1731 ( .A(u5__abc_78290_new_n1187_), .B(u5__abc_78290_new_n2031_), .Y(u5__abc_78290_new_n2032_));
NAND2X1 NAND2X1_1732 ( .A(u5__abc_78290_new_n1440_), .B(u5__abc_78290_new_n2032_), .Y(u5__abc_78290_new_n2033_));
NAND2X1 NAND2X1_1733 ( .A(u5__abc_78290_new_n1550_), .B(u5__abc_78290_new_n2038_), .Y(u5__abc_78290_new_n2039_));
NAND2X1 NAND2X1_1734 ( .A(u5__abc_78290_new_n2041_), .B(u5__abc_78290_new_n2045_), .Y(u5__abc_78290_new_n2046_));
NAND2X1 NAND2X1_1735 ( .A(u5__abc_78290_new_n2053_), .B(u5__abc_78290_new_n2051_), .Y(u5__abc_78290_new_n2054_));
NAND2X1 NAND2X1_1736 ( .A(u5__abc_78290_new_n594_), .B(u5__abc_78290_new_n607_), .Y(u5__abc_78290_new_n2062_));
NAND2X1 NAND2X1_1737 ( .A(u5__abc_78290_new_n1214_), .B(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n2076_));
NAND2X1 NAND2X1_1738 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1829_), .Y(u5__abc_78290_new_n2091_));
NAND2X1 NAND2X1_1739 ( .A(u5__abc_78290_new_n2091_), .B(u5__abc_78290_new_n1711_), .Y(u5__abc_78290_new_n2092_));
NAND2X1 NAND2X1_174 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1548_));
NAND2X1 NAND2X1_1740 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1790_), .Y(u5__abc_78290_new_n2096_));
NAND2X1 NAND2X1_1741 ( .A(u5__abc_78290_new_n1034_), .B(u5__abc_78290_new_n2096_), .Y(u5__abc_78290_new_n2097_));
NAND2X1 NAND2X1_1742 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1794_), .Y(u5__abc_78290_new_n2102_));
NAND2X1 NAND2X1_1743 ( .A(u5__abc_78290_new_n2101_), .B(u5__abc_78290_new_n2102_), .Y(u5__abc_78290_new_n2103_));
NAND2X1 NAND2X1_1744 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1720_), .Y(u5__abc_78290_new_n2106_));
NAND2X1 NAND2X1_1745 ( .A(u5__abc_78290_new_n1717_), .B(u5__abc_78290_new_n2106_), .Y(u5__abc_78290_new_n2112_));
NAND2X1 NAND2X1_1746 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1722_), .Y(u5__abc_78290_new_n2113_));
NAND2X1 NAND2X1_1747 ( .A(u5__abc_78290_new_n2135_), .B(u5__abc_78290_new_n1007_), .Y(u5__abc_78290_new_n2136_));
NAND2X1 NAND2X1_1748 ( .A(u5__abc_78290_new_n2148_), .B(u5__abc_78290_new_n1345_), .Y(u5__abc_78290_new_n2149_));
NAND2X1 NAND2X1_1749 ( .A(u5__abc_78290_new_n455_), .B(u5__abc_78290_new_n982_), .Y(u5__abc_78290_new_n2157_));
NAND2X1 NAND2X1_175 ( .A(u0__abc_74894_new_n1536_), .B(u0__abc_74894_new_n1554_), .Y(u0__0sp_tms_31_0__19_));
NAND2X1 NAND2X1_1750 ( .A(u5__abc_78290_new_n1651_), .B(u5__abc_78290_new_n1632_), .Y(u5__abc_78290_new_n2167_));
NAND2X1 NAND2X1_1751 ( .A(u5__abc_78290_new_n580_), .B(u5__abc_78290_new_n2173_), .Y(u5__abc_78290_new_n2174_));
NAND2X1 NAND2X1_1752 ( .A(u5__abc_78290_new_n2169_), .B(u5__abc_78290_new_n2175_), .Y(u5__abc_78290_new_n2176_));
NAND2X1 NAND2X1_1753 ( .A(u5__abc_78290_new_n1390_), .B(u5__abc_78290_new_n1641_), .Y(u5__abc_78290_new_n2179_));
NAND2X1 NAND2X1_1754 ( .A(u5__abc_78290_new_n1039_), .B(u5__abc_78290_new_n1089_), .Y(u5__abc_78290_new_n2180_));
NAND2X1 NAND2X1_1755 ( .A(u5__abc_78290_new_n1051_), .B(u5__abc_78290_new_n1045_), .Y(u5__abc_78290_new_n2196_));
NAND2X1 NAND2X1_1756 ( .A(u5__abc_78290_new_n1070_), .B(u5__abc_78290_new_n2196_), .Y(u5__abc_78290_new_n2197_));
NAND2X1 NAND2X1_1757 ( .A(u5__abc_78290_new_n1095_), .B(u5__abc_78290_new_n2201_), .Y(u5__abc_78290_new_n2202_));
NAND2X1 NAND2X1_1758 ( .A(u5__abc_78290_new_n2079_), .B(u5__abc_78290_new_n2028_), .Y(u5__abc_78290_new_n2206_));
NAND2X1 NAND2X1_1759 ( .A(u5__abc_78290_new_n2231_), .B(u5__abc_78290_new_n2045_), .Y(u5__abc_78290_new_n2232_));
NAND2X1 NAND2X1_176 ( .A(sp_tms_20_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1556_));
NAND2X1 NAND2X1_1760 ( .A(u5__abc_78290_new_n2165_), .B(u5__abc_78290_new_n2254_), .Y(u5__abc_78290_new_n2255_));
NAND2X1 NAND2X1_1761 ( .A(u5__abc_78290_new_n2249_), .B(u5__abc_78290_new_n1632_), .Y(u5__abc_78290_new_n2268_));
NAND2X1 NAND2X1_1762 ( .A(u5__abc_78290_new_n1072_), .B(u5__abc_78290_new_n1117_), .Y(u5__abc_78290_new_n2276_));
NAND2X1 NAND2X1_1763 ( .A(u5__abc_78290_new_n1363_), .B(u5__abc_78290_new_n2278_), .Y(u5__abc_78290_new_n2279_));
NAND2X1 NAND2X1_1764 ( .A(u5__abc_78290_new_n2288_), .B(u5__abc_78290_new_n2281_), .Y(u5__abc_78290_new_n2333_));
NAND2X1 NAND2X1_1765 ( .A(u5__abc_78290_new_n2356_), .B(u5__abc_78290_new_n2341_), .Y(u5__abc_78290_new_n2357_));
NAND2X1 NAND2X1_1766 ( .A(u5__abc_78290_new_n2358_), .B(u5__abc_78290_new_n2350_), .Y(u5__abc_78290_new_n2359_));
NAND2X1 NAND2X1_1767 ( .A(u5__abc_78290_new_n786_), .B(u5__abc_78290_new_n2056_), .Y(u5__abc_78290_new_n2370_));
NAND2X1 NAND2X1_1768 ( .A(u5__abc_78290_new_n2377_), .B(u5__abc_78290_new_n2371_), .Y(u5__abc_78290_new_n2378_));
NAND2X1 NAND2X1_1769 ( .A(u5__abc_78290_new_n2381_), .B(u5__abc_78290_new_n2277_), .Y(u5__abc_78290_new_n2382_));
NAND2X1 NAND2X1_177 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1557_), .Y(u0__abc_74894_new_n1558_));
NAND2X1 NAND2X1_1770 ( .A(u5__abc_78290_new_n2395_), .B(u5__abc_78290_new_n2400_), .Y(u5__abc_78290_new_n2401_));
NAND2X1 NAND2X1_1771 ( .A(u5__abc_78290_new_n2394_), .B(u5__abc_78290_new_n2402_), .Y(u5__abc_78290_new_n2403_));
NAND2X1 NAND2X1_1772 ( .A(u5__abc_78290_new_n2393_), .B(u5__abc_78290_new_n2406_), .Y(u5__abc_78290_new_n2407_));
NAND2X1 NAND2X1_1773 ( .A(u5__abc_78290_new_n1647_), .B(u5__abc_78290_new_n2178_), .Y(u5__abc_78290_new_n2428_));
NAND2X1 NAND2X1_1774 ( .A(u5_timer2_1_), .B(u5_timer2_0_), .Y(u5__abc_78290_new_n2452_));
NAND2X1 NAND2X1_1775 ( .A(u5__abc_78290_new_n2259_), .B(u5__abc_78290_new_n2437_), .Y(u5__abc_78290_new_n2468_));
NAND2X1 NAND2X1_1776 ( .A(u5__abc_78290_new_n2469_), .B(u5__abc_78290_new_n2472_), .Y(u5__abc_78290_new_n2473_));
NAND2X1 NAND2X1_1777 ( .A(u5__abc_78290_new_n2476_), .B(u5__abc_78290_new_n2475_), .Y(u5__abc_78290_new_n2477_));
NAND2X1 NAND2X1_1778 ( .A(u5__abc_78290_new_n2450_), .B(u5__abc_78290_new_n2041_), .Y(u5__abc_78290_new_n2510_));
NAND2X1 NAND2X1_1779 ( .A(u5__abc_78290_new_n2516_), .B(u5__abc_78290_new_n2379_), .Y(u5__abc_78290_new_n2517_));
NAND2X1 NAND2X1_178 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1559_), .Y(u0__abc_74894_new_n1560_));
NAND2X1 NAND2X1_1780 ( .A(u5__abc_78290_new_n2231_), .B(u5__abc_78290_new_n2413_), .Y(u5__abc_78290_new_n2522_));
NAND2X1 NAND2X1_1781 ( .A(u5__abc_78290_new_n2534_), .B(u5__abc_78290_new_n2536_), .Y(u5__abc_78290_new_n2537_));
NAND2X1 NAND2X1_1782 ( .A(u5_ack_cnt_1_), .B(u5_ack_cnt_0_), .Y(u5__abc_78290_new_n2541_));
NAND2X1 NAND2X1_1783 ( .A(u5__abc_78290_new_n2543_), .B(u5__abc_78290_new_n2535_), .Y(u5__abc_78290_new_n2544_));
NAND2X1 NAND2X1_1784 ( .A(u5_ack_cnt_2_), .B(u5__abc_78290_new_n2542_), .Y(u5__abc_78290_new_n2554_));
NAND2X1 NAND2X1_1785 ( .A(u5_mc_le), .B(u5_cmd_asserted2), .Y(u5__abc_78290_new_n2558_));
NAND2X1 NAND2X1_1786 ( .A(u5_mc_adv_r), .B(u5_mc_le), .Y(u5__abc_78290_new_n2563_));
NAND2X1 NAND2X1_1787 ( .A(u5__abc_78290_new_n2565_), .B(u5__abc_78290_new_n2157_), .Y(u5__abc_78290_new_n2566_));
NAND2X1 NAND2X1_1788 ( .A(u5__abc_78290_new_n2571_), .B(u5__abc_78290_new_n2208_), .Y(u5__abc_78290_new_n2572_));
NAND2X1 NAND2X1_1789 ( .A(u5__0mc_le_0_0_), .B(mc_adv_d), .Y(u5__abc_78290_new_n2574_));
NAND2X1 NAND2X1_179 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1561_));
NAND2X1 NAND2X1_1790 ( .A(u5__abc_78290_new_n1343_), .B(u5__abc_78290_new_n1478_), .Y(u5__abc_78290_new_n2577_));
NAND2X1 NAND2X1_1791 ( .A(u5__abc_78290_new_n1543_), .B(u5__abc_78290_new_n1492_), .Y(u5__abc_78290_new_n2618_));
NAND2X1 NAND2X1_1792 ( .A(u5_wb_cycle), .B(u5__abc_78290_new_n1609_), .Y(u5__abc_78290_new_n2636_));
NAND2X1 NAND2X1_1793 ( .A(u5__abc_78290_new_n2647_), .B(u5__abc_78290_new_n2648_), .Y(u5__abc_78290_new_n2649_));
NAND2X1 NAND2X1_1794 ( .A(u5_kro), .B(u5__abc_78290_new_n1414_), .Y(u5__abc_78290_new_n2650_));
NAND2X1 NAND2X1_1795 ( .A(u5_lookup_ready2), .B(bank_open), .Y(u5__abc_78290_new_n2651_));
NAND2X1 NAND2X1_1796 ( .A(u5__abc_78290_new_n2656_), .B(u5__abc_78290_new_n1478_), .Y(u5__abc_78290_new_n2657_));
NAND2X1 NAND2X1_1797 ( .A(u5__abc_78290_new_n1514_), .B(u5__abc_78290_new_n2666_), .Y(u5__abc_78290_new_n2667_));
NAND2X1 NAND2X1_1798 ( .A(u5_state_7_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2681_));
NAND2X1 NAND2X1_1799 ( .A(u5__abc_78290_new_n777_), .B(u5__abc_78290_new_n1990_), .Y(u5__abc_78290_new_n2682_));
NAND2X1 NAND2X1_18 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1159_), .Y(u0__abc_74894_new_n1160_));
NAND2X1 NAND2X1_180 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1562_));
NAND2X1 NAND2X1_1800 ( .A(u5__abc_78290_new_n2696_), .B(u5__abc_78290_new_n2698_), .Y(u5__abc_78290_new_n2699_));
NAND2X1 NAND2X1_1801 ( .A(u5__abc_78290_new_n2704_), .B(u5__abc_78290_new_n1262_), .Y(u5__abc_78290_new_n2705_));
NAND2X1 NAND2X1_1802 ( .A(u5_state_11_), .B(u5__abc_78290_new_n2605_), .Y(u5__abc_78290_new_n2712_));
NAND2X1 NAND2X1_1803 ( .A(u5_wb_cycle), .B(u1_wb_write_go), .Y(u5__abc_78290_new_n2714_));
NAND2X1 NAND2X1_1804 ( .A(u5__abc_78290_new_n492_), .B(u5__abc_78290_new_n1375_), .Y(u5__abc_78290_new_n2718_));
NAND2X1 NAND2X1_1805 ( .A(u5__abc_78290_new_n1325_), .B(u5__abc_78290_new_n1262_), .Y(u5__abc_78290_new_n2727_));
NAND2X1 NAND2X1_1806 ( .A(u5_state_14_), .B(u5__abc_78290_new_n2659_), .Y(u5__abc_78290_new_n2735_));
NAND2X1 NAND2X1_1807 ( .A(u5__abc_78290_new_n1420_), .B(u5__abc_78290_new_n2737_), .Y(u5__abc_78290_new_n2738_));
NAND2X1 NAND2X1_1808 ( .A(u5__abc_78290_new_n2653_), .B(u5__abc_78290_new_n2578_), .Y(u5__abc_78290_new_n2742_));
NAND2X1 NAND2X1_1809 ( .A(u5_state_15_), .B(u5_wb_wait), .Y(u5__abc_78290_new_n2743_));
NAND2X1 NAND2X1_181 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1565_));
NAND2X1 NAND2X1_1810 ( .A(u5__abc_78290_new_n1631_), .B(u5__abc_78290_new_n1609_), .Y(u5__abc_78290_new_n2766_));
NAND2X1 NAND2X1_1811 ( .A(u5__abc_78290_new_n571_), .B(u5__abc_78290_new_n1375_), .Y(u5__abc_78290_new_n2776_));
NAND2X1 NAND2X1_1812 ( .A(u5_state_19_), .B(u5__abc_78290_new_n1375_), .Y(u5__abc_78290_new_n2791_));
NAND2X1 NAND2X1_1813 ( .A(u5_state_22_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2804_));
NAND2X1 NAND2X1_1814 ( .A(u5_state_23_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2808_));
NAND2X1 NAND2X1_1815 ( .A(u5__abc_78290_new_n590_), .B(u5__abc_78290_new_n1990_), .Y(u5__abc_78290_new_n2809_));
NAND2X1 NAND2X1_1816 ( .A(u5_state_24_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2813_));
NAND2X1 NAND2X1_1817 ( .A(u5_tmr_done), .B(u5_ir_cnt_done), .Y(u5__abc_78290_new_n2815_));
NAND2X1 NAND2X1_1818 ( .A(u5_state_25_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2820_));
NAND2X1 NAND2X1_1819 ( .A(u5_state_26_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2825_));
NAND2X1 NAND2X1_182 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1568_));
NAND2X1 NAND2X1_1820 ( .A(u5_state_28_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2833_));
NAND2X1 NAND2X1_1821 ( .A(u5_state_29_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2839_));
NAND2X1 NAND2X1_1822 ( .A(u5__abc_78290_new_n2840_), .B(u5__abc_78290_new_n2841_), .Y(u5__abc_78290_new_n2842_));
NAND2X1 NAND2X1_1823 ( .A(u5_state_30_), .B(u5__abc_78290_new_n2680_), .Y(u5__abc_78290_new_n2844_));
NAND2X1 NAND2X1_1824 ( .A(u5__abc_78290_new_n2845_), .B(u5__abc_78290_new_n2846_), .Y(u5__abc_78290_new_n2847_));
NAND2X1 NAND2X1_1825 ( .A(u5_state_32_), .B(u5__abc_78290_new_n1375_), .Y(u5__abc_78290_new_n2852_));
NAND2X1 NAND2X1_1826 ( .A(u5_state_37_), .B(u5__abc_78290_new_n2565_), .Y(u5__abc_78290_new_n2869_));
NAND2X1 NAND2X1_1827 ( .A(u5__abc_78290_new_n698_), .B(u5__abc_78290_new_n2565_), .Y(u5__abc_78290_new_n2878_));
NAND2X1 NAND2X1_1828 ( .A(u5__abc_78290_new_n2897_), .B(u5__abc_78290_new_n2874_), .Y(u5__abc_78290_new_n2898_));
NAND2X1 NAND2X1_1829 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n2417_), .Y(u5__abc_78290_new_n2912_));
NAND2X1 NAND2X1_183 ( .A(u0__abc_74894_new_n1556_), .B(u0__abc_74894_new_n1574_), .Y(u0__0sp_tms_31_0__20_));
NAND2X1 NAND2X1_1830 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n2914_), .Y(u5__abc_78290_new_n2917_));
NAND2X1 NAND2X1_1831 ( .A(u5__abc_78290_new_n1482_), .B(u5__abc_78290_new_n1481_), .Y(u5__abc_78290_new_n2919_));
NAND2X1 NAND2X1_1832 ( .A(u5__abc_78290_new_n2920_), .B(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2921_));
NAND2X1 NAND2X1_1833 ( .A(u5__abc_78290_new_n938_), .B(u5__abc_78290_new_n1990_), .Y(u5__abc_78290_new_n2927_));
NAND2X1 NAND2X1_1834 ( .A(u3_wb_read_go), .B(u5__abc_78290_new_n2605_), .Y(u5__abc_78290_new_n2930_));
NAND2X1 NAND2X1_1835 ( .A(u5_state_55_), .B(u5_wb_wait), .Y(u5__abc_78290_new_n2935_));
NAND2X1 NAND2X1_1836 ( .A(u5__abc_78290_new_n2945_), .B(u5__abc_78290_new_n2942_), .Y(u5_next_state_56_));
NAND2X1 NAND2X1_1837 ( .A(u5__abc_78290_new_n2961_), .B(u5__abc_78290_new_n2958_), .Y(u5_next_state_58_));
NAND2X1 NAND2X1_1838 ( .A(u5__abc_78290_new_n1324_), .B(u5__abc_78290_new_n1487_), .Y(u5__abc_78290_new_n2967_));
NAND2X1 NAND2X1_1839 ( .A(u5__abc_78290_new_n2968_), .B(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2969_));
NAND2X1 NAND2X1_184 ( .A(sp_tms_21_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1576_));
NAND2X1 NAND2X1_1840 ( .A(u5_state_60_), .B(u5__abc_78290_new_n2970_), .Y(u5__abc_78290_new_n2971_));
NAND2X1 NAND2X1_1841 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n1616_), .Y(u5__abc_78290_new_n2979_));
NAND2X1 NAND2X1_1842 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1895_), .Y(u5__abc_78290_new_n2981_));
NAND2X1 NAND2X1_1843 ( .A(u5_state_63_), .B(u5__abc_78290_new_n2970_), .Y(u5__abc_78290_new_n2985_));
NAND2X1 NAND2X1_1844 ( .A(u5__abc_78290_new_n487_), .B(u5__abc_78290_new_n2605_), .Y(u5__abc_78290_new_n3003_));
NAND2X1 NAND2X1_1845 ( .A(u5__abc_78290_new_n3012_), .B(u5__abc_78290_new_n3008_), .Y(u5__abc_78290_new_n3013_));
NAND2X1 NAND2X1_1846 ( .A(u5__abc_78290_new_n1343_), .B(u5__abc_78290_new_n2782_), .Y(u5__abc_78290_new_n3017_));
NAND2X1 NAND2X1_1847 ( .A(u5__abc_78290_new_n1104_), .B(u5__abc_78290_new_n2568_), .Y(u5__abc_78290_new_n3023_));
NAND2X1 NAND2X1_1848 ( .A(u5__abc_78290_new_n1984_), .B(u5__abc_78290_new_n3029_), .Y(u5__abc_78290_new_n3030_));
NAND2X1 NAND2X1_1849 ( .A(u5__abc_78290_new_n3035_), .B(u5__abc_78290_new_n2795_), .Y(u5__abc_78290_new_n3036_));
NAND2X1 NAND2X1_185 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1577_), .Y(u0__abc_74894_new_n1578_));
NAND2X1 NAND2X1_1850 ( .A(u5_wb_stb_first), .B(u5__abc_78290_new_n1478_), .Y(u5__abc_78290_new_n3037_));
NAND2X1 NAND2X1_1851 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n1414_), .Y(u5__abc_78290_new_n3039_));
NAND2X1 NAND2X1_1852 ( .A(u5__abc_78290_new_n1363_), .B(u5__abc_78290_new_n1543_), .Y(u5__abc_78290_new_n3045_));
NAND2X1 NAND2X1_1853 ( .A(u5__abc_78290_new_n3051_), .B(u5__abc_78290_new_n3058_), .Y(u5_mc_c_oe_d));
NAND2X1 NAND2X1_1854 ( .A(u5__abc_78290_new_n3072_), .B(u5__abc_78290_new_n3080_), .Y(u5__abc_78290_new_n3081_));
NAND2X1 NAND2X1_1855 ( .A(u5__abc_78290_new_n2181_), .B(u5__abc_78290_new_n3087_), .Y(u5__abc_78290_new_n3088_));
NAND2X1 NAND2X1_1856 ( .A(u5__abc_78290_new_n3123_), .B(u5__abc_78290_new_n3072_), .Y(u5__abc_78290_new_n3124_));
NAND2X1 NAND2X1_1857 ( .A(u5__abc_78290_new_n3126_), .B(u5__abc_78290_new_n2221_), .Y(u5__abc_78290_new_n3127_));
NAND2X1 NAND2X1_1858 ( .A(u5__abc_78290_new_n3129_), .B(u5__abc_78290_new_n2280_), .Y(u5__abc_78290_new_n3130_));
NAND2X1 NAND2X1_1859 ( .A(u5__abc_78290_new_n2422_), .B(u5__abc_78290_new_n2391_), .Y(u5__abc_78290_new_n3147_));
NAND2X1 NAND2X1_186 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1579_), .Y(u0__abc_74894_new_n1580_));
NAND2X1 NAND2X1_1860 ( .A(u5_wb_cycle), .B(wb_cyc_i), .Y(u5__abc_78290_new_n3153_));
NAND2X1 NAND2X1_1861 ( .A(u5__abc_78290_new_n3155_), .B(u5__abc_78290_new_n3156_), .Y(u5__abc_78290_new_n3157_));
NAND2X1 NAND2X1_1862 ( .A(u6__abc_81318_new_n133_), .B(u6__abc_81318_new_n134_), .Y(u6__abc_81318_new_n135_));
NAND2X1 NAND2X1_1863 ( .A(mem_ack), .B(u6__abc_81318_new_n140_), .Y(u6__abc_81318_new_n141_));
NAND2X1 NAND2X1_1864 ( .A(rf_dout_0_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n147_));
NAND2X1 NAND2X1_1865 ( .A(rf_dout_1_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n150_));
NAND2X1 NAND2X1_1866 ( .A(rf_dout_2_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n153_));
NAND2X1 NAND2X1_1867 ( .A(rf_dout_3_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n156_));
NAND2X1 NAND2X1_1868 ( .A(rf_dout_4_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n159_));
NAND2X1 NAND2X1_1869 ( .A(rf_dout_5_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n162_));
NAND2X1 NAND2X1_187 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1581_));
NAND2X1 NAND2X1_1870 ( .A(rf_dout_6_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n165_));
NAND2X1 NAND2X1_1871 ( .A(rf_dout_7_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n168_));
NAND2X1 NAND2X1_1872 ( .A(rf_dout_8_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n171_));
NAND2X1 NAND2X1_1873 ( .A(rf_dout_9_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n174_));
NAND2X1 NAND2X1_1874 ( .A(rf_dout_10_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n177_));
NAND2X1 NAND2X1_1875 ( .A(rf_dout_11_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n180_));
NAND2X1 NAND2X1_1876 ( .A(rf_dout_12_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n183_));
NAND2X1 NAND2X1_1877 ( .A(rf_dout_13_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n186_));
NAND2X1 NAND2X1_1878 ( .A(rf_dout_14_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n189_));
NAND2X1 NAND2X1_1879 ( .A(rf_dout_15_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n192_));
NAND2X1 NAND2X1_188 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1582_));
NAND2X1 NAND2X1_1880 ( .A(rf_dout_16_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n195_));
NAND2X1 NAND2X1_1881 ( .A(rf_dout_17_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n198_));
NAND2X1 NAND2X1_1882 ( .A(rf_dout_18_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n201_));
NAND2X1 NAND2X1_1883 ( .A(rf_dout_19_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n204_));
NAND2X1 NAND2X1_1884 ( .A(rf_dout_20_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n207_));
NAND2X1 NAND2X1_1885 ( .A(rf_dout_21_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n210_));
NAND2X1 NAND2X1_1886 ( .A(rf_dout_22_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n213_));
NAND2X1 NAND2X1_1887 ( .A(rf_dout_23_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n216_));
NAND2X1 NAND2X1_1888 ( .A(rf_dout_24_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n219_));
NAND2X1 NAND2X1_1889 ( .A(rf_dout_25_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n222_));
NAND2X1 NAND2X1_189 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1585_));
NAND2X1 NAND2X1_1890 ( .A(rf_dout_26_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n225_));
NAND2X1 NAND2X1_1891 ( .A(rf_dout_27_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n228_));
NAND2X1 NAND2X1_1892 ( .A(rf_dout_28_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n231_));
NAND2X1 NAND2X1_1893 ( .A(rf_dout_29_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n234_));
NAND2X1 NAND2X1_1894 ( .A(rf_dout_30_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n237_));
NAND2X1 NAND2X1_1895 ( .A(rf_dout_31_), .B(u6__abc_81318_new_n135_), .Y(u6__abc_81318_new_n240_));
NAND2X1 NAND2X1_1896 ( .A(u6_rmw_en), .B(u6__abc_81318_new_n242_), .Y(u6__abc_81318_new_n245_));
NAND2X1 NAND2X1_1897 ( .A(u6__abc_81318_new_n254_), .B(u6__abc_81318_new_n252_), .Y(u6__abc_81318_new_n255_));
NAND2X1 NAND2X1_1898 ( .A(wb_cyc_i), .B(u6_read_go_r1), .Y(u6__abc_81318_new_n258_));
NAND2X1 NAND2X1_1899 ( .A(wb_cyc_i), .B(u6_write_go_r1), .Y(u6__abc_81318_new_n265_));
NAND2X1 NAND2X1_19 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1161_));
NAND2X1 NAND2X1_190 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1588_));
NAND2X1 NAND2X1_1900 ( .A(u6__abc_81318_new_n270_), .B(u6__abc_81318_new_n249_), .Y(u6__abc_81318_new_n273_));
NAND2X1 NAND2X1_1901 ( .A(wb_cyc_i), .B(u6__abc_81318_new_n137_), .Y(u6__abc_81318_new_n275_));
NAND2X1 NAND2X1_1902 ( .A(wb_stb_i), .B(wb_cyc_i), .Y(u7__abc_73829_new_n88_));
NAND2X1 NAND2X1_1903 ( .A(u7_mc_dqm_r_0_), .B(u7__abc_73829_new_n88_), .Y(u7__abc_73829_new_n89_));
NAND2X1 NAND2X1_1904 ( .A(u7_mc_dqm_r_1_), .B(u7__abc_73829_new_n88_), .Y(u7__abc_73829_new_n92_));
NAND2X1 NAND2X1_1905 ( .A(u7_mc_dqm_r_2_), .B(u7__abc_73829_new_n88_), .Y(u7__abc_73829_new_n95_));
NAND2X1 NAND2X1_1906 ( .A(u7_mc_dqm_r_3_), .B(u7__abc_73829_new_n88_), .Y(u7__abc_73829_new_n98_));
NAND2X1 NAND2X1_1907 ( .A(cs_0_), .B(u7__abc_73829_new_n101_), .Y(u7__abc_73829_new_n102_));
NAND2X1 NAND2X1_1908 ( .A(spec_req_cs_0_), .B(lmr_sel), .Y(u7__abc_73829_new_n103_));
NAND2X1 NAND2X1_1909 ( .A(u7__abc_73829_new_n104_), .B(u7__abc_73829_new_n108_), .Y(u7__0mc_cs__0_0_));
NAND2X1 NAND2X1_191 ( .A(u0__abc_74894_new_n1576_), .B(u0__abc_74894_new_n1594_), .Y(u0__0sp_tms_31_0__21_));
NAND2X1 NAND2X1_1910 ( .A(cs_1_), .B(u7__abc_73829_new_n101_), .Y(u7__abc_73829_new_n110_));
NAND2X1 NAND2X1_1911 ( .A(lmr_sel), .B(spec_req_cs_1_), .Y(u7__abc_73829_new_n111_));
NAND2X1 NAND2X1_1912 ( .A(u7__abc_73829_new_n112_), .B(u7__abc_73829_new_n114_), .Y(u7__0mc_cs__1_1_));
NAND2X1 NAND2X1_1913 ( .A(cs_2_), .B(u7__abc_73829_new_n101_), .Y(u7__abc_73829_new_n116_));
NAND2X1 NAND2X1_1914 ( .A(lmr_sel), .B(spec_req_cs_2_), .Y(u7__abc_73829_new_n117_));
NAND2X1 NAND2X1_1915 ( .A(u7__abc_73829_new_n118_), .B(u7__abc_73829_new_n120_), .Y(u7__0mc_cs__2_2_));
NAND2X1 NAND2X1_1916 ( .A(cs_3_), .B(u7__abc_73829_new_n101_), .Y(u7__abc_73829_new_n122_));
NAND2X1 NAND2X1_1917 ( .A(lmr_sel), .B(spec_req_cs_3_), .Y(u7__abc_73829_new_n123_));
NAND2X1 NAND2X1_1918 ( .A(u7__abc_73829_new_n124_), .B(u7__abc_73829_new_n126_), .Y(u7__0mc_cs__3_3_));
NAND2X1 NAND2X1_1919 ( .A(cs_4_), .B(u7__abc_73829_new_n101_), .Y(u7__abc_73829_new_n128_));
NAND2X1 NAND2X1_192 ( .A(sp_tms_22_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1596_));
NAND2X1 NAND2X1_1920 ( .A(lmr_sel), .B(spec_req_cs_4_), .Y(u7__abc_73829_new_n129_));
NAND2X1 NAND2X1_1921 ( .A(u7__abc_73829_new_n130_), .B(u7__abc_73829_new_n132_), .Y(u7__0mc_cs__4_4_));
NAND2X1 NAND2X1_1922 ( .A(cs_5_), .B(u7__abc_73829_new_n101_), .Y(u7__abc_73829_new_n134_));
NAND2X1 NAND2X1_1923 ( .A(lmr_sel), .B(spec_req_cs_5_), .Y(u7__abc_73829_new_n135_));
NAND2X1 NAND2X1_1924 ( .A(u7__abc_73829_new_n136_), .B(u7__abc_73829_new_n138_), .Y(u7__0mc_cs__5_5_));
NAND2X1 NAND2X1_1925 ( .A(cs_6_), .B(u7__abc_73829_new_n101_), .Y(u7__abc_73829_new_n140_));
NAND2X1 NAND2X1_1926 ( .A(lmr_sel), .B(spec_req_cs_6_), .Y(u7__abc_73829_new_n141_));
NAND2X1 NAND2X1_1927 ( .A(u7__abc_73829_new_n142_), .B(u7__abc_73829_new_n144_), .Y(u7__0mc_cs__6_6_));
NAND2X1 NAND2X1_1928 ( .A(cs_7_), .B(u7__abc_73829_new_n101_), .Y(u7__abc_73829_new_n146_));
NAND2X1 NAND2X1_1929 ( .A(lmr_sel), .B(spec_req_cs_7_), .Y(u7__abc_73829_new_n147_));
NAND2X1 NAND2X1_193 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1597_), .Y(u0__abc_74894_new_n1598_));
NAND2X1 NAND2X1_1930 ( .A(u7__abc_73829_new_n148_), .B(u7__abc_73829_new_n150_), .Y(u7__0mc_cs__7_7_));
NAND2X1 NAND2X1_1931 ( .A(data_oe), .B(mc_c_oe_d), .Y(u7__abc_73829_new_n155_));
NAND2X1 NAND2X1_194 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1599_), .Y(u0__abc_74894_new_n1600_));
NAND2X1 NAND2X1_195 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1601_));
NAND2X1 NAND2X1_196 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1602_));
NAND2X1 NAND2X1_197 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1605_));
NAND2X1 NAND2X1_198 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1608_));
NAND2X1 NAND2X1_199 ( .A(u0__abc_74894_new_n1596_), .B(u0__abc_74894_new_n1614_), .Y(u0__0sp_tms_31_0__22_));
NAND2X1 NAND2X1_2 ( .A(u0__abc_74894_new_n1102_), .B(u0__abc_74894_new_n1101_), .Y(u0__abc_74894_new_n1103_));
NAND2X1 NAND2X1_20 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1162_));
NAND2X1 NAND2X1_200 ( .A(sp_tms_23_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1616_));
NAND2X1 NAND2X1_201 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1617_), .Y(u0__abc_74894_new_n1618_));
NAND2X1 NAND2X1_202 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1619_), .Y(u0__abc_74894_new_n1620_));
NAND2X1 NAND2X1_203 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1621_));
NAND2X1 NAND2X1_204 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1622_));
NAND2X1 NAND2X1_205 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1625_));
NAND2X1 NAND2X1_206 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1628_));
NAND2X1 NAND2X1_207 ( .A(u0__abc_74894_new_n1616_), .B(u0__abc_74894_new_n1634_), .Y(u0__0sp_tms_31_0__23_));
NAND2X1 NAND2X1_208 ( .A(sp_tms_24_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1636_));
NAND2X1 NAND2X1_209 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1637_), .Y(u0__abc_74894_new_n1638_));
NAND2X1 NAND2X1_21 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1165_));
NAND2X1 NAND2X1_210 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1639_), .Y(u0__abc_74894_new_n1640_));
NAND2X1 NAND2X1_211 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1641_));
NAND2X1 NAND2X1_212 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1642_));
NAND2X1 NAND2X1_213 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1645_));
NAND2X1 NAND2X1_214 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1648_));
NAND2X1 NAND2X1_215 ( .A(u0__abc_74894_new_n1636_), .B(u0__abc_74894_new_n1654_), .Y(u0__0sp_tms_31_0__24_));
NAND2X1 NAND2X1_216 ( .A(sp_tms_25_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1656_));
NAND2X1 NAND2X1_217 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1657_), .Y(u0__abc_74894_new_n1658_));
NAND2X1 NAND2X1_218 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1659_), .Y(u0__abc_74894_new_n1660_));
NAND2X1 NAND2X1_219 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1661_));
NAND2X1 NAND2X1_22 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1168_));
NAND2X1 NAND2X1_220 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1662_));
NAND2X1 NAND2X1_221 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1665_));
NAND2X1 NAND2X1_222 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1668_));
NAND2X1 NAND2X1_223 ( .A(u0__abc_74894_new_n1656_), .B(u0__abc_74894_new_n1674_), .Y(u0__0sp_tms_31_0__25_));
NAND2X1 NAND2X1_224 ( .A(sp_tms_26_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1676_));
NAND2X1 NAND2X1_225 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1677_), .Y(u0__abc_74894_new_n1678_));
NAND2X1 NAND2X1_226 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1679_), .Y(u0__abc_74894_new_n1680_));
NAND2X1 NAND2X1_227 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1681_));
NAND2X1 NAND2X1_228 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1682_));
NAND2X1 NAND2X1_229 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1685_));
NAND2X1 NAND2X1_23 ( .A(u0__abc_74894_new_n1156_), .B(u0__abc_74894_new_n1174_), .Y(u0__0sp_tms_31_0__0_));
NAND2X1 NAND2X1_230 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1688_));
NAND2X1 NAND2X1_231 ( .A(u0__abc_74894_new_n1676_), .B(u0__abc_74894_new_n1694_), .Y(u0__0sp_tms_31_0__26_));
NAND2X1 NAND2X1_232 ( .A(sp_tms_27_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1696_));
NAND2X1 NAND2X1_233 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1697_), .Y(u0__abc_74894_new_n1698_));
NAND2X1 NAND2X1_234 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1699_), .Y(u0__abc_74894_new_n1700_));
NAND2X1 NAND2X1_235 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1701_));
NAND2X1 NAND2X1_236 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1702_));
NAND2X1 NAND2X1_237 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1705_));
NAND2X1 NAND2X1_238 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1708_));
NAND2X1 NAND2X1_239 ( .A(u0__abc_74894_new_n1696_), .B(u0__abc_74894_new_n1714_), .Y(u0__0sp_tms_31_0__27_));
NAND2X1 NAND2X1_24 ( .A(sp_tms_1_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1176_));
NAND2X1 NAND2X1_240 ( .A(cs_le_d), .B(u0__abc_74894_new_n1154_), .Y(u0__abc_74894_new_n1796_));
NAND2X1 NAND2X1_241 ( .A(sp_csc_1_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1817_));
NAND2X1 NAND2X1_242 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1818_), .Y(u0__abc_74894_new_n1819_));
NAND2X1 NAND2X1_243 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1820_), .Y(u0__abc_74894_new_n1821_));
NAND2X1 NAND2X1_244 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1822_));
NAND2X1 NAND2X1_245 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1823_));
NAND2X1 NAND2X1_246 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1826_));
NAND2X1 NAND2X1_247 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1829_));
NAND2X1 NAND2X1_248 ( .A(u0__abc_74894_new_n1817_), .B(u0__abc_74894_new_n1835_), .Y(u0__0sp_csc_31_0__1_));
NAND2X1 NAND2X1_249 ( .A(sp_csc_2_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1837_));
NAND2X1 NAND2X1_25 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1177_), .Y(u0__abc_74894_new_n1178_));
NAND2X1 NAND2X1_250 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1838_), .Y(u0__abc_74894_new_n1839_));
NAND2X1 NAND2X1_251 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1840_), .Y(u0__abc_74894_new_n1841_));
NAND2X1 NAND2X1_252 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1842_));
NAND2X1 NAND2X1_253 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1843_));
NAND2X1 NAND2X1_254 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1846_));
NAND2X1 NAND2X1_255 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1849_));
NAND2X1 NAND2X1_256 ( .A(u0__abc_74894_new_n1837_), .B(u0__abc_74894_new_n1855_), .Y(u0__0sp_csc_31_0__2_));
NAND2X1 NAND2X1_257 ( .A(sp_csc_3_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1857_));
NAND2X1 NAND2X1_258 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1858_), .Y(u0__abc_74894_new_n1859_));
NAND2X1 NAND2X1_259 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1860_), .Y(u0__abc_74894_new_n1861_));
NAND2X1 NAND2X1_26 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1179_), .Y(u0__abc_74894_new_n1180_));
NAND2X1 NAND2X1_260 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1862_));
NAND2X1 NAND2X1_261 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1863_));
NAND2X1 NAND2X1_262 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1866_));
NAND2X1 NAND2X1_263 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1869_));
NAND2X1 NAND2X1_264 ( .A(u0__abc_74894_new_n1857_), .B(u0__abc_74894_new_n1875_), .Y(u0__0sp_csc_31_0__3_));
NAND2X1 NAND2X1_265 ( .A(sp_csc_4_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1877_));
NAND2X1 NAND2X1_266 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1878_), .Y(u0__abc_74894_new_n1879_));
NAND2X1 NAND2X1_267 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1880_), .Y(u0__abc_74894_new_n1881_));
NAND2X1 NAND2X1_268 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1882_));
NAND2X1 NAND2X1_269 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1883_));
NAND2X1 NAND2X1_27 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1181_));
NAND2X1 NAND2X1_270 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1886_));
NAND2X1 NAND2X1_271 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1889_));
NAND2X1 NAND2X1_272 ( .A(u0__abc_74894_new_n1877_), .B(u0__abc_74894_new_n1895_), .Y(u0__0sp_csc_31_0__4_));
NAND2X1 NAND2X1_273 ( .A(sp_csc_5_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1897_));
NAND2X1 NAND2X1_274 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1898_), .Y(u0__abc_74894_new_n1899_));
NAND2X1 NAND2X1_275 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1900_), .Y(u0__abc_74894_new_n1901_));
NAND2X1 NAND2X1_276 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1902_));
NAND2X1 NAND2X1_277 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1903_));
NAND2X1 NAND2X1_278 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1906_));
NAND2X1 NAND2X1_279 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1909_));
NAND2X1 NAND2X1_28 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1182_));
NAND2X1 NAND2X1_280 ( .A(u0__abc_74894_new_n1897_), .B(u0__abc_74894_new_n1915_), .Y(u0__0sp_csc_31_0__5_));
NAND2X1 NAND2X1_281 ( .A(sp_csc_6_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1917_));
NAND2X1 NAND2X1_282 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1918_), .Y(u0__abc_74894_new_n1919_));
NAND2X1 NAND2X1_283 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1920_), .Y(u0__abc_74894_new_n1921_));
NAND2X1 NAND2X1_284 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1922_));
NAND2X1 NAND2X1_285 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1923_));
NAND2X1 NAND2X1_286 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1926_));
NAND2X1 NAND2X1_287 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1929_));
NAND2X1 NAND2X1_288 ( .A(u0__abc_74894_new_n1917_), .B(u0__abc_74894_new_n1935_), .Y(u0__0sp_csc_31_0__6_));
NAND2X1 NAND2X1_289 ( .A(sp_csc_7_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1937_));
NAND2X1 NAND2X1_29 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1185_));
NAND2X1 NAND2X1_290 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1938_), .Y(u0__abc_74894_new_n1939_));
NAND2X1 NAND2X1_291 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1940_), .Y(u0__abc_74894_new_n1941_));
NAND2X1 NAND2X1_292 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1942_));
NAND2X1 NAND2X1_293 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1943_));
NAND2X1 NAND2X1_294 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1946_));
NAND2X1 NAND2X1_295 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1949_));
NAND2X1 NAND2X1_296 ( .A(u0__abc_74894_new_n1937_), .B(u0__abc_74894_new_n1955_), .Y(u0__0sp_csc_31_0__7_));
NAND2X1 NAND2X1_297 ( .A(sp_csc_9_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1977_));
NAND2X1 NAND2X1_298 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1978_), .Y(u0__abc_74894_new_n1979_));
NAND2X1 NAND2X1_299 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1980_), .Y(u0__abc_74894_new_n1981_));
NAND2X1 NAND2X1_3 ( .A(u0_sreq_cs_le), .B(u0__abc_74894_new_n1104_), .Y(u0__abc_74894_new_n1107_));
NAND2X1 NAND2X1_30 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1188_));
NAND2X1 NAND2X1_300 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1982_));
NAND2X1 NAND2X1_301 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1983_));
NAND2X1 NAND2X1_302 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1986_));
NAND2X1 NAND2X1_303 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1989_));
NAND2X1 NAND2X1_304 ( .A(u0__abc_74894_new_n1977_), .B(u0__abc_74894_new_n1995_), .Y(u0__0sp_csc_31_0__9_));
NAND2X1 NAND2X1_305 ( .A(sp_csc_10_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n1997_));
NAND2X1 NAND2X1_306 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1998_), .Y(u0__abc_74894_new_n1999_));
NAND2X1 NAND2X1_307 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n2000_), .Y(u0__abc_74894_new_n2001_));
NAND2X1 NAND2X1_308 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n2002_));
NAND2X1 NAND2X1_309 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n2003_));
NAND2X1 NAND2X1_31 ( .A(u0__abc_74894_new_n1176_), .B(u0__abc_74894_new_n1194_), .Y(u0__0sp_tms_31_0__1_));
NAND2X1 NAND2X1_310 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n2006_));
NAND2X1 NAND2X1_311 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n2009_));
NAND2X1 NAND2X1_312 ( .A(u0__abc_74894_new_n1997_), .B(u0__abc_74894_new_n2015_), .Y(u0__0sp_csc_31_0__10_));
NAND2X1 NAND2X1_313 ( .A(tms_0_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2437_));
NAND2X1 NAND2X1_314 ( .A(1'h0), .B(u0__abc_74894_new_n1157_), .Y(u0__abc_74894_new_n2439_));
NAND2X1 NAND2X1_315 ( .A(1'h0), .B(u0__abc_74894_new_n1159_), .Y(u0__abc_74894_new_n2442_));
NAND2X1 NAND2X1_316 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2445_));
NAND2X1 NAND2X1_317 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2446_));
NAND2X1 NAND2X1_318 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2449_));
NAND2X1 NAND2X1_319 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2452_));
NAND2X1 NAND2X1_32 ( .A(sp_tms_2_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1196_));
NAND2X1 NAND2X1_320 ( .A(u0__abc_74894_new_n2437_), .B(u0__abc_74894_new_n2458_), .Y(u0__0tms_31_0__0_));
NAND2X1 NAND2X1_321 ( .A(tms_1_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2460_));
NAND2X1 NAND2X1_322 ( .A(1'h0), .B(u0__abc_74894_new_n1177_), .Y(u0__abc_74894_new_n2461_));
NAND2X1 NAND2X1_323 ( .A(1'h0), .B(u0__abc_74894_new_n1179_), .Y(u0__abc_74894_new_n2462_));
NAND2X1 NAND2X1_324 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2463_));
NAND2X1 NAND2X1_325 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2464_));
NAND2X1 NAND2X1_326 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2467_));
NAND2X1 NAND2X1_327 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2470_));
NAND2X1 NAND2X1_328 ( .A(u0__abc_74894_new_n2460_), .B(u0__abc_74894_new_n2474_), .Y(u0__0tms_31_0__1_));
NAND2X1 NAND2X1_329 ( .A(tms_2_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2476_));
NAND2X1 NAND2X1_33 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1197_), .Y(u0__abc_74894_new_n1198_));
NAND2X1 NAND2X1_330 ( .A(1'h0), .B(u0__abc_74894_new_n1197_), .Y(u0__abc_74894_new_n2477_));
NAND2X1 NAND2X1_331 ( .A(1'h0), .B(u0__abc_74894_new_n1199_), .Y(u0__abc_74894_new_n2478_));
NAND2X1 NAND2X1_332 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2479_));
NAND2X1 NAND2X1_333 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2480_));
NAND2X1 NAND2X1_334 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2483_));
NAND2X1 NAND2X1_335 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2486_));
NAND2X1 NAND2X1_336 ( .A(u0__abc_74894_new_n2476_), .B(u0__abc_74894_new_n2490_), .Y(u0__0tms_31_0__2_));
NAND2X1 NAND2X1_337 ( .A(tms_3_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2492_));
NAND2X1 NAND2X1_338 ( .A(1'h0), .B(u0__abc_74894_new_n1217_), .Y(u0__abc_74894_new_n2493_));
NAND2X1 NAND2X1_339 ( .A(1'h0), .B(u0__abc_74894_new_n1219_), .Y(u0__abc_74894_new_n2494_));
NAND2X1 NAND2X1_34 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1199_), .Y(u0__abc_74894_new_n1200_));
NAND2X1 NAND2X1_340 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2495_));
NAND2X1 NAND2X1_341 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2496_));
NAND2X1 NAND2X1_342 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2499_));
NAND2X1 NAND2X1_343 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2502_));
NAND2X1 NAND2X1_344 ( .A(u0__abc_74894_new_n2492_), .B(u0__abc_74894_new_n2506_), .Y(u0__0tms_31_0__3_));
NAND2X1 NAND2X1_345 ( .A(tms_4_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2508_));
NAND2X1 NAND2X1_346 ( .A(1'h0), .B(u0__abc_74894_new_n1237_), .Y(u0__abc_74894_new_n2509_));
NAND2X1 NAND2X1_347 ( .A(1'h0), .B(u0__abc_74894_new_n1239_), .Y(u0__abc_74894_new_n2510_));
NAND2X1 NAND2X1_348 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2511_));
NAND2X1 NAND2X1_349 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2512_));
NAND2X1 NAND2X1_35 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1201_));
NAND2X1 NAND2X1_350 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2515_));
NAND2X1 NAND2X1_351 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2518_));
NAND2X1 NAND2X1_352 ( .A(u0__abc_74894_new_n2508_), .B(u0__abc_74894_new_n2522_), .Y(u0__0tms_31_0__4_));
NAND2X1 NAND2X1_353 ( .A(tms_5_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2524_));
NAND2X1 NAND2X1_354 ( .A(1'h0), .B(u0__abc_74894_new_n1257_), .Y(u0__abc_74894_new_n2525_));
NAND2X1 NAND2X1_355 ( .A(1'h0), .B(u0__abc_74894_new_n1259_), .Y(u0__abc_74894_new_n2526_));
NAND2X1 NAND2X1_356 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2527_));
NAND2X1 NAND2X1_357 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2528_));
NAND2X1 NAND2X1_358 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2531_));
NAND2X1 NAND2X1_359 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2534_));
NAND2X1 NAND2X1_36 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1202_));
NAND2X1 NAND2X1_360 ( .A(u0__abc_74894_new_n2524_), .B(u0__abc_74894_new_n2538_), .Y(u0__0tms_31_0__5_));
NAND2X1 NAND2X1_361 ( .A(tms_6_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2540_));
NAND2X1 NAND2X1_362 ( .A(1'h0), .B(u0__abc_74894_new_n1277_), .Y(u0__abc_74894_new_n2541_));
NAND2X1 NAND2X1_363 ( .A(1'h0), .B(u0__abc_74894_new_n1279_), .Y(u0__abc_74894_new_n2542_));
NAND2X1 NAND2X1_364 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2543_));
NAND2X1 NAND2X1_365 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2544_));
NAND2X1 NAND2X1_366 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2547_));
NAND2X1 NAND2X1_367 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2550_));
NAND2X1 NAND2X1_368 ( .A(u0__abc_74894_new_n2540_), .B(u0__abc_74894_new_n2554_), .Y(u0__0tms_31_0__6_));
NAND2X1 NAND2X1_369 ( .A(tms_7_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2556_));
NAND2X1 NAND2X1_37 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1205_));
NAND2X1 NAND2X1_370 ( .A(1'h0), .B(u0__abc_74894_new_n1297_), .Y(u0__abc_74894_new_n2557_));
NAND2X1 NAND2X1_371 ( .A(1'h0), .B(u0__abc_74894_new_n1299_), .Y(u0__abc_74894_new_n2558_));
NAND2X1 NAND2X1_372 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2559_));
NAND2X1 NAND2X1_373 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2560_));
NAND2X1 NAND2X1_374 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2563_));
NAND2X1 NAND2X1_375 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2566_));
NAND2X1 NAND2X1_376 ( .A(u0__abc_74894_new_n2556_), .B(u0__abc_74894_new_n2570_), .Y(u0__0tms_31_0__7_));
NAND2X1 NAND2X1_377 ( .A(tms_8_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2572_));
NAND2X1 NAND2X1_378 ( .A(1'h0), .B(u0__abc_74894_new_n1317_), .Y(u0__abc_74894_new_n2573_));
NAND2X1 NAND2X1_379 ( .A(1'h0), .B(u0__abc_74894_new_n1319_), .Y(u0__abc_74894_new_n2574_));
NAND2X1 NAND2X1_38 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1208_));
NAND2X1 NAND2X1_380 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2575_));
NAND2X1 NAND2X1_381 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2576_));
NAND2X1 NAND2X1_382 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2579_));
NAND2X1 NAND2X1_383 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2582_));
NAND2X1 NAND2X1_384 ( .A(u0__abc_74894_new_n2572_), .B(u0__abc_74894_new_n2586_), .Y(u0__0tms_31_0__8_));
NAND2X1 NAND2X1_385 ( .A(tms_9_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2588_));
NAND2X1 NAND2X1_386 ( .A(1'h0), .B(u0__abc_74894_new_n1337_), .Y(u0__abc_74894_new_n2589_));
NAND2X1 NAND2X1_387 ( .A(1'h0), .B(u0__abc_74894_new_n1339_), .Y(u0__abc_74894_new_n2590_));
NAND2X1 NAND2X1_388 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2591_));
NAND2X1 NAND2X1_389 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2592_));
NAND2X1 NAND2X1_39 ( .A(u0__abc_74894_new_n1196_), .B(u0__abc_74894_new_n1214_), .Y(u0__0sp_tms_31_0__2_));
NAND2X1 NAND2X1_390 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2595_));
NAND2X1 NAND2X1_391 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2598_));
NAND2X1 NAND2X1_392 ( .A(u0__abc_74894_new_n2588_), .B(u0__abc_74894_new_n2602_), .Y(u0__0tms_31_0__9_));
NAND2X1 NAND2X1_393 ( .A(tms_10_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2604_));
NAND2X1 NAND2X1_394 ( .A(1'h0), .B(u0__abc_74894_new_n1357_), .Y(u0__abc_74894_new_n2605_));
NAND2X1 NAND2X1_395 ( .A(1'h0), .B(u0__abc_74894_new_n1359_), .Y(u0__abc_74894_new_n2606_));
NAND2X1 NAND2X1_396 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2607_));
NAND2X1 NAND2X1_397 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2608_));
NAND2X1 NAND2X1_398 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2611_));
NAND2X1 NAND2X1_399 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2614_));
NAND2X1 NAND2X1_4 ( .A(u0__abc_74894_new_n1101_), .B(u0__abc_74894_new_n1108_), .Y(u0__abc_74894_new_n1109_));
NAND2X1 NAND2X1_40 ( .A(sp_tms_3_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1216_));
NAND2X1 NAND2X1_400 ( .A(u0__abc_74894_new_n2604_), .B(u0__abc_74894_new_n2618_), .Y(u0__0tms_31_0__10_));
NAND2X1 NAND2X1_401 ( .A(tms_11_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2620_));
NAND2X1 NAND2X1_402 ( .A(1'h0), .B(u0__abc_74894_new_n1377_), .Y(u0__abc_74894_new_n2621_));
NAND2X1 NAND2X1_403 ( .A(1'h0), .B(u0__abc_74894_new_n1379_), .Y(u0__abc_74894_new_n2622_));
NAND2X1 NAND2X1_404 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2623_));
NAND2X1 NAND2X1_405 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2624_));
NAND2X1 NAND2X1_406 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2627_));
NAND2X1 NAND2X1_407 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2630_));
NAND2X1 NAND2X1_408 ( .A(u0__abc_74894_new_n2620_), .B(u0__abc_74894_new_n2634_), .Y(u0__0tms_31_0__11_));
NAND2X1 NAND2X1_409 ( .A(tms_12_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2636_));
NAND2X1 NAND2X1_41 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1217_), .Y(u0__abc_74894_new_n1218_));
NAND2X1 NAND2X1_410 ( .A(1'h0), .B(u0__abc_74894_new_n1397_), .Y(u0__abc_74894_new_n2637_));
NAND2X1 NAND2X1_411 ( .A(1'h0), .B(u0__abc_74894_new_n1399_), .Y(u0__abc_74894_new_n2638_));
NAND2X1 NAND2X1_412 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2639_));
NAND2X1 NAND2X1_413 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2640_));
NAND2X1 NAND2X1_414 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2643_));
NAND2X1 NAND2X1_415 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2646_));
NAND2X1 NAND2X1_416 ( .A(u0__abc_74894_new_n2636_), .B(u0__abc_74894_new_n2650_), .Y(u0__0tms_31_0__12_));
NAND2X1 NAND2X1_417 ( .A(tms_13_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2652_));
NAND2X1 NAND2X1_418 ( .A(1'h0), .B(u0__abc_74894_new_n1417_), .Y(u0__abc_74894_new_n2653_));
NAND2X1 NAND2X1_419 ( .A(1'h0), .B(u0__abc_74894_new_n1419_), .Y(u0__abc_74894_new_n2654_));
NAND2X1 NAND2X1_42 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1219_), .Y(u0__abc_74894_new_n1220_));
NAND2X1 NAND2X1_420 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2655_));
NAND2X1 NAND2X1_421 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2656_));
NAND2X1 NAND2X1_422 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2659_));
NAND2X1 NAND2X1_423 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2662_));
NAND2X1 NAND2X1_424 ( .A(u0__abc_74894_new_n2652_), .B(u0__abc_74894_new_n2666_), .Y(u0__0tms_31_0__13_));
NAND2X1 NAND2X1_425 ( .A(tms_14_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2668_));
NAND2X1 NAND2X1_426 ( .A(1'h0), .B(u0__abc_74894_new_n1437_), .Y(u0__abc_74894_new_n2669_));
NAND2X1 NAND2X1_427 ( .A(1'h0), .B(u0__abc_74894_new_n1439_), .Y(u0__abc_74894_new_n2670_));
NAND2X1 NAND2X1_428 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2671_));
NAND2X1 NAND2X1_429 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2672_));
NAND2X1 NAND2X1_43 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1221_));
NAND2X1 NAND2X1_430 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2675_));
NAND2X1 NAND2X1_431 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2678_));
NAND2X1 NAND2X1_432 ( .A(u0__abc_74894_new_n2668_), .B(u0__abc_74894_new_n2682_), .Y(u0__0tms_31_0__14_));
NAND2X1 NAND2X1_433 ( .A(tms_15_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2684_));
NAND2X1 NAND2X1_434 ( .A(1'h0), .B(u0__abc_74894_new_n1457_), .Y(u0__abc_74894_new_n2685_));
NAND2X1 NAND2X1_435 ( .A(1'h0), .B(u0__abc_74894_new_n1459_), .Y(u0__abc_74894_new_n2686_));
NAND2X1 NAND2X1_436 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2687_));
NAND2X1 NAND2X1_437 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2688_));
NAND2X1 NAND2X1_438 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2691_));
NAND2X1 NAND2X1_439 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2694_));
NAND2X1 NAND2X1_44 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1222_));
NAND2X1 NAND2X1_440 ( .A(u0__abc_74894_new_n2684_), .B(u0__abc_74894_new_n2698_), .Y(u0__0tms_31_0__15_));
NAND2X1 NAND2X1_441 ( .A(tms_16_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2700_));
NAND2X1 NAND2X1_442 ( .A(1'h0), .B(u0__abc_74894_new_n1477_), .Y(u0__abc_74894_new_n2701_));
NAND2X1 NAND2X1_443 ( .A(1'h0), .B(u0__abc_74894_new_n1479_), .Y(u0__abc_74894_new_n2702_));
NAND2X1 NAND2X1_444 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2703_));
NAND2X1 NAND2X1_445 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2704_));
NAND2X1 NAND2X1_446 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2707_));
NAND2X1 NAND2X1_447 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2710_));
NAND2X1 NAND2X1_448 ( .A(u0__abc_74894_new_n2700_), .B(u0__abc_74894_new_n2714_), .Y(u0__0tms_31_0__16_));
NAND2X1 NAND2X1_449 ( .A(tms_17_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2716_));
NAND2X1 NAND2X1_45 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1225_));
NAND2X1 NAND2X1_450 ( .A(1'h0), .B(u0__abc_74894_new_n1497_), .Y(u0__abc_74894_new_n2717_));
NAND2X1 NAND2X1_451 ( .A(1'h0), .B(u0__abc_74894_new_n1499_), .Y(u0__abc_74894_new_n2718_));
NAND2X1 NAND2X1_452 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2719_));
NAND2X1 NAND2X1_453 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2720_));
NAND2X1 NAND2X1_454 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2723_));
NAND2X1 NAND2X1_455 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2726_));
NAND2X1 NAND2X1_456 ( .A(u0__abc_74894_new_n2716_), .B(u0__abc_74894_new_n2730_), .Y(u0__0tms_31_0__17_));
NAND2X1 NAND2X1_457 ( .A(tms_18_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2732_));
NAND2X1 NAND2X1_458 ( .A(1'h0), .B(u0__abc_74894_new_n1517_), .Y(u0__abc_74894_new_n2733_));
NAND2X1 NAND2X1_459 ( .A(1'h0), .B(u0__abc_74894_new_n1519_), .Y(u0__abc_74894_new_n2734_));
NAND2X1 NAND2X1_46 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1228_));
NAND2X1 NAND2X1_460 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2735_));
NAND2X1 NAND2X1_461 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2736_));
NAND2X1 NAND2X1_462 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2739_));
NAND2X1 NAND2X1_463 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2742_));
NAND2X1 NAND2X1_464 ( .A(u0__abc_74894_new_n2732_), .B(u0__abc_74894_new_n2746_), .Y(u0__0tms_31_0__18_));
NAND2X1 NAND2X1_465 ( .A(tms_19_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2748_));
NAND2X1 NAND2X1_466 ( .A(1'h0), .B(u0__abc_74894_new_n1537_), .Y(u0__abc_74894_new_n2749_));
NAND2X1 NAND2X1_467 ( .A(1'h0), .B(u0__abc_74894_new_n1539_), .Y(u0__abc_74894_new_n2750_));
NAND2X1 NAND2X1_468 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2751_));
NAND2X1 NAND2X1_469 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2752_));
NAND2X1 NAND2X1_47 ( .A(u0__abc_74894_new_n1216_), .B(u0__abc_74894_new_n1234_), .Y(u0__0sp_tms_31_0__3_));
NAND2X1 NAND2X1_470 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2755_));
NAND2X1 NAND2X1_471 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2758_));
NAND2X1 NAND2X1_472 ( .A(u0__abc_74894_new_n2748_), .B(u0__abc_74894_new_n2762_), .Y(u0__0tms_31_0__19_));
NAND2X1 NAND2X1_473 ( .A(tms_20_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2764_));
NAND2X1 NAND2X1_474 ( .A(1'h0), .B(u0__abc_74894_new_n1557_), .Y(u0__abc_74894_new_n2765_));
NAND2X1 NAND2X1_475 ( .A(1'h0), .B(u0__abc_74894_new_n1559_), .Y(u0__abc_74894_new_n2766_));
NAND2X1 NAND2X1_476 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2767_));
NAND2X1 NAND2X1_477 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2768_));
NAND2X1 NAND2X1_478 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2771_));
NAND2X1 NAND2X1_479 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2774_));
NAND2X1 NAND2X1_48 ( .A(sp_tms_4_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1236_));
NAND2X1 NAND2X1_480 ( .A(u0__abc_74894_new_n2764_), .B(u0__abc_74894_new_n2778_), .Y(u0__0tms_31_0__20_));
NAND2X1 NAND2X1_481 ( .A(tms_21_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2780_));
NAND2X1 NAND2X1_482 ( .A(1'h0), .B(u0__abc_74894_new_n1577_), .Y(u0__abc_74894_new_n2781_));
NAND2X1 NAND2X1_483 ( .A(1'h0), .B(u0__abc_74894_new_n1579_), .Y(u0__abc_74894_new_n2782_));
NAND2X1 NAND2X1_484 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2783_));
NAND2X1 NAND2X1_485 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2784_));
NAND2X1 NAND2X1_486 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2787_));
NAND2X1 NAND2X1_487 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2790_));
NAND2X1 NAND2X1_488 ( .A(u0__abc_74894_new_n2780_), .B(u0__abc_74894_new_n2794_), .Y(u0__0tms_31_0__21_));
NAND2X1 NAND2X1_489 ( .A(tms_22_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2796_));
NAND2X1 NAND2X1_49 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1237_), .Y(u0__abc_74894_new_n1238_));
NAND2X1 NAND2X1_490 ( .A(1'h0), .B(u0__abc_74894_new_n1597_), .Y(u0__abc_74894_new_n2797_));
NAND2X1 NAND2X1_491 ( .A(1'h0), .B(u0__abc_74894_new_n1599_), .Y(u0__abc_74894_new_n2798_));
NAND2X1 NAND2X1_492 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2799_));
NAND2X1 NAND2X1_493 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2800_));
NAND2X1 NAND2X1_494 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2803_));
NAND2X1 NAND2X1_495 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2806_));
NAND2X1 NAND2X1_496 ( .A(u0__abc_74894_new_n2796_), .B(u0__abc_74894_new_n2810_), .Y(u0__0tms_31_0__22_));
NAND2X1 NAND2X1_497 ( .A(tms_23_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2812_));
NAND2X1 NAND2X1_498 ( .A(1'h0), .B(u0__abc_74894_new_n1617_), .Y(u0__abc_74894_new_n2813_));
NAND2X1 NAND2X1_499 ( .A(1'h0), .B(u0__abc_74894_new_n1619_), .Y(u0__abc_74894_new_n2814_));
NAND2X1 NAND2X1_5 ( .A(u0__abc_74894_new_n1101_), .B(u0__abc_74894_new_n1113_), .Y(u0__abc_74894_new_n1114_));
NAND2X1 NAND2X1_50 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1239_), .Y(u0__abc_74894_new_n1240_));
NAND2X1 NAND2X1_500 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2815_));
NAND2X1 NAND2X1_501 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2816_));
NAND2X1 NAND2X1_502 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2819_));
NAND2X1 NAND2X1_503 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2822_));
NAND2X1 NAND2X1_504 ( .A(u0__abc_74894_new_n2812_), .B(u0__abc_74894_new_n2826_), .Y(u0__0tms_31_0__23_));
NAND2X1 NAND2X1_505 ( .A(tms_24_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2828_));
NAND2X1 NAND2X1_506 ( .A(1'h0), .B(u0__abc_74894_new_n1637_), .Y(u0__abc_74894_new_n2829_));
NAND2X1 NAND2X1_507 ( .A(1'h0), .B(u0__abc_74894_new_n1639_), .Y(u0__abc_74894_new_n2830_));
NAND2X1 NAND2X1_508 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2831_));
NAND2X1 NAND2X1_509 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2832_));
NAND2X1 NAND2X1_51 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1241_));
NAND2X1 NAND2X1_510 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2835_));
NAND2X1 NAND2X1_511 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2838_));
NAND2X1 NAND2X1_512 ( .A(u0__abc_74894_new_n2828_), .B(u0__abc_74894_new_n2842_), .Y(u0__0tms_31_0__24_));
NAND2X1 NAND2X1_513 ( .A(tms_25_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2844_));
NAND2X1 NAND2X1_514 ( .A(1'h0), .B(u0__abc_74894_new_n1657_), .Y(u0__abc_74894_new_n2845_));
NAND2X1 NAND2X1_515 ( .A(1'h0), .B(u0__abc_74894_new_n1659_), .Y(u0__abc_74894_new_n2846_));
NAND2X1 NAND2X1_516 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2847_));
NAND2X1 NAND2X1_517 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2848_));
NAND2X1 NAND2X1_518 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2851_));
NAND2X1 NAND2X1_519 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2854_));
NAND2X1 NAND2X1_52 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1242_));
NAND2X1 NAND2X1_520 ( .A(u0__abc_74894_new_n2844_), .B(u0__abc_74894_new_n2858_), .Y(u0__0tms_31_0__25_));
NAND2X1 NAND2X1_521 ( .A(tms_26_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2860_));
NAND2X1 NAND2X1_522 ( .A(1'h0), .B(u0__abc_74894_new_n1677_), .Y(u0__abc_74894_new_n2861_));
NAND2X1 NAND2X1_523 ( .A(1'h0), .B(u0__abc_74894_new_n1679_), .Y(u0__abc_74894_new_n2862_));
NAND2X1 NAND2X1_524 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2863_));
NAND2X1 NAND2X1_525 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2864_));
NAND2X1 NAND2X1_526 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2867_));
NAND2X1 NAND2X1_527 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2870_));
NAND2X1 NAND2X1_528 ( .A(u0__abc_74894_new_n2860_), .B(u0__abc_74894_new_n2874_), .Y(u0__0tms_31_0__26_));
NAND2X1 NAND2X1_529 ( .A(tms_27_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n2876_));
NAND2X1 NAND2X1_53 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1245_));
NAND2X1 NAND2X1_530 ( .A(1'h0), .B(u0__abc_74894_new_n1697_), .Y(u0__abc_74894_new_n2877_));
NAND2X1 NAND2X1_531 ( .A(1'h0), .B(u0__abc_74894_new_n1699_), .Y(u0__abc_74894_new_n2878_));
NAND2X1 NAND2X1_532 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2879_));
NAND2X1 NAND2X1_533 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2880_));
NAND2X1 NAND2X1_534 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2883_));
NAND2X1 NAND2X1_535 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2886_));
NAND2X1 NAND2X1_536 ( .A(u0__abc_74894_new_n2876_), .B(u0__abc_74894_new_n2890_), .Y(u0__0tms_31_0__27_));
NAND2X1 NAND2X1_537 ( .A(csc_1_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n2973_));
NAND2X1 NAND2X1_538 ( .A(1'h0), .B(u0__abc_74894_new_n1818_), .Y(u0__abc_74894_new_n2974_));
NAND2X1 NAND2X1_539 ( .A(1'h0), .B(u0__abc_74894_new_n1820_), .Y(u0__abc_74894_new_n2975_));
NAND2X1 NAND2X1_54 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1248_));
NAND2X1 NAND2X1_540 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2976_));
NAND2X1 NAND2X1_541 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2977_));
NAND2X1 NAND2X1_542 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2980_));
NAND2X1 NAND2X1_543 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2983_));
NAND2X1 NAND2X1_544 ( .A(u0__abc_74894_new_n2983_), .B(u0__abc_74894_new_n2982_), .Y(u0__abc_74894_new_n2984_));
NAND2X1 NAND2X1_545 ( .A(csc_2_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n2989_));
NAND2X1 NAND2X1_546 ( .A(1'h0), .B(u0__abc_74894_new_n1838_), .Y(u0__abc_74894_new_n2990_));
NAND2X1 NAND2X1_547 ( .A(1'h0), .B(u0__abc_74894_new_n1840_), .Y(u0__abc_74894_new_n2991_));
NAND2X1 NAND2X1_548 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n2992_));
NAND2X1 NAND2X1_549 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2993_));
NAND2X1 NAND2X1_55 ( .A(u0__abc_74894_new_n1236_), .B(u0__abc_74894_new_n1254_), .Y(u0__0sp_tms_31_0__4_));
NAND2X1 NAND2X1_550 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2996_));
NAND2X1 NAND2X1_551 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n2999_));
NAND2X1 NAND2X1_552 ( .A(u0__abc_74894_new_n2999_), .B(u0__abc_74894_new_n2998_), .Y(u0__abc_74894_new_n3000_));
NAND2X1 NAND2X1_553 ( .A(csc_3_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n3005_));
NAND2X1 NAND2X1_554 ( .A(1'h0), .B(u0__abc_74894_new_n1858_), .Y(u0__abc_74894_new_n3006_));
NAND2X1 NAND2X1_555 ( .A(1'h0), .B(u0__abc_74894_new_n1860_), .Y(u0__abc_74894_new_n3007_));
NAND2X1 NAND2X1_556 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n3008_));
NAND2X1 NAND2X1_557 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3009_));
NAND2X1 NAND2X1_558 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3012_));
NAND2X1 NAND2X1_559 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3015_));
NAND2X1 NAND2X1_56 ( .A(sp_tms_5_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1256_));
NAND2X1 NAND2X1_560 ( .A(u0__abc_74894_new_n3015_), .B(u0__abc_74894_new_n3014_), .Y(u0__abc_74894_new_n3016_));
NAND2X1 NAND2X1_561 ( .A(csc_4_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n3021_));
NAND2X1 NAND2X1_562 ( .A(1'h0), .B(u0__abc_74894_new_n1878_), .Y(u0__abc_74894_new_n3022_));
NAND2X1 NAND2X1_563 ( .A(1'h0), .B(u0__abc_74894_new_n1880_), .Y(u0__abc_74894_new_n3023_));
NAND2X1 NAND2X1_564 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n3024_));
NAND2X1 NAND2X1_565 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3025_));
NAND2X1 NAND2X1_566 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3028_));
NAND2X1 NAND2X1_567 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3031_));
NAND2X1 NAND2X1_568 ( .A(u0__abc_74894_new_n3031_), .B(u0__abc_74894_new_n3030_), .Y(u0__abc_74894_new_n3032_));
NAND2X1 NAND2X1_569 ( .A(csc_5_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n3037_));
NAND2X1 NAND2X1_57 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1257_), .Y(u0__abc_74894_new_n1258_));
NAND2X1 NAND2X1_570 ( .A(1'h0), .B(u0__abc_74894_new_n1898_), .Y(u0__abc_74894_new_n3038_));
NAND2X1 NAND2X1_571 ( .A(1'h0), .B(u0__abc_74894_new_n1900_), .Y(u0__abc_74894_new_n3039_));
NAND2X1 NAND2X1_572 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n3040_));
NAND2X1 NAND2X1_573 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3041_));
NAND2X1 NAND2X1_574 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3044_));
NAND2X1 NAND2X1_575 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3047_));
NAND2X1 NAND2X1_576 ( .A(u0__abc_74894_new_n3047_), .B(u0__abc_74894_new_n3046_), .Y(u0__abc_74894_new_n3048_));
NAND2X1 NAND2X1_577 ( .A(csc_6_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n3053_));
NAND2X1 NAND2X1_578 ( .A(1'h0), .B(u0__abc_74894_new_n1918_), .Y(u0__abc_74894_new_n3054_));
NAND2X1 NAND2X1_579 ( .A(1'h0), .B(u0__abc_74894_new_n1920_), .Y(u0__abc_74894_new_n3055_));
NAND2X1 NAND2X1_58 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1259_), .Y(u0__abc_74894_new_n1260_));
NAND2X1 NAND2X1_580 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n3056_));
NAND2X1 NAND2X1_581 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3057_));
NAND2X1 NAND2X1_582 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3060_));
NAND2X1 NAND2X1_583 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3063_));
NAND2X1 NAND2X1_584 ( .A(u0__abc_74894_new_n3063_), .B(u0__abc_74894_new_n3062_), .Y(u0__abc_74894_new_n3064_));
NAND2X1 NAND2X1_585 ( .A(csc_7_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n3069_));
NAND2X1 NAND2X1_586 ( .A(1'h0), .B(u0__abc_74894_new_n1938_), .Y(u0__abc_74894_new_n3070_));
NAND2X1 NAND2X1_587 ( .A(1'h0), .B(u0__abc_74894_new_n1940_), .Y(u0__abc_74894_new_n3071_));
NAND2X1 NAND2X1_588 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n3072_));
NAND2X1 NAND2X1_589 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3073_));
NAND2X1 NAND2X1_59 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1261_));
NAND2X1 NAND2X1_590 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3076_));
NAND2X1 NAND2X1_591 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3079_));
NAND2X1 NAND2X1_592 ( .A(u0__abc_74894_new_n3079_), .B(u0__abc_74894_new_n3078_), .Y(u0__abc_74894_new_n3080_));
NAND2X1 NAND2X1_593 ( .A(csc_9_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n3101_));
NAND2X1 NAND2X1_594 ( .A(1'h0), .B(u0__abc_74894_new_n1978_), .Y(u0__abc_74894_new_n3102_));
NAND2X1 NAND2X1_595 ( .A(1'h0), .B(u0__abc_74894_new_n1980_), .Y(u0__abc_74894_new_n3103_));
NAND2X1 NAND2X1_596 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n3104_));
NAND2X1 NAND2X1_597 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3105_));
NAND2X1 NAND2X1_598 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3108_));
NAND2X1 NAND2X1_599 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3111_));
NAND2X1 NAND2X1_6 ( .A(u0__abc_74894_new_n1110_), .B(u0__abc_74894_new_n1116_), .Y(u0__abc_74894_new_n1117_));
NAND2X1 NAND2X1_60 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1262_));
NAND2X1 NAND2X1_600 ( .A(u0__abc_74894_new_n3111_), .B(u0__abc_74894_new_n3110_), .Y(u0__abc_74894_new_n3112_));
NAND2X1 NAND2X1_601 ( .A(csc_10_), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n3117_));
NAND2X1 NAND2X1_602 ( .A(1'h0), .B(u0__abc_74894_new_n1998_), .Y(u0__abc_74894_new_n3118_));
NAND2X1 NAND2X1_603 ( .A(1'h0), .B(u0__abc_74894_new_n2000_), .Y(u0__abc_74894_new_n3119_));
NAND2X1 NAND2X1_604 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n3120_));
NAND2X1 NAND2X1_605 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3121_));
NAND2X1 NAND2X1_606 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3124_));
NAND2X1 NAND2X1_607 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3127_));
NAND2X1 NAND2X1_608 ( .A(u0__abc_74894_new_n3127_), .B(u0__abc_74894_new_n3126_), .Y(u0__abc_74894_new_n3128_));
NAND2X1 NAND2X1_609 ( .A(u3_pen), .B(u0__abc_74894_new_n1796_), .Y(u0__abc_74894_new_n3133_));
NAND2X1 NAND2X1_61 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1265_));
NAND2X1 NAND2X1_610 ( .A(1'h0), .B(u0__abc_74894_new_n2018_), .Y(u0__abc_74894_new_n3134_));
NAND2X1 NAND2X1_611 ( .A(1'h0), .B(u0__abc_74894_new_n2020_), .Y(u0__abc_74894_new_n3135_));
NAND2X1 NAND2X1_612 ( .A(1'h0), .B(u0__abc_74894_new_n2444_), .Y(u0__abc_74894_new_n3136_));
NAND2X1 NAND2X1_613 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3137_));
NAND2X1 NAND2X1_614 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3140_));
NAND2X1 NAND2X1_615 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3143_));
NAND2X1 NAND2X1_616 ( .A(u0__abc_74894_new_n3143_), .B(u0__abc_74894_new_n3142_), .Y(u0__abc_74894_new_n3144_));
NAND2X1 NAND2X1_617 ( .A(cs_le), .B(u0__abc_74894_new_n1154_), .Y(u0__abc_74894_new_n3469_));
NAND2X1 NAND2X1_618 ( .A(wb_cyc_i), .B(u0_wp_err), .Y(u0__abc_74894_new_n3477_));
NAND2X1 NAND2X1_619 ( .A(cs_le), .B(1'h0), .Y(u0__abc_74894_new_n3494_));
NAND2X1 NAND2X1_62 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1268_));
NAND2X1 NAND2X1_620 ( .A(mc_data_ir_0_), .B(u0_rst_r3), .Y(u0__abc_74894_new_n3497_));
NAND2X1 NAND2X1_621 ( .A(u0_rst_r3), .B(mc_data_ir_1_), .Y(u0__abc_74894_new_n3500_));
NAND2X1 NAND2X1_622 ( .A(u0_rst_r3), .B(mc_data_ir_2_), .Y(u0__abc_74894_new_n3503_));
NAND2X1 NAND2X1_623 ( .A(u0_rst_r3), .B(mc_data_ir_3_), .Y(u0__abc_74894_new_n3506_));
NAND2X1 NAND2X1_624 ( .A(u0_rst_r3), .B(mc_data_ir_4_), .Y(u0__abc_74894_new_n3509_));
NAND2X1 NAND2X1_625 ( .A(u0_rst_r3), .B(mc_data_ir_5_), .Y(u0__abc_74894_new_n3512_));
NAND2X1 NAND2X1_626 ( .A(u0_rst_r3), .B(mc_data_ir_6_), .Y(u0__abc_74894_new_n3515_));
NAND2X1 NAND2X1_627 ( .A(u0_rst_r3), .B(mc_data_ir_7_), .Y(u0__abc_74894_new_n3518_));
NAND2X1 NAND2X1_628 ( .A(u0_rst_r3), .B(mc_data_ir_8_), .Y(u0__abc_74894_new_n3521_));
NAND2X1 NAND2X1_629 ( .A(u0_rst_r3), .B(mc_data_ir_9_), .Y(u0__abc_74894_new_n3524_));
NAND2X1 NAND2X1_63 ( .A(u0__abc_74894_new_n1256_), .B(u0__abc_74894_new_n1274_), .Y(u0__0sp_tms_31_0__5_));
NAND2X1 NAND2X1_630 ( .A(u0_rst_r3), .B(mc_data_ir_10_), .Y(u0__abc_74894_new_n3527_));
NAND2X1 NAND2X1_631 ( .A(u0_rst_r3), .B(mc_data_ir_11_), .Y(u0__abc_74894_new_n3530_));
NAND2X1 NAND2X1_632 ( .A(u0_rst_r3), .B(mc_data_ir_12_), .Y(u0__abc_74894_new_n3533_));
NAND2X1 NAND2X1_633 ( .A(u0_rst_r3), .B(mc_data_ir_13_), .Y(u0__abc_74894_new_n3536_));
NAND2X1 NAND2X1_634 ( .A(u0_rst_r3), .B(mc_data_ir_14_), .Y(u0__abc_74894_new_n3539_));
NAND2X1 NAND2X1_635 ( .A(u0_rst_r3), .B(mc_data_ir_15_), .Y(u0__abc_74894_new_n3542_));
NAND2X1 NAND2X1_636 ( .A(u0_rst_r3), .B(mc_data_ir_16_), .Y(u0__abc_74894_new_n3545_));
NAND2X1 NAND2X1_637 ( .A(u0_rst_r3), .B(mc_data_ir_17_), .Y(u0__abc_74894_new_n3548_));
NAND2X1 NAND2X1_638 ( .A(u0_rst_r3), .B(mc_data_ir_18_), .Y(u0__abc_74894_new_n3551_));
NAND2X1 NAND2X1_639 ( .A(u0_rst_r3), .B(mc_data_ir_19_), .Y(u0__abc_74894_new_n3554_));
NAND2X1 NAND2X1_64 ( .A(sp_tms_6_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1276_));
NAND2X1 NAND2X1_640 ( .A(u0_rst_r3), .B(mc_data_ir_20_), .Y(u0__abc_74894_new_n3557_));
NAND2X1 NAND2X1_641 ( .A(u0_rst_r3), .B(mc_data_ir_21_), .Y(u0__abc_74894_new_n3560_));
NAND2X1 NAND2X1_642 ( .A(u0_rst_r3), .B(mc_data_ir_22_), .Y(u0__abc_74894_new_n3563_));
NAND2X1 NAND2X1_643 ( .A(u0_rst_r3), .B(mc_data_ir_23_), .Y(u0__abc_74894_new_n3566_));
NAND2X1 NAND2X1_644 ( .A(u0_rst_r3), .B(mc_data_ir_24_), .Y(u0__abc_74894_new_n3569_));
NAND2X1 NAND2X1_645 ( .A(u0_rst_r3), .B(mc_data_ir_25_), .Y(u0__abc_74894_new_n3572_));
NAND2X1 NAND2X1_646 ( .A(u0_rst_r3), .B(mc_data_ir_26_), .Y(u0__abc_74894_new_n3575_));
NAND2X1 NAND2X1_647 ( .A(u0_rst_r3), .B(mc_data_ir_27_), .Y(u0__abc_74894_new_n3578_));
NAND2X1 NAND2X1_648 ( .A(u0_rst_r3), .B(mc_data_ir_28_), .Y(u0__abc_74894_new_n3581_));
NAND2X1 NAND2X1_649 ( .A(u0_rst_r3), .B(mc_data_ir_29_), .Y(u0__abc_74894_new_n3584_));
NAND2X1 NAND2X1_65 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1277_), .Y(u0__abc_74894_new_n1278_));
NAND2X1 NAND2X1_650 ( .A(u0_rst_r3), .B(mc_data_ir_30_), .Y(u0__abc_74894_new_n3587_));
NAND2X1 NAND2X1_651 ( .A(u0_rst_r3), .B(mc_data_ir_31_), .Y(u0__abc_74894_new_n3590_));
NAND2X1 NAND2X1_652 ( .A(u0__abc_74894_new_n3593_), .B(u0__abc_74894_new_n3594_), .Y(u0__abc_74894_new_n3595_));
NAND2X1 NAND2X1_653 ( .A(\wb_data_i[0] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3599_));
NAND2X1 NAND2X1_654 ( .A(\wb_data_i[1] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3602_));
NAND2X1 NAND2X1_655 ( .A(\wb_data_i[2] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3605_));
NAND2X1 NAND2X1_656 ( .A(\wb_data_i[3] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3608_));
NAND2X1 NAND2X1_657 ( .A(\wb_data_i[4] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3611_));
NAND2X1 NAND2X1_658 ( .A(\wb_data_i[5] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3614_));
NAND2X1 NAND2X1_659 ( .A(\wb_data_i[6] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3617_));
NAND2X1 NAND2X1_66 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1279_), .Y(u0__abc_74894_new_n1280_));
NAND2X1 NAND2X1_660 ( .A(\wb_data_i[7] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3620_));
NAND2X1 NAND2X1_661 ( .A(\wb_data_i[8] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3623_));
NAND2X1 NAND2X1_662 ( .A(\wb_data_i[9] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3626_));
NAND2X1 NAND2X1_663 ( .A(\wb_data_i[10] ), .B(u0__abc_74894_new_n3598_), .Y(u0__abc_74894_new_n3629_));
NAND2X1 NAND2X1_664 ( .A(\wb_data_i[1] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3635_));
NAND2X1 NAND2X1_665 ( .A(\wb_data_i[2] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3638_));
NAND2X1 NAND2X1_666 ( .A(\wb_data_i[3] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3641_));
NAND2X1 NAND2X1_667 ( .A(\wb_data_i[4] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3644_));
NAND2X1 NAND2X1_668 ( .A(\wb_data_i[5] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3647_));
NAND2X1 NAND2X1_669 ( .A(\wb_data_i[6] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3650_));
NAND2X1 NAND2X1_67 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1281_));
NAND2X1 NAND2X1_670 ( .A(\wb_data_i[7] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3653_));
NAND2X1 NAND2X1_671 ( .A(\wb_data_i[8] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3656_));
NAND2X1 NAND2X1_672 ( .A(\wb_data_i[9] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3659_));
NAND2X1 NAND2X1_673 ( .A(\wb_data_i[10] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3662_));
NAND2X1 NAND2X1_674 ( .A(\wb_data_i[24] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3665_));
NAND2X1 NAND2X1_675 ( .A(\wb_data_i[25] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3668_));
NAND2X1 NAND2X1_676 ( .A(\wb_data_i[26] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3671_));
NAND2X1 NAND2X1_677 ( .A(\wb_data_i[27] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3674_));
NAND2X1 NAND2X1_678 ( .A(\wb_data_i[28] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3677_));
NAND2X1 NAND2X1_679 ( .A(\wb_data_i[29] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3680_));
NAND2X1 NAND2X1_68 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1282_));
NAND2X1 NAND2X1_680 ( .A(\wb_data_i[30] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3683_));
NAND2X1 NAND2X1_681 ( .A(\wb_data_i[31] ), .B(u0__abc_74894_new_n3634_), .Y(u0__abc_74894_new_n3686_));
NAND2X1 NAND2X1_682 ( .A(\wb_addr_i[6] ), .B(u0__abc_74894_new_n3688_), .Y(u0__abc_74894_new_n3689_));
NAND2X1 NAND2X1_683 ( .A(u0__abc_74894_new_n3690_), .B(u0__abc_74894_new_n3691_), .Y(u0__abc_74894_new_n3692_));
NAND2X1 NAND2X1_684 ( .A(1'h0), .B(u0__abc_74894_new_n3693_), .Y(u0__abc_74894_new_n3694_));
NAND2X1 NAND2X1_685 ( .A(\wb_addr_i[2] ), .B(u0__abc_74894_new_n3690_), .Y(u0__abc_74894_new_n3695_));
NAND2X1 NAND2X1_686 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n3697_));
NAND2X1 NAND2X1_687 ( .A(\wb_addr_i[3] ), .B(\wb_addr_i[2] ), .Y(u0__abc_74894_new_n3698_));
NAND2X1 NAND2X1_688 ( .A(\wb_addr_i[3] ), .B(u0__abc_74894_new_n3691_), .Y(u0__abc_74894_new_n3700_));
NAND2X1 NAND2X1_689 ( .A(u0__abc_74894_new_n3705_), .B(u0__abc_74894_new_n3706_), .Y(u0__abc_74894_new_n3707_));
NAND2X1 NAND2X1_69 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1285_));
NAND2X1 NAND2X1_690 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n3709_));
NAND2X1 NAND2X1_691 ( .A(u0__abc_74894_new_n3705_), .B(u0__abc_74894_new_n3715_), .Y(u0__abc_74894_new_n3716_));
NAND2X1 NAND2X1_692 ( .A(u0__abc_74894_new_n3718_), .B(u0__abc_74894_new_n3715_), .Y(u0__abc_74894_new_n3719_));
NAND2X1 NAND2X1_693 ( .A(\wb_addr_i[4] ), .B(u0__abc_74894_new_n3704_), .Y(u0__abc_74894_new_n3730_));
NAND2X1 NAND2X1_694 ( .A(u0__abc_74894_new_n3726_), .B(u0__abc_74894_new_n3731_), .Y(u0__abc_74894_new_n3733_));
NAND2X1 NAND2X1_695 ( .A(u0__abc_74894_new_n3735_), .B(u0__abc_74894_new_n3731_), .Y(u0__abc_74894_new_n3736_));
NAND2X1 NAND2X1_696 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n3742_));
NAND2X1 NAND2X1_697 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3744_));
NAND2X1 NAND2X1_698 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3746_));
NAND2X1 NAND2X1_699 ( .A(u0__abc_74894_new_n3725_), .B(u0__abc_74894_new_n3731_), .Y(u0__abc_74894_new_n3748_));
NAND2X1 NAND2X1_7 ( .A(init_req), .B(1'h0), .Y(u0__abc_74894_new_n1121_));
NAND2X1 NAND2X1_70 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1288_));
NAND2X1 NAND2X1_700 ( .A(u0__abc_74894_new_n3688_), .B(u0__abc_74894_new_n3712_), .Y(u0__abc_74894_new_n3750_));
NAND2X1 NAND2X1_701 ( .A(u0__abc_74894_new_n3756_), .B(u0__abc_74894_new_n3757_), .Y(u0__abc_74894_new_n3758_));
NAND2X1 NAND2X1_702 ( .A(u0__abc_74894_new_n3760_), .B(u0__abc_74894_new_n3759_), .Y(u0__abc_74894_new_n3761_));
NAND2X1 NAND2X1_703 ( .A(u0__abc_74894_new_n3705_), .B(u0__abc_74894_new_n3710_), .Y(u0__abc_74894_new_n3765_));
NAND2X1 NAND2X1_704 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n3766_));
NAND2X1 NAND2X1_705 ( .A(u0__abc_74894_new_n3778_), .B(u0__abc_74894_new_n3779_), .Y(u0__abc_74894_new_n3780_));
NAND2X1 NAND2X1_706 ( .A(u0__abc_74894_new_n3782_), .B(u0__abc_74894_new_n3781_), .Y(u0__abc_74894_new_n3783_));
NAND2X1 NAND2X1_707 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n3786_));
NAND2X1 NAND2X1_708 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3799_));
NAND2X1 NAND2X1_709 ( .A(u0__abc_74894_new_n3803_), .B(u0__abc_74894_new_n3801_), .Y(u0__abc_74894_new_n3804_));
NAND2X1 NAND2X1_71 ( .A(u0__abc_74894_new_n1276_), .B(u0__abc_74894_new_n1294_), .Y(u0__0sp_tms_31_0__6_));
NAND2X1 NAND2X1_710 ( .A(\poc_o[3] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3806_));
NAND2X1 NAND2X1_711 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n3807_));
NAND2X1 NAND2X1_712 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3811_));
NAND2X1 NAND2X1_713 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3812_));
NAND2X1 NAND2X1_714 ( .A(u0__abc_74894_new_n3818_), .B(u0__abc_74894_new_n3817_), .Y(u0__abc_74894_new_n3819_));
NAND2X1 NAND2X1_715 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3822_));
NAND2X1 NAND2X1_716 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3823_));
NAND2X1 NAND2X1_717 ( .A(u0__abc_74894_new_n3827_), .B(u0__abc_74894_new_n3826_), .Y(u0__abc_74894_new_n3828_));
NAND2X1 NAND2X1_718 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3841_));
NAND2X1 NAND2X1_719 ( .A(1'h0), .B(u0__abc_74894_new_n3693_), .Y(u0__abc_74894_new_n3843_));
NAND2X1 NAND2X1_72 ( .A(sp_tms_7_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1296_));
NAND2X1 NAND2X1_720 ( .A(u0__abc_74894_new_n3688_), .B(u0__abc_74894_new_n3706_), .Y(u0__abc_74894_new_n3845_));
NAND2X1 NAND2X1_721 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3846_));
NAND2X1 NAND2X1_722 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3849_));
NAND2X1 NAND2X1_723 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3850_));
NAND2X1 NAND2X1_724 ( .A(u0_tms0_5_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n3854_));
NAND2X1 NAND2X1_725 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .Y(u0__abc_74894_new_n3855_));
NAND2X1 NAND2X1_726 ( .A(u0__abc_74894_new_n3858_), .B(u0__abc_74894_new_n3859_), .Y(u0__abc_74894_new_n3860_));
NAND2X1 NAND2X1_727 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3863_));
NAND2X1 NAND2X1_728 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3864_));
NAND2X1 NAND2X1_729 ( .A(u0__abc_74894_new_n3868_), .B(u0__abc_74894_new_n3867_), .Y(u0__abc_74894_new_n3869_));
NAND2X1 NAND2X1_73 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1297_), .Y(u0__abc_74894_new_n1298_));
NAND2X1 NAND2X1_730 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n3885_));
NAND2X1 NAND2X1_731 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n3886_));
NAND2X1 NAND2X1_732 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3887_));
NAND2X1 NAND2X1_733 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3893_));
NAND2X1 NAND2X1_734 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3900_));
NAND2X1 NAND2X1_735 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3901_));
NAND2X1 NAND2X1_736 ( .A(u0__abc_74894_new_n3905_), .B(u0__abc_74894_new_n3904_), .Y(u0__abc_74894_new_n3906_));
NAND2X1 NAND2X1_737 ( .A(ref_int_0_), .B(u0__abc_74894_new_n3729_), .Y(u0__abc_74894_new_n3911_));
NAND2X1 NAND2X1_738 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3919_));
NAND2X1 NAND2X1_739 ( .A(u0__abc_74894_new_n3921_), .B(u0__abc_74894_new_n3922_), .Y(u0__abc_74894_new_n3923_));
NAND2X1 NAND2X1_74 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1299_), .Y(u0__abc_74894_new_n1300_));
NAND2X1 NAND2X1_740 ( .A(u0_csc_mask_9_), .B(u0__abc_74894_new_n3749_), .Y(u0__abc_74894_new_n3925_));
NAND2X1 NAND2X1_741 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n3926_));
NAND2X1 NAND2X1_742 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n3930_));
NAND2X1 NAND2X1_743 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3931_));
NAND2X1 NAND2X1_744 ( .A(u0__abc_74894_new_n3935_), .B(u0__abc_74894_new_n3934_), .Y(u0__abc_74894_new_n3936_));
NAND2X1 NAND2X1_745 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3939_));
NAND2X1 NAND2X1_746 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3940_));
NAND2X1 NAND2X1_747 ( .A(u0__abc_74894_new_n3944_), .B(u0__abc_74894_new_n3943_), .Y(u0__abc_74894_new_n3945_));
NAND2X1 NAND2X1_748 ( .A(\poc_o[11] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3957_));
NAND2X1 NAND2X1_749 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3958_));
NAND2X1 NAND2X1_75 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1301_));
NAND2X1 NAND2X1_750 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3959_));
NAND2X1 NAND2X1_751 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3962_));
NAND2X1 NAND2X1_752 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n3963_));
NAND2X1 NAND2X1_753 ( .A(u0__abc_74894_new_n3968_), .B(u0__abc_74894_new_n3967_), .Y(u0__abc_74894_new_n3969_));
NAND2X1 NAND2X1_754 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3970_));
NAND2X1 NAND2X1_755 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n3971_));
NAND2X1 NAND2X1_756 ( .A(\poc_o[12] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n3976_));
NAND2X1 NAND2X1_757 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n3977_));
NAND2X1 NAND2X1_758 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n3978_));
NAND2X1 NAND2X1_759 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3981_));
NAND2X1 NAND2X1_76 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1302_));
NAND2X1 NAND2X1_760 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n3982_));
NAND2X1 NAND2X1_761 ( .A(u0__abc_74894_new_n3987_), .B(u0__abc_74894_new_n3986_), .Y(u0__abc_74894_new_n3988_));
NAND2X1 NAND2X1_762 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n3989_));
NAND2X1 NAND2X1_763 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n3990_));
NAND2X1 NAND2X1_764 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n3995_));
NAND2X1 NAND2X1_765 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n3996_));
NAND2X1 NAND2X1_766 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n3997_));
NAND2X1 NAND2X1_767 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4002_));
NAND2X1 NAND2X1_768 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4005_));
NAND2X1 NAND2X1_769 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4011_));
NAND2X1 NAND2X1_77 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1305_));
NAND2X1 NAND2X1_770 ( .A(u0_tms0_13_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4012_));
NAND2X1 NAND2X1_771 ( .A(u0_csc1_13_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4013_));
NAND2X1 NAND2X1_772 ( .A(u0_csc0_14_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4017_));
NAND2X1 NAND2X1_773 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4018_));
NAND2X1 NAND2X1_774 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4019_));
NAND2X1 NAND2X1_775 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4024_));
NAND2X1 NAND2X1_776 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4027_));
NAND2X1 NAND2X1_777 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4033_));
NAND2X1 NAND2X1_778 ( .A(u0_tms0_14_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4034_));
NAND2X1 NAND2X1_779 ( .A(u0_csc1_14_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4035_));
NAND2X1 NAND2X1_78 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1308_));
NAND2X1 NAND2X1_780 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4039_));
NAND2X1 NAND2X1_781 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4043_));
NAND2X1 NAND2X1_782 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4047_));
NAND2X1 NAND2X1_783 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4048_));
NAND2X1 NAND2X1_784 ( .A(u0_csc0_15_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4049_));
NAND2X1 NAND2X1_785 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4053_));
NAND2X1 NAND2X1_786 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4056_));
NAND2X1 NAND2X1_787 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4061_));
NAND2X1 NAND2X1_788 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4064_));
NAND2X1 NAND2X1_789 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4065_));
NAND2X1 NAND2X1_79 ( .A(u0__abc_74894_new_n1296_), .B(u0__abc_74894_new_n1314_), .Y(u0__0sp_tms_31_0__7_));
NAND2X1 NAND2X1_790 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4068_));
NAND2X1 NAND2X1_791 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4072_));
NAND2X1 NAND2X1_792 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .Y(u0__abc_74894_new_n4073_));
NAND2X1 NAND2X1_793 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4076_));
NAND2X1 NAND2X1_794 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4077_));
NAND2X1 NAND2X1_795 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4081_));
NAND2X1 NAND2X1_796 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4085_));
NAND2X1 NAND2X1_797 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4089_));
NAND2X1 NAND2X1_798 ( .A(u0_csc0_17_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4090_));
NAND2X1 NAND2X1_799 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4091_));
NAND2X1 NAND2X1_8 ( .A(u0__abc_74894_new_n1122_), .B(u0__abc_74894_new_n1115_), .Y(u0__abc_74894_new_n1123_));
NAND2X1 NAND2X1_80 ( .A(sp_tms_8_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1316_));
NAND2X1 NAND2X1_800 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4095_));
NAND2X1 NAND2X1_801 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4098_));
NAND2X1 NAND2X1_802 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4103_));
NAND2X1 NAND2X1_803 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4107_));
NAND2X1 NAND2X1_804 ( .A(u0_csc0_18_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4111_));
NAND2X1 NAND2X1_805 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4112_));
NAND2X1 NAND2X1_806 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4113_));
NAND2X1 NAND2X1_807 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4117_));
NAND2X1 NAND2X1_808 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4120_));
NAND2X1 NAND2X1_809 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4125_));
NAND2X1 NAND2X1_81 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1317_), .Y(u0__abc_74894_new_n1318_));
NAND2X1 NAND2X1_810 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4126_));
NAND2X1 NAND2X1_811 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4127_));
NAND2X1 NAND2X1_812 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4132_));
NAND2X1 NAND2X1_813 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4135_));
NAND2X1 NAND2X1_814 ( .A(u0_csc1_19_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4141_));
NAND2X1 NAND2X1_815 ( .A(u0_tms0_19_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4142_));
NAND2X1 NAND2X1_816 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4143_));
NAND2X1 NAND2X1_817 ( .A(\poc_o[20] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4147_));
NAND2X1 NAND2X1_818 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4148_));
NAND2X1 NAND2X1_819 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4149_));
NAND2X1 NAND2X1_82 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1319_), .Y(u0__abc_74894_new_n1320_));
NAND2X1 NAND2X1_820 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4152_));
NAND2X1 NAND2X1_821 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4153_));
NAND2X1 NAND2X1_822 ( .A(u0__abc_74894_new_n4158_), .B(u0__abc_74894_new_n4157_), .Y(u0__abc_74894_new_n4159_));
NAND2X1 NAND2X1_823 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4160_));
NAND2X1 NAND2X1_824 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4161_));
NAND2X1 NAND2X1_825 ( .A(u0_csc0_21_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4166_));
NAND2X1 NAND2X1_826 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4167_));
NAND2X1 NAND2X1_827 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4168_));
NAND2X1 NAND2X1_828 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4170_));
NAND2X1 NAND2X1_829 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4174_));
NAND2X1 NAND2X1_83 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1321_));
NAND2X1 NAND2X1_830 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4177_));
NAND2X1 NAND2X1_831 ( .A(u0_tms1_21_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4183_));
NAND2X1 NAND2X1_832 ( .A(u0_tms0_21_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4184_));
NAND2X1 NAND2X1_833 ( .A(u0_csc1_21_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4185_));
NAND2X1 NAND2X1_834 ( .A(\poc_o[22] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4189_));
NAND2X1 NAND2X1_835 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4190_));
NAND2X1 NAND2X1_836 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4191_));
NAND2X1 NAND2X1_837 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4194_));
NAND2X1 NAND2X1_838 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4195_));
NAND2X1 NAND2X1_839 ( .A(u0__abc_74894_new_n4200_), .B(u0__abc_74894_new_n4199_), .Y(u0__abc_74894_new_n4201_));
NAND2X1 NAND2X1_84 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1322_));
NAND2X1 NAND2X1_840 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4202_));
NAND2X1 NAND2X1_841 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4203_));
NAND2X1 NAND2X1_842 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4208_));
NAND2X1 NAND2X1_843 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4211_));
NAND2X1 NAND2X1_844 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4212_));
NAND2X1 NAND2X1_845 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4215_));
NAND2X1 NAND2X1_846 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4219_));
NAND2X1 NAND2X1_847 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .Y(u0__abc_74894_new_n4220_));
NAND2X1 NAND2X1_848 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4223_));
NAND2X1 NAND2X1_849 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4224_));
NAND2X1 NAND2X1_85 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1325_));
NAND2X1 NAND2X1_850 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4228_));
NAND2X1 NAND2X1_851 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4229_));
NAND2X1 NAND2X1_852 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4230_));
NAND2X1 NAND2X1_853 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4232_));
NAND2X1 NAND2X1_854 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4233_));
NAND2X1 NAND2X1_855 ( .A(1'h0), .B(u0__abc_74894_new_n3693_), .Y(u0__abc_74894_new_n4234_));
NAND2X1 NAND2X1_856 ( .A(u0_csc1_24_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4237_));
NAND2X1 NAND2X1_857 ( .A(u0_tms0_24_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4238_));
NAND2X1 NAND2X1_858 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4239_));
NAND2X1 NAND2X1_859 ( .A(u0_tms1_24_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4242_));
NAND2X1 NAND2X1_86 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1328_));
NAND2X1 NAND2X1_860 ( .A(\poc_o[24] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4243_));
NAND2X1 NAND2X1_861 ( .A(u0_csc0_24_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4244_));
NAND2X1 NAND2X1_862 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4246_));
NAND2X1 NAND2X1_863 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4247_));
NAND2X1 NAND2X1_864 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4248_));
NAND2X1 NAND2X1_865 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4250_));
NAND2X1 NAND2X1_866 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4254_));
NAND2X1 NAND2X1_867 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4255_));
NAND2X1 NAND2X1_868 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4256_));
NAND2X1 NAND2X1_869 ( .A(1'h0), .B(u0__abc_74894_new_n3693_), .Y(u0__abc_74894_new_n4258_));
NAND2X1 NAND2X1_87 ( .A(u0__abc_74894_new_n1316_), .B(u0__abc_74894_new_n1334_), .Y(u0__0sp_tms_31_0__8_));
NAND2X1 NAND2X1_870 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4259_));
NAND2X1 NAND2X1_871 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4260_));
NAND2X1 NAND2X1_872 ( .A(u0_tms1_25_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4263_));
NAND2X1 NAND2X1_873 ( .A(u0_tms0_25_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4264_));
NAND2X1 NAND2X1_874 ( .A(u0_csc1_25_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4265_));
NAND2X1 NAND2X1_875 ( .A(\poc_o[25] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4268_));
NAND2X1 NAND2X1_876 ( .A(u0_csc0_25_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4269_));
NAND2X1 NAND2X1_877 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4270_));
NAND2X1 NAND2X1_878 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4276_));
NAND2X1 NAND2X1_879 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4280_));
NAND2X1 NAND2X1_88 ( .A(sp_tms_9_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1336_));
NAND2X1 NAND2X1_880 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4281_));
NAND2X1 NAND2X1_881 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4282_));
NAND2X1 NAND2X1_882 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4284_));
NAND2X1 NAND2X1_883 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4285_));
NAND2X1 NAND2X1_884 ( .A(1'h0), .B(u0__abc_74894_new_n3693_), .Y(u0__abc_74894_new_n4286_));
NAND2X1 NAND2X1_885 ( .A(u0_tms0_26_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4289_));
NAND2X1 NAND2X1_886 ( .A(u0_csc1_26_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4290_));
NAND2X1 NAND2X1_887 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4291_));
NAND2X1 NAND2X1_888 ( .A(u0_tms1_26_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4294_));
NAND2X1 NAND2X1_889 ( .A(\poc_o[26] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4295_));
NAND2X1 NAND2X1_89 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1337_), .Y(u0__abc_74894_new_n1338_));
NAND2X1 NAND2X1_890 ( .A(u0_csc0_26_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4296_));
NAND2X1 NAND2X1_891 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4298_));
NAND2X1 NAND2X1_892 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4299_));
NAND2X1 NAND2X1_893 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4300_));
NAND2X1 NAND2X1_894 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4302_));
NAND2X1 NAND2X1_895 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4306_));
NAND2X1 NAND2X1_896 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4307_));
NAND2X1 NAND2X1_897 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4308_));
NAND2X1 NAND2X1_898 ( .A(1'h0), .B(u0__abc_74894_new_n3693_), .Y(u0__abc_74894_new_n4310_));
NAND2X1 NAND2X1_899 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4311_));
NAND2X1 NAND2X1_9 ( .A(init_req), .B(1'h0), .Y(u0__abc_74894_new_n1127_));
NAND2X1 NAND2X1_90 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1339_), .Y(u0__abc_74894_new_n1340_));
NAND2X1 NAND2X1_900 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4312_));
NAND2X1 NAND2X1_901 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4315_));
NAND2X1 NAND2X1_902 ( .A(u0_tms0_27_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4316_));
NAND2X1 NAND2X1_903 ( .A(u0_csc1_27_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4317_));
NAND2X1 NAND2X1_904 ( .A(u0_tms1_27_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4320_));
NAND2X1 NAND2X1_905 ( .A(\poc_o[27] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4321_));
NAND2X1 NAND2X1_906 ( .A(u0_csc0_27_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4322_));
NAND2X1 NAND2X1_907 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4324_));
NAND2X1 NAND2X1_908 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .Y(u0__abc_74894_new_n4325_));
NAND2X1 NAND2X1_909 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4326_));
NAND2X1 NAND2X1_91 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1341_));
NAND2X1 NAND2X1_910 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4329_));
NAND2X1 NAND2X1_911 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4333_));
NAND2X1 NAND2X1_912 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4334_));
NAND2X1 NAND2X1_913 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4335_));
NAND2X1 NAND2X1_914 ( .A(1'h0), .B(u0__abc_74894_new_n3699_), .Y(u0__abc_74894_new_n4337_));
NAND2X1 NAND2X1_915 ( .A(1'h0), .B(u0__abc_74894_new_n3745_), .Y(u0__abc_74894_new_n4338_));
NAND2X1 NAND2X1_916 ( .A(1'h0), .B(u0__abc_74894_new_n3693_), .Y(u0__abc_74894_new_n4339_));
NAND2X1 NAND2X1_917 ( .A(u0_tms0_28_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4342_));
NAND2X1 NAND2X1_918 ( .A(u0_csc1_28_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4343_));
NAND2X1 NAND2X1_919 ( .A(u0_tms1_28_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4344_));
NAND2X1 NAND2X1_92 ( .A(spec_req_cs_6_), .B(1'h0), .Y(u0__abc_74894_new_n1342_));
NAND2X1 NAND2X1_920 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4347_));
NAND2X1 NAND2X1_921 ( .A(\poc_o[28] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4348_));
NAND2X1 NAND2X1_922 ( .A(u0_csc0_28_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4349_));
NAND2X1 NAND2X1_923 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4351_));
NAND2X1 NAND2X1_924 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4352_));
NAND2X1 NAND2X1_925 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4353_));
NAND2X1 NAND2X1_926 ( .A(1'h0), .B(u0__abc_74894_new_n3696_), .Y(u0__abc_74894_new_n4355_));
NAND2X1 NAND2X1_927 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4359_));
NAND2X1 NAND2X1_928 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4360_));
NAND2X1 NAND2X1_929 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4361_));
NAND2X1 NAND2X1_93 ( .A(spec_req_cs_4_), .B(1'h0), .Y(u0__abc_74894_new_n1345_));
NAND2X1 NAND2X1_930 ( .A(u0__abc_74894_new_n4363_), .B(u0__abc_74894_new_n4364_), .Y(u0__abc_74894_new_n4365_));
NAND2X1 NAND2X1_931 ( .A(u0_tms0_29_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4367_));
NAND2X1 NAND2X1_932 ( .A(u0_csc1_29_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4368_));
NAND2X1 NAND2X1_933 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4369_));
NAND2X1 NAND2X1_934 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4373_));
NAND2X1 NAND2X1_935 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4374_));
NAND2X1 NAND2X1_936 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4375_));
NAND2X1 NAND2X1_937 ( .A(u0_csc0_29_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4377_));
NAND2X1 NAND2X1_938 ( .A(\poc_o[29] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4378_));
NAND2X1 NAND2X1_939 ( .A(u0_tms1_29_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4379_));
NAND2X1 NAND2X1_94 ( .A(spec_req_cs_2_), .B(1'h0), .Y(u0__abc_74894_new_n1348_));
NAND2X1 NAND2X1_940 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4383_));
NAND2X1 NAND2X1_941 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4384_));
NAND2X1 NAND2X1_942 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4385_));
NAND2X1 NAND2X1_943 ( .A(u0__abc_74894_new_n4387_), .B(u0__abc_74894_new_n4388_), .Y(u0__abc_74894_new_n4389_));
NAND2X1 NAND2X1_944 ( .A(u0_tms0_30_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4391_));
NAND2X1 NAND2X1_945 ( .A(u0_csc1_30_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4392_));
NAND2X1 NAND2X1_946 ( .A(u0_tms1_30_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4393_));
NAND2X1 NAND2X1_947 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4397_));
NAND2X1 NAND2X1_948 ( .A(1'h0), .B(u0__abc_74894_new_n3701_), .Y(u0__abc_74894_new_n4398_));
NAND2X1 NAND2X1_949 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4399_));
NAND2X1 NAND2X1_95 ( .A(u0__abc_74894_new_n1336_), .B(u0__abc_74894_new_n1354_), .Y(u0__0sp_tms_31_0__9_));
NAND2X1 NAND2X1_950 ( .A(u0_csc0_30_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4401_));
NAND2X1 NAND2X1_951 ( .A(\poc_o[30] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4402_));
NAND2X1 NAND2X1_952 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4403_));
NAND2X1 NAND2X1_953 ( .A(1'h0), .B(u0__abc_74894_new_n3741_), .Y(u0__abc_74894_new_n4407_));
NAND2X1 NAND2X1_954 ( .A(1'h0), .B(u0__abc_74894_new_n3720_), .Y(u0__abc_74894_new_n4408_));
NAND2X1 NAND2X1_955 ( .A(1'h0), .B(u0__abc_74894_new_n3743_), .Y(u0__abc_74894_new_n4409_));
NAND2X1 NAND2X1_956 ( .A(u0__abc_74894_new_n4411_), .B(u0__abc_74894_new_n4412_), .Y(u0__abc_74894_new_n4413_));
NAND2X1 NAND2X1_957 ( .A(u0_tms0_31_), .B(u0__abc_74894_new_n3737_), .Y(u0__abc_74894_new_n4415_));
NAND2X1 NAND2X1_958 ( .A(u0_csc1_31_), .B(u0__abc_74894_new_n3816_), .Y(u0__abc_74894_new_n4416_));
NAND2X1 NAND2X1_959 ( .A(u0_tms1_31_), .B(u0__abc_74894_new_n3802_), .Y(u0__abc_74894_new_n4417_));
NAND2X1 NAND2X1_96 ( .A(sp_tms_10_), .B(u0__abc_74894_new_n1155_), .Y(u0__abc_74894_new_n1356_));
NAND2X1 NAND2X1_960 ( .A(1'h0), .B(u0__abc_74894_new_n3708_), .Y(u0__abc_74894_new_n4421_));
NAND2X1 NAND2X1_961 ( .A(1'h0), .B(u0__abc_74894_new_n3717_), .Y(u0__abc_74894_new_n4422_));
NAND2X1 NAND2X1_962 ( .A(1'h0), .B(u0__abc_74894_new_n3713_), .Y(u0__abc_74894_new_n4423_));
NAND2X1 NAND2X1_963 ( .A(u0_csc0_31_), .B(u0__abc_74894_new_n3734_), .Y(u0__abc_74894_new_n4425_));
NAND2X1 NAND2X1_964 ( .A(\poc_o[31] ), .B(u0__abc_74894_new_n3751_), .Y(u0__abc_74894_new_n4426_));
NAND2X1 NAND2X1_965 ( .A(1'h0), .B(u0__abc_74894_new_n3711_), .Y(u0__abc_74894_new_n4427_));
NAND2X1 NAND2X1_966 ( .A(\wb_addr_i[30] ), .B(\wb_addr_i[29] ), .Y(u0__abc_74894_new_n4431_));
NAND2X1 NAND2X1_967 ( .A(u0__abc_74894_new_n1833_), .B(u0__abc_74894_new_n1853_), .Y(u0__abc_74894_new_n4437_));
NAND2X1 NAND2X1_968 ( .A(u0_csc0_0_), .B(u0__abc_74894_new_n1873_), .Y(u0__abc_74894_new_n4438_));
NAND2X1 NAND2X1_969 ( .A(u0__abc_74894_new_n1831_), .B(u0__abc_74894_new_n1851_), .Y(u0__abc_74894_new_n4440_));
NAND2X1 NAND2X1_97 ( .A(spec_req_cs_3_), .B(u0__abc_74894_new_n1357_), .Y(u0__abc_74894_new_n1358_));
NAND2X1 NAND2X1_970 ( .A(u0_csc1_0_), .B(u0__abc_74894_new_n1871_), .Y(u0__abc_74894_new_n4441_));
NAND2X1 NAND2X1_971 ( .A(u0__abc_74894_new_n3764_), .B(u0__abc_74894_new_n3785_), .Y(u0__abc_74894_new_n4443_));
NAND2X1 NAND2X1_972 ( .A(u0__abc_74894_new_n1818_), .B(u0__abc_74894_new_n1838_), .Y(u0__abc_74894_new_n4446_));
NAND2X1 NAND2X1_973 ( .A(1'h0), .B(u0__abc_74894_new_n1858_), .Y(u0__abc_74894_new_n4447_));
NAND2X1 NAND2X1_974 ( .A(u0__abc_74894_new_n1820_), .B(u0__abc_74894_new_n1840_), .Y(u0__abc_74894_new_n4452_));
NAND2X1 NAND2X1_975 ( .A(1'h0), .B(u0__abc_74894_new_n1860_), .Y(u0__abc_74894_new_n4453_));
NAND2X1 NAND2X1_976 ( .A(1'h0), .B(u0__abc_74894_new_n3797_), .Y(u0__abc_74894_new_n4456_));
NAND2X1 NAND2X1_977 ( .A(u0_lmr_ack_r), .B(u0__abc_74894_new_n4461_), .Y(u0__abc_74894_new_n4462_));
NAND2X1 NAND2X1_978 ( .A(u0_init_ack_r), .B(u0__abc_74894_new_n4463_), .Y(u0__abc_74894_new_n4464_));
NAND2X1 NAND2X1_979 ( .A(u0_u0__abc_72207_new_n206_), .B(u0_u0__abc_72207_new_n207_), .Y(u0_u0__abc_72207_new_n208_));
NAND2X1 NAND2X1_98 ( .A(spec_req_cs_5_), .B(u0__abc_74894_new_n1359_), .Y(u0__abc_74894_new_n1360_));
NAND2X1 NAND2X1_980 ( .A(u0_u0_inited), .B(u0_u0__abc_72207_new_n209_), .Y(u0_u0__abc_72207_new_n210_));
NAND2X1 NAND2X1_981 ( .A(u0_lmr_req0), .B(u0_u0__abc_72207_new_n211_), .Y(u0_u0__abc_72207_new_n212_));
NAND2X1 NAND2X1_982 ( .A(u0_u0_addr_r_4_), .B(u0_u0__abc_72207_new_n214_), .Y(u0_u0__abc_72207_new_n215_));
NAND2X1 NAND2X1_983 ( .A(u0_u0_addr_r_2_), .B(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n220_));
NAND2X1 NAND2X1_984 ( .A(u0_u0__abc_72207_new_n222_), .B(u0_u0__abc_72207_new_n223_), .Y(u0_u0__0tms_31_0__0_));
NAND2X1 NAND2X1_985 ( .A(u0_u0__abc_72207_new_n225_), .B(u0_u0__abc_72207_new_n226_), .Y(u0_u0__0tms_31_0__1_));
NAND2X1 NAND2X1_986 ( .A(u0_u0__abc_72207_new_n228_), .B(u0_u0__abc_72207_new_n229_), .Y(u0_u0__0tms_31_0__2_));
NAND2X1 NAND2X1_987 ( .A(u0_u0__abc_72207_new_n231_), .B(u0_u0__abc_72207_new_n232_), .Y(u0_u0__0tms_31_0__3_));
NAND2X1 NAND2X1_988 ( .A(u0_u0__abc_72207_new_n234_), .B(u0_u0__abc_72207_new_n235_), .Y(u0_u0__0tms_31_0__4_));
NAND2X1 NAND2X1_989 ( .A(u0_u0__abc_72207_new_n237_), .B(u0_u0__abc_72207_new_n238_), .Y(u0_u0__0tms_31_0__5_));
NAND2X1 NAND2X1_99 ( .A(1'h0), .B(u0__abc_74894_new_n1140_), .Y(u0__abc_74894_new_n1361_));
NAND2X1 NAND2X1_990 ( .A(u0_u0__abc_72207_new_n240_), .B(u0_u0__abc_72207_new_n241_), .Y(u0_u0__0tms_31_0__6_));
NAND2X1 NAND2X1_991 ( .A(u0_u0__abc_72207_new_n243_), .B(u0_u0__abc_72207_new_n244_), .Y(u0_u0__0tms_31_0__7_));
NAND2X1 NAND2X1_992 ( .A(u0_u0__abc_72207_new_n246_), .B(u0_u0__abc_72207_new_n247_), .Y(u0_u0__0tms_31_0__8_));
NAND2X1 NAND2X1_993 ( .A(u0_u0__abc_72207_new_n249_), .B(u0_u0__abc_72207_new_n250_), .Y(u0_u0__0tms_31_0__9_));
NAND2X1 NAND2X1_994 ( .A(u0_u0__abc_72207_new_n252_), .B(u0_u0__abc_72207_new_n253_), .Y(u0_u0__0tms_31_0__10_));
NAND2X1 NAND2X1_995 ( .A(u0_u0__abc_72207_new_n255_), .B(u0_u0__abc_72207_new_n256_), .Y(u0_u0__0tms_31_0__11_));
NAND2X1 NAND2X1_996 ( .A(u0_u0__abc_72207_new_n258_), .B(u0_u0__abc_72207_new_n259_), .Y(u0_u0__0tms_31_0__12_));
NAND2X1 NAND2X1_997 ( .A(u0_u0__abc_72207_new_n261_), .B(u0_u0__abc_72207_new_n262_), .Y(u0_u0__0tms_31_0__13_));
NAND2X1 NAND2X1_998 ( .A(u0_u0__abc_72207_new_n264_), .B(u0_u0__abc_72207_new_n265_), .Y(u0_u0__0tms_31_0__14_));
NAND2X1 NAND2X1_999 ( .A(u0_u0__abc_72207_new_n267_), .B(u0_u0__abc_72207_new_n268_), .Y(u0_u0__0tms_31_0__15_));
NAND3X1 NAND3X1_1 ( .A(u0__abc_74894_new_n1148_), .B(u0__abc_74894_new_n1151_), .C(u0__abc_74894_new_n1144_), .Y(u0__abc_74894_new_n1152_));
NAND3X1 NAND3X1_10 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1202_), .C(u0__abc_74894_new_n1201_), .Y(u0__abc_74894_new_n1203_));
NAND3X1 NAND3X1_100 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1645_), .C(u0__abc_74894_new_n1644_), .Y(u0__abc_74894_new_n1646_));
NAND3X1 NAND3X1_1000 ( .A(u5__abc_78290_new_n2061_), .B(u5__abc_78290_new_n2066_), .C(u5__abc_78290_new_n2060_), .Y(u5__abc_78290_new_n2067_));
NAND3X1 NAND3X1_1001 ( .A(u5__abc_78290_new_n2068_), .B(u5__abc_78290_new_n2070_), .C(u5__abc_78290_new_n2072_), .Y(u5__abc_78290_new_n2073_));
NAND3X1 NAND3X1_1002 ( .A(u5__abc_78290_new_n997_), .B(u5__abc_78290_new_n2056_), .C(u5__abc_78290_new_n2074_), .Y(u5__abc_78290_new_n2075_));
NAND3X1 NAND3X1_1003 ( .A(u5__abc_78290_new_n472_), .B(u5__abc_78290_new_n2076_), .C(u5__abc_78290_new_n1533_), .Y(u5__abc_78290_new_n2077_));
NAND3X1 NAND3X1_1004 ( .A(u5__abc_78290_new_n1996_), .B(u5__abc_78290_new_n1558_), .C(u5__abc_78290_new_n2079_), .Y(u5__abc_78290_new_n2080_));
NAND3X1 NAND3X1_1005 ( .A(u5__abc_78290_new_n2078_), .B(u5__abc_78290_new_n1549_), .C(u5__abc_78290_new_n2081_), .Y(u5__abc_78290_new_n2082_));
NAND3X1 NAND3X1_1006 ( .A(u5__abc_78290_new_n418_), .B(u5__abc_78290_new_n2098_), .C(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n2099_));
NAND3X1 NAND3X1_1007 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n2100_), .Y(u5__abc_78290_new_n2101_));
NAND3X1 NAND3X1_1008 ( .A(u5__abc_78290_new_n2106_), .B(u5__abc_78290_new_n1031_), .C(u5__abc_78290_new_n2107_), .Y(u5__abc_78290_new_n2108_));
NAND3X1 NAND3X1_1009 ( .A(u5__abc_78290_new_n2105_), .B(u5__abc_78290_new_n2109_), .C(u5__abc_78290_new_n2095_), .Y(u5__abc_78290_new_n2110_));
NAND3X1 NAND3X1_101 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1638_), .C(u0__abc_74894_new_n1646_), .Y(u0__abc_74894_new_n1647_));
NAND3X1 NAND3X1_1010 ( .A(u5__abc_78290_new_n1031_), .B(u5__abc_78290_new_n2113_), .C(u5__abc_78290_new_n1250_), .Y(u5__abc_78290_new_n2114_));
NAND3X1 NAND3X1_1011 ( .A(u5__abc_78290_new_n2115_), .B(u5__abc_78290_new_n2122_), .C(u5__abc_78290_new_n2095_), .Y(u5__abc_78290_new_n2123_));
NAND3X1 NAND3X1_1012 ( .A(u5__abc_78290_new_n2075_), .B(u5__abc_78290_new_n2127_), .C(u5__abc_78290_new_n2126_), .Y(u5__abc_78290_new_n2128_));
NAND3X1 NAND3X1_1013 ( .A(u5__abc_78290_new_n2040_), .B(u5__abc_78290_new_n2046_), .C(u5__abc_78290_new_n2128_), .Y(u5__abc_78290_new_n2129_));
NAND3X1 NAND3X1_1014 ( .A(u5__abc_78290_new_n786_), .B(u5__abc_78290_new_n612_), .C(u5__abc_78290_new_n2056_), .Y(u5__abc_78290_new_n2151_));
NAND3X1 NAND3X1_1015 ( .A(u5__abc_78290_new_n937_), .B(u5__abc_78290_new_n2157_), .C(u5__abc_78290_new_n2156_), .Y(u5__abc_78290_new_n2158_));
NAND3X1 NAND3X1_1016 ( .A(u5__abc_78290_new_n1039_), .B(u5__abc_78290_new_n882_), .C(u5__abc_78290_new_n2160_), .Y(u5__abc_78290_new_n2161_));
NAND3X1 NAND3X1_1017 ( .A(u5__abc_78290_new_n2154_), .B(u5__abc_78290_new_n2162_), .C(u5__abc_78290_new_n724_), .Y(u5__abc_78290_new_n2163_));
NAND3X1 NAND3X1_1018 ( .A(u5__abc_78290_new_n1193_), .B(u5__abc_78290_new_n1491_), .C(u5__abc_78290_new_n2171_), .Y(u5__abc_78290_new_n2172_));
NAND3X1 NAND3X1_1019 ( .A(u5__abc_78290_new_n2181_), .B(u5__abc_78290_new_n2184_), .C(u5__abc_78290_new_n1645_), .Y(u5__abc_78290_new_n2185_));
NAND3X1 NAND3X1_102 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1662_), .C(u0__abc_74894_new_n1661_), .Y(u0__abc_74894_new_n1663_));
NAND3X1 NAND3X1_1020 ( .A(u5__abc_78290_new_n1167_), .B(u5__abc_78290_new_n2193_), .C(u5__abc_78290_new_n2192_), .Y(u5__abc_78290_new_n2194_));
NAND3X1 NAND3X1_1021 ( .A(u5__abc_78290_new_n2195_), .B(u5__abc_78290_new_n2198_), .C(u5__abc_78290_new_n2203_), .Y(u5__abc_78290_new_n2204_));
NAND3X1 NAND3X1_1022 ( .A(u5__abc_78290_new_n2217_), .B(u5__abc_78290_new_n2219_), .C(u5__abc_78290_new_n1645_), .Y(u5__abc_78290_new_n2220_));
NAND3X1 NAND3X1_1023 ( .A(u5__abc_78290_new_n2216_), .B(u5__abc_78290_new_n2221_), .C(u5__abc_78290_new_n2178_), .Y(u5__abc_78290_new_n2222_));
NAND3X1 NAND3X1_1024 ( .A(u5__abc_78290_new_n2075_), .B(u5__abc_78290_new_n2239_), .C(u5__abc_78290_new_n2238_), .Y(u5__abc_78290_new_n2240_));
NAND3X1 NAND3X1_1025 ( .A(u5__abc_78290_new_n2040_), .B(u5__abc_78290_new_n2232_), .C(u5__abc_78290_new_n2240_), .Y(u5__abc_78290_new_n2241_));
NAND3X1 NAND3X1_1026 ( .A(u5__abc_78290_new_n2284_), .B(u5__abc_78290_new_n2286_), .C(u5__abc_78290_new_n2283_), .Y(u5__abc_78290_new_n2287_));
NAND3X1 NAND3X1_1027 ( .A(u5__abc_78290_new_n2278_), .B(u5__abc_78290_new_n1209_), .C(u5__abc_78290_new_n1988_), .Y(u5__abc_78290_new_n2289_));
NAND3X1 NAND3X1_1028 ( .A(u5__abc_78290_new_n2210_), .B(u5__abc_78290_new_n2263_), .C(u5__abc_78290_new_n2301_), .Y(u5__abc_78290_new_n2302_));
NAND3X1 NAND3X1_1029 ( .A(u5__abc_78290_new_n2265_), .B(u5__abc_78290_new_n2308_), .C(u5__abc_78290_new_n2270_), .Y(u5__abc_78290_new_n2309_));
NAND3X1 NAND3X1_103 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1660_), .C(u0__abc_74894_new_n1663_), .Y(u0__abc_74894_new_n1664_));
NAND3X1 NAND3X1_1030 ( .A(u5__abc_78290_new_n1996_), .B(u5__abc_78290_new_n1573_), .C(u5__abc_78290_new_n2329_), .Y(u5__abc_78290_new_n2330_));
NAND3X1 NAND3X1_1031 ( .A(u5__abc_78290_new_n2336_), .B(u5__abc_78290_new_n2338_), .C(u5__abc_78290_new_n2344_), .Y(u5__abc_78290_new_n2345_));
NAND3X1 NAND3X1_1032 ( .A(u5_timer_7_), .B(u5__abc_78290_new_n2357_), .C(u5__abc_78290_new_n2350_), .Y(u5__abc_78290_new_n2363_));
NAND3X1 NAND3X1_1033 ( .A(u5__abc_78290_new_n992_), .B(u5__abc_78290_new_n995_), .C(u5__abc_78290_new_n1525_), .Y(u5__abc_78290_new_n2369_));
NAND3X1 NAND3X1_1034 ( .A(u5__abc_78290_new_n666_), .B(u5__abc_78290_new_n702_), .C(u5__abc_78290_new_n2372_), .Y(u5__abc_78290_new_n2373_));
NAND3X1 NAND3X1_1035 ( .A(u5__abc_78290_new_n987_), .B(u5__abc_78290_new_n2375_), .C(u5__abc_78290_new_n2374_), .Y(u5__abc_78290_new_n2376_));
NAND3X1 NAND3X1_1036 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n1133_), .C(u5__abc_78290_new_n1637_), .Y(u5__abc_78290_new_n2383_));
NAND3X1 NAND3X1_1037 ( .A(u5__abc_78290_new_n1146_), .B(u5__abc_78290_new_n2386_), .C(u5__abc_78290_new_n1133_), .Y(u5__abc_78290_new_n2387_));
NAND3X1 NAND3X1_1038 ( .A(u5__abc_78290_new_n1386_), .B(u5__abc_78290_new_n1639_), .C(u5__abc_78290_new_n1637_), .Y(u5__abc_78290_new_n2389_));
NAND3X1 NAND3X1_1039 ( .A(u5__abc_78290_new_n1211_), .B(u5__abc_78290_new_n2283_), .C(u5__abc_78290_new_n2411_), .Y(u5__abc_78290_new_n2412_));
NAND3X1 NAND3X1_104 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1665_), .C(u0__abc_74894_new_n1664_), .Y(u0__abc_74894_new_n1666_));
NAND3X1 NAND3X1_1040 ( .A(u5__abc_78290_new_n2418_), .B(u5__abc_78290_new_n2419_), .C(u5__abc_78290_new_n2381_), .Y(u5__abc_78290_new_n2420_));
NAND3X1 NAND3X1_1041 ( .A(u5__abc_78290_new_n536_), .B(u5__abc_78290_new_n702_), .C(u5__abc_78290_new_n641_), .Y(u5__abc_78290_new_n2434_));
NAND3X1 NAND3X1_1042 ( .A(u5__abc_78290_new_n569_), .B(u5__abc_78290_new_n798_), .C(u5__abc_78290_new_n2061_), .Y(u5__abc_78290_new_n2439_));
NAND3X1 NAND3X1_1043 ( .A(u5__abc_78290_new_n1004_), .B(u5__abc_78290_new_n2438_), .C(u5__abc_78290_new_n2441_), .Y(u5__abc_78290_new_n2442_));
NAND3X1 NAND3X1_1044 ( .A(u5__abc_78290_new_n2053_), .B(u5__abc_78290_new_n2444_), .C(u5__abc_78290_new_n2445_), .Y(u5__abc_78290_new_n2446_));
NAND3X1 NAND3X1_1045 ( .A(u5__abc_78290_new_n1012_), .B(u5__abc_78290_new_n1015_), .C(u5__abc_78290_new_n990_), .Y(u5__abc_78290_new_n2448_));
NAND3X1 NAND3X1_1046 ( .A(u5__abc_78290_new_n2380_), .B(u5__abc_78290_new_n2498_), .C(u5__abc_78290_new_n2504_), .Y(u5__abc_78290_new_n2505_));
NAND3X1 NAND3X1_1047 ( .A(u5__abc_78290_new_n2465_), .B(u5__abc_78290_new_n2517_), .C(u5__abc_78290_new_n2479_), .Y(u5__abc_78290_new_n2518_));
NAND3X1 NAND3X1_1048 ( .A(u5__abc_78290_new_n2465_), .B(u5__abc_78290_new_n2391_), .C(u5__abc_78290_new_n2479_), .Y(u5__abc_78290_new_n2524_));
NAND3X1 NAND3X1_1049 ( .A(u5__abc_78290_new_n2199_), .B(u5__abc_78290_new_n2569_), .C(u5__abc_78290_new_n1072_), .Y(u5__abc_78290_new_n2570_));
NAND3X1 NAND3X1_105 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1658_), .C(u0__abc_74894_new_n1666_), .Y(u0__abc_74894_new_n1667_));
NAND3X1 NAND3X1_1050 ( .A(u5__abc_78290_new_n2597_), .B(u5__abc_78290_new_n2603_), .C(u5__abc_78290_new_n2596_), .Y(u5_next_state_1_));
NAND3X1 NAND3X1_1051 ( .A(u5__abc_78290_new_n2619_), .B(u5__abc_78290_new_n2634_), .C(u5__abc_78290_new_n2617_), .Y(u5__abc_78290_new_n2635_));
NAND3X1 NAND3X1_1052 ( .A(u5__abc_78290_new_n1324_), .B(u5_ap_en), .C(u5__abc_78290_new_n1412_), .Y(u5__abc_78290_new_n2637_));
NAND3X1 NAND3X1_1053 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n2637_), .C(u5__abc_78290_new_n2636_), .Y(u5__abc_78290_new_n2638_));
NAND3X1 NAND3X1_1054 ( .A(u5__abc_78290_new_n2665_), .B(u5__abc_78290_new_n2668_), .C(u5__abc_78290_new_n2663_), .Y(u5__abc_78290_new_n2669_));
NAND3X1 NAND3X1_1055 ( .A(u5_kro), .B(u5_wb_wait_r), .C(u5__abc_78290_new_n726_), .Y(u5__abc_78290_new_n2700_));
NAND3X1 NAND3X1_1056 ( .A(u5__abc_78290_new_n1257_), .B(u5__abc_78290_new_n2733_), .C(u5__abc_78290_new_n2731_), .Y(u5__abc_78290_new_n2734_));
NAND3X1 NAND3X1_1057 ( .A(u5__abc_78290_new_n2735_), .B(u5__abc_78290_new_n2738_), .C(u5__abc_78290_new_n2734_), .Y(u5_next_state_14_));
NAND3X1 NAND3X1_1058 ( .A(u5__abc_78290_new_n1324_), .B(u5__abc_78290_new_n1631_), .C(u5__abc_78290_new_n1412_), .Y(u5__abc_78290_new_n2756_));
NAND3X1 NAND3X1_1059 ( .A(u5_state_17_), .B(u5__abc_78290_new_n2592_), .C(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2772_));
NAND3X1 NAND3X1_106 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1682_), .C(u0__abc_74894_new_n1681_), .Y(u0__abc_74894_new_n1683_));
NAND3X1 NAND3X1_1060 ( .A(u5__abc_78290_new_n2775_), .B(u5__abc_78290_new_n2780_), .C(u5__abc_78290_new_n2772_), .Y(u5_next_state_17_));
NAND3X1 NAND3X1_1061 ( .A(u5_state_19_), .B(u5__abc_78290_new_n1342_), .C(u5__abc_78290_new_n2788_), .Y(u5__abc_78290_new_n2789_));
NAND3X1 NAND3X1_1062 ( .A(u5_state_20_), .B(u5__abc_78290_new_n2647_), .C(u5__abc_78290_new_n2788_), .Y(u5__abc_78290_new_n2797_));
NAND3X1 NAND3X1_1063 ( .A(u5_state_31_), .B(u5__abc_78290_new_n2680_), .C(u5__abc_78290_new_n2783_), .Y(u5__abc_78290_new_n2849_));
NAND3X1 NAND3X1_1064 ( .A(u5_state_52_), .B(u5__abc_78290_new_n1990_), .C(u5__abc_78290_new_n2218_), .Y(u5__abc_78290_new_n2924_));
NAND3X1 NAND3X1_1065 ( .A(u5__abc_78290_new_n2923_), .B(u5__abc_78290_new_n2924_), .C(u5__abc_78290_new_n2921_), .Y(u5_next_state_52_));
NAND3X1 NAND3X1_1066 ( .A(u5__abc_78290_new_n2192_), .B(u5__abc_78290_new_n2999_), .C(u5__abc_78290_new_n2277_), .Y(u5__abc_78290_new_n3000_));
NAND3X1 NAND3X1_1067 ( .A(u5__abc_78290_new_n767_), .B(u5__abc_78290_new_n2140_), .C(u5__abc_78290_new_n3006_), .Y(u5__abc_78290_new_n3007_));
NAND3X1 NAND3X1_1068 ( .A(u5__abc_78290_new_n1348_), .B(u5__abc_78290_new_n3010_), .C(u5__abc_78290_new_n2169_), .Y(u5__abc_78290_new_n3011_));
NAND3X1 NAND3X1_1069 ( .A(u5__abc_78290_new_n1193_), .B(u5__abc_78290_new_n1312_), .C(u5__abc_78290_new_n3018_), .Y(u5__abc_78290_new_n3019_));
NAND3X1 NAND3X1_107 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1680_), .C(u0__abc_74894_new_n1683_), .Y(u0__abc_74894_new_n1684_));
NAND3X1 NAND3X1_1070 ( .A(u5__abc_78290_new_n2283_), .B(u5__abc_78290_new_n3020_), .C(u5__abc_78290_new_n2280_), .Y(u5__abc_78290_new_n3021_));
NAND3X1 NAND3X1_1071 ( .A(u5__abc_78290_new_n2948_), .B(u5__abc_78290_new_n3024_), .C(u5__abc_78290_new_n1485_), .Y(mc_adsc_d));
NAND3X1 NAND3X1_1072 ( .A(u5__0no_wb_cycle_0_0_), .B(u5__abc_78290_new_n1343_), .C(u5__abc_78290_new_n3026_), .Y(u5__abc_78290_new_n3027_));
NAND3X1 NAND3X1_1073 ( .A(u5__abc_78290_new_n2175_), .B(u5__abc_78290_new_n2283_), .C(u5__abc_78290_new_n3032_), .Y(u5__abc_78290_new_n3033_));
NAND3X1 NAND3X1_1074 ( .A(u5__abc_78290_new_n2599_), .B(u5__abc_78290_new_n3042_), .C(u5__abc_78290_new_n574_), .Y(u5__abc_78290_new_n3043_));
NAND3X1 NAND3X1_1075 ( .A(u5__abc_78290_new_n2923_), .B(u5__abc_78290_new_n3043_), .C(u5__abc_78290_new_n3046_), .Y(u5__abc_78290_new_n3047_));
NAND3X1 NAND3X1_1076 ( .A(u5__abc_78290_new_n3037_), .B(u5__abc_78290_new_n3048_), .C(u5__abc_78290_new_n3036_), .Y(cs_le_d));
NAND3X1 NAND3X1_1077 ( .A(u5__abc_78290_new_n1312_), .B(u5__abc_78290_new_n3052_), .C(u5__abc_78290_new_n3029_), .Y(u5__abc_78290_new_n3053_));
NAND3X1 NAND3X1_1078 ( .A(u5__abc_78290_new_n1578_), .B(u5__abc_78290_new_n3055_), .C(u5__abc_78290_new_n3056_), .Y(u5__abc_78290_new_n3057_));
NAND3X1 NAND3X1_1079 ( .A(rfr_ack), .B(u5__abc_78290_new_n505_), .C(u5__abc_78290_new_n521_), .Y(u5__abc_78290_new_n3061_));
NAND3X1 NAND3X1_108 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1685_), .C(u0__abc_74894_new_n1684_), .Y(u0__abc_74894_new_n1686_));
NAND3X1 NAND3X1_1080 ( .A(u5__abc_78290_new_n2024_), .B(u5__abc_78290_new_n3063_), .C(u5__abc_78290_new_n3064_), .Y(u5__abc_78290_new_n3065_));
NAND3X1 NAND3X1_1081 ( .A(u5__abc_78290_new_n3060_), .B(u5__abc_78290_new_n1492_), .C(u5__abc_78290_new_n3065_), .Y(bank_clr_all));
NAND3X1 NAND3X1_1082 ( .A(u5__abc_78290_new_n2672_), .B(u5__abc_78290_new_n1437_), .C(u5__abc_78290_new_n1582_), .Y(u5__abc_78290_new_n3067_));
NAND3X1 NAND3X1_1083 ( .A(u5__abc_78290_new_n2173_), .B(u5__abc_78290_new_n3069_), .C(u5__abc_78290_new_n3064_), .Y(u5__abc_78290_new_n3070_));
NAND3X1 NAND3X1_1084 ( .A(u5__abc_78290_new_n3074_), .B(u5__abc_78290_new_n3076_), .C(u5__abc_78290_new_n1553_), .Y(u5__abc_78290_new_n3077_));
NAND3X1 NAND3X1_1085 ( .A(u5__abc_78290_new_n1528_), .B(u5__abc_78290_new_n3078_), .C(u5__abc_78290_new_n1117_), .Y(u5__abc_78290_new_n3079_));
NAND3X1 NAND3X1_1086 ( .A(u5__abc_78290_new_n2035_), .B(u5__abc_78290_new_n3084_), .C(u5__abc_78290_new_n2329_), .Y(u5__abc_78290_new_n3085_));
NAND3X1 NAND3X1_1087 ( .A(u5__abc_78290_new_n3091_), .B(u5__abc_78290_new_n3093_), .C(u5__abc_78290_new_n3092_), .Y(u5__abc_78290_new_n3094_));
NAND3X1 NAND3X1_1088 ( .A(u5__abc_78290_new_n3060_), .B(u5__abc_78290_new_n3100_), .C(u5__abc_78290_new_n3101_), .Y(u5__abc_78290_new_n3102_));
NAND3X1 NAND3X1_1089 ( .A(u5__abc_78290_new_n1291_), .B(u5__abc_78290_new_n3108_), .C(u5__abc_78290_new_n1460_), .Y(u5__abc_78290_new_n3109_));
NAND3X1 NAND3X1_109 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1678_), .C(u0__abc_74894_new_n1686_), .Y(u0__abc_74894_new_n1687_));
NAND3X1 NAND3X1_1090 ( .A(u5__abc_78290_new_n1384_), .B(u5__abc_78290_new_n1183_), .C(u5__abc_78290_new_n3121_), .Y(u5__abc_78290_new_n3122_));
NAND3X1 NAND3X1_1091 ( .A(u5__abc_78290_new_n1549_), .B(u5__abc_78290_new_n2078_), .C(u5__abc_78290_new_n3137_), .Y(u5__abc_78290_new_n3138_));
NAND3X1 NAND3X1_1092 ( .A(wb_stb_i), .B(cs_le), .C(wb_cyc_i), .Y(u5__abc_78290_new_n3141_));
NAND3X1 NAND3X1_1093 ( .A(wb_stb_i), .B(wb_cyc_i), .C(u5_lookup_ready1), .Y(u5__abc_78290_new_n3143_));
NAND3X1 NAND3X1_1094 ( .A(u5__abc_78290_new_n2425_), .B(u5__abc_78290_new_n3145_), .C(u5__abc_78290_new_n2465_), .Y(u5__abc_78290_new_n3146_));
NAND3X1 NAND3X1_1095 ( .A(u5__abc_78290_new_n1547_), .B(u5__abc_78290_new_n1992_), .C(u5__abc_78290_new_n2284_), .Y(u5__abc_78290_new_n3149_));
NAND3X1 NAND3X1_1096 ( .A(\wb_addr_i[30] ), .B(u6__abc_81318_new_n143_), .C(u6__abc_81318_new_n138_), .Y(u6__abc_81318_new_n144_));
NAND3X1 NAND3X1_1097 ( .A(wb_cyc_i), .B(wb_stb_i), .C(wb_we_i), .Y(u6__abc_81318_new_n243_));
NAND3X1 NAND3X1_1098 ( .A(wb_stb_i), .B(u6__abc_81318_new_n248_), .C(u6__abc_81318_new_n249_), .Y(u6__abc_81318_new_n250_));
NAND3X1 NAND3X1_1099 ( .A(wb_cyc_i), .B(u6__abc_81318_new_n251_), .C(u6__abc_81318_new_n255_), .Y(u6__abc_81318_new_n256_));
NAND3X1 NAND3X1_11 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1200_), .C(u0__abc_74894_new_n1203_), .Y(u0__abc_74894_new_n1204_));
NAND3X1 NAND3X1_110 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1702_), .C(u0__abc_74894_new_n1701_), .Y(u0__abc_74894_new_n1703_));
NAND3X1 NAND3X1_1100 ( .A(u6__abc_81318_new_n251_), .B(u6__0read_go_r_0_0_), .C(u6__abc_81318_new_n255_), .Y(u6__abc_81318_new_n260_));
NAND3X1 NAND3X1_1101 ( .A(wb_stb_i), .B(wb_we_i), .C(u6__abc_81318_new_n249_), .Y(u6__abc_81318_new_n263_));
NAND3X1 NAND3X1_1102 ( .A(u6__abc_81318_new_n251_), .B(u6__0write_go_r_0_0_), .C(u6__abc_81318_new_n255_), .Y(u6__abc_81318_new_n267_));
NAND3X1 NAND3X1_1103 ( .A(u6__abc_81318_new_n247_), .B(u6__abc_81318_new_n262_), .C(u6__abc_81318_new_n138_), .Y(u6__abc_81318_new_n269_));
NAND3X1 NAND3X1_1104 ( .A(u6_wb_first_r), .B(u6__abc_81318_new_n143_), .C(u6__abc_81318_new_n270_), .Y(u6__abc_81318_new_n271_));
NAND3X1 NAND3X1_1105 ( .A(u7__abc_73829_new_n75_), .B(u7__abc_73829_new_n79_), .C(u7__abc_73829_new_n77_), .Y(u7__0mc_dqm_3_0__0_));
NAND3X1 NAND3X1_1106 ( .A(u7__abc_73829_new_n75_), .B(u7__abc_73829_new_n79_), .C(u7__abc_73829_new_n81_), .Y(u7__0mc_dqm_3_0__1_));
NAND3X1 NAND3X1_1107 ( .A(u7__abc_73829_new_n75_), .B(u7__abc_73829_new_n79_), .C(u7__abc_73829_new_n83_), .Y(u7__0mc_dqm_3_0__2_));
NAND3X1 NAND3X1_1108 ( .A(u7__abc_73829_new_n75_), .B(u7__abc_73829_new_n79_), .C(u7__abc_73829_new_n85_), .Y(u7__0mc_dqm_3_0__3_));
NAND3X1 NAND3X1_1109 ( .A(u7__abc_73829_new_n100_), .B(u7__abc_73829_new_n103_), .C(u7__abc_73829_new_n102_), .Y(u7__abc_73829_new_n104_));
NAND3X1 NAND3X1_111 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1700_), .C(u0__abc_74894_new_n1703_), .Y(u0__abc_74894_new_n1704_));
NAND3X1 NAND3X1_1110 ( .A(u7__abc_73829_new_n100_), .B(u7__abc_73829_new_n111_), .C(u7__abc_73829_new_n110_), .Y(u7__abc_73829_new_n112_));
NAND3X1 NAND3X1_1111 ( .A(u7__abc_73829_new_n100_), .B(u7__abc_73829_new_n117_), .C(u7__abc_73829_new_n116_), .Y(u7__abc_73829_new_n118_));
NAND3X1 NAND3X1_1112 ( .A(u7__abc_73829_new_n100_), .B(u7__abc_73829_new_n123_), .C(u7__abc_73829_new_n122_), .Y(u7__abc_73829_new_n124_));
NAND3X1 NAND3X1_1113 ( .A(u7__abc_73829_new_n100_), .B(u7__abc_73829_new_n129_), .C(u7__abc_73829_new_n128_), .Y(u7__abc_73829_new_n130_));
NAND3X1 NAND3X1_1114 ( .A(u7__abc_73829_new_n100_), .B(u7__abc_73829_new_n135_), .C(u7__abc_73829_new_n134_), .Y(u7__abc_73829_new_n136_));
NAND3X1 NAND3X1_1115 ( .A(u7__abc_73829_new_n100_), .B(u7__abc_73829_new_n141_), .C(u7__abc_73829_new_n140_), .Y(u7__abc_73829_new_n142_));
NAND3X1 NAND3X1_1116 ( .A(u7__abc_73829_new_n100_), .B(u7__abc_73829_new_n147_), .C(u7__abc_73829_new_n146_), .Y(u7__abc_73829_new_n148_));
NAND3X1 NAND3X1_112 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1705_), .C(u0__abc_74894_new_n1704_), .Y(u0__abc_74894_new_n1706_));
NAND3X1 NAND3X1_113 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1698_), .C(u0__abc_74894_new_n1706_), .Y(u0__abc_74894_new_n1707_));
NAND3X1 NAND3X1_114 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1823_), .C(u0__abc_74894_new_n1822_), .Y(u0__abc_74894_new_n1824_));
NAND3X1 NAND3X1_115 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1821_), .C(u0__abc_74894_new_n1824_), .Y(u0__abc_74894_new_n1825_));
NAND3X1 NAND3X1_116 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1826_), .C(u0__abc_74894_new_n1825_), .Y(u0__abc_74894_new_n1827_));
NAND3X1 NAND3X1_117 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1819_), .C(u0__abc_74894_new_n1827_), .Y(u0__abc_74894_new_n1828_));
NAND3X1 NAND3X1_118 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1843_), .C(u0__abc_74894_new_n1842_), .Y(u0__abc_74894_new_n1844_));
NAND3X1 NAND3X1_119 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1841_), .C(u0__abc_74894_new_n1844_), .Y(u0__abc_74894_new_n1845_));
NAND3X1 NAND3X1_12 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1205_), .C(u0__abc_74894_new_n1204_), .Y(u0__abc_74894_new_n1206_));
NAND3X1 NAND3X1_120 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1846_), .C(u0__abc_74894_new_n1845_), .Y(u0__abc_74894_new_n1847_));
NAND3X1 NAND3X1_121 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1839_), .C(u0__abc_74894_new_n1847_), .Y(u0__abc_74894_new_n1848_));
NAND3X1 NAND3X1_122 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1863_), .C(u0__abc_74894_new_n1862_), .Y(u0__abc_74894_new_n1864_));
NAND3X1 NAND3X1_123 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1861_), .C(u0__abc_74894_new_n1864_), .Y(u0__abc_74894_new_n1865_));
NAND3X1 NAND3X1_124 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1866_), .C(u0__abc_74894_new_n1865_), .Y(u0__abc_74894_new_n1867_));
NAND3X1 NAND3X1_125 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1859_), .C(u0__abc_74894_new_n1867_), .Y(u0__abc_74894_new_n1868_));
NAND3X1 NAND3X1_126 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1883_), .C(u0__abc_74894_new_n1882_), .Y(u0__abc_74894_new_n1884_));
NAND3X1 NAND3X1_127 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1881_), .C(u0__abc_74894_new_n1884_), .Y(u0__abc_74894_new_n1885_));
NAND3X1 NAND3X1_128 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1886_), .C(u0__abc_74894_new_n1885_), .Y(u0__abc_74894_new_n1887_));
NAND3X1 NAND3X1_129 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1879_), .C(u0__abc_74894_new_n1887_), .Y(u0__abc_74894_new_n1888_));
NAND3X1 NAND3X1_13 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1198_), .C(u0__abc_74894_new_n1206_), .Y(u0__abc_74894_new_n1207_));
NAND3X1 NAND3X1_130 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1903_), .C(u0__abc_74894_new_n1902_), .Y(u0__abc_74894_new_n1904_));
NAND3X1 NAND3X1_131 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1901_), .C(u0__abc_74894_new_n1904_), .Y(u0__abc_74894_new_n1905_));
NAND3X1 NAND3X1_132 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1906_), .C(u0__abc_74894_new_n1905_), .Y(u0__abc_74894_new_n1907_));
NAND3X1 NAND3X1_133 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1899_), .C(u0__abc_74894_new_n1907_), .Y(u0__abc_74894_new_n1908_));
NAND3X1 NAND3X1_134 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1923_), .C(u0__abc_74894_new_n1922_), .Y(u0__abc_74894_new_n1924_));
NAND3X1 NAND3X1_135 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1921_), .C(u0__abc_74894_new_n1924_), .Y(u0__abc_74894_new_n1925_));
NAND3X1 NAND3X1_136 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1926_), .C(u0__abc_74894_new_n1925_), .Y(u0__abc_74894_new_n1927_));
NAND3X1 NAND3X1_137 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1919_), .C(u0__abc_74894_new_n1927_), .Y(u0__abc_74894_new_n1928_));
NAND3X1 NAND3X1_138 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1943_), .C(u0__abc_74894_new_n1942_), .Y(u0__abc_74894_new_n1944_));
NAND3X1 NAND3X1_139 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1941_), .C(u0__abc_74894_new_n1944_), .Y(u0__abc_74894_new_n1945_));
NAND3X1 NAND3X1_14 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1222_), .C(u0__abc_74894_new_n1221_), .Y(u0__abc_74894_new_n1223_));
NAND3X1 NAND3X1_140 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1946_), .C(u0__abc_74894_new_n1945_), .Y(u0__abc_74894_new_n1947_));
NAND3X1 NAND3X1_141 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1939_), .C(u0__abc_74894_new_n1947_), .Y(u0__abc_74894_new_n1948_));
NAND3X1 NAND3X1_142 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1983_), .C(u0__abc_74894_new_n1982_), .Y(u0__abc_74894_new_n1984_));
NAND3X1 NAND3X1_143 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1981_), .C(u0__abc_74894_new_n1984_), .Y(u0__abc_74894_new_n1985_));
NAND3X1 NAND3X1_144 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1986_), .C(u0__abc_74894_new_n1985_), .Y(u0__abc_74894_new_n1987_));
NAND3X1 NAND3X1_145 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1979_), .C(u0__abc_74894_new_n1987_), .Y(u0__abc_74894_new_n1988_));
NAND3X1 NAND3X1_146 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n2003_), .C(u0__abc_74894_new_n2002_), .Y(u0__abc_74894_new_n2004_));
NAND3X1 NAND3X1_147 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n2001_), .C(u0__abc_74894_new_n2004_), .Y(u0__abc_74894_new_n2005_));
NAND3X1 NAND3X1_148 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n2006_), .C(u0__abc_74894_new_n2005_), .Y(u0__abc_74894_new_n2007_));
NAND3X1 NAND3X1_149 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1999_), .C(u0__abc_74894_new_n2007_), .Y(u0__abc_74894_new_n2008_));
NAND3X1 NAND3X1_15 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1220_), .C(u0__abc_74894_new_n1223_), .Y(u0__abc_74894_new_n1224_));
NAND3X1 NAND3X1_150 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2446_), .C(u0__abc_74894_new_n2445_), .Y(u0__abc_74894_new_n2447_));
NAND3X1 NAND3X1_151 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2442_), .C(u0__abc_74894_new_n2447_), .Y(u0__abc_74894_new_n2448_));
NAND3X1 NAND3X1_152 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2449_), .C(u0__abc_74894_new_n2448_), .Y(u0__abc_74894_new_n2450_));
NAND3X1 NAND3X1_153 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2439_), .C(u0__abc_74894_new_n2450_), .Y(u0__abc_74894_new_n2451_));
NAND3X1 NAND3X1_154 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2464_), .C(u0__abc_74894_new_n2463_), .Y(u0__abc_74894_new_n2465_));
NAND3X1 NAND3X1_155 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2462_), .C(u0__abc_74894_new_n2465_), .Y(u0__abc_74894_new_n2466_));
NAND3X1 NAND3X1_156 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2467_), .C(u0__abc_74894_new_n2466_), .Y(u0__abc_74894_new_n2468_));
NAND3X1 NAND3X1_157 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2461_), .C(u0__abc_74894_new_n2468_), .Y(u0__abc_74894_new_n2469_));
NAND3X1 NAND3X1_158 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2480_), .C(u0__abc_74894_new_n2479_), .Y(u0__abc_74894_new_n2481_));
NAND3X1 NAND3X1_159 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2478_), .C(u0__abc_74894_new_n2481_), .Y(u0__abc_74894_new_n2482_));
NAND3X1 NAND3X1_16 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1225_), .C(u0__abc_74894_new_n1224_), .Y(u0__abc_74894_new_n1226_));
NAND3X1 NAND3X1_160 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2483_), .C(u0__abc_74894_new_n2482_), .Y(u0__abc_74894_new_n2484_));
NAND3X1 NAND3X1_161 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2477_), .C(u0__abc_74894_new_n2484_), .Y(u0__abc_74894_new_n2485_));
NAND3X1 NAND3X1_162 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2496_), .C(u0__abc_74894_new_n2495_), .Y(u0__abc_74894_new_n2497_));
NAND3X1 NAND3X1_163 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2494_), .C(u0__abc_74894_new_n2497_), .Y(u0__abc_74894_new_n2498_));
NAND3X1 NAND3X1_164 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2499_), .C(u0__abc_74894_new_n2498_), .Y(u0__abc_74894_new_n2500_));
NAND3X1 NAND3X1_165 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2493_), .C(u0__abc_74894_new_n2500_), .Y(u0__abc_74894_new_n2501_));
NAND3X1 NAND3X1_166 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2512_), .C(u0__abc_74894_new_n2511_), .Y(u0__abc_74894_new_n2513_));
NAND3X1 NAND3X1_167 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2510_), .C(u0__abc_74894_new_n2513_), .Y(u0__abc_74894_new_n2514_));
NAND3X1 NAND3X1_168 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2515_), .C(u0__abc_74894_new_n2514_), .Y(u0__abc_74894_new_n2516_));
NAND3X1 NAND3X1_169 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2509_), .C(u0__abc_74894_new_n2516_), .Y(u0__abc_74894_new_n2517_));
NAND3X1 NAND3X1_17 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1218_), .C(u0__abc_74894_new_n1226_), .Y(u0__abc_74894_new_n1227_));
NAND3X1 NAND3X1_170 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2528_), .C(u0__abc_74894_new_n2527_), .Y(u0__abc_74894_new_n2529_));
NAND3X1 NAND3X1_171 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2526_), .C(u0__abc_74894_new_n2529_), .Y(u0__abc_74894_new_n2530_));
NAND3X1 NAND3X1_172 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2531_), .C(u0__abc_74894_new_n2530_), .Y(u0__abc_74894_new_n2532_));
NAND3X1 NAND3X1_173 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2525_), .C(u0__abc_74894_new_n2532_), .Y(u0__abc_74894_new_n2533_));
NAND3X1 NAND3X1_174 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2544_), .C(u0__abc_74894_new_n2543_), .Y(u0__abc_74894_new_n2545_));
NAND3X1 NAND3X1_175 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2542_), .C(u0__abc_74894_new_n2545_), .Y(u0__abc_74894_new_n2546_));
NAND3X1 NAND3X1_176 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2547_), .C(u0__abc_74894_new_n2546_), .Y(u0__abc_74894_new_n2548_));
NAND3X1 NAND3X1_177 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2541_), .C(u0__abc_74894_new_n2548_), .Y(u0__abc_74894_new_n2549_));
NAND3X1 NAND3X1_178 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2560_), .C(u0__abc_74894_new_n2559_), .Y(u0__abc_74894_new_n2561_));
NAND3X1 NAND3X1_179 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2558_), .C(u0__abc_74894_new_n2561_), .Y(u0__abc_74894_new_n2562_));
NAND3X1 NAND3X1_18 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1242_), .C(u0__abc_74894_new_n1241_), .Y(u0__abc_74894_new_n1243_));
NAND3X1 NAND3X1_180 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2563_), .C(u0__abc_74894_new_n2562_), .Y(u0__abc_74894_new_n2564_));
NAND3X1 NAND3X1_181 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2557_), .C(u0__abc_74894_new_n2564_), .Y(u0__abc_74894_new_n2565_));
NAND3X1 NAND3X1_182 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2576_), .C(u0__abc_74894_new_n2575_), .Y(u0__abc_74894_new_n2577_));
NAND3X1 NAND3X1_183 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2574_), .C(u0__abc_74894_new_n2577_), .Y(u0__abc_74894_new_n2578_));
NAND3X1 NAND3X1_184 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2579_), .C(u0__abc_74894_new_n2578_), .Y(u0__abc_74894_new_n2580_));
NAND3X1 NAND3X1_185 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2573_), .C(u0__abc_74894_new_n2580_), .Y(u0__abc_74894_new_n2581_));
NAND3X1 NAND3X1_186 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2592_), .C(u0__abc_74894_new_n2591_), .Y(u0__abc_74894_new_n2593_));
NAND3X1 NAND3X1_187 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2590_), .C(u0__abc_74894_new_n2593_), .Y(u0__abc_74894_new_n2594_));
NAND3X1 NAND3X1_188 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2595_), .C(u0__abc_74894_new_n2594_), .Y(u0__abc_74894_new_n2596_));
NAND3X1 NAND3X1_189 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2589_), .C(u0__abc_74894_new_n2596_), .Y(u0__abc_74894_new_n2597_));
NAND3X1 NAND3X1_19 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1240_), .C(u0__abc_74894_new_n1243_), .Y(u0__abc_74894_new_n1244_));
NAND3X1 NAND3X1_190 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2608_), .C(u0__abc_74894_new_n2607_), .Y(u0__abc_74894_new_n2609_));
NAND3X1 NAND3X1_191 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2606_), .C(u0__abc_74894_new_n2609_), .Y(u0__abc_74894_new_n2610_));
NAND3X1 NAND3X1_192 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2611_), .C(u0__abc_74894_new_n2610_), .Y(u0__abc_74894_new_n2612_));
NAND3X1 NAND3X1_193 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2605_), .C(u0__abc_74894_new_n2612_), .Y(u0__abc_74894_new_n2613_));
NAND3X1 NAND3X1_194 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2624_), .C(u0__abc_74894_new_n2623_), .Y(u0__abc_74894_new_n2625_));
NAND3X1 NAND3X1_195 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2622_), .C(u0__abc_74894_new_n2625_), .Y(u0__abc_74894_new_n2626_));
NAND3X1 NAND3X1_196 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2627_), .C(u0__abc_74894_new_n2626_), .Y(u0__abc_74894_new_n2628_));
NAND3X1 NAND3X1_197 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2621_), .C(u0__abc_74894_new_n2628_), .Y(u0__abc_74894_new_n2629_));
NAND3X1 NAND3X1_198 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2640_), .C(u0__abc_74894_new_n2639_), .Y(u0__abc_74894_new_n2641_));
NAND3X1 NAND3X1_199 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2638_), .C(u0__abc_74894_new_n2641_), .Y(u0__abc_74894_new_n2642_));
NAND3X1 NAND3X1_2 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1162_), .C(u0__abc_74894_new_n1161_), .Y(u0__abc_74894_new_n1163_));
NAND3X1 NAND3X1_20 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1245_), .C(u0__abc_74894_new_n1244_), .Y(u0__abc_74894_new_n1246_));
NAND3X1 NAND3X1_200 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2643_), .C(u0__abc_74894_new_n2642_), .Y(u0__abc_74894_new_n2644_));
NAND3X1 NAND3X1_201 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2637_), .C(u0__abc_74894_new_n2644_), .Y(u0__abc_74894_new_n2645_));
NAND3X1 NAND3X1_202 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2656_), .C(u0__abc_74894_new_n2655_), .Y(u0__abc_74894_new_n2657_));
NAND3X1 NAND3X1_203 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2654_), .C(u0__abc_74894_new_n2657_), .Y(u0__abc_74894_new_n2658_));
NAND3X1 NAND3X1_204 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2659_), .C(u0__abc_74894_new_n2658_), .Y(u0__abc_74894_new_n2660_));
NAND3X1 NAND3X1_205 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2653_), .C(u0__abc_74894_new_n2660_), .Y(u0__abc_74894_new_n2661_));
NAND3X1 NAND3X1_206 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2672_), .C(u0__abc_74894_new_n2671_), .Y(u0__abc_74894_new_n2673_));
NAND3X1 NAND3X1_207 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2670_), .C(u0__abc_74894_new_n2673_), .Y(u0__abc_74894_new_n2674_));
NAND3X1 NAND3X1_208 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2675_), .C(u0__abc_74894_new_n2674_), .Y(u0__abc_74894_new_n2676_));
NAND3X1 NAND3X1_209 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2669_), .C(u0__abc_74894_new_n2676_), .Y(u0__abc_74894_new_n2677_));
NAND3X1 NAND3X1_21 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1238_), .C(u0__abc_74894_new_n1246_), .Y(u0__abc_74894_new_n1247_));
NAND3X1 NAND3X1_210 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2688_), .C(u0__abc_74894_new_n2687_), .Y(u0__abc_74894_new_n2689_));
NAND3X1 NAND3X1_211 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2686_), .C(u0__abc_74894_new_n2689_), .Y(u0__abc_74894_new_n2690_));
NAND3X1 NAND3X1_212 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2691_), .C(u0__abc_74894_new_n2690_), .Y(u0__abc_74894_new_n2692_));
NAND3X1 NAND3X1_213 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2685_), .C(u0__abc_74894_new_n2692_), .Y(u0__abc_74894_new_n2693_));
NAND3X1 NAND3X1_214 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2704_), .C(u0__abc_74894_new_n2703_), .Y(u0__abc_74894_new_n2705_));
NAND3X1 NAND3X1_215 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2702_), .C(u0__abc_74894_new_n2705_), .Y(u0__abc_74894_new_n2706_));
NAND3X1 NAND3X1_216 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2707_), .C(u0__abc_74894_new_n2706_), .Y(u0__abc_74894_new_n2708_));
NAND3X1 NAND3X1_217 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2701_), .C(u0__abc_74894_new_n2708_), .Y(u0__abc_74894_new_n2709_));
NAND3X1 NAND3X1_218 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2720_), .C(u0__abc_74894_new_n2719_), .Y(u0__abc_74894_new_n2721_));
NAND3X1 NAND3X1_219 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2718_), .C(u0__abc_74894_new_n2721_), .Y(u0__abc_74894_new_n2722_));
NAND3X1 NAND3X1_22 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1262_), .C(u0__abc_74894_new_n1261_), .Y(u0__abc_74894_new_n1263_));
NAND3X1 NAND3X1_220 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2723_), .C(u0__abc_74894_new_n2722_), .Y(u0__abc_74894_new_n2724_));
NAND3X1 NAND3X1_221 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2717_), .C(u0__abc_74894_new_n2724_), .Y(u0__abc_74894_new_n2725_));
NAND3X1 NAND3X1_222 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2736_), .C(u0__abc_74894_new_n2735_), .Y(u0__abc_74894_new_n2737_));
NAND3X1 NAND3X1_223 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2734_), .C(u0__abc_74894_new_n2737_), .Y(u0__abc_74894_new_n2738_));
NAND3X1 NAND3X1_224 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2739_), .C(u0__abc_74894_new_n2738_), .Y(u0__abc_74894_new_n2740_));
NAND3X1 NAND3X1_225 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2733_), .C(u0__abc_74894_new_n2740_), .Y(u0__abc_74894_new_n2741_));
NAND3X1 NAND3X1_226 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2752_), .C(u0__abc_74894_new_n2751_), .Y(u0__abc_74894_new_n2753_));
NAND3X1 NAND3X1_227 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2750_), .C(u0__abc_74894_new_n2753_), .Y(u0__abc_74894_new_n2754_));
NAND3X1 NAND3X1_228 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2755_), .C(u0__abc_74894_new_n2754_), .Y(u0__abc_74894_new_n2756_));
NAND3X1 NAND3X1_229 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2749_), .C(u0__abc_74894_new_n2756_), .Y(u0__abc_74894_new_n2757_));
NAND3X1 NAND3X1_23 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1260_), .C(u0__abc_74894_new_n1263_), .Y(u0__abc_74894_new_n1264_));
NAND3X1 NAND3X1_230 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2768_), .C(u0__abc_74894_new_n2767_), .Y(u0__abc_74894_new_n2769_));
NAND3X1 NAND3X1_231 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2766_), .C(u0__abc_74894_new_n2769_), .Y(u0__abc_74894_new_n2770_));
NAND3X1 NAND3X1_232 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2771_), .C(u0__abc_74894_new_n2770_), .Y(u0__abc_74894_new_n2772_));
NAND3X1 NAND3X1_233 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2765_), .C(u0__abc_74894_new_n2772_), .Y(u0__abc_74894_new_n2773_));
NAND3X1 NAND3X1_234 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2784_), .C(u0__abc_74894_new_n2783_), .Y(u0__abc_74894_new_n2785_));
NAND3X1 NAND3X1_235 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2782_), .C(u0__abc_74894_new_n2785_), .Y(u0__abc_74894_new_n2786_));
NAND3X1 NAND3X1_236 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2787_), .C(u0__abc_74894_new_n2786_), .Y(u0__abc_74894_new_n2788_));
NAND3X1 NAND3X1_237 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2781_), .C(u0__abc_74894_new_n2788_), .Y(u0__abc_74894_new_n2789_));
NAND3X1 NAND3X1_238 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2800_), .C(u0__abc_74894_new_n2799_), .Y(u0__abc_74894_new_n2801_));
NAND3X1 NAND3X1_239 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2798_), .C(u0__abc_74894_new_n2801_), .Y(u0__abc_74894_new_n2802_));
NAND3X1 NAND3X1_24 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1265_), .C(u0__abc_74894_new_n1264_), .Y(u0__abc_74894_new_n1266_));
NAND3X1 NAND3X1_240 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2803_), .C(u0__abc_74894_new_n2802_), .Y(u0__abc_74894_new_n2804_));
NAND3X1 NAND3X1_241 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2797_), .C(u0__abc_74894_new_n2804_), .Y(u0__abc_74894_new_n2805_));
NAND3X1 NAND3X1_242 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2816_), .C(u0__abc_74894_new_n2815_), .Y(u0__abc_74894_new_n2817_));
NAND3X1 NAND3X1_243 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2814_), .C(u0__abc_74894_new_n2817_), .Y(u0__abc_74894_new_n2818_));
NAND3X1 NAND3X1_244 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2819_), .C(u0__abc_74894_new_n2818_), .Y(u0__abc_74894_new_n2820_));
NAND3X1 NAND3X1_245 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2813_), .C(u0__abc_74894_new_n2820_), .Y(u0__abc_74894_new_n2821_));
NAND3X1 NAND3X1_246 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2832_), .C(u0__abc_74894_new_n2831_), .Y(u0__abc_74894_new_n2833_));
NAND3X1 NAND3X1_247 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2830_), .C(u0__abc_74894_new_n2833_), .Y(u0__abc_74894_new_n2834_));
NAND3X1 NAND3X1_248 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2835_), .C(u0__abc_74894_new_n2834_), .Y(u0__abc_74894_new_n2836_));
NAND3X1 NAND3X1_249 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2829_), .C(u0__abc_74894_new_n2836_), .Y(u0__abc_74894_new_n2837_));
NAND3X1 NAND3X1_25 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1258_), .C(u0__abc_74894_new_n1266_), .Y(u0__abc_74894_new_n1267_));
NAND3X1 NAND3X1_250 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2848_), .C(u0__abc_74894_new_n2847_), .Y(u0__abc_74894_new_n2849_));
NAND3X1 NAND3X1_251 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2846_), .C(u0__abc_74894_new_n2849_), .Y(u0__abc_74894_new_n2850_));
NAND3X1 NAND3X1_252 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2851_), .C(u0__abc_74894_new_n2850_), .Y(u0__abc_74894_new_n2852_));
NAND3X1 NAND3X1_253 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2845_), .C(u0__abc_74894_new_n2852_), .Y(u0__abc_74894_new_n2853_));
NAND3X1 NAND3X1_254 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2864_), .C(u0__abc_74894_new_n2863_), .Y(u0__abc_74894_new_n2865_));
NAND3X1 NAND3X1_255 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2862_), .C(u0__abc_74894_new_n2865_), .Y(u0__abc_74894_new_n2866_));
NAND3X1 NAND3X1_256 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2867_), .C(u0__abc_74894_new_n2866_), .Y(u0__abc_74894_new_n2868_));
NAND3X1 NAND3X1_257 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2861_), .C(u0__abc_74894_new_n2868_), .Y(u0__abc_74894_new_n2869_));
NAND3X1 NAND3X1_258 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2880_), .C(u0__abc_74894_new_n2879_), .Y(u0__abc_74894_new_n2881_));
NAND3X1 NAND3X1_259 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2878_), .C(u0__abc_74894_new_n2881_), .Y(u0__abc_74894_new_n2882_));
NAND3X1 NAND3X1_26 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1282_), .C(u0__abc_74894_new_n1281_), .Y(u0__abc_74894_new_n1283_));
NAND3X1 NAND3X1_260 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2883_), .C(u0__abc_74894_new_n2882_), .Y(u0__abc_74894_new_n2884_));
NAND3X1 NAND3X1_261 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2877_), .C(u0__abc_74894_new_n2884_), .Y(u0__abc_74894_new_n2885_));
NAND3X1 NAND3X1_262 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2977_), .C(u0__abc_74894_new_n2976_), .Y(u0__abc_74894_new_n2978_));
NAND3X1 NAND3X1_263 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2975_), .C(u0__abc_74894_new_n2978_), .Y(u0__abc_74894_new_n2979_));
NAND3X1 NAND3X1_264 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2980_), .C(u0__abc_74894_new_n2979_), .Y(u0__abc_74894_new_n2981_));
NAND3X1 NAND3X1_265 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2974_), .C(u0__abc_74894_new_n2981_), .Y(u0__abc_74894_new_n2982_));
NAND3X1 NAND3X1_266 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n2993_), .C(u0__abc_74894_new_n2992_), .Y(u0__abc_74894_new_n2994_));
NAND3X1 NAND3X1_267 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n2991_), .C(u0__abc_74894_new_n2994_), .Y(u0__abc_74894_new_n2995_));
NAND3X1 NAND3X1_268 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n2996_), .C(u0__abc_74894_new_n2995_), .Y(u0__abc_74894_new_n2997_));
NAND3X1 NAND3X1_269 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n2990_), .C(u0__abc_74894_new_n2997_), .Y(u0__abc_74894_new_n2998_));
NAND3X1 NAND3X1_27 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1280_), .C(u0__abc_74894_new_n1283_), .Y(u0__abc_74894_new_n1284_));
NAND3X1 NAND3X1_270 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n3009_), .C(u0__abc_74894_new_n3008_), .Y(u0__abc_74894_new_n3010_));
NAND3X1 NAND3X1_271 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n3007_), .C(u0__abc_74894_new_n3010_), .Y(u0__abc_74894_new_n3011_));
NAND3X1 NAND3X1_272 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n3012_), .C(u0__abc_74894_new_n3011_), .Y(u0__abc_74894_new_n3013_));
NAND3X1 NAND3X1_273 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n3006_), .C(u0__abc_74894_new_n3013_), .Y(u0__abc_74894_new_n3014_));
NAND3X1 NAND3X1_274 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n3025_), .C(u0__abc_74894_new_n3024_), .Y(u0__abc_74894_new_n3026_));
NAND3X1 NAND3X1_275 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n3023_), .C(u0__abc_74894_new_n3026_), .Y(u0__abc_74894_new_n3027_));
NAND3X1 NAND3X1_276 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n3028_), .C(u0__abc_74894_new_n3027_), .Y(u0__abc_74894_new_n3029_));
NAND3X1 NAND3X1_277 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n3022_), .C(u0__abc_74894_new_n3029_), .Y(u0__abc_74894_new_n3030_));
NAND3X1 NAND3X1_278 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n3041_), .C(u0__abc_74894_new_n3040_), .Y(u0__abc_74894_new_n3042_));
NAND3X1 NAND3X1_279 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n3039_), .C(u0__abc_74894_new_n3042_), .Y(u0__abc_74894_new_n3043_));
NAND3X1 NAND3X1_28 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1285_), .C(u0__abc_74894_new_n1284_), .Y(u0__abc_74894_new_n1286_));
NAND3X1 NAND3X1_280 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n3044_), .C(u0__abc_74894_new_n3043_), .Y(u0__abc_74894_new_n3045_));
NAND3X1 NAND3X1_281 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n3038_), .C(u0__abc_74894_new_n3045_), .Y(u0__abc_74894_new_n3046_));
NAND3X1 NAND3X1_282 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n3057_), .C(u0__abc_74894_new_n3056_), .Y(u0__abc_74894_new_n3058_));
NAND3X1 NAND3X1_283 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n3055_), .C(u0__abc_74894_new_n3058_), .Y(u0__abc_74894_new_n3059_));
NAND3X1 NAND3X1_284 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n3060_), .C(u0__abc_74894_new_n3059_), .Y(u0__abc_74894_new_n3061_));
NAND3X1 NAND3X1_285 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n3054_), .C(u0__abc_74894_new_n3061_), .Y(u0__abc_74894_new_n3062_));
NAND3X1 NAND3X1_286 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n3073_), .C(u0__abc_74894_new_n3072_), .Y(u0__abc_74894_new_n3074_));
NAND3X1 NAND3X1_287 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n3071_), .C(u0__abc_74894_new_n3074_), .Y(u0__abc_74894_new_n3075_));
NAND3X1 NAND3X1_288 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n3076_), .C(u0__abc_74894_new_n3075_), .Y(u0__abc_74894_new_n3077_));
NAND3X1 NAND3X1_289 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n3070_), .C(u0__abc_74894_new_n3077_), .Y(u0__abc_74894_new_n3078_));
NAND3X1 NAND3X1_29 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1278_), .C(u0__abc_74894_new_n1286_), .Y(u0__abc_74894_new_n1287_));
NAND3X1 NAND3X1_290 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n3105_), .C(u0__abc_74894_new_n3104_), .Y(u0__abc_74894_new_n3106_));
NAND3X1 NAND3X1_291 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n3103_), .C(u0__abc_74894_new_n3106_), .Y(u0__abc_74894_new_n3107_));
NAND3X1 NAND3X1_292 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n3108_), .C(u0__abc_74894_new_n3107_), .Y(u0__abc_74894_new_n3109_));
NAND3X1 NAND3X1_293 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n3102_), .C(u0__abc_74894_new_n3109_), .Y(u0__abc_74894_new_n3110_));
NAND3X1 NAND3X1_294 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n3121_), .C(u0__abc_74894_new_n3120_), .Y(u0__abc_74894_new_n3122_));
NAND3X1 NAND3X1_295 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n3119_), .C(u0__abc_74894_new_n3122_), .Y(u0__abc_74894_new_n3123_));
NAND3X1 NAND3X1_296 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n3124_), .C(u0__abc_74894_new_n3123_), .Y(u0__abc_74894_new_n3125_));
NAND3X1 NAND3X1_297 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n3118_), .C(u0__abc_74894_new_n3125_), .Y(u0__abc_74894_new_n3126_));
NAND3X1 NAND3X1_298 ( .A(u0__abc_74894_new_n2443_), .B(u0__abc_74894_new_n3137_), .C(u0__abc_74894_new_n3136_), .Y(u0__abc_74894_new_n3138_));
NAND3X1 NAND3X1_299 ( .A(u0__abc_74894_new_n2441_), .B(u0__abc_74894_new_n3135_), .C(u0__abc_74894_new_n3138_), .Y(u0__abc_74894_new_n3139_));
NAND3X1 NAND3X1_3 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1160_), .C(u0__abc_74894_new_n1163_), .Y(u0__abc_74894_new_n1164_));
NAND3X1 NAND3X1_30 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1302_), .C(u0__abc_74894_new_n1301_), .Y(u0__abc_74894_new_n1303_));
NAND3X1 NAND3X1_300 ( .A(u0__abc_74894_new_n2440_), .B(u0__abc_74894_new_n3140_), .C(u0__abc_74894_new_n3139_), .Y(u0__abc_74894_new_n3141_));
NAND3X1 NAND3X1_301 ( .A(u0__abc_74894_new_n2438_), .B(u0__abc_74894_new_n3134_), .C(u0__abc_74894_new_n3141_), .Y(u0__abc_74894_new_n3142_));
NAND3X1 NAND3X1_302 ( .A(u0__abc_74894_new_n3472_), .B(u0__abc_74894_new_n3473_), .C(u0__abc_74894_new_n3474_), .Y(u0__abc_74894_new_n3475_));
NAND3X1 NAND3X1_303 ( .A(u0_rf_we), .B(u0_wb_addr_r_3_), .C(u0__abc_74894_new_n3596_), .Y(u0__abc_74894_new_n3597_));
NAND3X1 NAND3X1_304 ( .A(u0_rf_we), .B(u0__abc_74894_new_n3596_), .C(u0__abc_74894_new_n3632_), .Y(u0__abc_74894_new_n3633_));
NAND3X1 NAND3X1_305 ( .A(u0__abc_74894_new_n3694_), .B(u0__abc_74894_new_n3697_), .C(u0__abc_74894_new_n3702_), .Y(u0__abc_74894_new_n3703_));
NAND3X1 NAND3X1_306 ( .A(u0__abc_74894_new_n3721_), .B(u0__abc_74894_new_n3709_), .C(u0__abc_74894_new_n3714_), .Y(u0__abc_74894_new_n3722_));
NAND3X1 NAND3X1_307 ( .A(\wb_addr_i[3] ), .B(u0__abc_74894_new_n3691_), .C(u0__abc_74894_new_n3731_), .Y(u0__abc_74894_new_n3732_));
NAND3X1 NAND3X1_308 ( .A(u0__abc_74894_new_n3742_), .B(u0__abc_74894_new_n3744_), .C(u0__abc_74894_new_n3746_), .Y(u0__abc_74894_new_n3747_));
NAND3X1 NAND3X1_309 ( .A(u0__abc_74894_new_n3754_), .B(u0__abc_74894_new_n3723_), .C(u0__abc_74894_new_n3740_), .Y(rf_dout_0_));
NAND3X1 NAND3X1_31 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1300_), .C(u0__abc_74894_new_n1303_), .Y(u0__abc_74894_new_n1304_));
NAND3X1 NAND3X1_310 ( .A(u0__abc_74894_new_n3768_), .B(u0__abc_74894_new_n3762_), .C(u0__abc_74894_new_n3776_), .Y(rf_dout_1_));
NAND3X1 NAND3X1_311 ( .A(u0__abc_74894_new_n3789_), .B(u0__abc_74894_new_n3784_), .C(u0__abc_74894_new_n3795_), .Y(rf_dout_2_));
NAND3X1 NAND3X1_312 ( .A(u0__abc_74894_new_n3807_), .B(u0__abc_74894_new_n3808_), .C(u0__abc_74894_new_n3806_), .Y(u0__abc_74894_new_n3809_));
NAND3X1 NAND3X1_313 ( .A(u0__abc_74894_new_n3811_), .B(u0__abc_74894_new_n3812_), .C(u0__abc_74894_new_n3810_), .Y(u0__abc_74894_new_n3813_));
NAND3X1 NAND3X1_314 ( .A(u0__abc_74894_new_n3820_), .B(u0__abc_74894_new_n3814_), .C(u0__abc_74894_new_n3805_), .Y(rf_dout_3_));
NAND3X1 NAND3X1_315 ( .A(u0__abc_74894_new_n3822_), .B(u0__abc_74894_new_n3823_), .C(u0__abc_74894_new_n3824_), .Y(u0__abc_74894_new_n3825_));
NAND3X1 NAND3X1_316 ( .A(u0__abc_74894_new_n3829_), .B(u0__abc_74894_new_n3832_), .C(u0__abc_74894_new_n3838_), .Y(rf_dout_4_));
NAND3X1 NAND3X1_317 ( .A(u0__abc_74894_new_n3849_), .B(u0__abc_74894_new_n3850_), .C(u0__abc_74894_new_n3851_), .Y(u0__abc_74894_new_n3852_));
NAND3X1 NAND3X1_318 ( .A(u0__abc_74894_new_n3855_), .B(u0__abc_74894_new_n3854_), .C(u0__abc_74894_new_n3853_), .Y(u0__abc_74894_new_n3856_));
NAND3X1 NAND3X1_319 ( .A(u0__abc_74894_new_n3848_), .B(u0__abc_74894_new_n3861_), .C(u0__abc_74894_new_n3857_), .Y(rf_dout_5_));
NAND3X1 NAND3X1_32 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1305_), .C(u0__abc_74894_new_n1304_), .Y(u0__abc_74894_new_n1306_));
NAND3X1 NAND3X1_320 ( .A(u0__abc_74894_new_n3863_), .B(u0__abc_74894_new_n3864_), .C(u0__abc_74894_new_n3865_), .Y(u0__abc_74894_new_n3866_));
NAND3X1 NAND3X1_321 ( .A(u0__abc_74894_new_n3870_), .B(u0__abc_74894_new_n3873_), .C(u0__abc_74894_new_n3879_), .Y(rf_dout_6_));
NAND3X1 NAND3X1_322 ( .A(u0__abc_74894_new_n3885_), .B(u0__abc_74894_new_n3887_), .C(u0__abc_74894_new_n3886_), .Y(u0__abc_74894_new_n3888_));
NAND3X1 NAND3X1_323 ( .A(u0__abc_74894_new_n3893_), .B(u0__abc_74894_new_n3894_), .C(u0__abc_74894_new_n3896_), .Y(u0__abc_74894_new_n3897_));
NAND3X1 NAND3X1_324 ( .A(u0__abc_74894_new_n3883_), .B(u0__abc_74894_new_n3889_), .C(u0__abc_74894_new_n3898_), .Y(rf_dout_7_));
NAND3X1 NAND3X1_325 ( .A(u0__abc_74894_new_n3900_), .B(u0__abc_74894_new_n3901_), .C(u0__abc_74894_new_n3902_), .Y(u0__abc_74894_new_n3903_));
NAND3X1 NAND3X1_326 ( .A(u0__abc_74894_new_n3911_), .B(u0__abc_74894_new_n3912_), .C(u0__abc_74894_new_n3914_), .Y(u0__abc_74894_new_n3915_));
NAND3X1 NAND3X1_327 ( .A(u0__abc_74894_new_n3907_), .B(u0__abc_74894_new_n3910_), .C(u0__abc_74894_new_n3916_), .Y(rf_dout_8_));
NAND3X1 NAND3X1_328 ( .A(u0__abc_74894_new_n3925_), .B(u0__abc_74894_new_n3926_), .C(u0__abc_74894_new_n3927_), .Y(u0__abc_74894_new_n3928_));
NAND3X1 NAND3X1_329 ( .A(u0__abc_74894_new_n3930_), .B(u0__abc_74894_new_n3931_), .C(u0__abc_74894_new_n3929_), .Y(u0__abc_74894_new_n3932_));
NAND3X1 NAND3X1_33 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1298_), .C(u0__abc_74894_new_n1306_), .Y(u0__abc_74894_new_n1307_));
NAND3X1 NAND3X1_330 ( .A(u0__abc_74894_new_n3937_), .B(u0__abc_74894_new_n3933_), .C(u0__abc_74894_new_n3924_), .Y(rf_dout_9_));
NAND3X1 NAND3X1_331 ( .A(u0__abc_74894_new_n3939_), .B(u0__abc_74894_new_n3940_), .C(u0__abc_74894_new_n3941_), .Y(u0__abc_74894_new_n3942_));
NAND3X1 NAND3X1_332 ( .A(u0__abc_74894_new_n3946_), .B(u0__abc_74894_new_n3949_), .C(u0__abc_74894_new_n3955_), .Y(rf_dout_10_));
NAND3X1 NAND3X1_333 ( .A(u0__abc_74894_new_n3958_), .B(u0__abc_74894_new_n3959_), .C(u0__abc_74894_new_n3960_), .Y(u0__abc_74894_new_n3961_));
NAND3X1 NAND3X1_334 ( .A(u0__abc_74894_new_n3962_), .B(u0__abc_74894_new_n3963_), .C(u0__abc_74894_new_n3964_), .Y(u0__abc_74894_new_n3965_));
NAND3X1 NAND3X1_335 ( .A(u0__abc_74894_new_n3970_), .B(u0__abc_74894_new_n3971_), .C(u0__abc_74894_new_n3972_), .Y(u0__abc_74894_new_n3973_));
NAND3X1 NAND3X1_336 ( .A(u0__abc_74894_new_n3957_), .B(u0__abc_74894_new_n3966_), .C(u0__abc_74894_new_n3974_), .Y(rf_dout_11_));
NAND3X1 NAND3X1_337 ( .A(u0__abc_74894_new_n3977_), .B(u0__abc_74894_new_n3978_), .C(u0__abc_74894_new_n3979_), .Y(u0__abc_74894_new_n3980_));
NAND3X1 NAND3X1_338 ( .A(u0__abc_74894_new_n3981_), .B(u0__abc_74894_new_n3982_), .C(u0__abc_74894_new_n3983_), .Y(u0__abc_74894_new_n3984_));
NAND3X1 NAND3X1_339 ( .A(u0__abc_74894_new_n3989_), .B(u0__abc_74894_new_n3990_), .C(u0__abc_74894_new_n3991_), .Y(u0__abc_74894_new_n3992_));
NAND3X1 NAND3X1_34 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1322_), .C(u0__abc_74894_new_n1321_), .Y(u0__abc_74894_new_n1323_));
NAND3X1 NAND3X1_340 ( .A(u0__abc_74894_new_n3976_), .B(u0__abc_74894_new_n3985_), .C(u0__abc_74894_new_n3993_), .Y(rf_dout_12_));
NAND3X1 NAND3X1_341 ( .A(u0__abc_74894_new_n3995_), .B(u0__abc_74894_new_n3996_), .C(u0__abc_74894_new_n3997_), .Y(u0__abc_74894_new_n3998_));
NAND3X1 NAND3X1_342 ( .A(u0__abc_74894_new_n4011_), .B(u0__abc_74894_new_n4013_), .C(u0__abc_74894_new_n4012_), .Y(u0__abc_74894_new_n4014_));
NAND3X1 NAND3X1_343 ( .A(u0__abc_74894_new_n4000_), .B(u0__abc_74894_new_n4015_), .C(u0__abc_74894_new_n4008_), .Y(rf_dout_13_));
NAND3X1 NAND3X1_344 ( .A(u0__abc_74894_new_n4018_), .B(u0__abc_74894_new_n4019_), .C(u0__abc_74894_new_n4017_), .Y(u0__abc_74894_new_n4020_));
NAND3X1 NAND3X1_345 ( .A(u0__abc_74894_new_n4033_), .B(u0__abc_74894_new_n4035_), .C(u0__abc_74894_new_n4034_), .Y(u0__abc_74894_new_n4036_));
NAND3X1 NAND3X1_346 ( .A(u0__abc_74894_new_n4022_), .B(u0__abc_74894_new_n4037_), .C(u0__abc_74894_new_n4030_), .Y(rf_dout_14_));
NAND3X1 NAND3X1_347 ( .A(u0__abc_74894_new_n4047_), .B(u0__abc_74894_new_n4048_), .C(u0__abc_74894_new_n4049_), .Y(u0__abc_74894_new_n4050_));
NAND3X1 NAND3X1_348 ( .A(u0__abc_74894_new_n4051_), .B(u0__abc_74894_new_n4059_), .C(u0__abc_74894_new_n4046_), .Y(rf_dout_15_));
NAND3X1 NAND3X1_349 ( .A(u0__abc_74894_new_n4064_), .B(u0__abc_74894_new_n4065_), .C(u0__abc_74894_new_n4063_), .Y(u0__abc_74894_new_n4066_));
NAND3X1 NAND3X1_35 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1320_), .C(u0__abc_74894_new_n1323_), .Y(u0__abc_74894_new_n1324_));
NAND3X1 NAND3X1_350 ( .A(u0__abc_74894_new_n4072_), .B(u0__abc_74894_new_n4073_), .C(u0__abc_74894_new_n4071_), .Y(u0__abc_74894_new_n4074_));
NAND3X1 NAND3X1_351 ( .A(u0__abc_74894_new_n4076_), .B(u0__abc_74894_new_n4077_), .C(u0__abc_74894_new_n4075_), .Y(u0__abc_74894_new_n4078_));
NAND3X1 NAND3X1_352 ( .A(u0__abc_74894_new_n4070_), .B(u0__abc_74894_new_n4067_), .C(u0__abc_74894_new_n4079_), .Y(rf_dout_16_));
NAND3X1 NAND3X1_353 ( .A(u0__abc_74894_new_n4089_), .B(u0__abc_74894_new_n4091_), .C(u0__abc_74894_new_n4090_), .Y(u0__abc_74894_new_n4092_));
NAND3X1 NAND3X1_354 ( .A(u0__abc_74894_new_n4093_), .B(u0__abc_74894_new_n4101_), .C(u0__abc_74894_new_n4088_), .Y(rf_dout_17_));
NAND3X1 NAND3X1_355 ( .A(u0__abc_74894_new_n4112_), .B(u0__abc_74894_new_n4113_), .C(u0__abc_74894_new_n4111_), .Y(u0__abc_74894_new_n4114_));
NAND3X1 NAND3X1_356 ( .A(u0__abc_74894_new_n4115_), .B(u0__abc_74894_new_n4123_), .C(u0__abc_74894_new_n4110_), .Y(rf_dout_18_));
NAND3X1 NAND3X1_357 ( .A(u0__abc_74894_new_n4125_), .B(u0__abc_74894_new_n4126_), .C(u0__abc_74894_new_n4127_), .Y(u0__abc_74894_new_n4128_));
NAND3X1 NAND3X1_358 ( .A(u0__abc_74894_new_n4143_), .B(u0__abc_74894_new_n4141_), .C(u0__abc_74894_new_n4142_), .Y(u0__abc_74894_new_n4144_));
NAND3X1 NAND3X1_359 ( .A(u0__abc_74894_new_n4130_), .B(u0__abc_74894_new_n4145_), .C(u0__abc_74894_new_n4138_), .Y(rf_dout_19_));
NAND3X1 NAND3X1_36 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1325_), .C(u0__abc_74894_new_n1324_), .Y(u0__abc_74894_new_n1326_));
NAND3X1 NAND3X1_360 ( .A(u0__abc_74894_new_n4148_), .B(u0__abc_74894_new_n4149_), .C(u0__abc_74894_new_n4150_), .Y(u0__abc_74894_new_n4151_));
NAND3X1 NAND3X1_361 ( .A(u0__abc_74894_new_n4152_), .B(u0__abc_74894_new_n4153_), .C(u0__abc_74894_new_n4154_), .Y(u0__abc_74894_new_n4155_));
NAND3X1 NAND3X1_362 ( .A(u0__abc_74894_new_n4160_), .B(u0__abc_74894_new_n4161_), .C(u0__abc_74894_new_n4162_), .Y(u0__abc_74894_new_n4163_));
NAND3X1 NAND3X1_363 ( .A(u0__abc_74894_new_n4147_), .B(u0__abc_74894_new_n4156_), .C(u0__abc_74894_new_n4164_), .Y(rf_dout_20_));
NAND3X1 NAND3X1_364 ( .A(u0__abc_74894_new_n4167_), .B(u0__abc_74894_new_n4168_), .C(u0__abc_74894_new_n4166_), .Y(u0__abc_74894_new_n4169_));
NAND3X1 NAND3X1_365 ( .A(u0__abc_74894_new_n4185_), .B(u0__abc_74894_new_n4183_), .C(u0__abc_74894_new_n4184_), .Y(u0__abc_74894_new_n4186_));
NAND3X1 NAND3X1_366 ( .A(u0__abc_74894_new_n4172_), .B(u0__abc_74894_new_n4187_), .C(u0__abc_74894_new_n4180_), .Y(rf_dout_21_));
NAND3X1 NAND3X1_367 ( .A(u0__abc_74894_new_n4190_), .B(u0__abc_74894_new_n4191_), .C(u0__abc_74894_new_n4192_), .Y(u0__abc_74894_new_n4193_));
NAND3X1 NAND3X1_368 ( .A(u0__abc_74894_new_n4194_), .B(u0__abc_74894_new_n4195_), .C(u0__abc_74894_new_n4196_), .Y(u0__abc_74894_new_n4197_));
NAND3X1 NAND3X1_369 ( .A(u0__abc_74894_new_n4202_), .B(u0__abc_74894_new_n4203_), .C(u0__abc_74894_new_n4204_), .Y(u0__abc_74894_new_n4205_));
NAND3X1 NAND3X1_37 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1318_), .C(u0__abc_74894_new_n1326_), .Y(u0__abc_74894_new_n1327_));
NAND3X1 NAND3X1_370 ( .A(u0__abc_74894_new_n4189_), .B(u0__abc_74894_new_n4198_), .C(u0__abc_74894_new_n4206_), .Y(rf_dout_22_));
NAND3X1 NAND3X1_371 ( .A(u0__abc_74894_new_n4211_), .B(u0__abc_74894_new_n4212_), .C(u0__abc_74894_new_n4210_), .Y(u0__abc_74894_new_n4213_));
NAND3X1 NAND3X1_372 ( .A(u0__abc_74894_new_n4219_), .B(u0__abc_74894_new_n4220_), .C(u0__abc_74894_new_n4218_), .Y(u0__abc_74894_new_n4221_));
NAND3X1 NAND3X1_373 ( .A(u0__abc_74894_new_n4223_), .B(u0__abc_74894_new_n4224_), .C(u0__abc_74894_new_n4222_), .Y(u0__abc_74894_new_n4225_));
NAND3X1 NAND3X1_374 ( .A(u0__abc_74894_new_n4217_), .B(u0__abc_74894_new_n4214_), .C(u0__abc_74894_new_n4226_), .Y(rf_dout_23_));
NAND3X1 NAND3X1_375 ( .A(u0__abc_74894_new_n4229_), .B(u0__abc_74894_new_n4228_), .C(u0__abc_74894_new_n4230_), .Y(u0__abc_74894_new_n4231_));
NAND3X1 NAND3X1_376 ( .A(u0__abc_74894_new_n4232_), .B(u0__abc_74894_new_n4233_), .C(u0__abc_74894_new_n4234_), .Y(u0__abc_74894_new_n4235_));
NAND3X1 NAND3X1_377 ( .A(u0__abc_74894_new_n4239_), .B(u0__abc_74894_new_n4237_), .C(u0__abc_74894_new_n4238_), .Y(u0__abc_74894_new_n4240_));
NAND3X1 NAND3X1_378 ( .A(u0__abc_74894_new_n4243_), .B(u0__abc_74894_new_n4242_), .C(u0__abc_74894_new_n4244_), .Y(u0__abc_74894_new_n4245_));
NAND3X1 NAND3X1_379 ( .A(u0__abc_74894_new_n4246_), .B(u0__abc_74894_new_n4248_), .C(u0__abc_74894_new_n4247_), .Y(u0__abc_74894_new_n4249_));
NAND3X1 NAND3X1_38 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1342_), .C(u0__abc_74894_new_n1341_), .Y(u0__abc_74894_new_n1343_));
NAND3X1 NAND3X1_380 ( .A(u0__abc_74894_new_n4236_), .B(u0__abc_74894_new_n4241_), .C(u0__abc_74894_new_n4252_), .Y(rf_dout_24_));
NAND3X1 NAND3X1_381 ( .A(u0__abc_74894_new_n4255_), .B(u0__abc_74894_new_n4254_), .C(u0__abc_74894_new_n4256_), .Y(u0__abc_74894_new_n4257_));
NAND3X1 NAND3X1_382 ( .A(u0__abc_74894_new_n4258_), .B(u0__abc_74894_new_n4260_), .C(u0__abc_74894_new_n4259_), .Y(u0__abc_74894_new_n4261_));
NAND3X1 NAND3X1_383 ( .A(u0__abc_74894_new_n4265_), .B(u0__abc_74894_new_n4263_), .C(u0__abc_74894_new_n4264_), .Y(u0__abc_74894_new_n4266_));
NAND3X1 NAND3X1_384 ( .A(u0__abc_74894_new_n4270_), .B(u0__abc_74894_new_n4268_), .C(u0__abc_74894_new_n4269_), .Y(u0__abc_74894_new_n4271_));
NAND3X1 NAND3X1_385 ( .A(u0__abc_74894_new_n4262_), .B(u0__abc_74894_new_n4267_), .C(u0__abc_74894_new_n4278_), .Y(rf_dout_25_));
NAND3X1 NAND3X1_386 ( .A(u0__abc_74894_new_n4281_), .B(u0__abc_74894_new_n4280_), .C(u0__abc_74894_new_n4282_), .Y(u0__abc_74894_new_n4283_));
NAND3X1 NAND3X1_387 ( .A(u0__abc_74894_new_n4284_), .B(u0__abc_74894_new_n4286_), .C(u0__abc_74894_new_n4285_), .Y(u0__abc_74894_new_n4287_));
NAND3X1 NAND3X1_388 ( .A(u0__abc_74894_new_n4290_), .B(u0__abc_74894_new_n4291_), .C(u0__abc_74894_new_n4289_), .Y(u0__abc_74894_new_n4292_));
NAND3X1 NAND3X1_389 ( .A(u0__abc_74894_new_n4295_), .B(u0__abc_74894_new_n4294_), .C(u0__abc_74894_new_n4296_), .Y(u0__abc_74894_new_n4297_));
NAND3X1 NAND3X1_39 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1340_), .C(u0__abc_74894_new_n1343_), .Y(u0__abc_74894_new_n1344_));
NAND3X1 NAND3X1_390 ( .A(u0__abc_74894_new_n4299_), .B(u0__abc_74894_new_n4300_), .C(u0__abc_74894_new_n4298_), .Y(u0__abc_74894_new_n4301_));
NAND3X1 NAND3X1_391 ( .A(u0__abc_74894_new_n4288_), .B(u0__abc_74894_new_n4293_), .C(u0__abc_74894_new_n4304_), .Y(rf_dout_26_));
NAND3X1 NAND3X1_392 ( .A(u0__abc_74894_new_n4307_), .B(u0__abc_74894_new_n4306_), .C(u0__abc_74894_new_n4308_), .Y(u0__abc_74894_new_n4309_));
NAND3X1 NAND3X1_393 ( .A(u0__abc_74894_new_n4310_), .B(u0__abc_74894_new_n4312_), .C(u0__abc_74894_new_n4311_), .Y(u0__abc_74894_new_n4313_));
NAND3X1 NAND3X1_394 ( .A(u0__abc_74894_new_n4315_), .B(u0__abc_74894_new_n4317_), .C(u0__abc_74894_new_n4316_), .Y(u0__abc_74894_new_n4318_));
NAND3X1 NAND3X1_395 ( .A(u0__abc_74894_new_n4321_), .B(u0__abc_74894_new_n4320_), .C(u0__abc_74894_new_n4322_), .Y(u0__abc_74894_new_n4323_));
NAND3X1 NAND3X1_396 ( .A(u0__abc_74894_new_n4325_), .B(u0__abc_74894_new_n4324_), .C(u0__abc_74894_new_n4326_), .Y(u0__abc_74894_new_n4327_));
NAND3X1 NAND3X1_397 ( .A(u0__abc_74894_new_n4314_), .B(u0__abc_74894_new_n4319_), .C(u0__abc_74894_new_n4331_), .Y(rf_dout_27_));
NAND3X1 NAND3X1_398 ( .A(u0__abc_74894_new_n4334_), .B(u0__abc_74894_new_n4333_), .C(u0__abc_74894_new_n4335_), .Y(u0__abc_74894_new_n4336_));
NAND3X1 NAND3X1_399 ( .A(u0__abc_74894_new_n4337_), .B(u0__abc_74894_new_n4339_), .C(u0__abc_74894_new_n4338_), .Y(u0__abc_74894_new_n4340_));
NAND3X1 NAND3X1_4 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1165_), .C(u0__abc_74894_new_n1164_), .Y(u0__abc_74894_new_n1166_));
NAND3X1 NAND3X1_40 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1345_), .C(u0__abc_74894_new_n1344_), .Y(u0__abc_74894_new_n1346_));
NAND3X1 NAND3X1_400 ( .A(u0__abc_74894_new_n4343_), .B(u0__abc_74894_new_n4342_), .C(u0__abc_74894_new_n4344_), .Y(u0__abc_74894_new_n4345_));
NAND3X1 NAND3X1_401 ( .A(u0__abc_74894_new_n4347_), .B(u0__abc_74894_new_n4348_), .C(u0__abc_74894_new_n4349_), .Y(u0__abc_74894_new_n4350_));
NAND3X1 NAND3X1_402 ( .A(u0__abc_74894_new_n4352_), .B(u0__abc_74894_new_n4353_), .C(u0__abc_74894_new_n4351_), .Y(u0__abc_74894_new_n4354_));
NAND3X1 NAND3X1_403 ( .A(u0__abc_74894_new_n4341_), .B(u0__abc_74894_new_n4346_), .C(u0__abc_74894_new_n4357_), .Y(rf_dout_28_));
NAND3X1 NAND3X1_404 ( .A(u0__abc_74894_new_n4360_), .B(u0__abc_74894_new_n4359_), .C(u0__abc_74894_new_n4361_), .Y(u0__abc_74894_new_n4362_));
NAND3X1 NAND3X1_405 ( .A(u0__abc_74894_new_n4368_), .B(u0__abc_74894_new_n4369_), .C(u0__abc_74894_new_n4367_), .Y(u0__abc_74894_new_n4370_));
NAND3X1 NAND3X1_406 ( .A(u0__abc_74894_new_n4374_), .B(u0__abc_74894_new_n4375_), .C(u0__abc_74894_new_n4373_), .Y(u0__abc_74894_new_n4376_));
NAND3X1 NAND3X1_407 ( .A(u0__abc_74894_new_n4378_), .B(u0__abc_74894_new_n4377_), .C(u0__abc_74894_new_n4379_), .Y(u0__abc_74894_new_n4380_));
NAND3X1 NAND3X1_408 ( .A(u0__abc_74894_new_n4371_), .B(u0__abc_74894_new_n4366_), .C(u0__abc_74894_new_n4381_), .Y(rf_dout_29_));
NAND3X1 NAND3X1_409 ( .A(u0__abc_74894_new_n4384_), .B(u0__abc_74894_new_n4383_), .C(u0__abc_74894_new_n4385_), .Y(u0__abc_74894_new_n4386_));
NAND3X1 NAND3X1_41 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1338_), .C(u0__abc_74894_new_n1346_), .Y(u0__abc_74894_new_n1347_));
NAND3X1 NAND3X1_410 ( .A(u0__abc_74894_new_n4392_), .B(u0__abc_74894_new_n4391_), .C(u0__abc_74894_new_n4393_), .Y(u0__abc_74894_new_n4394_));
NAND3X1 NAND3X1_411 ( .A(u0__abc_74894_new_n4398_), .B(u0__abc_74894_new_n4399_), .C(u0__abc_74894_new_n4397_), .Y(u0__abc_74894_new_n4400_));
NAND3X1 NAND3X1_412 ( .A(u0__abc_74894_new_n4403_), .B(u0__abc_74894_new_n4401_), .C(u0__abc_74894_new_n4402_), .Y(u0__abc_74894_new_n4404_));
NAND3X1 NAND3X1_413 ( .A(u0__abc_74894_new_n4395_), .B(u0__abc_74894_new_n4390_), .C(u0__abc_74894_new_n4405_), .Y(rf_dout_30_));
NAND3X1 NAND3X1_414 ( .A(u0__abc_74894_new_n4408_), .B(u0__abc_74894_new_n4407_), .C(u0__abc_74894_new_n4409_), .Y(u0__abc_74894_new_n4410_));
NAND3X1 NAND3X1_415 ( .A(u0__abc_74894_new_n4416_), .B(u0__abc_74894_new_n4415_), .C(u0__abc_74894_new_n4417_), .Y(u0__abc_74894_new_n4418_));
NAND3X1 NAND3X1_416 ( .A(u0__abc_74894_new_n4422_), .B(u0__abc_74894_new_n4423_), .C(u0__abc_74894_new_n4421_), .Y(u0__abc_74894_new_n4424_));
NAND3X1 NAND3X1_417 ( .A(u0__abc_74894_new_n4427_), .B(u0__abc_74894_new_n4425_), .C(u0__abc_74894_new_n4426_), .Y(u0__abc_74894_new_n4428_));
NAND3X1 NAND3X1_418 ( .A(u0__abc_74894_new_n4419_), .B(u0__abc_74894_new_n4414_), .C(u0__abc_74894_new_n4429_), .Y(rf_dout_31_));
NAND3X1 NAND3X1_419 ( .A(wb_we_i), .B(u0__abc_74894_new_n1154_), .C(u0__abc_74894_new_n4432_), .Y(u0__abc_74894_new_n4433_));
NAND3X1 NAND3X1_42 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1362_), .C(u0__abc_74894_new_n1361_), .Y(u0__abc_74894_new_n1363_));
NAND3X1 NAND3X1_420 ( .A(u0__abc_74894_new_n4465_), .B(u0__abc_74894_new_n4462_), .C(u0__abc_74894_new_n4464_), .Y(u0__0sreq_cs_le_0_0_));
NAND3X1 NAND3X1_421 ( .A(u0__abc_74894_new_n4470_), .B(u0__abc_74894_new_n4471_), .C(u0__abc_74894_new_n4469_), .Y(u0__0init_req_0_0_));
NAND3X1 NAND3X1_422 ( .A(u0__abc_74894_new_n1102_), .B(u0__abc_74894_new_n1108_), .C(u0__abc_74894_new_n1113_), .Y(u0__abc_74894_new_n4473_));
NAND3X1 NAND3X1_423 ( .A(u0__abc_74894_new_n4475_), .B(u0__abc_74894_new_n4476_), .C(u0__abc_74894_new_n4474_), .Y(u0__0lmr_req_0_0_));
NAND3X1 NAND3X1_424 ( .A(u0_rf_we), .B(u0_u0__abc_72207_new_n216_), .C(u0_u0__abc_72207_new_n217_), .Y(u0_u0__abc_72207_new_n218_));
NAND3X1 NAND3X1_425 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[0] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n222_));
NAND3X1 NAND3X1_426 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[1] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n225_));
NAND3X1 NAND3X1_427 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[2] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n228_));
NAND3X1 NAND3X1_428 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[3] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n231_));
NAND3X1 NAND3X1_429 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[4] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n234_));
NAND3X1 NAND3X1_43 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1360_), .C(u0__abc_74894_new_n1363_), .Y(u0__abc_74894_new_n1364_));
NAND3X1 NAND3X1_430 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[5] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n237_));
NAND3X1 NAND3X1_431 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[6] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n240_));
NAND3X1 NAND3X1_432 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[7] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n243_));
NAND3X1 NAND3X1_433 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[8] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n246_));
NAND3X1 NAND3X1_434 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[9] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n249_));
NAND3X1 NAND3X1_435 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[10] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n252_));
NAND3X1 NAND3X1_436 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[11] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n255_));
NAND3X1 NAND3X1_437 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[12] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n258_));
NAND3X1 NAND3X1_438 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[13] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n261_));
NAND3X1 NAND3X1_439 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[14] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n264_));
NAND3X1 NAND3X1_44 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1365_), .C(u0__abc_74894_new_n1364_), .Y(u0__abc_74894_new_n1366_));
NAND3X1 NAND3X1_440 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[15] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n267_));
NAND3X1 NAND3X1_441 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[16] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n270_));
NAND3X1 NAND3X1_442 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[17] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n273_));
NAND3X1 NAND3X1_443 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[18] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n276_));
NAND3X1 NAND3X1_444 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[19] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n279_));
NAND3X1 NAND3X1_445 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[20] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n282_));
NAND3X1 NAND3X1_446 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[21] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n285_));
NAND3X1 NAND3X1_447 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[22] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n288_));
NAND3X1 NAND3X1_448 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[23] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n291_));
NAND3X1 NAND3X1_449 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[24] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n294_));
NAND3X1 NAND3X1_45 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1358_), .C(u0__abc_74894_new_n1366_), .Y(u0__abc_74894_new_n1367_));
NAND3X1 NAND3X1_450 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[25] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n297_));
NAND3X1 NAND3X1_451 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[26] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n300_));
NAND3X1 NAND3X1_452 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[27] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n303_));
NAND3X1 NAND3X1_453 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[28] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n306_));
NAND3X1 NAND3X1_454 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[29] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n309_));
NAND3X1 NAND3X1_455 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[30] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n312_));
NAND3X1 NAND3X1_456 ( .A(u0_u0_addr_r_2_), .B(\wb_data_i[31] ), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n315_));
NAND3X1 NAND3X1_457 ( .A(u0_u0__abc_72207_new_n318_), .B(u0_u0__abc_72207_new_n319_), .C(u0_u0__abc_72207_new_n321_), .Y(u0_u0__abc_72207_new_n322_));
NAND3X1 NAND3X1_458 ( .A(u0_u0__abc_72207_new_n318_), .B(u0_u0__abc_72207_new_n327_), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n328_));
NAND3X1 NAND3X1_459 ( .A(u0_u0__abc_72207_new_n324_), .B(u0_u0__abc_72207_new_n328_), .C(u0_u0__abc_72207_new_n326_), .Y(u0_u0__abc_72207_new_n329_));
NAND3X1 NAND3X1_46 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1382_), .C(u0__abc_74894_new_n1381_), .Y(u0__abc_74894_new_n1383_));
NAND3X1 NAND3X1_460 ( .A(u0_u0__abc_72207_new_n318_), .B(u0_u0__abc_72207_new_n345_), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n346_));
NAND3X1 NAND3X1_461 ( .A(u0_u0__abc_72207_new_n324_), .B(u0_u0__abc_72207_new_n346_), .C(u0_u0__abc_72207_new_n344_), .Y(u0_u0__abc_72207_new_n347_));
NAND3X1 NAND3X1_462 ( .A(u0_u0__abc_72207_new_n318_), .B(u0_u0__abc_72207_new_n352_), .C(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n353_));
NAND3X1 NAND3X1_463 ( .A(u0_u0__abc_72207_new_n324_), .B(u0_u0__abc_72207_new_n353_), .C(u0_u0__abc_72207_new_n351_), .Y(u0_u0__abc_72207_new_n354_));
NAND3X1 NAND3X1_464 ( .A(u0_u0__abc_72207_new_n440_), .B(u0_u0__abc_72207_new_n448_), .C(u0_u0__abc_72207_new_n457_), .Y(u0_u0__abc_72207_new_n458_));
NAND3X1 NAND3X1_465 ( .A(u0_u1_addr_r_4_), .B(u0_u1_addr_r_3_), .C(u0_u1__abc_72470_new_n213_), .Y(u0_u1__abc_72470_new_n214_));
NAND3X1 NAND3X1_466 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[0] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n218_));
NAND3X1 NAND3X1_467 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[1] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n221_));
NAND3X1 NAND3X1_468 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[2] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n224_));
NAND3X1 NAND3X1_469 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[3] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n227_));
NAND3X1 NAND3X1_47 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1380_), .C(u0__abc_74894_new_n1383_), .Y(u0__abc_74894_new_n1384_));
NAND3X1 NAND3X1_470 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[4] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n230_));
NAND3X1 NAND3X1_471 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[5] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n233_));
NAND3X1 NAND3X1_472 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[6] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n236_));
NAND3X1 NAND3X1_473 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[7] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n239_));
NAND3X1 NAND3X1_474 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[8] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n242_));
NAND3X1 NAND3X1_475 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[9] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n245_));
NAND3X1 NAND3X1_476 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[10] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n248_));
NAND3X1 NAND3X1_477 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[11] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n251_));
NAND3X1 NAND3X1_478 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[12] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n254_));
NAND3X1 NAND3X1_479 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[13] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n257_));
NAND3X1 NAND3X1_48 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1385_), .C(u0__abc_74894_new_n1384_), .Y(u0__abc_74894_new_n1386_));
NAND3X1 NAND3X1_480 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[14] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n260_));
NAND3X1 NAND3X1_481 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[15] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n263_));
NAND3X1 NAND3X1_482 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[16] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n266_));
NAND3X1 NAND3X1_483 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[17] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n269_));
NAND3X1 NAND3X1_484 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[18] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n272_));
NAND3X1 NAND3X1_485 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[19] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n275_));
NAND3X1 NAND3X1_486 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[20] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n278_));
NAND3X1 NAND3X1_487 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[21] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n281_));
NAND3X1 NAND3X1_488 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[22] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n284_));
NAND3X1 NAND3X1_489 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[23] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n287_));
NAND3X1 NAND3X1_49 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1378_), .C(u0__abc_74894_new_n1386_), .Y(u0__abc_74894_new_n1387_));
NAND3X1 NAND3X1_490 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[24] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n290_));
NAND3X1 NAND3X1_491 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[25] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n293_));
NAND3X1 NAND3X1_492 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[26] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n296_));
NAND3X1 NAND3X1_493 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[27] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n299_));
NAND3X1 NAND3X1_494 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[28] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n302_));
NAND3X1 NAND3X1_495 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[29] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n305_));
NAND3X1 NAND3X1_496 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[30] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n308_));
NAND3X1 NAND3X1_497 ( .A(u0_u1_addr_r_2_), .B(\wb_data_i[31] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n311_));
NAND3X1 NAND3X1_498 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[0] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n315_));
NAND3X1 NAND3X1_499 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[1] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n318_));
NAND3X1 NAND3X1_5 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1158_), .C(u0__abc_74894_new_n1166_), .Y(u0__abc_74894_new_n1167_));
NAND3X1 NAND3X1_50 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1402_), .C(u0__abc_74894_new_n1401_), .Y(u0__abc_74894_new_n1403_));
NAND3X1 NAND3X1_500 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[2] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n321_));
NAND3X1 NAND3X1_501 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[3] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n324_));
NAND3X1 NAND3X1_502 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[4] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n327_));
NAND3X1 NAND3X1_503 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[5] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n330_));
NAND3X1 NAND3X1_504 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[6] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n333_));
NAND3X1 NAND3X1_505 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[7] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n336_));
NAND3X1 NAND3X1_506 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[8] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n339_));
NAND3X1 NAND3X1_507 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[9] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n342_));
NAND3X1 NAND3X1_508 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[10] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n345_));
NAND3X1 NAND3X1_509 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[11] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n348_));
NAND3X1 NAND3X1_51 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1400_), .C(u0__abc_74894_new_n1403_), .Y(u0__abc_74894_new_n1404_));
NAND3X1 NAND3X1_510 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[12] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n351_));
NAND3X1 NAND3X1_511 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[13] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n354_));
NAND3X1 NAND3X1_512 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[14] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n357_));
NAND3X1 NAND3X1_513 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[15] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n360_));
NAND3X1 NAND3X1_514 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[16] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n363_));
NAND3X1 NAND3X1_515 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[17] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n366_));
NAND3X1 NAND3X1_516 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[18] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n369_));
NAND3X1 NAND3X1_517 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[19] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n372_));
NAND3X1 NAND3X1_518 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[20] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n375_));
NAND3X1 NAND3X1_519 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[21] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n378_));
NAND3X1 NAND3X1_52 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1405_), .C(u0__abc_74894_new_n1404_), .Y(u0__abc_74894_new_n1406_));
NAND3X1 NAND3X1_520 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[22] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n381_));
NAND3X1 NAND3X1_521 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[23] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n384_));
NAND3X1 NAND3X1_522 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[24] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n387_));
NAND3X1 NAND3X1_523 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[25] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n390_));
NAND3X1 NAND3X1_524 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[26] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n393_));
NAND3X1 NAND3X1_525 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[27] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n396_));
NAND3X1 NAND3X1_526 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[28] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n399_));
NAND3X1 NAND3X1_527 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[29] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n402_));
NAND3X1 NAND3X1_528 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[30] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n405_));
NAND3X1 NAND3X1_529 ( .A(u0_u1__abc_72470_new_n210_), .B(\wb_data_i[31] ), .C(u0_u1__abc_72470_new_n217_), .Y(u0_u1__abc_72470_new_n408_));
NAND3X1 NAND3X1_53 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1398_), .C(u0__abc_74894_new_n1406_), .Y(u0__abc_74894_new_n1407_));
NAND3X1 NAND3X1_530 ( .A(u0_u1__abc_72470_new_n417_), .B(u0_u1__abc_72470_new_n424_), .C(u0_u1__abc_72470_new_n433_), .Y(u0_u1__abc_72470_new_n434_));
NAND3X1 NAND3X1_531 ( .A(u0_csc1_0_), .B(u0_u1_init_req_we), .C(u0_u1__abc_72470_new_n439_), .Y(u0_u1__abc_72470_new_n440_));
NAND3X1 NAND3X1_532 ( .A(csc_s_5_), .B(u1__abc_72801_new_n269_), .C(u1__abc_72801_new_n270_), .Y(u1__abc_72801_new_n271_));
NAND3X1 NAND3X1_533 ( .A(u1__abc_72801_new_n291_), .B(u1__abc_72801_new_n293_), .C(u1__abc_72801_new_n290_), .Y(u1__abc_72801_new_n294_));
NAND3X1 NAND3X1_534 ( .A(u1__abc_72801_new_n298_), .B(u1__abc_72801_new_n296_), .C(u1__abc_72801_new_n303_), .Y(u1__abc_72801_new_n304_));
NAND3X1 NAND3X1_535 ( .A(csc_s_5_), .B(\wb_addr_i[22] ), .C(u1__abc_72801_new_n269_), .Y(u1__abc_72801_new_n316_));
NAND3X1 NAND3X1_536 ( .A(u1__abc_72801_new_n315_), .B(u1__abc_72801_new_n314_), .C(u1__abc_72801_new_n318_), .Y(u1__abc_72801_new_n319_));
NAND3X1 NAND3X1_537 ( .A(u1__abc_72801_new_n336_), .B(u1__abc_72801_new_n282_), .C(u1__abc_72801_new_n337_), .Y(u1__abc_72801_new_n338_));
NAND3X1 NAND3X1_538 ( .A(\wb_addr_i[14] ), .B(u1__abc_72801_new_n273_), .C(u1__abc_72801_new_n268_), .Y(u1__abc_72801_new_n347_));
NAND3X1 NAND3X1_539 ( .A(u1_bas), .B(u1__abc_72801_new_n347_), .C(u1__abc_72801_new_n325_), .Y(u1__abc_72801_new_n348_));
NAND3X1 NAND3X1_54 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1422_), .C(u0__abc_74894_new_n1421_), .Y(u0__abc_74894_new_n1423_));
NAND3X1 NAND3X1_540 ( .A(\wb_addr_i[16] ), .B(u1__abc_72801_new_n349_), .C(u1__abc_72801_new_n351_), .Y(u1__abc_72801_new_n352_));
NAND3X1 NAND3X1_541 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n355_), .C(u1__abc_72801_new_n352_), .Y(u1__abc_72801_new_n356_));
NAND3X1 NAND3X1_542 ( .A(cs_le), .B(u1__abc_72801_new_n348_), .C(u1__abc_72801_new_n356_), .Y(u1__abc_72801_new_n357_));
NAND3X1 NAND3X1_543 ( .A(\wb_addr_i[15] ), .B(u1__abc_72801_new_n349_), .C(u1__abc_72801_new_n351_), .Y(u1__abc_72801_new_n360_));
NAND3X1 NAND3X1_544 ( .A(u1_bas), .B(u1__abc_72801_new_n362_), .C(u1__abc_72801_new_n360_), .Y(u1__abc_72801_new_n363_));
NAND3X1 NAND3X1_545 ( .A(\wb_addr_i[17] ), .B(u1__abc_72801_new_n349_), .C(u1__abc_72801_new_n351_), .Y(u1__abc_72801_new_n364_));
NAND3X1 NAND3X1_546 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n367_), .C(u1__abc_72801_new_n364_), .Y(u1__abc_72801_new_n368_));
NAND3X1 NAND3X1_547 ( .A(cs_le), .B(u1__abc_72801_new_n363_), .C(u1__abc_72801_new_n368_), .Y(u1__abc_72801_new_n369_));
NAND3X1 NAND3X1_548 ( .A(\wb_addr_i[18] ), .B(u1__abc_72801_new_n349_), .C(u1__abc_72801_new_n351_), .Y(u1__abc_72801_new_n372_));
NAND3X1 NAND3X1_549 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n375_), .C(u1__abc_72801_new_n372_), .Y(u1__abc_72801_new_n376_));
NAND3X1 NAND3X1_55 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1420_), .C(u0__abc_74894_new_n1423_), .Y(u0__abc_74894_new_n1424_));
NAND3X1 NAND3X1_550 ( .A(u1_bas), .B(u1__abc_72801_new_n355_), .C(u1__abc_72801_new_n352_), .Y(u1__abc_72801_new_n377_));
NAND3X1 NAND3X1_551 ( .A(cs_le), .B(u1__abc_72801_new_n376_), .C(u1__abc_72801_new_n377_), .Y(u1__abc_72801_new_n378_));
NAND3X1 NAND3X1_552 ( .A(u1_bas), .B(u1__abc_72801_new_n367_), .C(u1__abc_72801_new_n364_), .Y(u1__abc_72801_new_n381_));
NAND3X1 NAND3X1_553 ( .A(\wb_addr_i[19] ), .B(u1__abc_72801_new_n349_), .C(u1__abc_72801_new_n351_), .Y(u1__abc_72801_new_n382_));
NAND3X1 NAND3X1_554 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n385_), .C(u1__abc_72801_new_n382_), .Y(u1__abc_72801_new_n386_));
NAND3X1 NAND3X1_555 ( .A(cs_le), .B(u1__abc_72801_new_n381_), .C(u1__abc_72801_new_n386_), .Y(u1__abc_72801_new_n387_));
NAND3X1 NAND3X1_556 ( .A(u1_bas), .B(u1__abc_72801_new_n375_), .C(u1__abc_72801_new_n372_), .Y(u1__abc_72801_new_n390_));
NAND3X1 NAND3X1_557 ( .A(\wb_addr_i[20] ), .B(u1__abc_72801_new_n349_), .C(u1__abc_72801_new_n351_), .Y(u1__abc_72801_new_n391_));
NAND3X1 NAND3X1_558 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n394_), .C(u1__abc_72801_new_n391_), .Y(u1__abc_72801_new_n395_));
NAND3X1 NAND3X1_559 ( .A(cs_le), .B(u1__abc_72801_new_n390_), .C(u1__abc_72801_new_n395_), .Y(u1__abc_72801_new_n396_));
NAND3X1 NAND3X1_56 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1425_), .C(u0__abc_74894_new_n1424_), .Y(u0__abc_74894_new_n1426_));
NAND3X1 NAND3X1_560 ( .A(\wb_addr_i[22] ), .B(u1__abc_72801_new_n273_), .C(u1__abc_72801_new_n268_), .Y(u1__abc_72801_new_n412_));
NAND3X1 NAND3X1_561 ( .A(\wb_addr_i[21] ), .B(u1__abc_72801_new_n273_), .C(u1__abc_72801_new_n268_), .Y(u1__abc_72801_new_n418_));
NAND3X1 NAND3X1_562 ( .A(u1_bas), .B(u1__abc_72801_new_n418_), .C(u1__abc_72801_new_n403_), .Y(u1__abc_72801_new_n419_));
NAND3X1 NAND3X1_563 ( .A(\wb_addr_i[23] ), .B(u1__abc_72801_new_n349_), .C(u1__abc_72801_new_n351_), .Y(u1__abc_72801_new_n420_));
NAND3X1 NAND3X1_564 ( .A(u1__abc_72801_new_n421_), .B(u1__abc_72801_new_n426_), .C(u1__abc_72801_new_n420_), .Y(u1__abc_72801_new_n427_));
NAND3X1 NAND3X1_565 ( .A(cs_le), .B(u1__abc_72801_new_n419_), .C(u1__abc_72801_new_n427_), .Y(u1__abc_72801_new_n428_));
NAND3X1 NAND3X1_566 ( .A(u1__abc_72801_new_n435_), .B(u1__abc_72801_new_n436_), .C(u1__abc_72801_new_n437_), .Y(u1__abc_72801_new_n438_));
NAND3X1 NAND3X1_567 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n448_), .C(u1__abc_72801_new_n449_), .Y(u1__abc_72801_new_n450_));
NAND3X1 NAND3X1_568 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n453_), .C(u1__abc_72801_new_n454_), .Y(u1__abc_72801_new_n455_));
NAND3X1 NAND3X1_569 ( .A(u1_acs_addr_0_), .B(u1_acs_addr_1_), .C(u1_acs_addr_2_), .Y(u1_u0__abc_72719_new_n54_));
NAND3X1 NAND3X1_57 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1418_), .C(u0__abc_74894_new_n1426_), .Y(u0__abc_74894_new_n1427_));
NAND3X1 NAND3X1_570 ( .A(u1_acs_addr_4_), .B(u1_acs_addr_5_), .C(u1_u0__abc_72719_new_n58_), .Y(u1_u0__abc_72719_new_n61_));
NAND3X1 NAND3X1_571 ( .A(u1_u0__abc_72719_new_n77_), .B(u1_u0__abc_72719_new_n58_), .C(u1_u0__abc_72719_new_n70_), .Y(u1_u0__abc_72719_new_n78_));
NAND3X1 NAND3X1_572 ( .A(u1_acs_addr_13_), .B(u1_u0_inc_next), .C(u1_acs_addr_12_), .Y(u1_u0__abc_72719_new_n91_));
NAND3X1 NAND3X1_573 ( .A(u1_acs_addr_13_), .B(u1_u0__abc_72719_new_n89_), .C(u1_u0__abc_72719_new_n96_), .Y(u1_u0__abc_72719_new_n97_));
NAND3X1 NAND3X1_574 ( .A(u1_acs_addr_20_), .B(u1_u0__abc_72719_new_n109_), .C(u1_u0__abc_72719_new_n100_), .Y(u1_u0__abc_72719_new_n111_));
NAND3X1 NAND3X1_575 ( .A(u1_u0__abc_72719_new_n109_), .B(u1_u0__abc_72719_new_n120_), .C(u1_u0__abc_72719_new_n100_), .Y(u1_u0__abc_72719_new_n121_));
NAND3X1 NAND3X1_576 ( .A(u1_acs_addr_22_), .B(u1_u0__abc_72719_new_n125_), .C(u1_u0__abc_72719_new_n126_), .Y(u1_u0__abc_72719_new_n127_));
NAND3X1 NAND3X1_577 ( .A(u2_u0__abc_73914_new_n270_), .B(u2_u0__abc_73914_new_n272_), .C(u2_u0__abc_73914_new_n269_), .Y(u2_u0__abc_73914_new_n273_));
NAND3X1 NAND3X1_578 ( .A(u2_u0__abc_73914_new_n274_), .B(u2_u0__abc_73914_new_n276_), .C(u2_u0__abc_73914_new_n281_), .Y(u2_u0__abc_73914_new_n282_));
NAND3X1 NAND3X1_579 ( .A(u2_u0__abc_73914_new_n311_), .B(u2_u0__abc_73914_new_n312_), .C(u2_u0__abc_73914_new_n310_), .Y(u2_u0__abc_73914_new_n313_));
NAND3X1 NAND3X1_58 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1442_), .C(u0__abc_74894_new_n1441_), .Y(u0__abc_74894_new_n1443_));
NAND3X1 NAND3X1_580 ( .A(u2_u0__abc_73914_new_n315_), .B(u2_u0__abc_73914_new_n316_), .C(u2_u0__abc_73914_new_n317_), .Y(u2_u0__abc_73914_new_n318_));
NAND3X1 NAND3X1_581 ( .A(u2_u0__abc_73914_new_n319_), .B(u2_u0__abc_73914_new_n320_), .C(u2_u0__abc_73914_new_n321_), .Y(u2_u0__abc_73914_new_n322_));
NAND3X1 NAND3X1_582 ( .A(u2_u0__abc_73914_new_n326_), .B(u2_u0__abc_73914_new_n325_), .C(u2_u0__abc_73914_new_n323_), .Y(u2_u0__abc_73914_new_n327_));
NAND3X1 NAND3X1_583 ( .A(u2_u0__abc_73914_new_n330_), .B(u2_u0__abc_73914_new_n331_), .C(u2_u0__abc_73914_new_n332_), .Y(u2_u0__abc_73914_new_n333_));
NAND3X1 NAND3X1_584 ( .A(u2_u0__abc_73914_new_n336_), .B(u2_u0__abc_73914_new_n335_), .C(u2_u0__abc_73914_new_n337_), .Y(u2_u0__abc_73914_new_n338_));
NAND3X1 NAND3X1_585 ( .A(u2_u0__abc_73914_new_n339_), .B(u2_u0__abc_73914_new_n340_), .C(u2_u0__abc_73914_new_n343_), .Y(u2_u0__abc_73914_new_n344_));
NAND3X1 NAND3X1_586 ( .A(u2_u0__abc_73914_new_n351_), .B(u2_u0__abc_73914_new_n352_), .C(u2_u0__abc_73914_new_n350_), .Y(u2_u0__abc_73914_new_n353_));
NAND3X1 NAND3X1_587 ( .A(u2_u0__abc_73914_new_n354_), .B(u2_u0__abc_73914_new_n357_), .C(u2_u0__abc_73914_new_n362_), .Y(u2_u0__abc_73914_new_n363_));
NAND3X1 NAND3X1_588 ( .A(u2_u0__abc_73914_new_n368_), .B(u2_u0__abc_73914_new_n370_), .C(u2_u0__abc_73914_new_n366_), .Y(u2_u0__abc_73914_new_n371_));
NAND3X1 NAND3X1_589 ( .A(u2_u0__abc_73914_new_n237_), .B(u2_u0__abc_73914_new_n392_), .C(u2_u0__abc_73914_new_n393_), .Y(u2_u0__abc_73914_new_n394_));
NAND3X1 NAND3X1_59 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1440_), .C(u0__abc_74894_new_n1443_), .Y(u0__abc_74894_new_n1444_));
NAND3X1 NAND3X1_590 ( .A(u2_u1__abc_73914_new_n270_), .B(u2_u1__abc_73914_new_n272_), .C(u2_u1__abc_73914_new_n269_), .Y(u2_u1__abc_73914_new_n273_));
NAND3X1 NAND3X1_591 ( .A(u2_u1__abc_73914_new_n274_), .B(u2_u1__abc_73914_new_n276_), .C(u2_u1__abc_73914_new_n281_), .Y(u2_u1__abc_73914_new_n282_));
NAND3X1 NAND3X1_592 ( .A(u2_u1__abc_73914_new_n311_), .B(u2_u1__abc_73914_new_n312_), .C(u2_u1__abc_73914_new_n310_), .Y(u2_u1__abc_73914_new_n313_));
NAND3X1 NAND3X1_593 ( .A(u2_u1__abc_73914_new_n315_), .B(u2_u1__abc_73914_new_n316_), .C(u2_u1__abc_73914_new_n317_), .Y(u2_u1__abc_73914_new_n318_));
NAND3X1 NAND3X1_594 ( .A(u2_u1__abc_73914_new_n319_), .B(u2_u1__abc_73914_new_n320_), .C(u2_u1__abc_73914_new_n321_), .Y(u2_u1__abc_73914_new_n322_));
NAND3X1 NAND3X1_595 ( .A(u2_u1__abc_73914_new_n326_), .B(u2_u1__abc_73914_new_n325_), .C(u2_u1__abc_73914_new_n323_), .Y(u2_u1__abc_73914_new_n327_));
NAND3X1 NAND3X1_596 ( .A(u2_u1__abc_73914_new_n330_), .B(u2_u1__abc_73914_new_n331_), .C(u2_u1__abc_73914_new_n332_), .Y(u2_u1__abc_73914_new_n333_));
NAND3X1 NAND3X1_597 ( .A(u2_u1__abc_73914_new_n336_), .B(u2_u1__abc_73914_new_n335_), .C(u2_u1__abc_73914_new_n337_), .Y(u2_u1__abc_73914_new_n338_));
NAND3X1 NAND3X1_598 ( .A(u2_u1__abc_73914_new_n339_), .B(u2_u1__abc_73914_new_n340_), .C(u2_u1__abc_73914_new_n343_), .Y(u2_u1__abc_73914_new_n344_));
NAND3X1 NAND3X1_599 ( .A(u2_u1__abc_73914_new_n351_), .B(u2_u1__abc_73914_new_n352_), .C(u2_u1__abc_73914_new_n350_), .Y(u2_u1__abc_73914_new_n353_));
NAND3X1 NAND3X1_6 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1182_), .C(u0__abc_74894_new_n1181_), .Y(u0__abc_74894_new_n1183_));
NAND3X1 NAND3X1_60 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1445_), .C(u0__abc_74894_new_n1444_), .Y(u0__abc_74894_new_n1446_));
NAND3X1 NAND3X1_600 ( .A(u2_u1__abc_73914_new_n354_), .B(u2_u1__abc_73914_new_n357_), .C(u2_u1__abc_73914_new_n362_), .Y(u2_u1__abc_73914_new_n363_));
NAND3X1 NAND3X1_601 ( .A(u2_u1__abc_73914_new_n368_), .B(u2_u1__abc_73914_new_n370_), .C(u2_u1__abc_73914_new_n366_), .Y(u2_u1__abc_73914_new_n371_));
NAND3X1 NAND3X1_602 ( .A(u2_u1__abc_73914_new_n237_), .B(u2_u1__abc_73914_new_n392_), .C(u2_u1__abc_73914_new_n393_), .Y(u2_u1__abc_73914_new_n394_));
NAND3X1 NAND3X1_603 ( .A(u3_rd_fifo_out_33_), .B(u3__abc_73372_new_n632_), .C(u3__abc_73372_new_n631_), .Y(u3__abc_73372_new_n633_));
NAND3X1 NAND3X1_604 ( .A(u3__abc_73372_new_n630_), .B(u3__abc_73372_new_n637_), .C(u3__abc_73372_new_n633_), .Y(u3__abc_73372_new_n638_));
NAND3X1 NAND3X1_605 ( .A(u3__abc_73372_new_n634_), .B(u3__abc_73372_new_n632_), .C(u3__abc_73372_new_n631_), .Y(u3__abc_73372_new_n641_));
NAND3X1 NAND3X1_606 ( .A(u3__abc_73372_new_n639_), .B(u3__abc_73372_new_n640_), .C(u3__abc_73372_new_n641_), .Y(u3__abc_73372_new_n642_));
NAND3X1 NAND3X1_607 ( .A(u3_rd_fifo_out_34_), .B(u3__abc_73372_new_n656_), .C(u3__abc_73372_new_n657_), .Y(u3__abc_73372_new_n660_));
NAND3X1 NAND3X1_608 ( .A(u3__abc_73372_new_n652_), .B(u3__abc_73372_new_n654_), .C(u3__abc_73372_new_n653_), .Y(u3__abc_73372_new_n661_));
NAND3X1 NAND3X1_609 ( .A(u3__abc_73372_new_n650_), .B(u3__abc_73372_new_n661_), .C(u3__abc_73372_new_n660_), .Y(u3__abc_73372_new_n662_));
NAND3X1 NAND3X1_61 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1438_), .C(u0__abc_74894_new_n1446_), .Y(u0__abc_74894_new_n1447_));
NAND3X1 NAND3X1_610 ( .A(u3__abc_73372_new_n668_), .B(u3__abc_73372_new_n673_), .C(u3__abc_73372_new_n663_), .Y(u3__abc_73372_new_n674_));
NAND3X1 NAND3X1_611 ( .A(u3__abc_73372_new_n662_), .B(u3__abc_73372_new_n675_), .C(u3__abc_73372_new_n659_), .Y(u3__abc_73372_new_n676_));
NAND3X1 NAND3X1_612 ( .A(u3_rd_fifo_out_32_), .B(u3__abc_73372_new_n682_), .C(u3__abc_73372_new_n681_), .Y(u3__abc_73372_new_n683_));
NAND3X1 NAND3X1_613 ( .A(u3__abc_73372_new_n679_), .B(u3__abc_73372_new_n686_), .C(u3__abc_73372_new_n683_), .Y(u3__abc_73372_new_n687_));
NAND3X1 NAND3X1_614 ( .A(u3__abc_73372_new_n684_), .B(u3__abc_73372_new_n682_), .C(u3__abc_73372_new_n681_), .Y(u3__abc_73372_new_n690_));
NAND3X1 NAND3X1_615 ( .A(u3__abc_73372_new_n688_), .B(u3__abc_73372_new_n689_), .C(u3__abc_73372_new_n690_), .Y(u3__abc_73372_new_n691_));
NAND3X1 NAND3X1_616 ( .A(u3__abc_73372_new_n687_), .B(u3__abc_73372_new_n691_), .C(u3__abc_73372_new_n694_), .Y(u3__abc_73372_new_n695_));
NAND3X1 NAND3X1_617 ( .A(u3_rd_fifo_out_35_), .B(u3__abc_73372_new_n706_), .C(u3__abc_73372_new_n707_), .Y(u3__abc_73372_new_n710_));
NAND3X1 NAND3X1_618 ( .A(u3__abc_73372_new_n702_), .B(u3__abc_73372_new_n704_), .C(u3__abc_73372_new_n703_), .Y(u3__abc_73372_new_n711_));
NAND3X1 NAND3X1_619 ( .A(u3__abc_73372_new_n700_), .B(u3__abc_73372_new_n711_), .C(u3__abc_73372_new_n710_), .Y(u3__abc_73372_new_n712_));
NAND3X1 NAND3X1_62 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1462_), .C(u0__abc_74894_new_n1461_), .Y(u0__abc_74894_new_n1463_));
NAND3X1 NAND3X1_620 ( .A(u3__abc_73372_new_n718_), .B(u3__abc_73372_new_n723_), .C(u3__abc_73372_new_n713_), .Y(u3__abc_73372_new_n724_));
NAND3X1 NAND3X1_621 ( .A(u3__abc_73372_new_n712_), .B(u3__abc_73372_new_n725_), .C(u3__abc_73372_new_n709_), .Y(u3__abc_73372_new_n726_));
NAND3X1 NAND3X1_622 ( .A(mem_ack), .B(u3_pen), .C(u3__abc_73372_new_n627_), .Y(u3__abc_73372_new_n729_));
NAND3X1 NAND3X1_623 ( .A(u3_u0_r0_0_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n741_));
NAND3X1 NAND3X1_624 ( .A(u3_u0__abc_74260_new_n743_), .B(u3_u0__abc_74260_new_n748_), .C(u3_u0__abc_74260_new_n741_), .Y(u3_rd_fifo_out_0_));
NAND3X1 NAND3X1_625 ( .A(u3_u0_r0_1_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n750_));
NAND3X1 NAND3X1_626 ( .A(u3_u0__abc_74260_new_n751_), .B(u3_u0__abc_74260_new_n752_), .C(u3_u0__abc_74260_new_n750_), .Y(u3_rd_fifo_out_1_));
NAND3X1 NAND3X1_627 ( .A(u3_u0_r0_2_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n754_));
NAND3X1 NAND3X1_628 ( .A(u3_u0__abc_74260_new_n755_), .B(u3_u0__abc_74260_new_n756_), .C(u3_u0__abc_74260_new_n754_), .Y(u3_rd_fifo_out_2_));
NAND3X1 NAND3X1_629 ( .A(u3_u0_r0_3_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n758_));
NAND3X1 NAND3X1_63 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1460_), .C(u0__abc_74894_new_n1463_), .Y(u0__abc_74894_new_n1464_));
NAND3X1 NAND3X1_630 ( .A(u3_u0__abc_74260_new_n759_), .B(u3_u0__abc_74260_new_n760_), .C(u3_u0__abc_74260_new_n758_), .Y(u3_rd_fifo_out_3_));
NAND3X1 NAND3X1_631 ( .A(u3_u0_r0_4_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n762_));
NAND3X1 NAND3X1_632 ( .A(u3_u0__abc_74260_new_n763_), .B(u3_u0__abc_74260_new_n764_), .C(u3_u0__abc_74260_new_n762_), .Y(u3_rd_fifo_out_4_));
NAND3X1 NAND3X1_633 ( .A(u3_u0_r0_5_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n766_));
NAND3X1 NAND3X1_634 ( .A(u3_u0__abc_74260_new_n767_), .B(u3_u0__abc_74260_new_n768_), .C(u3_u0__abc_74260_new_n766_), .Y(u3_rd_fifo_out_5_));
NAND3X1 NAND3X1_635 ( .A(u3_u0_r0_6_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n770_));
NAND3X1 NAND3X1_636 ( .A(u3_u0__abc_74260_new_n771_), .B(u3_u0__abc_74260_new_n772_), .C(u3_u0__abc_74260_new_n770_), .Y(u3_rd_fifo_out_6_));
NAND3X1 NAND3X1_637 ( .A(u3_u0_r0_7_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n774_));
NAND3X1 NAND3X1_638 ( .A(u3_u0__abc_74260_new_n775_), .B(u3_u0__abc_74260_new_n776_), .C(u3_u0__abc_74260_new_n774_), .Y(u3_rd_fifo_out_7_));
NAND3X1 NAND3X1_639 ( .A(u3_u0_r0_8_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n778_));
NAND3X1 NAND3X1_64 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1465_), .C(u0__abc_74894_new_n1464_), .Y(u0__abc_74894_new_n1466_));
NAND3X1 NAND3X1_640 ( .A(u3_u0__abc_74260_new_n779_), .B(u3_u0__abc_74260_new_n780_), .C(u3_u0__abc_74260_new_n778_), .Y(u3_rd_fifo_out_8_));
NAND3X1 NAND3X1_641 ( .A(u3_u0_r0_9_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n782_));
NAND3X1 NAND3X1_642 ( .A(u3_u0__abc_74260_new_n783_), .B(u3_u0__abc_74260_new_n784_), .C(u3_u0__abc_74260_new_n782_), .Y(u3_rd_fifo_out_9_));
NAND3X1 NAND3X1_643 ( .A(u3_u0_r0_10_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n786_));
NAND3X1 NAND3X1_644 ( .A(u3_u0__abc_74260_new_n787_), .B(u3_u0__abc_74260_new_n788_), .C(u3_u0__abc_74260_new_n786_), .Y(u3_rd_fifo_out_10_));
NAND3X1 NAND3X1_645 ( .A(u3_u0_r0_11_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n790_));
NAND3X1 NAND3X1_646 ( .A(u3_u0__abc_74260_new_n791_), .B(u3_u0__abc_74260_new_n792_), .C(u3_u0__abc_74260_new_n790_), .Y(u3_rd_fifo_out_11_));
NAND3X1 NAND3X1_647 ( .A(u3_u0_r0_12_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n794_));
NAND3X1 NAND3X1_648 ( .A(u3_u0__abc_74260_new_n795_), .B(u3_u0__abc_74260_new_n796_), .C(u3_u0__abc_74260_new_n794_), .Y(u3_rd_fifo_out_12_));
NAND3X1 NAND3X1_649 ( .A(u3_u0_r0_13_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n798_));
NAND3X1 NAND3X1_65 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1458_), .C(u0__abc_74894_new_n1466_), .Y(u0__abc_74894_new_n1467_));
NAND3X1 NAND3X1_650 ( .A(u3_u0__abc_74260_new_n799_), .B(u3_u0__abc_74260_new_n800_), .C(u3_u0__abc_74260_new_n798_), .Y(u3_rd_fifo_out_13_));
NAND3X1 NAND3X1_651 ( .A(u3_u0_r0_14_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n802_));
NAND3X1 NAND3X1_652 ( .A(u3_u0__abc_74260_new_n803_), .B(u3_u0__abc_74260_new_n804_), .C(u3_u0__abc_74260_new_n802_), .Y(u3_rd_fifo_out_14_));
NAND3X1 NAND3X1_653 ( .A(u3_u0_r0_15_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n806_));
NAND3X1 NAND3X1_654 ( .A(u3_u0__abc_74260_new_n807_), .B(u3_u0__abc_74260_new_n808_), .C(u3_u0__abc_74260_new_n806_), .Y(u3_rd_fifo_out_15_));
NAND3X1 NAND3X1_655 ( .A(u3_u0_r0_16_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n810_));
NAND3X1 NAND3X1_656 ( .A(u3_u0__abc_74260_new_n811_), .B(u3_u0__abc_74260_new_n812_), .C(u3_u0__abc_74260_new_n810_), .Y(u3_rd_fifo_out_16_));
NAND3X1 NAND3X1_657 ( .A(u3_u0_r0_17_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n814_));
NAND3X1 NAND3X1_658 ( .A(u3_u0__abc_74260_new_n815_), .B(u3_u0__abc_74260_new_n816_), .C(u3_u0__abc_74260_new_n814_), .Y(u3_rd_fifo_out_17_));
NAND3X1 NAND3X1_659 ( .A(u3_u0_r0_18_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n818_));
NAND3X1 NAND3X1_66 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1482_), .C(u0__abc_74894_new_n1481_), .Y(u0__abc_74894_new_n1483_));
NAND3X1 NAND3X1_660 ( .A(u3_u0__abc_74260_new_n819_), .B(u3_u0__abc_74260_new_n820_), .C(u3_u0__abc_74260_new_n818_), .Y(u3_rd_fifo_out_18_));
NAND3X1 NAND3X1_661 ( .A(u3_u0_r0_19_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n822_));
NAND3X1 NAND3X1_662 ( .A(u3_u0__abc_74260_new_n823_), .B(u3_u0__abc_74260_new_n824_), .C(u3_u0__abc_74260_new_n822_), .Y(u3_rd_fifo_out_19_));
NAND3X1 NAND3X1_663 ( .A(u3_u0_r0_20_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n826_));
NAND3X1 NAND3X1_664 ( .A(u3_u0__abc_74260_new_n827_), .B(u3_u0__abc_74260_new_n828_), .C(u3_u0__abc_74260_new_n826_), .Y(u3_rd_fifo_out_20_));
NAND3X1 NAND3X1_665 ( .A(u3_u0_r0_21_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n830_));
NAND3X1 NAND3X1_666 ( .A(u3_u0__abc_74260_new_n831_), .B(u3_u0__abc_74260_new_n832_), .C(u3_u0__abc_74260_new_n830_), .Y(u3_rd_fifo_out_21_));
NAND3X1 NAND3X1_667 ( .A(u3_u0_r0_22_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n834_));
NAND3X1 NAND3X1_668 ( .A(u3_u0__abc_74260_new_n835_), .B(u3_u0__abc_74260_new_n836_), .C(u3_u0__abc_74260_new_n834_), .Y(u3_rd_fifo_out_22_));
NAND3X1 NAND3X1_669 ( .A(u3_u0_r0_23_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n838_));
NAND3X1 NAND3X1_67 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1480_), .C(u0__abc_74894_new_n1483_), .Y(u0__abc_74894_new_n1484_));
NAND3X1 NAND3X1_670 ( .A(u3_u0__abc_74260_new_n839_), .B(u3_u0__abc_74260_new_n840_), .C(u3_u0__abc_74260_new_n838_), .Y(u3_rd_fifo_out_23_));
NAND3X1 NAND3X1_671 ( .A(u3_u0_r0_24_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n842_));
NAND3X1 NAND3X1_672 ( .A(u3_u0__abc_74260_new_n843_), .B(u3_u0__abc_74260_new_n844_), .C(u3_u0__abc_74260_new_n842_), .Y(u3_rd_fifo_out_24_));
NAND3X1 NAND3X1_673 ( .A(u3_u0_r0_25_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n846_));
NAND3X1 NAND3X1_674 ( .A(u3_u0__abc_74260_new_n847_), .B(u3_u0__abc_74260_new_n848_), .C(u3_u0__abc_74260_new_n846_), .Y(u3_rd_fifo_out_25_));
NAND3X1 NAND3X1_675 ( .A(u3_u0_r0_26_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n850_));
NAND3X1 NAND3X1_676 ( .A(u3_u0__abc_74260_new_n851_), .B(u3_u0__abc_74260_new_n852_), .C(u3_u0__abc_74260_new_n850_), .Y(u3_rd_fifo_out_26_));
NAND3X1 NAND3X1_677 ( .A(u3_u0_r0_27_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n854_));
NAND3X1 NAND3X1_678 ( .A(u3_u0__abc_74260_new_n855_), .B(u3_u0__abc_74260_new_n856_), .C(u3_u0__abc_74260_new_n854_), .Y(u3_rd_fifo_out_27_));
NAND3X1 NAND3X1_679 ( .A(u3_u0_r0_28_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n858_));
NAND3X1 NAND3X1_68 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1485_), .C(u0__abc_74894_new_n1484_), .Y(u0__abc_74894_new_n1486_));
NAND3X1 NAND3X1_680 ( .A(u3_u0__abc_74260_new_n859_), .B(u3_u0__abc_74260_new_n860_), .C(u3_u0__abc_74260_new_n858_), .Y(u3_rd_fifo_out_28_));
NAND3X1 NAND3X1_681 ( .A(u3_u0_r0_29_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n862_));
NAND3X1 NAND3X1_682 ( .A(u3_u0__abc_74260_new_n863_), .B(u3_u0__abc_74260_new_n864_), .C(u3_u0__abc_74260_new_n862_), .Y(u3_rd_fifo_out_29_));
NAND3X1 NAND3X1_683 ( .A(u3_u0_r0_30_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n866_));
NAND3X1 NAND3X1_684 ( .A(u3_u0__abc_74260_new_n867_), .B(u3_u0__abc_74260_new_n868_), .C(u3_u0__abc_74260_new_n866_), .Y(u3_rd_fifo_out_30_));
NAND3X1 NAND3X1_685 ( .A(u3_u0_r0_31_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n870_));
NAND3X1 NAND3X1_686 ( .A(u3_u0__abc_74260_new_n871_), .B(u3_u0__abc_74260_new_n872_), .C(u3_u0__abc_74260_new_n870_), .Y(u3_rd_fifo_out_31_));
NAND3X1 NAND3X1_687 ( .A(u3_u0_r0_32_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n874_));
NAND3X1 NAND3X1_688 ( .A(u3_u0__abc_74260_new_n875_), .B(u3_u0__abc_74260_new_n876_), .C(u3_u0__abc_74260_new_n874_), .Y(u3_rd_fifo_out_32_));
NAND3X1 NAND3X1_689 ( .A(u3_u0_r0_33_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n878_));
NAND3X1 NAND3X1_69 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1478_), .C(u0__abc_74894_new_n1486_), .Y(u0__abc_74894_new_n1487_));
NAND3X1 NAND3X1_690 ( .A(u3_u0__abc_74260_new_n879_), .B(u3_u0__abc_74260_new_n880_), .C(u3_u0__abc_74260_new_n878_), .Y(u3_rd_fifo_out_33_));
NAND3X1 NAND3X1_691 ( .A(u3_u0_r0_34_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n882_));
NAND3X1 NAND3X1_692 ( .A(u3_u0__abc_74260_new_n883_), .B(u3_u0__abc_74260_new_n884_), .C(u3_u0__abc_74260_new_n882_), .Y(u3_rd_fifo_out_34_));
NAND3X1 NAND3X1_693 ( .A(u3_u0_r0_35_), .B(u3_u0__abc_74260_new_n736_), .C(u3_u0__abc_74260_new_n740_), .Y(u3_u0__abc_74260_new_n886_));
NAND3X1 NAND3X1_694 ( .A(u3_u0__abc_74260_new_n887_), .B(u3_u0__abc_74260_new_n888_), .C(u3_u0__abc_74260_new_n886_), .Y(u3_rd_fifo_out_35_));
NAND3X1 NAND3X1_695 ( .A(u4__abc_74770_new_n68_), .B(u4__abc_74770_new_n69_), .C(u4__abc_74770_new_n67_), .Y(u4__0rfr_en_0_0_));
NAND3X1 NAND3X1_696 ( .A(u4__abc_74770_new_n82_), .B(u4__abc_74770_new_n83_), .C(u4__abc_74770_new_n88_), .Y(u4__abc_74770_new_n89_));
NAND3X1 NAND3X1_697 ( .A(u4_rfr_cnt_0_), .B(u4_rfr_cnt_1_), .C(u4_rfr_cnt_2_), .Y(u4__abc_74770_new_n102_));
NAND3X1 NAND3X1_698 ( .A(u4__abc_74770_new_n122_), .B(u4__abc_74770_new_n124_), .C(u4__abc_74770_new_n112_), .Y(u4__abc_74770_new_n125_));
NAND3X1 NAND3X1_699 ( .A(u4__abc_74770_new_n130_), .B(u4__abc_74770_new_n131_), .C(u4__abc_74770_new_n129_), .Y(u4__abc_74770_new_n132_));
NAND3X1 NAND3X1_7 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1180_), .C(u0__abc_74894_new_n1183_), .Y(u0__abc_74894_new_n1184_));
NAND3X1 NAND3X1_70 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1502_), .C(u0__abc_74894_new_n1501_), .Y(u0__abc_74894_new_n1503_));
NAND3X1 NAND3X1_700 ( .A(u4_ps_cnt_0_), .B(u4_ps_cnt_1_), .C(u4_rfr_en), .Y(u4__abc_74770_new_n139_));
NAND3X1 NAND3X1_701 ( .A(u4_ps_cnt_3_), .B(u4_ps_cnt_4_), .C(u4_ps_cnt_5_), .Y(u4__abc_74770_new_n154_));
NAND3X1 NAND3X1_702 ( .A(u4_ps_cnt_3_), .B(u4_ps_cnt_4_), .C(u4__abc_74770_new_n148_), .Y(u4__abc_74770_new_n158_));
NAND3X1 NAND3X1_703 ( .A(u4_ps_cnt_6_), .B(u4_ps_cnt_7_), .C(u4__abc_74770_new_n165_), .Y(u4__abc_74770_new_n166_));
NAND3X1 NAND3X1_704 ( .A(u4_ps_cnt_6_), .B(u4__abc_74770_new_n155_), .C(u4__abc_74770_new_n148_), .Y(u4__abc_74770_new_n168_));
NAND3X1 NAND3X1_705 ( .A(ref_int_2_), .B(u4__abc_74770_new_n181_), .C(u4__abc_74770_new_n184_), .Y(u4__abc_74770_new_n185_));
NAND3X1 NAND3X1_706 ( .A(u5__abc_78290_new_n427_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n429_), .Y(u5__abc_78290_new_n430_));
NAND3X1 NAND3X1_707 ( .A(u5_state_30_), .B(u5__abc_78290_new_n437_), .C(u5__abc_78290_new_n438_), .Y(u5__abc_78290_new_n439_));
NAND3X1 NAND3X1_708 ( .A(u5_state_32_), .B(u5__abc_78290_new_n467_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n468_));
NAND3X1 NAND3X1_709 ( .A(u5__abc_78290_new_n402_), .B(u5__abc_78290_new_n465_), .C(u5__abc_78290_new_n469_), .Y(u5__abc_78290_new_n470_));
NAND3X1 NAND3X1_71 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1500_), .C(u0__abc_74894_new_n1503_), .Y(u0__abc_74894_new_n1504_));
NAND3X1 NAND3X1_710 ( .A(u5__abc_78290_new_n481_), .B(u5_state_31_), .C(u5__abc_78290_new_n438_), .Y(u5__abc_78290_new_n482_));
NAND3X1 NAND3X1_711 ( .A(u5__abc_78290_new_n473_), .B(u5__abc_78290_new_n483_), .C(u5__abc_78290_new_n480_), .Y(u5__abc_78290_new_n484_));
NAND3X1 NAND3X1_712 ( .A(u5__abc_78290_new_n472_), .B(u5__abc_78290_new_n441_), .C(u5__abc_78290_new_n484_), .Y(u5_suspended_d));
NAND3X1 NAND3X1_713 ( .A(u5_burst_act_rd), .B(u5_cke_o_del), .C(u5__abc_78290_new_n487_), .Y(u5__abc_78290_new_n488_));
NAND3X1 NAND3X1_714 ( .A(u5__abc_78290_new_n411_), .B(u5__abc_78290_new_n494_), .C(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n495_));
NAND3X1 NAND3X1_715 ( .A(u5__abc_78290_new_n434_), .B(u5__abc_78290_new_n502_), .C(u5__abc_78290_new_n450_), .Y(u5__abc_78290_new_n503_));
NAND3X1 NAND3X1_716 ( .A(u5__abc_78290_new_n499_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n504_), .Y(u5__abc_78290_new_n505_));
NAND3X1 NAND3X1_717 ( .A(u5__abc_78290_new_n435_), .B(u5__abc_78290_new_n508_), .C(u5__abc_78290_new_n450_), .Y(u5__abc_78290_new_n509_));
NAND3X1 NAND3X1_718 ( .A(u5__abc_78290_new_n499_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n510_), .Y(u5__abc_78290_new_n511_));
NAND3X1 NAND3X1_719 ( .A(u5__abc_78290_new_n465_), .B(u5__abc_78290_new_n518_), .C(u5__abc_78290_new_n392_), .Y(u5__abc_78290_new_n519_));
NAND3X1 NAND3X1_72 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1505_), .C(u0__abc_74894_new_n1504_), .Y(u0__abc_74894_new_n1506_));
NAND3X1 NAND3X1_720 ( .A(u5__abc_78290_new_n473_), .B(u5__abc_78290_new_n525_), .C(u5__abc_78290_new_n526_), .Y(u5__abc_78290_new_n527_));
NAND3X1 NAND3X1_721 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n528_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n529_));
NAND3X1 NAND3X1_722 ( .A(u5__abc_78290_new_n531_), .B(u5__abc_78290_new_n533_), .C(u5__abc_78290_new_n465_), .Y(u5__abc_78290_new_n534_));
NAND3X1 NAND3X1_723 ( .A(u5_state_28_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n540_), .Y(u5__abc_78290_new_n541_));
NAND3X1 NAND3X1_724 ( .A(u5__abc_78290_new_n536_), .B(u5__abc_78290_new_n529_), .C(u5__abc_78290_new_n541_), .Y(u5__abc_78290_new_n542_));
NAND3X1 NAND3X1_725 ( .A(u5_state_29_), .B(u5__abc_78290_new_n523_), .C(u5__abc_78290_new_n451_), .Y(u5__abc_78290_new_n544_));
NAND3X1 NAND3X1_726 ( .A(u5__abc_78290_new_n423_), .B(u5__abc_78290_new_n546_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n547_));
NAND3X1 NAND3X1_727 ( .A(u5__abc_78290_new_n550_), .B(u5__abc_78290_new_n431_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n551_));
NAND3X1 NAND3X1_728 ( .A(u5_state_27_), .B(u5__abc_78290_new_n392_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n552_));
NAND3X1 NAND3X1_729 ( .A(u5__abc_78290_new_n521_), .B(u5__abc_78290_new_n543_), .C(u5__abc_78290_new_n554_), .Y(u5__abc_78290_new_n555_));
NAND3X1 NAND3X1_73 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1498_), .C(u0__abc_74894_new_n1506_), .Y(u0__abc_74894_new_n1507_));
NAND3X1 NAND3X1_730 ( .A(u5_state_19_), .B(u5__abc_78290_new_n558_), .C(u5__abc_78290_new_n425_), .Y(u5__abc_78290_new_n559_));
NAND3X1 NAND3X1_731 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n562_), .C(u5__abc_78290_new_n566_), .Y(u5__abc_78290_new_n567_));
NAND3X1 NAND3X1_732 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n568_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n569_));
NAND3X1 NAND3X1_733 ( .A(u5__abc_78290_new_n571_), .B(u5_state_16_), .C(u5__abc_78290_new_n424_), .Y(u5__abc_78290_new_n572_));
NAND3X1 NAND3X1_734 ( .A(u5__abc_78290_new_n582_), .B(u5_state_24_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n583_));
NAND3X1 NAND3X1_735 ( .A(u5__abc_78290_new_n499_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n586_), .Y(u5__abc_78290_new_n587_));
NAND3X1 NAND3X1_736 ( .A(u5__abc_78290_new_n591_), .B(u5__abc_78290_new_n588_), .C(u5__abc_78290_new_n589_), .Y(u5__abc_78290_new_n592_));
NAND3X1 NAND3X1_737 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n593_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n594_));
NAND3X1 NAND3X1_738 ( .A(u5__abc_78290_new_n597_), .B(u5__abc_78290_new_n588_), .C(u5__abc_78290_new_n589_), .Y(u5__abc_78290_new_n598_));
NAND3X1 NAND3X1_739 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n599_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n600_));
NAND3X1 NAND3X1_74 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1522_), .C(u0__abc_74894_new_n1521_), .Y(u0__abc_74894_new_n1523_));
NAND3X1 NAND3X1_740 ( .A(u5__abc_78290_new_n604_), .B(u5__abc_78290_new_n588_), .C(u5__abc_78290_new_n602_), .Y(u5__abc_78290_new_n605_));
NAND3X1 NAND3X1_741 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n606_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n607_));
NAND3X1 NAND3X1_742 ( .A(u5__abc_78290_new_n561_), .B(u5__abc_78290_new_n569_), .C(u5__abc_78290_new_n610_), .Y(u5__abc_78290_new_n611_));
NAND3X1 NAND3X1_743 ( .A(u5__abc_78290_new_n387_), .B(u5__abc_78290_new_n616_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n617_));
NAND3X1 NAND3X1_744 ( .A(u5__abc_78290_new_n387_), .B(u5__abc_78290_new_n389_), .C(u5__abc_78290_new_n621_), .Y(u5__abc_78290_new_n622_));
NAND3X1 NAND3X1_745 ( .A(u5__abc_78290_new_n628_), .B(u5__abc_78290_new_n421_), .C(u5__abc_78290_new_n626_), .Y(u5__abc_78290_new_n629_));
NAND3X1 NAND3X1_746 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n630_), .Y(u5__abc_78290_new_n631_));
NAND3X1 NAND3X1_747 ( .A(u5__abc_78290_new_n633_), .B(u5__abc_78290_new_n636_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n637_));
NAND3X1 NAND3X1_748 ( .A(u5__abc_78290_new_n643_), .B(u5__abc_78290_new_n396_), .C(u5__abc_78290_new_n645_), .Y(u5__abc_78290_new_n646_));
NAND3X1 NAND3X1_749 ( .A(u5__abc_78290_new_n647_), .B(u5__abc_78290_new_n642_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n648_));
NAND3X1 NAND3X1_75 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1520_), .C(u0__abc_74894_new_n1523_), .Y(u0__abc_74894_new_n1524_));
NAND3X1 NAND3X1_750 ( .A(u5__abc_78290_new_n649_), .B(u5__abc_78290_new_n651_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n652_));
NAND3X1 NAND3X1_751 ( .A(u5_state_47_), .B(u5__abc_78290_new_n394_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n657_));
NAND3X1 NAND3X1_752 ( .A(u5__abc_78290_new_n658_), .B(u5__abc_78290_new_n642_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n659_));
NAND3X1 NAND3X1_753 ( .A(u5_state_39_), .B(u5__abc_78290_new_n401_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n664_));
NAND3X1 NAND3X1_754 ( .A(u5__abc_78290_new_n665_), .B(u5__abc_78290_new_n661_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n666_));
NAND3X1 NAND3X1_755 ( .A(u5__abc_78290_new_n648_), .B(u5__abc_78290_new_n668_), .C(u5__abc_78290_new_n641_), .Y(u5__abc_78290_new_n669_));
NAND3X1 NAND3X1_756 ( .A(u5_state_42_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n673_), .Y(u5__abc_78290_new_n674_));
NAND3X1 NAND3X1_757 ( .A(u5_state_37_), .B(u5__abc_78290_new_n400_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n679_));
NAND3X1 NAND3X1_758 ( .A(u5_state_46_), .B(u5__abc_78290_new_n394_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n689_));
NAND3X1 NAND3X1_759 ( .A(u5__abc_78290_new_n688_), .B(u5__abc_78290_new_n690_), .C(u5__abc_78290_new_n392_), .Y(u5__abc_78290_new_n691_));
NAND3X1 NAND3X1_76 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1525_), .C(u0__abc_74894_new_n1524_), .Y(u0__abc_74894_new_n1526_));
NAND3X1 NAND3X1_760 ( .A(u5_state_45_), .B(u5__abc_78290_new_n393_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n694_));
NAND3X1 NAND3X1_761 ( .A(u5_state_38_), .B(u5__abc_78290_new_n401_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n700_));
NAND3X1 NAND3X1_762 ( .A(u5__abc_78290_new_n701_), .B(u5__abc_78290_new_n661_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n702_));
NAND3X1 NAND3X1_763 ( .A(u5_state_44_), .B(u5__abc_78290_new_n393_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n705_));
NAND3X1 NAND3X1_764 ( .A(u5__abc_78290_new_n711_), .B(u5__abc_78290_new_n397_), .C(u5__abc_78290_new_n395_), .Y(u5__abc_78290_new_n712_));
NAND3X1 NAND3X1_765 ( .A(u5__abc_78290_new_n644_), .B(u5__abc_78290_new_n396_), .C(u5__abc_78290_new_n395_), .Y(u5__abc_78290_new_n717_));
NAND3X1 NAND3X1_766 ( .A(u5__abc_78290_new_n716_), .B(u5__abc_78290_new_n392_), .C(u5__abc_78290_new_n718_), .Y(u5__abc_78290_new_n719_));
NAND3X1 NAND3X1_767 ( .A(u5__abc_78290_new_n725_), .B(u5__abc_78290_new_n411_), .C(u5__abc_78290_new_n727_), .Y(u5__abc_78290_new_n728_));
NAND3X1 NAND3X1_768 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n729_), .Y(u5__abc_78290_new_n730_));
NAND3X1 NAND3X1_769 ( .A(u5__abc_78290_new_n733_), .B(u5__abc_78290_new_n419_), .C(u5__abc_78290_new_n420_), .Y(u5__abc_78290_new_n734_));
NAND3X1 NAND3X1_77 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1518_), .C(u0__abc_74894_new_n1526_), .Y(u0__abc_74894_new_n1527_));
NAND3X1 NAND3X1_770 ( .A(u5_state_7_), .B(u5__abc_78290_new_n417_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n735_));
NAND3X1 NAND3X1_771 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n737_), .Y(u5__abc_78290_new_n738_));
NAND3X1 NAND3X1_772 ( .A(u5__abc_78290_new_n740_), .B(u5__abc_78290_new_n411_), .C(u5__abc_78290_new_n742_), .Y(u5__abc_78290_new_n743_));
NAND3X1 NAND3X1_773 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n744_), .Y(u5__abc_78290_new_n745_));
NAND3X1 NAND3X1_774 ( .A(u5__abc_78290_new_n749_), .B(u5__abc_78290_new_n750_), .C(u5__abc_78290_new_n684_), .Y(u5__abc_78290_new_n751_));
NAND3X1 NAND3X1_775 ( .A(u5__abc_78290_new_n447_), .B(u5__abc_78290_new_n755_), .C(u5__abc_78290_new_n684_), .Y(u5__abc_78290_new_n756_));
NAND3X1 NAND3X1_776 ( .A(u5__abc_78290_new_n758_), .B(u5__abc_78290_new_n392_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n759_));
NAND3X1 NAND3X1_777 ( .A(u5_state_14_), .B(u5__abc_78290_new_n410_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n760_));
NAND3X1 NAND3X1_778 ( .A(u5__abc_78290_new_n765_), .B(u5__abc_78290_new_n392_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n766_));
NAND3X1 NAND3X1_779 ( .A(u5__abc_78290_new_n419_), .B(u5__abc_78290_new_n420_), .C(u5__abc_78290_new_n772_), .Y(u5__abc_78290_new_n773_));
NAND3X1 NAND3X1_78 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1542_), .C(u0__abc_74894_new_n1541_), .Y(u0__abc_74894_new_n1543_));
NAND3X1 NAND3X1_780 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n774_), .Y(u5__abc_78290_new_n775_));
NAND3X1 NAND3X1_781 ( .A(u5_state_6_), .B(u5__abc_78290_new_n417_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n780_));
NAND3X1 NAND3X1_782 ( .A(u5__abc_78290_new_n779_), .B(u5__abc_78290_new_n781_), .C(u5__abc_78290_new_n684_), .Y(u5__abc_78290_new_n782_));
NAND3X1 NAND3X1_783 ( .A(u5__abc_78290_new_n787_), .B(u5__abc_78290_new_n419_), .C(u5__abc_78290_new_n418_), .Y(u5__abc_78290_new_n788_));
NAND3X1 NAND3X1_784 ( .A(u5_state_1_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n789_), .Y(u5__abc_78290_new_n790_));
NAND3X1 NAND3X1_785 ( .A(u5__abc_78290_new_n793_), .B(u5__abc_78290_new_n419_), .C(u5__abc_78290_new_n418_), .Y(u5__abc_78290_new_n794_));
NAND3X1 NAND3X1_786 ( .A(u5_state_0_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n795_), .Y(u5__abc_78290_new_n796_));
NAND3X1 NAND3X1_787 ( .A(u5__abc_78290_new_n473_), .B(u5__abc_78290_new_n800_), .C(u5__abc_78290_new_n801_), .Y(u5__abc_78290_new_n802_));
NAND3X1 NAND3X1_788 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n803_), .Y(u5__abc_78290_new_n804_));
NAND3X1 NAND3X1_789 ( .A(u5__abc_78290_new_n513_), .B(u5__abc_78290_new_n404_), .C(u5__abc_78290_new_n402_), .Y(u5__abc_78290_new_n806_));
NAND3X1 NAND3X1_79 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1540_), .C(u0__abc_74894_new_n1543_), .Y(u0__abc_74894_new_n1544_));
NAND3X1 NAND3X1_790 ( .A(u5__abc_78290_new_n423_), .B(u5__abc_78290_new_n684_), .C(u5__abc_78290_new_n807_), .Y(u5__abc_78290_new_n808_));
NAND3X1 NAND3X1_791 ( .A(u5__abc_78290_new_n811_), .B(u5__abc_78290_new_n813_), .C(u5__abc_78290_new_n465_), .Y(u5__abc_78290_new_n814_));
NAND3X1 NAND3X1_792 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n820_), .Y(u5__abc_78290_new_n821_));
NAND3X1 NAND3X1_793 ( .A(u5__abc_78290_new_n823_), .B(u5__abc_78290_new_n412_), .C(u5__abc_78290_new_n413_), .Y(u5__abc_78290_new_n824_));
NAND3X1 NAND3X1_794 ( .A(u5_state_12_), .B(u5__abc_78290_new_n409_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n825_));
NAND3X1 NAND3X1_795 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n827_), .Y(u5__abc_78290_new_n828_));
NAND3X1 NAND3X1_796 ( .A(u5__abc_78290_new_n829_), .B(u5__abc_78290_new_n412_), .C(u5__abc_78290_new_n413_), .Y(u5__abc_78290_new_n830_));
NAND3X1 NAND3X1_797 ( .A(u5_state_15_), .B(u5__abc_78290_new_n410_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n831_));
NAND3X1 NAND3X1_798 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n833_), .Y(u5__abc_78290_new_n834_));
NAND3X1 NAND3X1_799 ( .A(u5_state_62_), .B(u5__abc_78290_new_n379_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n841_));
NAND3X1 NAND3X1_8 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1185_), .C(u0__abc_74894_new_n1184_), .Y(u0__abc_74894_new_n1186_));
NAND3X1 NAND3X1_80 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1545_), .C(u0__abc_74894_new_n1544_), .Y(u0__abc_74894_new_n1546_));
NAND3X1 NAND3X1_800 ( .A(u5__abc_78290_new_n840_), .B(u5__abc_78290_new_n383_), .C(u5__abc_78290_new_n842_), .Y(u5__abc_78290_new_n843_));
NAND3X1 NAND3X1_801 ( .A(u5__abc_78290_new_n846_), .B(u5__abc_78290_new_n381_), .C(u5__abc_78290_new_n382_), .Y(u5__abc_78290_new_n847_));
NAND3X1 NAND3X1_802 ( .A(u5__abc_78290_new_n848_), .B(u5__abc_78290_new_n851_), .C(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n852_));
NAND3X1 NAND3X1_803 ( .A(u5__abc_78290_new_n854_), .B(u5__abc_78290_new_n381_), .C(u5__abc_78290_new_n382_), .Y(u5__abc_78290_new_n855_));
NAND3X1 NAND3X1_804 ( .A(u5__abc_78290_new_n856_), .B(u5__abc_78290_new_n858_), .C(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n859_));
NAND3X1 NAND3X1_805 ( .A(u5__abc_78290_new_n418_), .B(u5__abc_78290_new_n863_), .C(u5__abc_78290_new_n865_), .Y(u5__abc_78290_new_n866_));
NAND3X1 NAND3X1_806 ( .A(u5__abc_78290_new_n684_), .B(u5__abc_78290_new_n867_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n868_));
NAND3X1 NAND3X1_807 ( .A(u5__abc_78290_new_n862_), .B(u5__abc_78290_new_n420_), .C(u5__abc_78290_new_n870_), .Y(u5__abc_78290_new_n871_));
NAND3X1 NAND3X1_808 ( .A(u5__abc_78290_new_n684_), .B(u5__abc_78290_new_n873_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n874_));
NAND3X1 NAND3X1_809 ( .A(u5__abc_78290_new_n868_), .B(u5__abc_78290_new_n874_), .C(u5__abc_78290_new_n861_), .Y(u5__abc_78290_new_n875_));
NAND3X1 NAND3X1_81 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1538_), .C(u0__abc_74894_new_n1546_), .Y(u0__abc_74894_new_n1547_));
NAND3X1 NAND3X1_810 ( .A(u5__abc_78290_new_n876_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n877_));
NAND3X1 NAND3X1_811 ( .A(u5__abc_78290_new_n379_), .B(u5__abc_78290_new_n461_), .C(u5__abc_78290_new_n879_), .Y(u5__abc_78290_new_n880_));
NAND3X1 NAND3X1_812 ( .A(u5__abc_78290_new_n837_), .B(u5__abc_78290_new_n885_), .C(u5__abc_78290_new_n786_), .Y(u5__abc_78290_new_n886_));
NAND3X1 NAND3X1_813 ( .A(u5__abc_78290_new_n889_), .B(u5__abc_78290_new_n411_), .C(u5__abc_78290_new_n890_), .Y(u5__abc_78290_new_n891_));
NAND3X1 NAND3X1_814 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n407_), .C(u5__abc_78290_new_n892_), .Y(u5__abc_78290_new_n893_));
NAND3X1 NAND3X1_815 ( .A(u5_state_36_), .B(u5__abc_78290_new_n400_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n896_));
NAND3X1 NAND3X1_816 ( .A(u5__abc_78290_new_n897_), .B(u5__abc_78290_new_n900_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n901_));
NAND3X1 NAND3X1_817 ( .A(u5__abc_78290_new_n903_), .B(u5__abc_78290_new_n906_), .C(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n907_));
NAND3X1 NAND3X1_818 ( .A(u5__abc_78290_new_n910_), .B(u5__abc_78290_new_n913_), .C(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n914_));
NAND3X1 NAND3X1_819 ( .A(u5__abc_78290_new_n917_), .B(u5__abc_78290_new_n919_), .C(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n920_));
NAND3X1 NAND3X1_82 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1562_), .C(u0__abc_74894_new_n1561_), .Y(u0__abc_74894_new_n1563_));
NAND3X1 NAND3X1_820 ( .A(u5__abc_78290_new_n901_), .B(u5__abc_78290_new_n922_), .C(u5__abc_78290_new_n916_), .Y(u5__abc_78290_new_n923_));
NAND3X1 NAND3X1_821 ( .A(u5__abc_78290_new_n924_), .B(u5__abc_78290_new_n926_), .C(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n927_));
NAND3X1 NAND3X1_822 ( .A(u5__abc_78290_new_n929_), .B(u5__abc_78290_new_n388_), .C(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n930_));
NAND3X1 NAND3X1_823 ( .A(u5__abc_78290_new_n931_), .B(u5__abc_78290_new_n934_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n935_));
NAND3X1 NAND3X1_824 ( .A(u5__abc_78290_new_n938_), .B(u5__abc_78290_new_n388_), .C(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n939_));
NAND3X1 NAND3X1_825 ( .A(u5__abc_78290_new_n940_), .B(u5__abc_78290_new_n943_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n944_));
NAND3X1 NAND3X1_826 ( .A(u5__abc_78290_new_n946_), .B(u5__abc_78290_new_n388_), .C(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n947_));
NAND3X1 NAND3X1_827 ( .A(u5__abc_78290_new_n948_), .B(u5__abc_78290_new_n950_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n951_));
NAND3X1 NAND3X1_828 ( .A(u5__abc_78290_new_n888_), .B(u5__abc_78290_new_n895_), .C(u5__abc_78290_new_n955_), .Y(u5__abc_78290_new_n956_));
NAND3X1 NAND3X1_829 ( .A(u5__abc_78290_new_n612_), .B(u5__abc_78290_new_n724_), .C(u5__abc_78290_new_n957_), .Y(u5__abc_78290_new_n958_));
NAND3X1 NAND3X1_83 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1560_), .C(u0__abc_74894_new_n1563_), .Y(u0__abc_74894_new_n1564_));
NAND3X1 NAND3X1_830 ( .A(u5__abc_78290_new_n961_), .B(u5__abc_78290_new_n966_), .C(u5__abc_78290_new_n965_), .Y(u5__abc_78290_new_n967_));
NAND3X1 NAND3X1_831 ( .A(u5__abc_78290_new_n976_), .B(u5__abc_78290_new_n388_), .C(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n977_));
NAND3X1 NAND3X1_832 ( .A(u5__abc_78290_new_n978_), .B(u5__abc_78290_new_n980_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n981_));
NAND3X1 NAND3X1_833 ( .A(u5__abc_78290_new_n845_), .B(u5__abc_78290_new_n985_), .C(u5__abc_78290_new_n884_), .Y(u5__abc_78290_new_n986_));
NAND3X1 NAND3X1_834 ( .A(u5__abc_78290_new_n648_), .B(u5__abc_78290_new_n659_), .C(u5__abc_78290_new_n987_), .Y(u5__abc_78290_new_n988_));
NAND3X1 NAND3X1_835 ( .A(u5__abc_78290_new_n666_), .B(u5__abc_78290_new_n702_), .C(u5__abc_78290_new_n624_), .Y(u5__abc_78290_new_n989_));
NAND3X1 NAND3X1_836 ( .A(u5__abc_78290_new_n992_), .B(u5__abc_78290_new_n995_), .C(u5__abc_78290_new_n990_), .Y(u5__abc_78290_new_n996_));
NAND3X1 NAND3X1_837 ( .A(u5__abc_78290_new_n1004_), .B(u5__abc_78290_new_n1007_), .C(u5__abc_78290_new_n1010_), .Y(u5__abc_78290_new_n1011_));
NAND3X1 NAND3X1_838 ( .A(u5__abc_78290_new_n1016_), .B(u5__abc_78290_new_n1015_), .C(u5__abc_78290_new_n1012_), .Y(u5__abc_78290_new_n1017_));
NAND3X1 NAND3X1_839 ( .A(u5__abc_78290_new_n421_), .B(u5__abc_78290_new_n1020_), .C(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n1021_));
NAND3X1 NAND3X1_84 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1565_), .C(u0__abc_74894_new_n1564_), .Y(u0__abc_74894_new_n1566_));
NAND3X1 NAND3X1_840 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n1022_), .Y(u5__abc_78290_new_n1023_));
NAND3X1 NAND3X1_841 ( .A(u5__abc_78290_new_n421_), .B(u5__abc_78290_new_n1024_), .C(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n1025_));
NAND3X1 NAND3X1_842 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n1026_), .Y(u5__abc_78290_new_n1027_));
NAND3X1 NAND3X1_843 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n545_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1029_));
NAND3X1 NAND3X1_844 ( .A(u5__abc_78290_new_n562_), .B(u5__abc_78290_new_n566_), .C(u5__abc_78290_new_n453_), .Y(u5__abc_78290_new_n1032_));
NAND3X1 NAND3X1_845 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n1033_), .Y(u5__abc_78290_new_n1034_));
NAND3X1 NAND3X1_846 ( .A(u5__abc_78290_new_n839_), .B(u5__abc_78290_new_n478_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1039_));
NAND3X1 NAND3X1_847 ( .A(u5__abc_78290_new_n840_), .B(u5_state_62_), .C(u5__abc_78290_new_n379_), .Y(u5__abc_78290_new_n1040_));
NAND3X1 NAND3X1_848 ( .A(u5__abc_78290_new_n461_), .B(u5__abc_78290_new_n1041_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1042_));
NAND3X1 NAND3X1_849 ( .A(u5__abc_78290_new_n378_), .B(u5__abc_78290_new_n461_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1044_));
NAND3X1 NAND3X1_85 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1558_), .C(u0__abc_74894_new_n1566_), .Y(u0__abc_74894_new_n1567_));
NAND3X1 NAND3X1_850 ( .A(u5__abc_78290_new_n1056_), .B(u5__abc_78290_new_n444_), .C(u5__abc_78290_new_n1055_), .Y(u5__abc_78290_new_n1057_));
NAND3X1 NAND3X1_851 ( .A(u5__abc_78290_new_n1059_), .B(u5__abc_78290_new_n444_), .C(u5__abc_78290_new_n1055_), .Y(u5__abc_78290_new_n1060_));
NAND3X1 NAND3X1_852 ( .A(u5_state_63_), .B(u5__abc_78290_new_n1065_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1066_));
NAND3X1 NAND3X1_853 ( .A(u5__abc_78290_new_n383_), .B(u5__abc_78290_new_n461_), .C(u5__abc_78290_new_n1067_), .Y(u5__abc_78290_new_n1068_));
NAND3X1 NAND3X1_854 ( .A(u5__abc_78290_new_n381_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1075_), .Y(u5__abc_78290_new_n1076_));
NAND3X1 NAND3X1_855 ( .A(u5__abc_78290_new_n386_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1080_), .Y(u5__abc_78290_new_n1081_));
NAND3X1 NAND3X1_856 ( .A(u5__abc_78290_new_n1082_), .B(u5__abc_78290_new_n1079_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1083_));
NAND3X1 NAND3X1_857 ( .A(u5__abc_78290_new_n385_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1086_), .Y(u5__abc_78290_new_n1087_));
NAND3X1 NAND3X1_858 ( .A(u5__abc_78290_new_n385_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1090_), .Y(u5__abc_78290_new_n1091_));
NAND3X1 NAND3X1_859 ( .A(u5_state_59_), .B(u5__abc_78290_new_n904_), .C(u5__abc_78290_new_n382_), .Y(u5__abc_78290_new_n1097_));
NAND3X1 NAND3X1_86 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1582_), .C(u0__abc_74894_new_n1581_), .Y(u0__abc_74894_new_n1583_));
NAND3X1 NAND3X1_860 ( .A(u5__abc_78290_new_n382_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1100_), .Y(u5__abc_78290_new_n1101_));
NAND3X1 NAND3X1_861 ( .A(u5__abc_78290_new_n381_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1106_), .Y(u5__abc_78290_new_n1107_));
NAND3X1 NAND3X1_862 ( .A(u5__abc_78290_new_n386_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1110_), .Y(u5__abc_78290_new_n1111_));
NAND3X1 NAND3X1_863 ( .A(u5_state_39_), .B(u5__abc_78290_new_n662_), .C(u5__abc_78290_new_n401_), .Y(u5__abc_78290_new_n1118_));
NAND3X1 NAND3X1_864 ( .A(u5__abc_78290_new_n698_), .B(u5_state_38_), .C(u5__abc_78290_new_n401_), .Y(u5__abc_78290_new_n1121_));
NAND3X1 NAND3X1_865 ( .A(u5_state_40_), .B(u5__abc_78290_new_n643_), .C(u5__abc_78290_new_n396_), .Y(u5__abc_78290_new_n1125_));
NAND3X1 NAND3X1_866 ( .A(u5_state_47_), .B(u5__abc_78290_new_n655_), .C(u5__abc_78290_new_n394_), .Y(u5__abc_78290_new_n1129_));
NAND3X1 NAND3X1_867 ( .A(u5__abc_78290_new_n388_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1140_), .Y(u5__abc_78290_new_n1141_));
NAND3X1 NAND3X1_868 ( .A(u5__abc_78290_new_n388_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1143_), .Y(u5__abc_78290_new_n1144_));
NAND3X1 NAND3X1_869 ( .A(u5__abc_78290_new_n703_), .B(u5_state_44_), .C(u5__abc_78290_new_n393_), .Y(u5__abc_78290_new_n1150_));
NAND3X1 NAND3X1_87 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1580_), .C(u0__abc_74894_new_n1583_), .Y(u0__abc_74894_new_n1584_));
NAND3X1 NAND3X1_870 ( .A(u5_state_43_), .B(u5__abc_78290_new_n711_), .C(u5__abc_78290_new_n397_), .Y(u5__abc_78290_new_n1153_));
NAND3X1 NAND3X1_871 ( .A(u5__abc_78290_new_n686_), .B(u5_state_46_), .C(u5__abc_78290_new_n394_), .Y(u5__abc_78290_new_n1158_));
NAND3X1 NAND3X1_872 ( .A(u5_state_45_), .B(u5__abc_78290_new_n692_), .C(u5__abc_78290_new_n393_), .Y(u5__abc_78290_new_n1162_));
NAND3X1 NAND3X1_873 ( .A(u5__abc_78290_new_n644_), .B(u5_state_41_), .C(u5__abc_78290_new_n396_), .Y(u5__abc_78290_new_n1172_));
NAND3X1 NAND3X1_874 ( .A(u5_state_37_), .B(u5__abc_78290_new_n677_), .C(u5__abc_78290_new_n400_), .Y(u5__abc_78290_new_n1176_));
NAND3X1 NAND3X1_875 ( .A(u5__abc_78290_new_n898_), .B(u5_state_36_), .C(u5__abc_78290_new_n400_), .Y(u5__abc_78290_new_n1179_));
NAND3X1 NAND3X1_876 ( .A(u5__abc_78290_new_n1072_), .B(u5__abc_78290_new_n1117_), .C(u5__abc_78290_new_n1185_), .Y(u5__abc_78290_new_n1186_));
NAND3X1 NAND3X1_877 ( .A(u5__abc_78290_new_n506_), .B(u5_state_26_), .C(u5__abc_78290_new_n435_), .Y(u5__abc_78290_new_n1202_));
NAND3X1 NAND3X1_878 ( .A(u5__abc_78290_new_n522_), .B(u5_state_28_), .C(u5__abc_78290_new_n451_), .Y(u5__abc_78290_new_n1213_));
NAND3X1 NAND3X1_879 ( .A(u5__abc_78290_new_n530_), .B(u5_state_33_), .C(u5__abc_78290_new_n403_), .Y(u5__abc_78290_new_n1217_));
NAND3X1 NAND3X1_88 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1585_), .C(u0__abc_74894_new_n1584_), .Y(u0__abc_74894_new_n1586_));
NAND3X1 NAND3X1_880 ( .A(u5__abc_78290_new_n602_), .B(u5__abc_78290_new_n818_), .C(u5__abc_78290_new_n453_), .Y(u5__abc_78290_new_n1220_));
NAND3X1 NAND3X1_881 ( .A(u5__abc_78290_new_n447_), .B(u5__abc_78290_new_n1227_), .C(u5__abc_78290_new_n1225_), .Y(u5__abc_78290_new_n1228_));
NAND3X1 NAND3X1_882 ( .A(u5__abc_78290_new_n410_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1230_), .Y(u5__abc_78290_new_n1231_));
NAND3X1 NAND3X1_883 ( .A(u5__abc_78290_new_n513_), .B(u5_state_34_), .C(u5__abc_78290_new_n404_), .Y(u5__abc_78290_new_n1236_));
NAND3X1 NAND3X1_884 ( .A(u5_state_27_), .B(u5__abc_78290_new_n548_), .C(u5__abc_78290_new_n435_), .Y(u5__abc_78290_new_n1241_));
NAND3X1 NAND3X1_885 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n1242_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1243_));
NAND3X1 NAND3X1_886 ( .A(u5__abc_78290_new_n404_), .B(u5__abc_78290_new_n1245_), .C(u5__abc_78290_new_n402_), .Y(u5__abc_78290_new_n1246_));
NAND3X1 NAND3X1_887 ( .A(u5__abc_78290_new_n447_), .B(u5__abc_78290_new_n1255_), .C(u5__abc_78290_new_n1225_), .Y(u5__abc_78290_new_n1256_));
NAND3X1 NAND3X1_888 ( .A(u5__abc_78290_new_n412_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1259_), .Y(u5__abc_78290_new_n1260_));
NAND3X1 NAND3X1_889 ( .A(u5__abc_78290_new_n412_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1264_), .Y(u5__abc_78290_new_n1265_));
NAND3X1 NAND3X1_89 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1578_), .C(u0__abc_74894_new_n1586_), .Y(u0__abc_74894_new_n1587_));
NAND3X1 NAND3X1_890 ( .A(u5__abc_78290_new_n410_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1269_), .Y(u5__abc_78290_new_n1270_));
NAND3X1 NAND3X1_891 ( .A(u5__abc_78290_new_n413_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n493_), .Y(u5__abc_78290_new_n1276_));
NAND3X1 NAND3X1_892 ( .A(u5__abc_78290_new_n413_), .B(u5__abc_78290_new_n428_), .C(u5__abc_78290_new_n1279_), .Y(u5__abc_78290_new_n1280_));
NAND3X1 NAND3X1_893 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1285_), .C(u5__abc_78290_new_n421_), .Y(u5__abc_78290_new_n1286_));
NAND3X1 NAND3X1_894 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1288_), .C(u5__abc_78290_new_n421_), .Y(u5__abc_78290_new_n1289_));
NAND3X1 NAND3X1_895 ( .A(u5__abc_78290_new_n628_), .B(u5__abc_78290_new_n421_), .C(u5__abc_78290_new_n626_), .Y(u5__abc_78290_new_n1295_));
NAND3X1 NAND3X1_896 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1308_), .C(u5__abc_78290_new_n418_), .Y(u5__abc_78290_new_n1309_));
NAND3X1 NAND3X1_897 ( .A(u5__abc_78290_new_n1301_), .B(u5__abc_78290_new_n1312_), .C(u5__abc_78290_new_n1306_), .Y(u5__abc_78290_new_n1313_));
NAND3X1 NAND3X1_898 ( .A(u5__abc_78290_new_n1330_), .B(u5__abc_78290_new_n1331_), .C(u5__abc_78290_new_n1329_), .Y(u5__abc_78290_new_n1332_));
NAND3X1 NAND3X1_899 ( .A(u5__abc_78290_new_n1354_), .B(u5__abc_78290_new_n1348_), .C(u5__abc_78290_new_n1352_), .Y(u5__abc_78290_new_n1355_));
NAND3X1 NAND3X1_9 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1178_), .C(u0__abc_74894_new_n1186_), .Y(u0__abc_74894_new_n1187_));
NAND3X1 NAND3X1_90 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1602_), .C(u0__abc_74894_new_n1601_), .Y(u0__abc_74894_new_n1603_));
NAND3X1 NAND3X1_900 ( .A(u5__abc_78290_new_n1357_), .B(u5__abc_78290_new_n1359_), .C(u5__abc_78290_new_n1201_), .Y(u5__abc_78290_new_n1360_));
NAND3X1 NAND3X1_901 ( .A(u5__abc_78290_new_n1282_), .B(u5__abc_78290_new_n1109_), .C(u5__abc_78290_new_n1368_), .Y(u5__abc_78290_new_n1369_));
NAND3X1 NAND3X1_902 ( .A(u5__abc_78290_new_n1370_), .B(u5__abc_78290_new_n1366_), .C(u5__abc_78290_new_n1367_), .Y(u5__abc_78290_new_n1371_));
NAND3X1 NAND3X1_903 ( .A(u5__abc_78290_new_n1393_), .B(u5__abc_78290_new_n1089_), .C(u5__abc_78290_new_n1395_), .Y(u5__abc_78290_new_n1396_));
NAND3X1 NAND3X1_904 ( .A(u5__abc_78290_new_n1379_), .B(u5__abc_78290_new_n1426_), .C(u5__abc_78290_new_n1347_), .Y(u5_cmd_0_));
NAND3X1 NAND3X1_905 ( .A(u5__abc_78290_new_n1193_), .B(u5__abc_78290_new_n1436_), .C(u5__abc_78290_new_n1437_), .Y(u5__abc_78290_new_n1438_));
NAND3X1 NAND3X1_906 ( .A(u5__abc_78290_new_n1445_), .B(u5__abc_78290_new_n1448_), .C(u5__abc_78290_new_n1373_), .Y(u5__abc_78290_new_n1449_));
NAND3X1 NAND3X1_907 ( .A(u5__abc_78290_new_n1444_), .B(u5__abc_78290_new_n1462_), .C(u5__abc_78290_new_n1379_), .Y(u5__abc_78290_new_n1463_));
NAND3X1 NAND3X1_908 ( .A(rfr_req), .B(u5__abc_78290_new_n997_), .C(u5__abc_78290_new_n1018_), .Y(u5__abc_78290_new_n1468_));
NAND3X1 NAND3X1_909 ( .A(u5__abc_78290_new_n1036_), .B(u5__abc_78290_new_n1470_), .C(u5__abc_78290_new_n1468_), .Y(u5__abc_78290_new_n1471_));
NAND3X1 NAND3X1_91 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1600_), .C(u0__abc_74894_new_n1603_), .Y(u0__abc_74894_new_n1604_));
NAND3X1 NAND3X1_910 ( .A(u5__abc_78290_new_n1494_), .B(u5__abc_78290_new_n1503_), .C(u5__abc_78290_new_n1499_), .Y(u5__abc_78290_new_n1504_));
NAND3X1 NAND3X1_911 ( .A(u5__abc_78290_new_n1390_), .B(u5__abc_78290_new_n1397_), .C(u5__abc_78290_new_n1445_), .Y(u5__abc_78290_new_n1505_));
NAND3X1 NAND3X1_912 ( .A(u5__abc_78290_new_n1489_), .B(u5__abc_78290_new_n1506_), .C(u5__abc_78290_new_n1485_), .Y(u5__abc_78290_new_n1507_));
NAND3X1 NAND3X1_913 ( .A(u5__abc_78290_new_n1444_), .B(u5__abc_78290_new_n1518_), .C(u5__abc_78290_new_n1516_), .Y(u5__abc_78290_new_n1519_));
NAND3X1 NAND3X1_914 ( .A(u5__abc_78290_new_n1157_), .B(u5__abc_78290_new_n1526_), .C(u5__abc_78290_new_n1528_), .Y(u5__abc_78290_new_n1529_));
NAND3X1 NAND3X1_915 ( .A(u5__abc_78290_new_n1525_), .B(u5__abc_78290_new_n995_), .C(u5__abc_78290_new_n1530_), .Y(u5__abc_78290_new_n1531_));
NAND3X1 NAND3X1_916 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n1539_), .C(u5__abc_78290_new_n418_), .Y(u5__abc_78290_new_n1540_));
NAND3X1 NAND3X1_917 ( .A(u5__abc_78290_new_n1437_), .B(u5__abc_78290_new_n1543_), .C(u5__abc_78290_new_n1547_), .Y(u5__abc_78290_new_n1548_));
NAND3X1 NAND3X1_918 ( .A(u5__abc_78290_new_n1555_), .B(u5__abc_78290_new_n1357_), .C(u5__abc_78290_new_n1553_), .Y(u5__abc_78290_new_n1556_));
NAND3X1 NAND3X1_919 ( .A(u5__abc_78290_new_n997_), .B(u5__abc_78290_new_n1575_), .C(u5__abc_78290_new_n1573_), .Y(u5__abc_78290_new_n1576_));
NAND3X1 NAND3X1_92 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1605_), .C(u0__abc_74894_new_n1604_), .Y(u0__abc_74894_new_n1606_));
NAND3X1 NAND3X1_920 ( .A(u5__abc_78290_new_n1577_), .B(u5__abc_78290_new_n1578_), .C(u5__abc_78290_new_n1584_), .Y(u5__abc_78290_new_n1585_));
NAND3X1 NAND3X1_921 ( .A(u5__abc_78290_new_n536_), .B(u5__abc_78290_new_n1588_), .C(u5__abc_78290_new_n769_), .Y(u5__abc_78290_new_n1589_));
NAND3X1 NAND3X1_922 ( .A(u5__abc_78290_new_n1563_), .B(u5__abc_78290_new_n1590_), .C(u5__abc_78290_new_n1550_), .Y(u5__abc_78290_new_n1591_));
NAND3X1 NAND3X1_923 ( .A(u5__abc_78290_new_n1406_), .B(u5__abc_78290_new_n1633_), .C(u5__abc_78290_new_n1632_), .Y(u5__abc_78290_new_n1634_));
NAND3X1 NAND3X1_924 ( .A(u5__abc_78290_new_n1109_), .B(u5__abc_78290_new_n1395_), .C(u5__abc_78290_new_n1643_), .Y(u5__abc_78290_new_n1644_));
NAND3X1 NAND3X1_925 ( .A(tms_s_1_), .B(u5__abc_78290_new_n1404_), .C(u5__abc_78290_new_n1632_), .Y(u5__abc_78290_new_n1661_));
NAND3X1 NAND3X1_926 ( .A(u5__abc_78290_new_n1692_), .B(u5__abc_78290_new_n369_), .C(u5__abc_78290_new_n1673_), .Y(u5__abc_78290_new_n1694_));
NAND3X1 NAND3X1_927 ( .A(1'h0), .B(u5__abc_78290_new_n1318_), .C(u5__abc_78290_new_n1675_), .Y(u5__abc_78290_new_n1697_));
NAND3X1 NAND3X1_928 ( .A(u5_state_32_), .B(u5__abc_78290_new_n467_), .C(u5__abc_78290_new_n403_), .Y(u5__abc_78290_new_n1713_));
NAND3X1 NAND3X1_929 ( .A(u5__abc_78290_new_n428_), .B(u5__abc_78290_new_n455_), .C(u5__abc_78290_new_n1716_), .Y(u5__abc_78290_new_n1717_));
NAND3X1 NAND3X1_93 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1598_), .C(u0__abc_74894_new_n1606_), .Y(u0__abc_74894_new_n1607_));
NAND3X1 NAND3X1_930 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n440_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1719_));
NAND3X1 NAND3X1_931 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n1214_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1721_));
NAND3X1 NAND3X1_932 ( .A(u5__abc_78290_new_n450_), .B(u5__abc_78290_new_n1195_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1730_));
NAND3X1 NAND3X1_933 ( .A(u5__abc_78290_new_n582_), .B(u5_state_24_), .C(u5__abc_78290_new_n434_), .Y(u5__abc_78290_new_n1733_));
NAND3X1 NAND3X1_934 ( .A(u5__abc_78290_new_n423_), .B(u5__abc_78290_new_n1735_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n1736_));
NAND3X1 NAND3X1_935 ( .A(u5__abc_78290_new_n588_), .B(u5__abc_78290_new_n1738_), .C(u5__abc_78290_new_n453_), .Y(u5__abc_78290_new_n1739_));
NAND3X1 NAND3X1_936 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n1745_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1746_));
NAND3X1 NAND3X1_937 ( .A(u5__abc_78290_new_n588_), .B(u5__abc_78290_new_n1748_), .C(u5__abc_78290_new_n453_), .Y(u5__abc_78290_new_n1749_));
NAND3X1 NAND3X1_938 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n1754_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1755_));
NAND3X1 NAND3X1_939 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n1757_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1758_));
NAND3X1 NAND3X1_94 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1622_), .C(u0__abc_74894_new_n1621_), .Y(u0__abc_74894_new_n1623_));
NAND3X1 NAND3X1_940 ( .A(u5__abc_78290_new_n423_), .B(u5__abc_78290_new_n1764_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n1765_));
NAND3X1 NAND3X1_941 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n1766_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1767_));
NAND3X1 NAND3X1_942 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n1770_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1771_));
NAND3X1 NAND3X1_943 ( .A(u5__abc_78290_new_n603_), .B(u5_state_21_), .C(u5__abc_78290_new_n429_), .Y(u5__abc_78290_new_n1772_));
NAND3X1 NAND3X1_944 ( .A(u5__abc_78290_new_n423_), .B(u5__abc_78290_new_n1774_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n1775_));
NAND3X1 NAND3X1_945 ( .A(u5_state_12_), .B(u5__abc_78290_new_n823_), .C(u5__abc_78290_new_n409_), .Y(u5__abc_78290_new_n1777_));
NAND3X1 NAND3X1_946 ( .A(u5__abc_78290_new_n414_), .B(u5__abc_78290_new_n1782_), .C(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n1783_));
NAND3X1 NAND3X1_947 ( .A(u5__abc_78290_new_n453_), .B(u5__abc_78290_new_n1788_), .C(u5__abc_78290_new_n423_), .Y(u5__abc_78290_new_n1789_));
NAND3X1 NAND3X1_948 ( .A(u5__abc_78290_new_n418_), .B(u5__abc_78290_new_n1791_), .C(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n1792_));
NAND3X1 NAND3X1_949 ( .A(u5__abc_78290_new_n1769_), .B(u5__abc_78290_new_n1795_), .C(u5__abc_78290_new_n1787_), .Y(u5__abc_78290_new_n1796_));
NAND3X1 NAND3X1_95 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1620_), .C(u0__abc_74894_new_n1623_), .Y(u0__abc_74894_new_n1624_));
NAND3X1 NAND3X1_950 ( .A(u5__abc_78290_new_n411_), .B(u5__abc_78290_new_n1797_), .C(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n1798_));
NAND3X1 NAND3X1_951 ( .A(u5__abc_78290_new_n411_), .B(u5__abc_78290_new_n1803_), .C(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n1804_));
NAND3X1 NAND3X1_952 ( .A(u5__abc_78290_new_n414_), .B(u5__abc_78290_new_n1807_), .C(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n1808_));
NAND3X1 NAND3X1_953 ( .A(u5__abc_78290_new_n747_), .B(u5_state_13_), .C(u5__abc_78290_new_n409_), .Y(u5__abc_78290_new_n1813_));
NAND3X1 NAND3X1_954 ( .A(u5__abc_78290_new_n411_), .B(u5__abc_78290_new_n1817_), .C(u5__abc_78290_new_n447_), .Y(u5__abc_78290_new_n1818_));
NAND3X1 NAND3X1_955 ( .A(u5__abc_78290_new_n421_), .B(u5__abc_78290_new_n1822_), .C(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n1823_));
NAND3X1 NAND3X1_956 ( .A(u5__abc_78290_new_n421_), .B(u5__abc_78290_new_n1825_), .C(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n1826_));
NAND3X1 NAND3X1_957 ( .A(u5__abc_78290_new_n1812_), .B(u5__abc_78290_new_n1802_), .C(u5__abc_78290_new_n1830_), .Y(u5__abc_78290_new_n1831_));
NAND3X1 NAND3X1_958 ( .A(u5__abc_78290_new_n1725_), .B(u5__abc_78290_new_n1762_), .C(u5__abc_78290_new_n1832_), .Y(u5__abc_78290_new_n1833_));
NAND3X1 NAND3X1_959 ( .A(u5_state_51_), .B(u5__abc_78290_new_n614_), .C(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n1834_));
NAND3X1 NAND3X1_96 ( .A(u0__abc_74894_new_n1119_), .B(u0__abc_74894_new_n1625_), .C(u0__abc_74894_new_n1624_), .Y(u0__abc_74894_new_n1626_));
NAND3X1 NAND3X1_960 ( .A(u5__abc_78290_new_n619_), .B(u5_state_50_), .C(u5__abc_78290_new_n389_), .Y(u5__abc_78290_new_n1839_));
NAND3X1 NAND3X1_961 ( .A(u5__abc_78290_new_n458_), .B(u5__abc_78290_new_n1840_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1841_));
NAND3X1 NAND3X1_962 ( .A(u5__abc_78290_new_n387_), .B(u5__abc_78290_new_n1844_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n1845_));
NAND3X1 NAND3X1_963 ( .A(u5__abc_78290_new_n458_), .B(u5__abc_78290_new_n1849_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1850_));
NAND3X1 NAND3X1_964 ( .A(u5__abc_78290_new_n476_), .B(u5__abc_78290_new_n1126_), .C(u5__abc_78290_new_n392_), .Y(u5__abc_78290_new_n1857_));
NAND3X1 NAND3X1_965 ( .A(u5__abc_78290_new_n392_), .B(u5__abc_78290_new_n1860_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n1861_));
NAND3X1 NAND3X1_966 ( .A(u5__abc_78290_new_n476_), .B(u5__abc_78290_new_n1163_), .C(u5__abc_78290_new_n392_), .Y(u5__abc_78290_new_n1868_));
NAND3X1 NAND3X1_967 ( .A(u5__abc_78290_new_n476_), .B(u5__abc_78290_new_n1151_), .C(u5__abc_78290_new_n392_), .Y(u5__abc_78290_new_n1871_));
NAND3X1 NAND3X1_968 ( .A(u5__abc_78290_new_n476_), .B(u5__abc_78290_new_n1170_), .C(u5__abc_78290_new_n392_), .Y(u5__abc_78290_new_n1878_));
NAND3X1 NAND3X1_969 ( .A(u5__abc_78290_new_n476_), .B(u5__abc_78290_new_n1173_), .C(u5__abc_78290_new_n392_), .Y(u5__abc_78290_new_n1879_));
NAND3X1 NAND3X1_97 ( .A(u0__abc_74894_new_n1112_), .B(u0__abc_74894_new_n1618_), .C(u0__abc_74894_new_n1626_), .Y(u0__abc_74894_new_n1627_));
NAND3X1 NAND3X1_970 ( .A(u5__abc_78290_new_n465_), .B(u5__abc_78290_new_n1177_), .C(u5__abc_78290_new_n392_), .Y(u5__abc_78290_new_n1882_));
NAND3X1 NAND3X1_971 ( .A(u5_state_63_), .B(u5__abc_78290_new_n1065_), .C(u5__abc_78290_new_n379_), .Y(u5__abc_78290_new_n1892_));
NAND3X1 NAND3X1_972 ( .A(u5__abc_78290_new_n461_), .B(u5__abc_78290_new_n1893_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1894_));
NAND3X1 NAND3X1_973 ( .A(u5__abc_78290_new_n461_), .B(u5__abc_78290_new_n1898_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1899_));
NAND3X1 NAND3X1_974 ( .A(u5__abc_78290_new_n461_), .B(u5__abc_78290_new_n1901_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1902_));
NAND3X1 NAND3X1_975 ( .A(u5__abc_78290_new_n444_), .B(u5__abc_78290_new_n1906_), .C(u5__abc_78290_new_n684_), .Y(u5__abc_78290_new_n1907_));
NAND3X1 NAND3X1_976 ( .A(u5__abc_78290_new_n418_), .B(u5__abc_78290_new_n1909_), .C(u5__abc_78290_new_n444_), .Y(u5__abc_78290_new_n1910_));
NAND3X1 NAND3X1_977 ( .A(u5__abc_78290_new_n1890_), .B(u5__abc_78290_new_n1896_), .C(u5__abc_78290_new_n1914_), .Y(u5__abc_78290_new_n1915_));
NAND3X1 NAND3X1_978 ( .A(u5__abc_78290_new_n458_), .B(u5__abc_78290_new_n1917_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1918_));
NAND3X1 NAND3X1_979 ( .A(u5__abc_78290_new_n458_), .B(u5__abc_78290_new_n1920_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1921_));
NAND3X1 NAND3X1_98 ( .A(u0__abc_74894_new_n1134_), .B(u0__abc_74894_new_n1642_), .C(u0__abc_74894_new_n1641_), .Y(u0__abc_74894_new_n1643_));
NAND3X1 NAND3X1_980 ( .A(u5__abc_78290_new_n407_), .B(u5__abc_78290_new_n455_), .C(u5__abc_78290_new_n1925_), .Y(u5__abc_78290_new_n1926_));
NAND3X1 NAND3X1_981 ( .A(u5__abc_78290_new_n380_), .B(u5__abc_78290_new_n1927_), .C(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n1928_));
NAND3X1 NAND3X1_982 ( .A(u5__abc_78290_new_n380_), .B(u5__abc_78290_new_n1931_), .C(u5__abc_78290_new_n461_), .Y(u5__abc_78290_new_n1932_));
NAND3X1 NAND3X1_983 ( .A(u5__abc_78290_new_n461_), .B(u5__abc_78290_new_n1935_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1936_));
NAND3X1 NAND3X1_984 ( .A(u5__abc_78290_new_n458_), .B(u5__abc_78290_new_n1940_), .C(u5__abc_78290_new_n407_), .Y(u5__abc_78290_new_n1941_));
NAND3X1 NAND3X1_985 ( .A(u5__abc_78290_new_n390_), .B(u5__abc_78290_new_n1943_), .C(u5__abc_78290_new_n458_), .Y(u5__abc_78290_new_n1944_));
NAND3X1 NAND3X1_986 ( .A(u5__abc_78290_new_n1923_), .B(u5__abc_78290_new_n1947_), .C(u5__abc_78290_new_n1938_), .Y(u5__abc_78290_new_n1948_));
NAND3X1 NAND3X1_987 ( .A(u5__abc_78290_new_n1867_), .B(u5__abc_78290_new_n1889_), .C(u5__abc_78290_new_n1949_), .Y(u5__abc_78290_new_n1950_));
NAND3X1 NAND3X1_988 ( .A(u5__abc_78290_new_n1711_), .B(u5__abc_78290_new_n1712_), .C(u5__abc_78290_new_n1951_), .Y(u5__abc_78290_new_n1952_));
NAND3X1 NAND3X1_989 ( .A(u5__abc_78290_new_n1706_), .B(u5__abc_78290_new_n370_), .C(u5__abc_78290_new_n369_), .Y(u5__abc_78290_new_n1953_));
NAND3X1 NAND3X1_99 ( .A(u0__abc_74894_new_n1125_), .B(u0__abc_74894_new_n1640_), .C(u0__abc_74894_new_n1643_), .Y(u0__abc_74894_new_n1644_));
NAND3X1 NAND3X1_990 ( .A(u5__abc_78290_new_n1579_), .B(u5__abc_78290_new_n1994_), .C(u5__abc_78290_new_n1988_), .Y(u5__abc_78290_new_n1995_));
NAND3X1 NAND3X1_991 ( .A(u5__abc_78290_new_n1263_), .B(u5__abc_78290_new_n1274_), .C(u5__abc_78290_new_n1570_), .Y(u5__abc_78290_new_n1999_));
NAND3X1 NAND3X1_992 ( .A(u5__abc_78290_new_n1544_), .B(u5__abc_78290_new_n2007_), .C(u5__abc_78290_new_n1986_), .Y(u5__abc_78290_new_n2008_));
NAND3X1 NAND3X1_993 ( .A(u5__abc_78290_new_n2026_), .B(u5__abc_78290_new_n2024_), .C(u5__abc_78290_new_n2023_), .Y(u5__abc_78290_new_n2027_));
NAND3X1 NAND3X1_994 ( .A(u5__abc_78290_new_n1354_), .B(u5__abc_78290_new_n1376_), .C(u5__abc_78290_new_n2028_), .Y(u5__abc_78290_new_n2029_));
NAND3X1 NAND3X1_995 ( .A(u5__abc_78290_new_n769_), .B(u5__abc_78290_new_n2035_), .C(u5__abc_78290_new_n2036_), .Y(u5__abc_78290_new_n2037_));
NAND3X1 NAND3X1_996 ( .A(u5__abc_78290_new_n472_), .B(u5__abc_78290_new_n1263_), .C(u5__abc_78290_new_n1552_), .Y(u5__abc_78290_new_n2042_));
NAND3X1 NAND3X1_997 ( .A(u5__abc_78290_new_n1563_), .B(u5__abc_78290_new_n2043_), .C(u5__abc_78290_new_n1550_), .Y(u5__abc_78290_new_n2044_));
NAND3X1 NAND3X1_998 ( .A(u5__abc_78290_new_n529_), .B(u5__abc_78290_new_n541_), .C(u5__abc_78290_new_n554_), .Y(u5__abc_78290_new_n2057_));
NAND3X1 NAND3X1_999 ( .A(u5__abc_78290_new_n505_), .B(u5__abc_78290_new_n587_), .C(u5__abc_78290_new_n2058_), .Y(u5__abc_78290_new_n2059_));
NOR2X1 NOR2X1_1 ( .A(init_ack), .B(lmr_ack), .Y(_abc_81086_new_n236_));
NOR2X1 NOR2X1_10 ( .A(cs_le), .B(cs_2_), .Y(u0__abc_74894_new_n3483_));
NOR2X1 NOR2X1_100 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n4475_));
NOR2X1 NOR2X1_1000 ( .A(u5__abc_78290_new_n670_), .B(u5__abc_78290_new_n681_), .Y(u5__abc_78290_new_n2874_));
NOR2X1 NOR2X1_1001 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n643_), .Y(u5__abc_78290_new_n2882_));
NOR2X1 NOR2X1_1002 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n711_), .Y(u5__abc_78290_new_n2887_));
NOR2X1 NOR2X1_1003 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n692_), .Y(u5__abc_78290_new_n2893_));
NOR2X1 NOR2X1_1004 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n655_), .Y(u5__abc_78290_new_n2902_));
NOR2X1 NOR2X1_1005 ( .A(u5__abc_78290_new_n1512_), .B(u5__abc_78290_new_n2864_), .Y(u5__abc_78290_new_n2905_));
NOR2X1 NOR2X1_1006 ( .A(u5__abc_78290_new_n2906_), .B(u5__abc_78290_new_n2613_), .Y(u5_next_state_47_));
NOR2X1 NOR2X1_1007 ( .A(u5__abc_78290_new_n1131_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n2908_));
NOR2X1 NOR2X1_1008 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n634_), .Y(u5__abc_78290_new_n2909_));
NOR2X1 NOR2X1_1009 ( .A(u5__abc_78290_new_n1600_), .B(u5__abc_78290_new_n1078_), .Y(u5__abc_78290_new_n2922_));
NOR2X1 NOR2X1_101 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n4476_));
NOR2X1 NOR2X1_1010 ( .A(u5_state_55_), .B(u5__abc_78290_new_n2930_), .Y(u5__abc_78290_new_n2934_));
NOR2X1 NOR2X1_1011 ( .A(u5__abc_78290_new_n1597_), .B(u5__abc_78290_new_n1083_), .Y(u5__abc_78290_new_n2937_));
NOR2X1 NOR2X1_1012 ( .A(u5__abc_78290_new_n911_), .B(u5__abc_78290_new_n1414_), .Y(u5__abc_78290_new_n2940_));
NOR2X1 NOR2X1_1013 ( .A(u5__abc_78290_new_n2943_), .B(u5__abc_78290_new_n1083_), .Y(u5__abc_78290_new_n2944_));
NOR2X1 NOR2X1_1014 ( .A(u3_wb_read_go), .B(u5__abc_78290_new_n1349_), .Y(u5__abc_78290_new_n2947_));
NOR2X1 NOR2X1_1015 ( .A(u5__abc_78290_new_n1414_), .B(u5__abc_78290_new_n1990_), .Y(u5__abc_78290_new_n2950_));
NOR2X1 NOR2X1_1016 ( .A(u5__abc_78290_new_n2147_), .B(u5__abc_78290_new_n1368_), .Y(u5__abc_78290_new_n2952_));
NOR2X1 NOR2X1_1017 ( .A(u5__abc_78290_new_n1606_), .B(u5__abc_78290_new_n1335_), .Y(u5__abc_78290_new_n2956_));
NOR2X1 NOR2X1_1018 ( .A(u5__abc_78290_new_n904_), .B(u5__abc_78290_new_n2591_), .Y(u5__abc_78290_new_n2957_));
NOR2X1 NOR2X1_1019 ( .A(u5__abc_78290_new_n2950_), .B(u5__abc_78290_new_n2959_), .Y(u5__abc_78290_new_n2960_));
NOR2X1 NOR2X1_102 ( .A(u0__abc_74894_new_n1100_), .B(u0__abc_74894_new_n4462_), .Y(u0_lmr_ack0));
NOR2X1 NOR2X1_1020 ( .A(u5_tmr2_done), .B(mc_ack_r), .Y(u5__abc_78290_new_n2970_));
NOR2X1 NOR2X1_1021 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n854_), .Y(u5__abc_78290_new_n2974_));
NOR2X1 NOR2X1_1022 ( .A(u5__abc_78290_new_n1335_), .B(u5__abc_78290_new_n1326_), .Y(u5__abc_78290_new_n2982_));
NOR2X1 NOR2X1_1023 ( .A(u5__abc_78290_new_n840_), .B(u5__abc_78290_new_n2591_), .Y(u5__abc_78290_new_n2983_));
NOR2X1 NOR2X1_1024 ( .A(u5__abc_78290_new_n2996_), .B(u5__abc_78290_new_n2995_), .Y(u5__abc_78290_new_n2997_));
NOR2X1 NOR2X1_1025 ( .A(u5__abc_78290_new_n1124_), .B(u5__abc_78290_new_n1182_), .Y(u5__abc_78290_new_n2998_));
NOR2X1 NOR2X1_1026 ( .A(u5__abc_78290_new_n3000_), .B(u5__abc_78290_new_n2994_), .Y(u5__abc_78290_new_n3001_));
NOR2X1 NOR2X1_1027 ( .A(u5__abc_78290_new_n1414_), .B(u5__abc_78290_new_n3003_), .Y(u5__abc_78290_new_n3004_));
NOR2X1 NOR2X1_1028 ( .A(u5__abc_78290_new_n2174_), .B(u5__abc_78290_new_n3011_), .Y(u5__abc_78290_new_n3012_));
NOR2X1 NOR2X1_1029 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n3013_), .Y(u5__abc_78290_new_n3014_));
NOR2X1 NOR2X1_103 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n4462_), .Y(u0_lmr_ack1));
NOR2X1 NOR2X1_1030 ( .A(u5__abc_78290_new_n3017_), .B(u5__abc_78290_new_n1305_), .Y(u5__abc_78290_new_n3018_));
NOR2X1 NOR2X1_1031 ( .A(u5__abc_78290_new_n3019_), .B(u5__abc_78290_new_n3016_), .Y(u5__abc_78290_new_n3020_));
NOR2X1 NOR2X1_1032 ( .A(u5__abc_78290_new_n2952_), .B(u5__abc_78290_new_n3023_), .Y(u5__abc_78290_new_n3024_));
NOR2X1 NOR2X1_1033 ( .A(lmr_req), .B(u5_susp_req_r), .Y(u5__abc_78290_new_n3026_));
NOR2X1 NOR2X1_1034 ( .A(u5__abc_78290_new_n1283_), .B(u5__abc_78290_new_n1234_), .Y(u5__abc_78290_new_n3028_));
NOR2X1 NOR2X1_1035 ( .A(u5__abc_78290_new_n3030_), .B(u5__abc_78290_new_n1989_), .Y(u5__abc_78290_new_n3031_));
NOR2X1 NOR2X1_1036 ( .A(u5__0no_wb_cycle_0_0_), .B(u5__abc_78290_new_n2650_), .Y(u5__abc_78290_new_n3042_));
NOR2X1 NOR2X1_1037 ( .A(u5__abc_78290_new_n3044_), .B(u5__abc_78290_new_n3045_), .Y(u5__abc_78290_new_n3046_));
NOR2X1 NOR2X1_1038 ( .A(u5__abc_78290_new_n3053_), .B(u5__abc_78290_new_n3054_), .Y(u5__abc_78290_new_n3055_));
NOR2X1 NOR2X1_1039 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n3057_), .Y(u5__abc_78290_new_n3058_));
NOR2X1 NOR2X1_104 ( .A(u0__abc_74894_new_n1100_), .B(u0__abc_74894_new_n4464_), .Y(u0_init_ack0));
NOR2X1 NOR2X1_1040 ( .A(u5__abc_78290_new_n3061_), .B(u5__abc_78290_new_n1542_), .Y(u5__abc_78290_new_n3062_));
NOR2X1 NOR2X1_1041 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n2177_), .Y(u5__abc_78290_new_n3064_));
NOR2X1 NOR2X1_1042 ( .A(u5__abc_78290_new_n1989_), .B(u5__abc_78290_new_n3067_), .Y(u5__abc_78290_new_n3068_));
NOR2X1 NOR2X1_1043 ( .A(u5__abc_78290_new_n1394_), .B(u5__abc_78290_new_n3073_), .Y(u5__abc_78290_new_n3074_));
NOR2X1 NOR2X1_1044 ( .A(u5__abc_78290_new_n1388_), .B(u5__abc_78290_new_n3075_), .Y(u5__abc_78290_new_n3076_));
NOR2X1 NOR2X1_1045 ( .A(u5__abc_78290_new_n1356_), .B(u5__abc_78290_new_n1353_), .Y(u5__abc_78290_new_n3078_));
NOR2X1 NOR2X1_1046 ( .A(u5__abc_78290_new_n3077_), .B(u5__abc_78290_new_n3079_), .Y(u5__abc_78290_new_n3080_));
NOR2X1 NOR2X1_1047 ( .A(u5__abc_78290_new_n1283_), .B(u5__abc_78290_new_n1275_), .Y(u5__abc_78290_new_n3084_));
NOR2X1 NOR2X1_1048 ( .A(u5__abc_78290_new_n1640_), .B(u5__abc_78290_new_n2206_), .Y(u5__abc_78290_new_n3087_));
NOR2X1 NOR2X1_1049 ( .A(u5__abc_78290_new_n3089_), .B(u5__abc_78290_new_n3090_), .Y(u5__abc_78290_new_n3091_));
NOR2X1 NOR2X1_105 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n4464_), .Y(u0_init_ack1));
NOR2X1 NOR2X1_1050 ( .A(u5__abc_78290_new_n1401_), .B(u5__abc_78290_new_n3075_), .Y(u5__abc_78290_new_n3092_));
NOR2X1 NOR2X1_1051 ( .A(u5__abc_78290_new_n1283_), .B(u5__abc_78290_new_n2183_), .Y(u5__abc_78290_new_n3093_));
NOR2X1 NOR2X1_1052 ( .A(u5__abc_78290_new_n2027_), .B(u5__abc_78290_new_n3095_), .Y(u5__abc_78290_new_n3096_));
NOR2X1 NOR2X1_1053 ( .A(u5__abc_78290_new_n3099_), .B(u5__abc_78290_new_n574_), .Y(u5__abc_78290_new_n3100_));
NOR2X1 NOR2X1_1054 ( .A(u5__abc_78290_new_n1356_), .B(u5__abc_78290_new_n1459_), .Y(u5__abc_78290_new_n3101_));
NOR2X1 NOR2X1_1055 ( .A(u5__abc_78290_new_n1094_), .B(u5__abc_78290_new_n3116_), .Y(u5__abc_78290_new_n3117_));
NOR2X1 NOR2X1_1056 ( .A(u5__abc_78290_new_n1484_), .B(u5__abc_78290_new_n3119_), .Y(u5__0oe__0_0_));
NOR2X1 NOR2X1_1057 ( .A(u5__abc_78290_new_n1532_), .B(u5__abc_78290_new_n1387_), .Y(u5__abc_78290_new_n3121_));
NOR2X1 NOR2X1_1058 ( .A(u5__abc_78290_new_n1116_), .B(u5__abc_78290_new_n3122_), .Y(u5__abc_78290_new_n3123_));
NOR2X1 NOR2X1_1059 ( .A(u5__abc_78290_new_n3124_), .B(u5__abc_78290_new_n1566_), .Y(u5_pack_le1_d));
NOR2X1 NOR2X1_106 ( .A(u0_csc0_2_), .B(u0_csc0_1_), .Y(u0_u0__abc_72207_new_n207_));
NOR2X1 NOR2X1_1060 ( .A(u5__abc_78290_new_n3127_), .B(u5__abc_78290_new_n1568_), .Y(err));
NOR2X1 NOR2X1_1061 ( .A(u5__abc_78290_new_n1999_), .B(u5__abc_78290_new_n1987_), .Y(u5__abc_78290_new_n3129_));
NOR2X1 NOR2X1_1062 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n3130_), .Y(init_ack));
NOR2X1 NOR2X1_1063 ( .A(u5__abc_78290_new_n1609_), .B(u5__abc_78290_new_n3132_), .Y(u5__abc_78290_new_n3133_));
NOR2X1 NOR2X1_1064 ( .A(u5__abc_78290_new_n1574_), .B(u5__abc_78290_new_n1562_), .Y(u5__abc_78290_new_n3136_));
NOR2X1 NOR2X1_1065 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n3138_), .Y(u5__abc_78290_new_n3139_));
NOR2X1 NOR2X1_1066 ( .A(u5__abc_78290_new_n2407_), .B(u5__abc_78290_new_n2413_), .Y(u5__abc_78290_new_n3145_));
NOR2X1 NOR2X1_1067 ( .A(u5__abc_78290_new_n3147_), .B(u5__abc_78290_new_n3146_), .Y(u5__0tmr2_done_0_0_));
NOR2X1 NOR2X1_1068 ( .A(\wb_addr_i[30] ), .B(\wb_addr_i[31] ), .Y(u6__abc_81318_new_n134_));
NOR2X1 NOR2X1_1069 ( .A(u6__abc_81318_new_n136_), .B(u6__abc_81318_new_n137_), .Y(u6__abc_81318_new_n138_));
NOR2X1 NOR2X1_107 ( .A(u0_u0__abc_72207_new_n205_), .B(u0_u0__abc_72207_new_n208_), .Y(u0_u0__abc_72207_new_n209_));
NOR2X1 NOR2X1_1070 ( .A(u6__abc_81318_new_n243_), .B(u6__abc_81318_new_n245_), .Y(u6__0rmw_r_0_0_));
NOR2X1 NOR2X1_1071 ( .A(u1_wr_hold), .B(u6__abc_81318_new_n253_), .Y(u6__abc_81318_new_n254_));
NOR2X1 NOR2X1_1072 ( .A(u6__abc_81318_new_n140_), .B(u6__abc_81318_new_n273_), .Y(u6__0wb_err_0_0_));
NOR2X1 NOR2X1_1073 ( .A(susp_sel), .B(rfr_ack), .Y(u7__abc_73829_new_n100_));
NOR2X1 NOR2X1_1074 ( .A(fs), .B(suspended_o), .Y(u7__0mc_rp_0_0_));
NOR2X1 NOR2X1_1075 ( .A(susp_sel), .B(u7__abc_73829_new_n155_), .Y(u7__0mc_data_oe_0_0_));
NOR2X1 NOR2X1_108 ( .A(u0_u0__abc_72207_new_n215_), .B(u0_u0__abc_72207_new_n218_), .Y(u0_u0__abc_72207_new_n219_));
NOR2X1 NOR2X1_109 ( .A(u0_u0__abc_72207_new_n442_), .B(u0_u0__abc_72207_new_n447_), .Y(u0_u0__abc_72207_new_n448_));
NOR2X1 NOR2X1_11 ( .A(cs_le), .B(cs_3_), .Y(u0__abc_74894_new_n3485_));
NOR2X1 NOR2X1_110 ( .A(u0_u0__abc_72207_new_n451_), .B(u0_u0__abc_72207_new_n456_), .Y(u0_u0__abc_72207_new_n457_));
NOR2X1 NOR2X1_111 ( .A(u0_u0__abc_72207_new_n434_), .B(u0_u0__abc_72207_new_n458_), .Y(u0_u0_wp_err));
NOR2X1 NOR2X1_112 ( .A(u0_u0_inited), .B(u0_u0__abc_72207_new_n325_), .Y(u0_u0__abc_72207_new_n463_));
NOR2X1 NOR2X1_113 ( .A(u0_csc1_2_), .B(u0_csc1_1_), .Y(u0_u1__abc_72470_new_n203_));
NOR2X1 NOR2X1_114 ( .A(u0_u1__abc_72470_new_n201_), .B(u0_u1__abc_72470_new_n204_), .Y(u0_u1__abc_72470_new_n205_));
NOR2X1 NOR2X1_115 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .Y(u0_u1__0lmr_req_we_0_0_));
NOR2X1 NOR2X1_116 ( .A(u0_u1__abc_72470_new_n212_), .B(u0_u1__abc_72470_new_n214_), .Y(u0_u1__abc_72470_new_n217_));
NOR2X1 NOR2X1_117 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .Y(u0_u1__0init_req_we_0_0_));
NOR2X1 NOR2X1_118 ( .A(u0_u1__abc_72470_new_n427_), .B(u0_u1__abc_72470_new_n432_), .Y(u0_u1__abc_72470_new_n433_));
NOR2X1 NOR2X1_119 ( .A(u0_u1__abc_72470_new_n411_), .B(u0_u1__abc_72470_new_n434_), .Y(u0_u1_wp_err));
NOR2X1 NOR2X1_12 ( .A(cs_le), .B(cs_4_), .Y(u0__abc_74894_new_n3487_));
NOR2X1 NOR2X1_120 ( .A(u1__abc_72801_new_n261_), .B(u1__abc_72801_new_n266_), .Y(u1__abc_72801_new_n267_));
NOR2X1 NOR2X1_121 ( .A(u1__abc_72801_new_n267_), .B(u1__abc_72801_new_n264_), .Y(u1__abc_72801_new_n268_));
NOR2X1 NOR2X1_122 ( .A(csc_s_5_), .B(csc_s_4_), .Y(u1__abc_72801_new_n278_));
NOR2X1 NOR2X1_123 ( .A(csc_s_7_), .B(csc_s_6_), .Y(u1__abc_72801_new_n279_));
NOR2X1 NOR2X1_124 ( .A(csc_s_5_), .B(u1__abc_72801_new_n269_), .Y(u1__abc_72801_new_n280_));
NOR2X1 NOR2X1_125 ( .A(csc_s_7_), .B(u1__abc_72801_new_n265_), .Y(u1__abc_72801_new_n281_));
NOR2X1 NOR2X1_126 ( .A(u1_bas), .B(u1__abc_72801_new_n285_), .Y(u1__abc_72801_new_n286_));
NOR2X1 NOR2X1_127 ( .A(u1__abc_72801_new_n266_), .B(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n289_));
NOR2X1 NOR2X1_128 ( .A(u1__abc_72801_new_n289_), .B(u1__abc_72801_new_n264_), .Y(u1__abc_72801_new_n290_));
NOR2X1 NOR2X1_129 ( .A(csc_s_4_), .B(u1__abc_72801_new_n260_), .Y(u1__abc_72801_new_n292_));
NOR2X1 NOR2X1_13 ( .A(cs_le), .B(cs_5_), .Y(u0__abc_74894_new_n3489_));
NOR2X1 NOR2X1_130 ( .A(u1__abc_72801_new_n287_), .B(u1__abc_72801_new_n294_), .Y(u1__abc_72801_new_n295_));
NOR2X1 NOR2X1_131 ( .A(u1_bas), .B(u1__abc_72801_new_n310_), .Y(u1__abc_72801_new_n311_));
NOR2X1 NOR2X1_132 ( .A(u1__abc_72801_new_n312_), .B(u1__abc_72801_new_n294_), .Y(u1__abc_72801_new_n313_));
NOR2X1 NOR2X1_133 ( .A(u1_bas), .B(u1__abc_72801_new_n326_), .Y(u1__abc_72801_new_n327_));
NOR2X1 NOR2X1_134 ( .A(csc_s_6_), .B(u1__abc_72801_new_n262_), .Y(u1__abc_72801_new_n335_));
NOR2X1 NOR2X1_135 ( .A(u1__abc_72801_new_n258_), .B(u1__abc_72801_new_n266_), .Y(u1__abc_72801_new_n340_));
NOR2X1 NOR2X1_136 ( .A(u1__abc_72801_new_n289_), .B(u1__abc_72801_new_n299_), .Y(u1__abc_72801_new_n349_));
NOR2X1 NOR2X1_137 ( .A(u1__abc_72801_new_n425_), .B(u1__abc_72801_new_n424_), .Y(u1__abc_72801_new_n426_));
NOR2X1 NOR2X1_138 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n414_), .Y(u1__abc_72801_new_n431_));
NOR2X1 NOR2X1_139 ( .A(u1__abc_72801_new_n287_), .B(u1__abc_72801_new_n274_), .Y(u1__abc_72801_new_n447_));
NOR2X1 NOR2X1_14 ( .A(cs_le), .B(cs_6_), .Y(u0__abc_74894_new_n3491_));
NOR2X1 NOR2X1_140 ( .A(cs_le), .B(wb_we_i), .Y(u1__abc_72801_new_n491_));
NOR2X1 NOR2X1_141 ( .A(u1__abc_72801_new_n280_), .B(u1__abc_72801_new_n292_), .Y(u1__abc_72801_new_n493_));
NOR2X1 NOR2X1_142 ( .A(u1__abc_72801_new_n460_), .B(u1__abc_72801_new_n261_), .Y(u1__abc_72801_new_n500_));
NOR2X1 NOR2X1_143 ( .A(u1__abc_72801_new_n537_), .B(u1__abc_72801_new_n261_), .Y(u1__abc_72801_new_n542_));
NOR2X1 NOR2X1_144 ( .A(wb_stb_i), .B(u1_sram_addr_0_), .Y(u1__abc_72801_new_n620_));
NOR2X1 NOR2X1_145 ( .A(wb_stb_i), .B(u1_sram_addr_1_), .Y(u1__abc_72801_new_n622_));
NOR2X1 NOR2X1_146 ( .A(wb_stb_i), .B(u1_sram_addr_2_), .Y(u1__abc_72801_new_n624_));
NOR2X1 NOR2X1_147 ( .A(wb_stb_i), .B(u1_sram_addr_3_), .Y(u1__abc_72801_new_n626_));
NOR2X1 NOR2X1_148 ( .A(wb_stb_i), .B(u1_sram_addr_4_), .Y(u1__abc_72801_new_n628_));
NOR2X1 NOR2X1_149 ( .A(wb_stb_i), .B(u1_sram_addr_5_), .Y(u1__abc_72801_new_n630_));
NOR2X1 NOR2X1_15 ( .A(u0_wb_addr_r_5_), .B(u0_wb_addr_r_4_), .Y(u0__abc_74894_new_n3594_));
NOR2X1 NOR2X1_150 ( .A(wb_stb_i), .B(u1_sram_addr_6_), .Y(u1__abc_72801_new_n632_));
NOR2X1 NOR2X1_151 ( .A(wb_stb_i), .B(u1_sram_addr_7_), .Y(u1__abc_72801_new_n634_));
NOR2X1 NOR2X1_152 ( .A(wb_stb_i), .B(u1_sram_addr_8_), .Y(u1__abc_72801_new_n636_));
NOR2X1 NOR2X1_153 ( .A(wb_stb_i), .B(u1_sram_addr_9_), .Y(u1__abc_72801_new_n638_));
NOR2X1 NOR2X1_154 ( .A(wb_stb_i), .B(u1_sram_addr_10_), .Y(u1__abc_72801_new_n640_));
NOR2X1 NOR2X1_155 ( .A(wb_stb_i), .B(u1_sram_addr_11_), .Y(u1__abc_72801_new_n642_));
NOR2X1 NOR2X1_156 ( .A(wb_stb_i), .B(u1_sram_addr_12_), .Y(u1__abc_72801_new_n644_));
NOR2X1 NOR2X1_157 ( .A(wb_stb_i), .B(u1_sram_addr_13_), .Y(u1__abc_72801_new_n646_));
NOR2X1 NOR2X1_158 ( .A(wb_stb_i), .B(u1_sram_addr_17_), .Y(u1__abc_72801_new_n657_));
NOR2X1 NOR2X1_159 ( .A(wb_stb_i), .B(u1_sram_addr_18_), .Y(u1__abc_72801_new_n659_));
NOR2X1 NOR2X1_16 ( .A(u0__abc_74894_new_n3597_), .B(u0__abc_74894_new_n3595_), .Y(u0__abc_74894_new_n3598_));
NOR2X1 NOR2X1_160 ( .A(wb_stb_i), .B(u1_sram_addr_19_), .Y(u1__abc_72801_new_n661_));
NOR2X1 NOR2X1_161 ( .A(wb_stb_i), .B(u1_sram_addr_20_), .Y(u1__abc_72801_new_n663_));
NOR2X1 NOR2X1_162 ( .A(wb_stb_i), .B(u1_sram_addr_21_), .Y(u1__abc_72801_new_n665_));
NOR2X1 NOR2X1_163 ( .A(wb_stb_i), .B(u1_sram_addr_22_), .Y(u1__abc_72801_new_n667_));
NOR2X1 NOR2X1_164 ( .A(wb_stb_i), .B(u1_sram_addr_23_), .Y(u1__abc_72801_new_n669_));
NOR2X1 NOR2X1_165 ( .A(csc_s_1_), .B(u1__abc_72801_new_n671_), .Y(u1__abc_72801_new_n672_));
NOR2X1 NOR2X1_166 ( .A(csc_s_3_), .B(csc_s_1_), .Y(u1__abc_72801_new_n674_));
NOR2X1 NOR2X1_167 ( .A(u1__abc_72801_new_n677_), .B(u1__abc_72801_new_n671_), .Y(u1__abc_72801_new_n678_));
NOR2X1 NOR2X1_168 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n680_), .Y(u1__abc_72801_new_n681_));
NOR2X1 NOR2X1_169 ( .A(cas_), .B(u1__abc_72801_new_n682_), .Y(u1__abc_72801_new_n683_));
NOR2X1 NOR2X1_17 ( .A(u0__abc_74894_new_n3633_), .B(u0__abc_74894_new_n3595_), .Y(u0__abc_74894_new_n3634_));
NOR2X1 NOR2X1_170 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n691_), .Y(u1__abc_72801_new_n692_));
NOR2X1 NOR2X1_171 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n699_), .Y(u1__abc_72801_new_n700_));
NOR2X1 NOR2X1_172 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n708_), .Y(u1__abc_72801_new_n709_));
NOR2X1 NOR2X1_173 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n716_), .Y(u1__abc_72801_new_n717_));
NOR2X1 NOR2X1_174 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n724_), .Y(u1__abc_72801_new_n725_));
NOR2X1 NOR2X1_175 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n732_), .Y(u1__abc_72801_new_n733_));
NOR2X1 NOR2X1_176 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n740_), .Y(u1__abc_72801_new_n741_));
NOR2X1 NOR2X1_177 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n748_), .Y(u1__abc_72801_new_n749_));
NOR2X1 NOR2X1_178 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n756_), .Y(u1__abc_72801_new_n757_));
NOR2X1 NOR2X1_179 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n765_), .Y(u1__abc_72801_new_n766_));
NOR2X1 NOR2X1_18 ( .A(\wb_addr_i[5] ), .B(\wb_addr_i[4] ), .Y(u0__abc_74894_new_n3688_));
NOR2X1 NOR2X1_180 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n773_), .Y(u1__abc_72801_new_n774_));
NOR2X1 NOR2X1_181 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n781_), .Y(u1__abc_72801_new_n782_));
NOR2X1 NOR2X1_182 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n786_), .Y(u1__abc_72801_new_n787_));
NOR2X1 NOR2X1_183 ( .A(u1__abc_72801_new_n676_), .B(u1__abc_72801_new_n820_), .Y(u1__abc_72801_new_n821_));
NOR2X1 NOR2X1_184 ( .A(u1_u0__abc_72719_new_n52_), .B(u1_u0__abc_72719_new_n57_), .Y(u1_u0__abc_72719_new_n58_));
NOR2X1 NOR2X1_185 ( .A(u1_u0__abc_72719_new_n60_), .B(u1_u0__abc_72719_new_n62_), .Y(u1_u0__0out_r_12_0__5_));
NOR2X1 NOR2X1_186 ( .A(u1_u0__abc_72719_new_n68_), .B(u1_u0__abc_72719_new_n69_), .Y(u1_u0__abc_72719_new_n70_));
NOR2X1 NOR2X1_187 ( .A(u1_u0__abc_72719_new_n74_), .B(u1_u0__abc_72719_new_n75_), .Y(u1_u0__abc_72719_new_n77_));
NOR2X1 NOR2X1_188 ( .A(u1_u0__abc_72719_new_n81_), .B(u1_u0__abc_72719_new_n82_), .Y(u1_u0__abc_72719_new_n83_));
NOR2X1 NOR2X1_189 ( .A(u1_u0__abc_72719_new_n99_), .B(u1_u0__abc_72719_new_n91_), .Y(u1_u0__abc_72719_new_n100_));
NOR2X1 NOR2X1_19 ( .A(u0__abc_74894_new_n3692_), .B(u0__abc_74894_new_n3689_), .Y(u0__abc_74894_new_n3693_));
NOR2X1 NOR2X1_190 ( .A(u1_u0__abc_72719_new_n104_), .B(u1_u0__abc_72719_new_n102_), .Y(u1_acs_addr_pl1_17_));
NOR2X1 NOR2X1_191 ( .A(u1_u0__abc_72719_new_n103_), .B(u1_u0__abc_72719_new_n108_), .Y(u1_u0__abc_72719_new_n109_));
NOR2X1 NOR2X1_192 ( .A(u1_u0_inc_next), .B(u1_acs_addr_12_), .Y(u1_u0__abc_72719_new_n129_));
NOR2X1 NOR2X1_193 ( .A(u1_u0__abc_72719_new_n129_), .B(u1_u0__abc_72719_new_n89_), .Y(u1_acs_addr_pl1_12_));
NOR2X1 NOR2X1_194 ( .A(u2__abc_74202_new_n64_), .B(u2__abc_74202_new_n65_), .Y(u2_bank_set_0));
NOR2X1 NOR2X1_195 ( .A(u2__abc_74202_new_n64_), .B(u2__abc_74202_new_n67_), .Y(u2_bank_set_1));
NOR2X1 NOR2X1_196 ( .A(u2__abc_74202_new_n65_), .B(u2__abc_74202_new_n81_), .Y(u2_bank_clr_0));
NOR2X1 NOR2X1_197 ( .A(u2__abc_74202_new_n67_), .B(u2__abc_74202_new_n81_), .Y(u2_bank_clr_1));
NOR2X1 NOR2X1_198 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .Y(u2_u0__abc_73914_new_n180_));
NOR2X1 NOR2X1_199 ( .A(bank_adr_0_), .B(u2_u0__abc_73914_new_n208_), .Y(u2_u0__abc_73914_new_n237_));
NOR2X1 NOR2X1_2 ( .A(susp_sel), .B(rfr_ack), .Y(_abc_81086_new_n240_));
NOR2X1 NOR2X1_20 ( .A(u0__abc_74894_new_n3695_), .B(u0__abc_74894_new_n3689_), .Y(u0__abc_74894_new_n3696_));
NOR2X1 NOR2X1_200 ( .A(u2_u0__abc_73914_new_n282_), .B(u2_u0__abc_73914_new_n273_), .Y(u2_u0__abc_73914_new_n283_));
NOR2X1 NOR2X1_201 ( .A(u2_u0_b3_last_row_10_), .B(row_adr_10_), .Y(u2_u0__abc_73914_new_n286_));
NOR2X1 NOR2X1_202 ( .A(u2_u0_b3_last_row_3_), .B(row_adr_3_), .Y(u2_u0__abc_73914_new_n289_));
NOR2X1 NOR2X1_203 ( .A(u2_u0__abc_73914_new_n313_), .B(u2_u0__abc_73914_new_n305_), .Y(u2_u0__abc_73914_new_n314_));
NOR2X1 NOR2X1_204 ( .A(u2_u0__abc_73914_new_n353_), .B(u2_u0__abc_73914_new_n363_), .Y(u2_u0__abc_73914_new_n364_));
NOR2X1 NOR2X1_205 ( .A(u2_u0__abc_73914_new_n382_), .B(u2_u0__abc_73914_new_n371_), .Y(u2_u0__abc_73914_new_n383_));
NOR2X1 NOR2X1_206 ( .A(row_adr_10_), .B(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_73914_new_n386_));
NOR2X1 NOR2X1_207 ( .A(row_adr_5_), .B(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_73914_new_n390_));
NOR2X1 NOR2X1_208 ( .A(u2_bank_clr_all_0), .B(u2_u0__abc_73914_new_n405_), .Y(u2_u0__abc_73914_new_n406_));
NOR2X1 NOR2X1_209 ( .A(u2_bank_clr_all_0), .B(u2_u0__abc_73914_new_n409_), .Y(u2_u0__abc_73914_new_n410_));
NOR2X1 NOR2X1_21 ( .A(u0__abc_74894_new_n3698_), .B(u0__abc_74894_new_n3689_), .Y(u0__abc_74894_new_n3699_));
NOR2X1 NOR2X1_210 ( .A(u2_bank_clr_all_0), .B(u2_u0__abc_73914_new_n399_), .Y(u2_u0__abc_73914_new_n415_));
NOR2X1 NOR2X1_211 ( .A(u2_u0__abc_73914_new_n404_), .B(u2_u0__abc_73914_new_n179_), .Y(u2_u0__abc_73914_new_n418_));
NOR2X1 NOR2X1_212 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .Y(u2_u1__abc_73914_new_n180_));
NOR2X1 NOR2X1_213 ( .A(bank_adr_0_), .B(u2_u1__abc_73914_new_n208_), .Y(u2_u1__abc_73914_new_n237_));
NOR2X1 NOR2X1_214 ( .A(u2_u1__abc_73914_new_n282_), .B(u2_u1__abc_73914_new_n273_), .Y(u2_u1__abc_73914_new_n283_));
NOR2X1 NOR2X1_215 ( .A(u2_u1_b3_last_row_10_), .B(row_adr_10_), .Y(u2_u1__abc_73914_new_n286_));
NOR2X1 NOR2X1_216 ( .A(u2_u1_b3_last_row_3_), .B(row_adr_3_), .Y(u2_u1__abc_73914_new_n289_));
NOR2X1 NOR2X1_217 ( .A(u2_u1__abc_73914_new_n313_), .B(u2_u1__abc_73914_new_n305_), .Y(u2_u1__abc_73914_new_n314_));
NOR2X1 NOR2X1_218 ( .A(u2_u1__abc_73914_new_n353_), .B(u2_u1__abc_73914_new_n363_), .Y(u2_u1__abc_73914_new_n364_));
NOR2X1 NOR2X1_219 ( .A(u2_u1__abc_73914_new_n382_), .B(u2_u1__abc_73914_new_n371_), .Y(u2_u1__abc_73914_new_n383_));
NOR2X1 NOR2X1_22 ( .A(u0__abc_74894_new_n3700_), .B(u0__abc_74894_new_n3689_), .Y(u0__abc_74894_new_n3701_));
NOR2X1 NOR2X1_220 ( .A(row_adr_10_), .B(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_73914_new_n386_));
NOR2X1 NOR2X1_221 ( .A(row_adr_5_), .B(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_73914_new_n390_));
NOR2X1 NOR2X1_222 ( .A(u2_bank_clr_all_1), .B(u2_u1__abc_73914_new_n405_), .Y(u2_u1__abc_73914_new_n406_));
NOR2X1 NOR2X1_223 ( .A(u2_bank_clr_all_1), .B(u2_u1__abc_73914_new_n409_), .Y(u2_u1__abc_73914_new_n410_));
NOR2X1 NOR2X1_224 ( .A(u2_bank_clr_all_1), .B(u2_u1__abc_73914_new_n399_), .Y(u2_u1__abc_73914_new_n415_));
NOR2X1 NOR2X1_225 ( .A(u2_u1__abc_73914_new_n404_), .B(u2_u1__abc_73914_new_n179_), .Y(u2_u1__abc_73914_new_n418_));
NOR2X1 NOR2X1_226 ( .A(csc_2_), .B(csc_3_), .Y(u3__abc_73372_new_n275_));
NOR2X1 NOR2X1_227 ( .A(csc_1_), .B(mem_ack_r), .Y(u3__abc_73372_new_n276_));
NOR2X1 NOR2X1_228 ( .A(u3_byte2_0_), .B(pack_le2), .Y(u3__abc_73372_new_n316_));
NOR2X1 NOR2X1_229 ( .A(pack_le2), .B(u3_byte2_1_), .Y(u3__abc_73372_new_n319_));
NOR2X1 NOR2X1_23 ( .A(\wb_addr_i[4] ), .B(u0__abc_74894_new_n3704_), .Y(u0__abc_74894_new_n3705_));
NOR2X1 NOR2X1_230 ( .A(pack_le2), .B(u3_byte2_2_), .Y(u3__abc_73372_new_n322_));
NOR2X1 NOR2X1_231 ( .A(pack_le2), .B(u3_byte2_3_), .Y(u3__abc_73372_new_n325_));
NOR2X1 NOR2X1_232 ( .A(pack_le2), .B(u3_byte2_4_), .Y(u3__abc_73372_new_n328_));
NOR2X1 NOR2X1_233 ( .A(pack_le2), .B(u3_byte2_5_), .Y(u3__abc_73372_new_n331_));
NOR2X1 NOR2X1_234 ( .A(pack_le2), .B(u3_byte2_6_), .Y(u3__abc_73372_new_n334_));
NOR2X1 NOR2X1_235 ( .A(pack_le2), .B(u3_byte2_7_), .Y(u3__abc_73372_new_n337_));
NOR2X1 NOR2X1_236 ( .A(csc_4_), .B(csc_5_), .Y(u3__abc_73372_new_n339_));
NOR2X1 NOR2X1_237 ( .A(csc_5_), .B(u3__abc_73372_new_n344_), .Y(u3__abc_73372_new_n345_));
NOR2X1 NOR2X1_238 ( .A(pack_le0), .B(u3_byte0_0_), .Y(u3__abc_73372_new_n386_));
NOR2X1 NOR2X1_239 ( .A(pack_le0), .B(u3_byte0_1_), .Y(u3__abc_73372_new_n388_));
NOR2X1 NOR2X1_24 ( .A(\wb_addr_i[6] ), .B(u0__abc_74894_new_n3700_), .Y(u0__abc_74894_new_n3706_));
NOR2X1 NOR2X1_240 ( .A(pack_le0), .B(u3_byte0_2_), .Y(u3__abc_73372_new_n390_));
NOR2X1 NOR2X1_241 ( .A(pack_le0), .B(u3_byte0_3_), .Y(u3__abc_73372_new_n392_));
NOR2X1 NOR2X1_242 ( .A(pack_le0), .B(u3_byte0_4_), .Y(u3__abc_73372_new_n394_));
NOR2X1 NOR2X1_243 ( .A(pack_le0), .B(u3_byte0_5_), .Y(u3__abc_73372_new_n396_));
NOR2X1 NOR2X1_244 ( .A(pack_le0), .B(u3_byte0_6_), .Y(u3__abc_73372_new_n398_));
NOR2X1 NOR2X1_245 ( .A(pack_le0), .B(u3_byte0_7_), .Y(u3__abc_73372_new_n400_));
NOR2X1 NOR2X1_246 ( .A(u3_rd_fifo_out_8_), .B(u3_rd_fifo_out_9_), .Y(u3__abc_73372_new_n635_));
NOR2X1 NOR2X1_247 ( .A(u3_rd_fifo_out_20_), .B(u3_rd_fifo_out_21_), .Y(u3__abc_73372_new_n664_));
NOR2X1 NOR2X1_248 ( .A(u3_rd_fifo_out_19_), .B(u3__abc_73372_new_n570_), .Y(u3__abc_73372_new_n666_));
NOR2X1 NOR2X1_249 ( .A(u3_rd_fifo_out_18_), .B(u3__abc_73372_new_n574_), .Y(u3__abc_73372_new_n667_));
NOR2X1 NOR2X1_25 ( .A(\wb_addr_i[6] ), .B(u0__abc_74894_new_n3692_), .Y(u0__abc_74894_new_n3710_));
NOR2X1 NOR2X1_250 ( .A(u3_rd_fifo_out_21_), .B(u3__abc_73372_new_n578_), .Y(u3__abc_73372_new_n669_));
NOR2X1 NOR2X1_251 ( .A(u3_rd_fifo_out_20_), .B(u3__abc_73372_new_n582_), .Y(u3__abc_73372_new_n670_));
NOR2X1 NOR2X1_252 ( .A(u3_rd_fifo_out_18_), .B(u3_rd_fifo_out_19_), .Y(u3__abc_73372_new_n671_));
NOR2X1 NOR2X1_253 ( .A(u3_rd_fifo_out_0_), .B(u3_rd_fifo_out_1_), .Y(u3__abc_73372_new_n680_));
NOR2X1 NOR2X1_254 ( .A(u3_rd_fifo_out_28_), .B(u3_rd_fifo_out_29_), .Y(u3__abc_73372_new_n714_));
NOR2X1 NOR2X1_255 ( .A(u3_rd_fifo_out_27_), .B(u3__abc_73372_new_n602_), .Y(u3__abc_73372_new_n716_));
NOR2X1 NOR2X1_256 ( .A(u3_rd_fifo_out_26_), .B(u3__abc_73372_new_n606_), .Y(u3__abc_73372_new_n717_));
NOR2X1 NOR2X1_257 ( .A(u3_rd_fifo_out_29_), .B(u3__abc_73372_new_n610_), .Y(u3__abc_73372_new_n719_));
NOR2X1 NOR2X1_258 ( .A(u3_rd_fifo_out_28_), .B(u3__abc_73372_new_n614_), .Y(u3__abc_73372_new_n720_));
NOR2X1 NOR2X1_259 ( .A(u3_rd_fifo_out_26_), .B(u3_rd_fifo_out_27_), .Y(u3__abc_73372_new_n721_));
NOR2X1 NOR2X1_26 ( .A(\wb_addr_i[6] ), .B(u0__abc_74894_new_n3695_), .Y(u0__abc_74894_new_n3712_));
NOR2X1 NOR2X1_260 ( .A(u3_u0__abc_74260_new_n654_), .B(u3_u0__abc_74260_new_n651_), .Y(u3_u0__abc_74260_new_n655_));
NOR2X1 NOR2X1_261 ( .A(u3_rd_fifo_clr), .B(u3_u0__abc_74260_new_n656_), .Y(u3_u0__0wr_adr_3_0__1_));
NOR2X1 NOR2X1_262 ( .A(u3_u0_r0_0_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n662_));
NOR2X1 NOR2X1_263 ( .A(u3_u0_r0_1_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n664_));
NOR2X1 NOR2X1_264 ( .A(u3_u0_r0_2_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n666_));
NOR2X1 NOR2X1_265 ( .A(u3_u0_r0_3_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n668_));
NOR2X1 NOR2X1_266 ( .A(u3_u0_r0_4_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n670_));
NOR2X1 NOR2X1_267 ( .A(u3_u0_r0_5_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n672_));
NOR2X1 NOR2X1_268 ( .A(u3_u0_r0_6_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n674_));
NOR2X1 NOR2X1_269 ( .A(u3_u0_r0_7_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n676_));
NOR2X1 NOR2X1_27 ( .A(\wb_addr_i[6] ), .B(u0__abc_74894_new_n3698_), .Y(u0__abc_74894_new_n3715_));
NOR2X1 NOR2X1_270 ( .A(u3_u0_r0_8_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n678_));
NOR2X1 NOR2X1_271 ( .A(u3_u0_r0_9_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n680_));
NOR2X1 NOR2X1_272 ( .A(u3_u0_r0_10_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n682_));
NOR2X1 NOR2X1_273 ( .A(u3_u0_r0_11_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n684_));
NOR2X1 NOR2X1_274 ( .A(u3_u0_r0_12_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n686_));
NOR2X1 NOR2X1_275 ( .A(u3_u0_r0_13_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n688_));
NOR2X1 NOR2X1_276 ( .A(u3_u0_r0_14_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n690_));
NOR2X1 NOR2X1_277 ( .A(u3_u0_r0_15_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n692_));
NOR2X1 NOR2X1_278 ( .A(u3_u0_r0_16_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n694_));
NOR2X1 NOR2X1_279 ( .A(u3_u0_r0_17_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n696_));
NOR2X1 NOR2X1_28 ( .A(u0__abc_74894_new_n3703_), .B(u0__abc_74894_new_n3722_), .Y(u0__abc_74894_new_n3723_));
NOR2X1 NOR2X1_280 ( .A(u3_u0_r0_18_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n698_));
NOR2X1 NOR2X1_281 ( .A(u3_u0_r0_19_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n700_));
NOR2X1 NOR2X1_282 ( .A(u3_u0_r0_20_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n702_));
NOR2X1 NOR2X1_283 ( .A(u3_u0_r0_21_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n704_));
NOR2X1 NOR2X1_284 ( .A(u3_u0_r0_22_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n706_));
NOR2X1 NOR2X1_285 ( .A(u3_u0_r0_23_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n708_));
NOR2X1 NOR2X1_286 ( .A(u3_u0_r0_24_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n710_));
NOR2X1 NOR2X1_287 ( .A(u3_u0_r0_25_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n712_));
NOR2X1 NOR2X1_288 ( .A(u3_u0_r0_26_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n714_));
NOR2X1 NOR2X1_289 ( .A(u3_u0_r0_27_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n716_));
NOR2X1 NOR2X1_29 ( .A(\wb_addr_i[6] ), .B(u0__abc_74894_new_n3730_), .Y(u0__abc_74894_new_n3731_));
NOR2X1 NOR2X1_290 ( .A(u3_u0_r0_28_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n718_));
NOR2X1 NOR2X1_291 ( .A(u3_u0_r0_29_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n720_));
NOR2X1 NOR2X1_292 ( .A(u3_u0_r0_30_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n722_));
NOR2X1 NOR2X1_293 ( .A(u3_u0_r0_31_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n724_));
NOR2X1 NOR2X1_294 ( .A(u3_u0_r0_32_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n726_));
NOR2X1 NOR2X1_295 ( .A(u3_u0_r0_33_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n728_));
NOR2X1 NOR2X1_296 ( .A(u3_u0_r0_34_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n730_));
NOR2X1 NOR2X1_297 ( .A(u3_u0_r0_35_), .B(u3_u0__abc_74260_new_n655_), .Y(u3_u0__abc_74260_new_n732_));
NOR2X1 NOR2X1_298 ( .A(u3_u0_rd_adr_0_), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_74260_new_n737_));
NOR2X1 NOR2X1_299 ( .A(u3_u0_rd_adr_2_), .B(u3_u0__abc_74260_new_n648_), .Y(u3_u0__abc_74260_new_n738_));
NOR2X1 NOR2X1_3 ( .A(\wb_addr_i[30] ), .B(\wb_addr_i[29] ), .Y(_abc_81086_new_n464_));
NOR2X1 NOR2X1_30 ( .A(u0__abc_74894_new_n3747_), .B(u0__abc_74894_new_n3753_), .Y(u0__abc_74894_new_n3754_));
NOR2X1 NOR2X1_300 ( .A(u3_u0_rd_adr_3_), .B(u3_u0__abc_74260_new_n645_), .Y(u3_u0__abc_74260_new_n739_));
NOR2X1 NOR2X1_301 ( .A(u3_u0__abc_74260_new_n734_), .B(u3_u0__abc_74260_new_n735_), .Y(u3_u0__abc_74260_new_n744_));
NOR2X1 NOR2X1_302 ( .A(u3_u0__abc_74260_new_n746_), .B(u3_u0__abc_74260_new_n745_), .Y(u3_u0__abc_74260_new_n747_));
NOR2X1 NOR2X1_303 ( .A(cs_need_rfr_2_), .B(cs_need_rfr_3_), .Y(u4__abc_74770_new_n65_));
NOR2X1 NOR2X1_304 ( .A(cs_need_rfr_0_), .B(cs_need_rfr_1_), .Y(u4__abc_74770_new_n66_));
NOR2X1 NOR2X1_305 ( .A(cs_need_rfr_6_), .B(cs_need_rfr_7_), .Y(u4__abc_74770_new_n68_));
NOR2X1 NOR2X1_306 ( .A(cs_need_rfr_4_), .B(cs_need_rfr_5_), .Y(u4__abc_74770_new_n69_));
NOR2X1 NOR2X1_307 ( .A(u4__abc_74770_new_n81_), .B(u4__abc_74770_new_n89_), .Y(u4__0rfr_early_0_0_));
NOR2X1 NOR2X1_308 ( .A(u4_rfr_clr), .B(rfr_req), .Y(u4__abc_74770_new_n91_));
NOR2X1 NOR2X1_309 ( .A(rfr_ack), .B(u4__abc_74770_new_n91_), .Y(u4__0rfr_req_0_0_));
NOR2X1 NOR2X1_31 ( .A(u0__abc_74894_new_n3758_), .B(u0__abc_74894_new_n3761_), .Y(u0__abc_74894_new_n3762_));
NOR2X1 NOR2X1_310 ( .A(u4__abc_74770_new_n93_), .B(u4__abc_74770_new_n95_), .Y(u4__0rfr_cnt_7_0__0_));
NOR2X1 NOR2X1_311 ( .A(u4__abc_74770_new_n99_), .B(u4__abc_74770_new_n98_), .Y(u4__0rfr_cnt_7_0__1_));
NOR2X1 NOR2X1_312 ( .A(u4__abc_74770_new_n101_), .B(u4__abc_74770_new_n102_), .Y(u4__abc_74770_new_n103_));
NOR2X1 NOR2X1_313 ( .A(u4__abc_74770_new_n103_), .B(u4__abc_74770_new_n104_), .Y(u4__0rfr_cnt_7_0__2_));
NOR2X1 NOR2X1_314 ( .A(u4__abc_74770_new_n106_), .B(u4__abc_74770_new_n102_), .Y(u4__abc_74770_new_n107_));
NOR2X1 NOR2X1_315 ( .A(u4__abc_74770_new_n110_), .B(u4__abc_74770_new_n113_), .Y(u4__0rfr_cnt_7_0__4_));
NOR2X1 NOR2X1_316 ( .A(rfr_ps_val_4_), .B(rfr_ps_val_5_), .Y(u4__abc_74770_new_n127_));
NOR2X1 NOR2X1_317 ( .A(rfr_ps_val_6_), .B(rfr_ps_val_7_), .Y(u4__abc_74770_new_n128_));
NOR2X1 NOR2X1_318 ( .A(rfr_ps_val_0_), .B(rfr_ps_val_1_), .Y(u4__abc_74770_new_n130_));
NOR2X1 NOR2X1_319 ( .A(rfr_ps_val_2_), .B(rfr_ps_val_3_), .Y(u4__abc_74770_new_n131_));
NOR2X1 NOR2X1_32 ( .A(u0__abc_74894_new_n3763_), .B(u0__abc_74894_new_n3767_), .Y(u0__abc_74894_new_n3768_));
NOR2X1 NOR2X1_320 ( .A(u4__abc_74770_new_n147_), .B(u4__abc_74770_new_n139_), .Y(u4__abc_74770_new_n148_));
NOR2X1 NOR2X1_321 ( .A(u4_rfr_cnt_1_), .B(u4__abc_74770_new_n174_), .Y(u4__abc_74770_new_n176_));
NOR2X1 NOR2X1_322 ( .A(u4__abc_74770_new_n111_), .B(u4__abc_74770_new_n102_), .Y(u4__abc_74770_new_n181_));
NOR2X1 NOR2X1_323 ( .A(u5_burst_cnt_1_), .B(u5_burst_cnt_0_), .Y(u5__abc_78290_new_n367_));
NOR2X1 NOR2X1_324 ( .A(u5_burst_cnt_3_), .B(u5__abc_78290_new_n368_), .Y(u5__abc_78290_new_n369_));
NOR2X1 NOR2X1_325 ( .A(u5_burst_cnt_5_), .B(u5_burst_cnt_4_), .Y(u5__abc_78290_new_n370_));
NOR2X1 NOR2X1_326 ( .A(u5_burst_cnt_7_), .B(u5_burst_cnt_6_), .Y(u5__abc_78290_new_n371_));
NOR2X1 NOR2X1_327 ( .A(u5_burst_cnt_9_), .B(u5_burst_cnt_8_), .Y(u5__abc_78290_new_n374_));
NOR2X1 NOR2X1_328 ( .A(u5__abc_78290_new_n375_), .B(u5__abc_78290_new_n372_), .Y(u5__abc_78290_new_n376_));
NOR2X1 NOR2X1_329 ( .A(u5_state_63_), .B(u5_state_62_), .Y(u5__abc_78290_new_n378_));
NOR2X1 NOR2X1_33 ( .A(u0__abc_74894_new_n3631_), .B(u0__abc_74894_new_n3770_), .Y(u0__abc_74894_new_n3771_));
NOR2X1 NOR2X1_330 ( .A(u5_state_61_), .B(u5_state_60_), .Y(u5__abc_78290_new_n379_));
NOR2X1 NOR2X1_331 ( .A(u5_state_59_), .B(u5_state_58_), .Y(u5__abc_78290_new_n381_));
NOR2X1 NOR2X1_332 ( .A(u5_state_57_), .B(u5_state_56_), .Y(u5__abc_78290_new_n382_));
NOR2X1 NOR2X1_333 ( .A(u5_state_55_), .B(u5_state_54_), .Y(u5__abc_78290_new_n385_));
NOR2X1 NOR2X1_334 ( .A(u5_state_53_), .B(u5_state_52_), .Y(u5__abc_78290_new_n386_));
NOR2X1 NOR2X1_335 ( .A(u5_state_51_), .B(u5_state_50_), .Y(u5__abc_78290_new_n388_));
NOR2X1 NOR2X1_336 ( .A(u5_state_49_), .B(u5_state_48_), .Y(u5__abc_78290_new_n389_));
NOR2X1 NOR2X1_337 ( .A(u5__abc_78290_new_n384_), .B(u5__abc_78290_new_n391_), .Y(u5__abc_78290_new_n392_));
NOR2X1 NOR2X1_338 ( .A(u5_state_47_), .B(u5_state_46_), .Y(u5__abc_78290_new_n393_));
NOR2X1 NOR2X1_339 ( .A(u5_state_45_), .B(u5_state_44_), .Y(u5__abc_78290_new_n394_));
NOR2X1 NOR2X1_34 ( .A(u0__abc_74894_new_n3780_), .B(u0__abc_74894_new_n3783_), .Y(u0__abc_74894_new_n3784_));
NOR2X1 NOR2X1_340 ( .A(u5_state_43_), .B(u5_state_42_), .Y(u5__abc_78290_new_n396_));
NOR2X1 NOR2X1_341 ( .A(u5_state_40_), .B(u5_state_41_), .Y(u5__abc_78290_new_n397_));
NOR2X1 NOR2X1_342 ( .A(u5_state_39_), .B(u5_state_38_), .Y(u5__abc_78290_new_n400_));
NOR2X1 NOR2X1_343 ( .A(u5_state_37_), .B(u5_state_36_), .Y(u5__abc_78290_new_n401_));
NOR2X1 NOR2X1_344 ( .A(u5_state_35_), .B(u5_state_34_), .Y(u5__abc_78290_new_n403_));
NOR2X1 NOR2X1_345 ( .A(u5_state_32_), .B(u5_state_33_), .Y(u5__abc_78290_new_n404_));
NOR2X1 NOR2X1_346 ( .A(u5__abc_78290_new_n399_), .B(u5__abc_78290_new_n406_), .Y(u5__abc_78290_new_n407_));
NOR2X1 NOR2X1_347 ( .A(u5_state_15_), .B(u5_state_14_), .Y(u5__abc_78290_new_n409_));
NOR2X1 NOR2X1_348 ( .A(u5_state_12_), .B(u5_state_13_), .Y(u5__abc_78290_new_n410_));
NOR2X1 NOR2X1_349 ( .A(u5_state_11_), .B(u5_state_10_), .Y(u5__abc_78290_new_n412_));
NOR2X1 NOR2X1_35 ( .A(u0__abc_74894_new_n3788_), .B(u0__abc_74894_new_n3787_), .Y(u0__abc_74894_new_n3789_));
NOR2X1 NOR2X1_350 ( .A(u5_state_9_), .B(u5_state_8_), .Y(u5__abc_78290_new_n413_));
NOR2X1 NOR2X1_351 ( .A(u5_state_7_), .B(u5_state_6_), .Y(u5__abc_78290_new_n416_));
NOR2X1 NOR2X1_352 ( .A(u5_state_5_), .B(u5_state_4_), .Y(u5__abc_78290_new_n417_));
NOR2X1 NOR2X1_353 ( .A(u5_state_3_), .B(u5_state_2_), .Y(u5__abc_78290_new_n419_));
NOR2X1 NOR2X1_354 ( .A(u5_state_1_), .B(u5_state_0_), .Y(u5__abc_78290_new_n420_));
NOR2X1 NOR2X1_355 ( .A(u5__abc_78290_new_n415_), .B(u5__abc_78290_new_n422_), .Y(u5__abc_78290_new_n423_));
NOR2X1 NOR2X1_356 ( .A(u5_state_19_), .B(u5_state_18_), .Y(u5__abc_78290_new_n424_));
NOR2X1 NOR2X1_357 ( .A(u5_state_17_), .B(u5_state_16_), .Y(u5__abc_78290_new_n425_));
NOR2X1 NOR2X1_358 ( .A(u5_state_20_), .B(u5_state_21_), .Y(u5__abc_78290_new_n427_));
NOR2X1 NOR2X1_359 ( .A(u5_state_65_), .B(u5_state_64_), .Y(u5__abc_78290_new_n428_));
NOR2X1 NOR2X1_36 ( .A(u0__abc_74894_new_n3637_), .B(u0__abc_74894_new_n3770_), .Y(u0__abc_74894_new_n3790_));
NOR2X1 NOR2X1_360 ( .A(u5_state_23_), .B(u5_state_22_), .Y(u5__abc_78290_new_n429_));
NOR2X1 NOR2X1_361 ( .A(u5__abc_78290_new_n426_), .B(u5__abc_78290_new_n430_), .Y(u5__abc_78290_new_n431_));
NOR2X1 NOR2X1_362 ( .A(u5__abc_78290_new_n432_), .B(u5__abc_78290_new_n408_), .Y(u5__abc_78290_new_n433_));
NOR2X1 NOR2X1_363 ( .A(u5_state_27_), .B(u5_state_26_), .Y(u5__abc_78290_new_n434_));
NOR2X1 NOR2X1_364 ( .A(u5_state_25_), .B(u5_state_24_), .Y(u5__abc_78290_new_n435_));
NOR2X1 NOR2X1_365 ( .A(u5_state_29_), .B(u5_state_28_), .Y(u5__abc_78290_new_n438_));
NOR2X1 NOR2X1_366 ( .A(u5__abc_78290_new_n436_), .B(u5__abc_78290_new_n439_), .Y(u5__abc_78290_new_n440_));
NOR2X1 NOR2X1_367 ( .A(u5__abc_78290_new_n442_), .B(u5__abc_78290_new_n443_), .Y(u5__abc_78290_new_n444_));
NOR2X1 NOR2X1_368 ( .A(u5__abc_78290_new_n445_), .B(u5__abc_78290_new_n446_), .Y(u5__abc_78290_new_n447_));
NOR2X1 NOR2X1_369 ( .A(u5__abc_78290_new_n426_), .B(u5__abc_78290_new_n449_), .Y(u5__abc_78290_new_n450_));
NOR2X1 NOR2X1_37 ( .A(u0__abc_74894_new_n3800_), .B(u0__abc_74894_new_n3804_), .Y(u0__abc_74894_new_n3805_));
NOR2X1 NOR2X1_370 ( .A(u5_state_30_), .B(u5_state_31_), .Y(u5__abc_78290_new_n451_));
NOR2X1 NOR2X1_371 ( .A(u5__abc_78290_new_n436_), .B(u5__abc_78290_new_n452_), .Y(u5__abc_78290_new_n453_));
NOR2X1 NOR2X1_372 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n454_), .Y(u5__abc_78290_new_n455_));
NOR2X1 NOR2X1_373 ( .A(u5__abc_78290_new_n456_), .B(u5__abc_78290_new_n457_), .Y(u5__abc_78290_new_n458_));
NOR2X1 NOR2X1_374 ( .A(u5__abc_78290_new_n459_), .B(u5__abc_78290_new_n460_), .Y(u5__abc_78290_new_n461_));
NOR2X1 NOR2X1_375 ( .A(u5__abc_78290_new_n463_), .B(u5__abc_78290_new_n464_), .Y(u5__abc_78290_new_n465_));
NOR2X1 NOR2X1_376 ( .A(u5__abc_78290_new_n466_), .B(u5__abc_78290_new_n468_), .Y(u5__abc_78290_new_n469_));
NOR2X1 NOR2X1_377 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n470_), .Y(u5__abc_78290_new_n471_));
NOR2X1 NOR2X1_378 ( .A(u5__abc_78290_new_n474_), .B(u5__abc_78290_new_n475_), .Y(u5__abc_78290_new_n476_));
NOR2X1 NOR2X1_379 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n477_), .Y(u5__abc_78290_new_n478_));
NOR2X1 NOR2X1_38 ( .A(u0__abc_74894_new_n3809_), .B(u0__abc_74894_new_n3813_), .Y(u0__abc_74894_new_n3814_));
NOR2X1 NOR2X1_380 ( .A(u5__abc_78290_new_n430_), .B(u5__abc_78290_new_n448_), .Y(u5__abc_78290_new_n479_));
NOR2X1 NOR2X1_381 ( .A(u5__abc_78290_new_n426_), .B(u5__abc_78290_new_n482_), .Y(u5__abc_78290_new_n483_));
NOR2X1 NOR2X1_382 ( .A(u5_cnt), .B(u5__abc_78290_new_n486_), .Y(u5__abc_78290_new_n487_));
NOR2X1 NOR2X1_383 ( .A(u5_state_10_), .B(u5__abc_78290_new_n492_), .Y(u5__abc_78290_new_n493_));
NOR2X1 NOR2X1_384 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n495_), .Y(u5__abc_78290_new_n496_));
NOR2X1 NOR2X1_385 ( .A(u5__abc_78290_new_n501_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n502_));
NOR2X1 NOR2X1_386 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n503_), .Y(u5__abc_78290_new_n504_));
NOR2X1 NOR2X1_387 ( .A(u5__abc_78290_new_n507_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n508_));
NOR2X1 NOR2X1_388 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n509_), .Y(u5__abc_78290_new_n510_));
NOR2X1 NOR2X1_389 ( .A(u5__abc_78290_new_n513_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n514_));
NOR2X1 NOR2X1_39 ( .A(u0__abc_74894_new_n3700_), .B(u0__abc_74894_new_n3815_), .Y(u0__abc_74894_new_n3816_));
NOR2X1 NOR2X1_390 ( .A(u5__abc_78290_new_n516_), .B(u5__abc_78290_new_n474_), .Y(u5__abc_78290_new_n517_));
NOR2X1 NOR2X1_391 ( .A(u5_state_31_), .B(u5__abc_78290_new_n524_), .Y(u5__abc_78290_new_n525_));
NOR2X1 NOR2X1_392 ( .A(u5__abc_78290_new_n481_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n526_));
NOR2X1 NOR2X1_393 ( .A(u5__abc_78290_new_n527_), .B(u5__abc_78290_new_n448_), .Y(u5__abc_78290_new_n528_));
NOR2X1 NOR2X1_394 ( .A(u5__abc_78290_new_n530_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n531_));
NOR2X1 NOR2X1_395 ( .A(u5__abc_78290_new_n532_), .B(u5__abc_78290_new_n474_), .Y(u5__abc_78290_new_n533_));
NOR2X1 NOR2X1_396 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n534_), .Y(u5__abc_78290_new_n535_));
NOR2X1 NOR2X1_397 ( .A(u5__abc_78290_new_n537_), .B(u5__abc_78290_new_n436_), .Y(u5__abc_78290_new_n538_));
NOR2X1 NOR2X1_398 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n539_), .Y(u5__abc_78290_new_n540_));
NOR2X1 NOR2X1_399 ( .A(u5__abc_78290_new_n436_), .B(u5__abc_78290_new_n544_), .Y(u5__abc_78290_new_n545_));
NOR2X1 NOR2X1_4 ( .A(u0__abc_74894_new_n1128_), .B(u0__abc_74894_new_n1137_), .Y(u0__abc_74894_new_n1144_));
NOR2X1 NOR2X1_40 ( .A(u0__abc_74894_new_n3825_), .B(u0__abc_74894_new_n3828_), .Y(u0__abc_74894_new_n3829_));
NOR2X1 NOR2X1_400 ( .A(u5__abc_78290_new_n549_), .B(u5__abc_78290_new_n452_), .Y(u5__abc_78290_new_n550_));
NOR2X1 NOR2X1_401 ( .A(u5__abc_78290_new_n559_), .B(u5__abc_78290_new_n557_), .Y(u5__abc_78290_new_n560_));
NOR2X1 NOR2X1_402 ( .A(u5__abc_78290_new_n565_), .B(u5__abc_78290_new_n563_), .Y(u5__abc_78290_new_n566_));
NOR2X1 NOR2X1_403 ( .A(u5__abc_78290_new_n567_), .B(u5__abc_78290_new_n448_), .Y(u5__abc_78290_new_n568_));
NOR2X1 NOR2X1_404 ( .A(u5__abc_78290_new_n573_), .B(u5__abc_78290_new_n570_), .Y(u5__abc_78290_new_n574_));
NOR2X1 NOR2X1_405 ( .A(u5_state_19_), .B(u5__abc_78290_new_n558_), .Y(u5__abc_78290_new_n575_));
NOR2X1 NOR2X1_406 ( .A(u5__abc_78290_new_n576_), .B(u5__abc_78290_new_n557_), .Y(u5__abc_78290_new_n577_));
NOR2X1 NOR2X1_407 ( .A(u5__abc_78290_new_n578_), .B(u5__abc_78290_new_n570_), .Y(u5__abc_78290_new_n579_));
NOR2X1 NOR2X1_408 ( .A(u5__abc_78290_new_n574_), .B(u5__abc_78290_new_n579_), .Y(u5__abc_78290_new_n580_));
NOR2X1 NOR2X1_409 ( .A(u5__abc_78290_new_n581_), .B(u5__abc_78290_new_n583_), .Y(u5__abc_78290_new_n584_));
NOR2X1 NOR2X1_41 ( .A(u0__abc_74894_new_n3643_), .B(u0__abc_74894_new_n3770_), .Y(u0__abc_74894_new_n3833_));
NOR2X1 NOR2X1_410 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n585_), .Y(u5__abc_78290_new_n586_));
NOR2X1 NOR2X1_411 ( .A(u5_state_22_), .B(u5__abc_78290_new_n590_), .Y(u5__abc_78290_new_n591_));
NOR2X1 NOR2X1_412 ( .A(u5__abc_78290_new_n592_), .B(u5__abc_78290_new_n448_), .Y(u5__abc_78290_new_n593_));
NOR2X1 NOR2X1_413 ( .A(u5_state_23_), .B(u5__abc_78290_new_n596_), .Y(u5__abc_78290_new_n597_));
NOR2X1 NOR2X1_414 ( .A(u5__abc_78290_new_n598_), .B(u5__abc_78290_new_n448_), .Y(u5__abc_78290_new_n599_));
NOR2X1 NOR2X1_415 ( .A(u5_state_21_), .B(u5__abc_78290_new_n603_), .Y(u5__abc_78290_new_n604_));
NOR2X1 NOR2X1_416 ( .A(u5__abc_78290_new_n605_), .B(u5__abc_78290_new_n448_), .Y(u5__abc_78290_new_n606_));
NOR2X1 NOR2X1_417 ( .A(u5__abc_78290_new_n608_), .B(u5__abc_78290_new_n595_), .Y(u5__abc_78290_new_n609_));
NOR2X1 NOR2X1_418 ( .A(u5__abc_78290_new_n556_), .B(u5__abc_78290_new_n611_), .Y(u5__abc_78290_new_n612_));
NOR2X1 NOR2X1_419 ( .A(u5__abc_78290_new_n613_), .B(u5__abc_78290_new_n615_), .Y(u5__abc_78290_new_n616_));
NOR2X1 NOR2X1_42 ( .A(u0__abc_74894_new_n3856_), .B(u0__abc_74894_new_n3852_), .Y(u0__abc_74894_new_n3857_));
NOR2X1 NOR2X1_420 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n617_), .Y(u5__abc_78290_new_n618_));
NOR2X1 NOR2X1_421 ( .A(u5__abc_78290_new_n620_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n621_));
NOR2X1 NOR2X1_422 ( .A(u5_state_5_), .B(u5__abc_78290_new_n627_), .Y(u5__abc_78290_new_n628_));
NOR2X1 NOR2X1_423 ( .A(u5__abc_78290_new_n415_), .B(u5__abc_78290_new_n629_), .Y(u5__abc_78290_new_n630_));
NOR2X1 NOR2X1_424 ( .A(u5__abc_78290_new_n632_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n633_));
NOR2X1 NOR2X1_425 ( .A(u5__abc_78290_new_n635_), .B(u5__abc_78290_new_n459_), .Y(u5__abc_78290_new_n636_));
NOR2X1 NOR2X1_426 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n637_), .Y(u5__abc_78290_new_n638_));
NOR2X1 NOR2X1_427 ( .A(u5__abc_78290_new_n640_), .B(u5__abc_78290_new_n625_), .Y(u5__abc_78290_new_n641_));
NOR2X1 NOR2X1_428 ( .A(u5__abc_78290_new_n406_), .B(u5__abc_78290_new_n462_), .Y(u5__abc_78290_new_n642_));
NOR2X1 NOR2X1_429 ( .A(u5__abc_78290_new_n644_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n645_));
NOR2X1 NOR2X1_43 ( .A(u0__abc_74894_new_n3866_), .B(u0__abc_74894_new_n3869_), .Y(u0__abc_74894_new_n3870_));
NOR2X1 NOR2X1_430 ( .A(u5__abc_78290_new_n463_), .B(u5__abc_78290_new_n646_), .Y(u5__abc_78290_new_n647_));
NOR2X1 NOR2X1_431 ( .A(u5__abc_78290_new_n634_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n649_));
NOR2X1 NOR2X1_432 ( .A(u5__abc_78290_new_n650_), .B(u5__abc_78290_new_n459_), .Y(u5__abc_78290_new_n651_));
NOR2X1 NOR2X1_433 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n652_), .Y(u5__abc_78290_new_n653_));
NOR2X1 NOR2X1_434 ( .A(u5__abc_78290_new_n657_), .B(u5__abc_78290_new_n656_), .Y(u5__abc_78290_new_n658_));
NOR2X1 NOR2X1_435 ( .A(u5__abc_78290_new_n399_), .B(u5__abc_78290_new_n462_), .Y(u5__abc_78290_new_n661_));
NOR2X1 NOR2X1_436 ( .A(u5__abc_78290_new_n664_), .B(u5__abc_78290_new_n663_), .Y(u5__abc_78290_new_n665_));
NOR2X1 NOR2X1_437 ( .A(u5__abc_78290_new_n667_), .B(u5__abc_78290_new_n660_), .Y(u5__abc_78290_new_n668_));
NOR2X1 NOR2X1_438 ( .A(u5_state_43_), .B(u5__abc_78290_new_n672_), .Y(u5__abc_78290_new_n673_));
NOR2X1 NOR2X1_439 ( .A(u5__abc_78290_new_n463_), .B(u5__abc_78290_new_n674_), .Y(u5__abc_78290_new_n675_));
NOR2X1 NOR2X1_44 ( .A(u0__abc_74894_new_n3649_), .B(u0__abc_74894_new_n3770_), .Y(u0__abc_74894_new_n3874_));
NOR2X1 NOR2X1_440 ( .A(u5__abc_78290_new_n679_), .B(u5__abc_78290_new_n678_), .Y(u5__abc_78290_new_n680_));
NOR2X1 NOR2X1_441 ( .A(u5__abc_78290_new_n683_), .B(u5__abc_78290_new_n557_), .Y(u5__abc_78290_new_n684_));
NOR2X1 NOR2X1_442 ( .A(u5__abc_78290_new_n689_), .B(u5__abc_78290_new_n406_), .Y(u5__abc_78290_new_n690_));
NOR2X1 NOR2X1_443 ( .A(u5__abc_78290_new_n694_), .B(u5__abc_78290_new_n693_), .Y(u5__abc_78290_new_n695_));
NOR2X1 NOR2X1_444 ( .A(u5__abc_78290_new_n700_), .B(u5__abc_78290_new_n699_), .Y(u5__abc_78290_new_n701_));
NOR2X1 NOR2X1_445 ( .A(u5__abc_78290_new_n705_), .B(u5__abc_78290_new_n704_), .Y(u5__abc_78290_new_n706_));
NOR2X1 NOR2X1_446 ( .A(u5__abc_78290_new_n708_), .B(u5__abc_78290_new_n697_), .Y(u5__abc_78290_new_n709_));
NOR2X1 NOR2X1_447 ( .A(u5__abc_78290_new_n710_), .B(u5__abc_78290_new_n712_), .Y(u5__abc_78290_new_n713_));
NOR2X1 NOR2X1_448 ( .A(u5__abc_78290_new_n671_), .B(u5__abc_78290_new_n714_), .Y(u5__abc_78290_new_n715_));
NOR2X1 NOR2X1_449 ( .A(u5__abc_78290_new_n643_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n716_));
NOR2X1 NOR2X1_45 ( .A(u0__abc_74894_new_n3884_), .B(u0__abc_74894_new_n3888_), .Y(u0__abc_74894_new_n3889_));
NOR2X1 NOR2X1_450 ( .A(u5__abc_78290_new_n406_), .B(u5__abc_78290_new_n717_), .Y(u5__abc_78290_new_n718_));
NOR2X1 NOR2X1_451 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n719_), .Y(u5__abc_78290_new_n720_));
NOR2X1 NOR2X1_452 ( .A(u5__abc_78290_new_n720_), .B(u5__abc_78290_new_n715_), .Y(u5__abc_78290_new_n721_));
NOR2X1 NOR2X1_453 ( .A(u5__abc_78290_new_n669_), .B(u5__abc_78290_new_n723_), .Y(u5__abc_78290_new_n724_));
NOR2X1 NOR2X1_454 ( .A(u5__abc_78290_new_n422_), .B(u5__abc_78290_new_n728_), .Y(u5__abc_78290_new_n729_));
NOR2X1 NOR2X1_455 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n730_), .Y(u5__abc_78290_new_n731_));
NOR2X1 NOR2X1_456 ( .A(u5__abc_78290_new_n734_), .B(u5__abc_78290_new_n735_), .Y(u5__abc_78290_new_n736_));
NOR2X1 NOR2X1_457 ( .A(u5__abc_78290_new_n422_), .B(u5__abc_78290_new_n743_), .Y(u5__abc_78290_new_n744_));
NOR2X1 NOR2X1_458 ( .A(u5__abc_78290_new_n746_), .B(u5__abc_78290_new_n748_), .Y(u5__abc_78290_new_n749_));
NOR2X1 NOR2X1_459 ( .A(u5__abc_78290_new_n754_), .B(u5__abc_78290_new_n442_), .Y(u5__abc_78290_new_n755_));
NOR2X1 NOR2X1_46 ( .A(u0__abc_74894_new_n3892_), .B(u0__abc_74894_new_n3897_), .Y(u0__abc_74894_new_n3898_));
NOR2X1 NOR2X1_460 ( .A(u5__abc_78290_new_n757_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n758_));
NOR2X1 NOR2X1_461 ( .A(u5__abc_78290_new_n760_), .B(u5__abc_78290_new_n422_), .Y(u5__abc_78290_new_n761_));
NOR2X1 NOR2X1_462 ( .A(u5__abc_78290_new_n753_), .B(u5__abc_78290_new_n768_), .Y(u5__abc_78290_new_n769_));
NOR2X1 NOR2X1_463 ( .A(u5_state_4_), .B(u5__abc_78290_new_n771_), .Y(u5__abc_78290_new_n772_));
NOR2X1 NOR2X1_464 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n775_), .Y(u5__abc_78290_new_n776_));
NOR2X1 NOR2X1_465 ( .A(u5__abc_78290_new_n780_), .B(u5__abc_78290_new_n415_), .Y(u5__abc_78290_new_n781_));
NOR2X1 NOR2X1_466 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n782_), .Y(u5__abc_78290_new_n783_));
NOR2X1 NOR2X1_467 ( .A(u5__abc_78290_new_n783_), .B(u5__abc_78290_new_n776_), .Y(u5__abc_78290_new_n784_));
NOR2X1 NOR2X1_468 ( .A(u5__abc_78290_new_n739_), .B(u5__abc_78290_new_n785_), .Y(u5__abc_78290_new_n786_));
NOR2X1 NOR2X1_469 ( .A(u5__abc_78290_new_n415_), .B(u5__abc_78290_new_n788_), .Y(u5__abc_78290_new_n789_));
NOR2X1 NOR2X1_47 ( .A(u0__abc_74894_new_n3903_), .B(u0__abc_74894_new_n3906_), .Y(u0__abc_74894_new_n3907_));
NOR2X1 NOR2X1_470 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n790_), .Y(u5__abc_78290_new_n791_));
NOR2X1 NOR2X1_471 ( .A(u5__abc_78290_new_n415_), .B(u5__abc_78290_new_n794_), .Y(u5__abc_78290_new_n795_));
NOR2X1 NOR2X1_472 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n796_), .Y(u5__abc_78290_new_n797_));
NOR2X1 NOR2X1_473 ( .A(u5_state_30_), .B(u5__abc_78290_new_n524_), .Y(u5__abc_78290_new_n800_));
NOR2X1 NOR2X1_474 ( .A(u5__abc_78290_new_n437_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n801_));
NOR2X1 NOR2X1_475 ( .A(u5__abc_78290_new_n683_), .B(u5__abc_78290_new_n802_), .Y(u5__abc_78290_new_n803_));
NOR2X1 NOR2X1_476 ( .A(u5__abc_78290_new_n805_), .B(u5__abc_78290_new_n806_), .Y(u5__abc_78290_new_n807_));
NOR2X1 NOR2X1_477 ( .A(u5__abc_78290_new_n809_), .B(u5__abc_78290_new_n799_), .Y(u5__abc_78290_new_n810_));
NOR2X1 NOR2X1_478 ( .A(u5__abc_78290_new_n467_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n811_));
NOR2X1 NOR2X1_479 ( .A(u5__abc_78290_new_n812_), .B(u5__abc_78290_new_n474_), .Y(u5__abc_78290_new_n813_));
NOR2X1 NOR2X1_48 ( .A(u0__abc_74894_new_n3920_), .B(u0__abc_74894_new_n3923_), .Y(u0__abc_74894_new_n3924_));
NOR2X1 NOR2X1_480 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n814_), .Y(u5__abc_78290_new_n815_));
NOR2X1 NOR2X1_481 ( .A(u5__abc_78290_new_n817_), .B(u5__abc_78290_new_n426_), .Y(u5__abc_78290_new_n818_));
NOR2X1 NOR2X1_482 ( .A(u5__abc_78290_new_n824_), .B(u5__abc_78290_new_n825_), .Y(u5__abc_78290_new_n826_));
NOR2X1 NOR2X1_483 ( .A(u5__abc_78290_new_n830_), .B(u5__abc_78290_new_n831_), .Y(u5__abc_78290_new_n832_));
NOR2X1 NOR2X1_484 ( .A(u5__abc_78290_new_n835_), .B(u5__abc_78290_new_n822_), .Y(u5__abc_78290_new_n836_));
NOR2X1 NOR2X1_485 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n685_), .Y(u5__abc_78290_new_n838_));
NOR2X1 NOR2X1_486 ( .A(u5_state_64_), .B(u5__abc_78290_new_n489_), .Y(u5__abc_78290_new_n839_));
NOR2X1 NOR2X1_487 ( .A(u5__abc_78290_new_n841_), .B(u5__abc_78290_new_n391_), .Y(u5__abc_78290_new_n842_));
NOR2X1 NOR2X1_488 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n843_), .Y(u5__abc_78290_new_n844_));
NOR2X1 NOR2X1_489 ( .A(u5__abc_78290_new_n849_), .B(u5__abc_78290_new_n850_), .Y(u5__abc_78290_new_n851_));
NOR2X1 NOR2X1_49 ( .A(u0__abc_74894_new_n3928_), .B(u0__abc_74894_new_n3932_), .Y(u0__abc_74894_new_n3933_));
NOR2X1 NOR2X1_490 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n852_), .Y(u5__abc_78290_new_n853_));
NOR2X1 NOR2X1_491 ( .A(u5__abc_78290_new_n849_), .B(u5__abc_78290_new_n857_), .Y(u5__abc_78290_new_n858_));
NOR2X1 NOR2X1_492 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n859_), .Y(u5__abc_78290_new_n860_));
NOR2X1 NOR2X1_493 ( .A(u5__abc_78290_new_n862_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n863_));
NOR2X1 NOR2X1_494 ( .A(u5_state_3_), .B(u5__abc_78290_new_n864_), .Y(u5__abc_78290_new_n865_));
NOR2X1 NOR2X1_495 ( .A(u5__abc_78290_new_n415_), .B(u5__abc_78290_new_n866_), .Y(u5__abc_78290_new_n867_));
NOR2X1 NOR2X1_496 ( .A(u5__abc_78290_new_n869_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n870_));
NOR2X1 NOR2X1_497 ( .A(u5__abc_78290_new_n871_), .B(u5__abc_78290_new_n872_), .Y(u5__abc_78290_new_n873_));
NOR2X1 NOR2X1_498 ( .A(u5_state_65_), .B(u5__abc_78290_new_n490_), .Y(u5__abc_78290_new_n876_));
NOR2X1 NOR2X1_499 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n880_), .Y(u5__abc_78290_new_n881_));
NOR2X1 NOR2X1_5 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3472_));
NOR2X1 NOR2X1_50 ( .A(u0__abc_74894_new_n3942_), .B(u0__abc_74894_new_n3945_), .Y(u0__abc_74894_new_n3946_));
NOR2X1 NOR2X1_500 ( .A(u5__abc_78290_new_n883_), .B(u5__abc_78290_new_n875_), .Y(u5__abc_78290_new_n884_));
NOR2X1 NOR2X1_501 ( .A(u5_dv_r), .B(u5__abc_78290_new_n887_), .Y(u5__abc_78290_new_n888_));
NOR2X1 NOR2X1_502 ( .A(u5__abc_78290_new_n422_), .B(u5__abc_78290_new_n891_), .Y(u5__abc_78290_new_n892_));
NOR2X1 NOR2X1_503 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n893_), .Y(u5__abc_78290_new_n894_));
NOR2X1 NOR2X1_504 ( .A(u5__abc_78290_new_n896_), .B(u5__abc_78290_new_n399_), .Y(u5__abc_78290_new_n897_));
NOR2X1 NOR2X1_505 ( .A(u5__abc_78290_new_n899_), .B(u5__abc_78290_new_n462_), .Y(u5__abc_78290_new_n900_));
NOR2X1 NOR2X1_506 ( .A(u5__abc_78290_new_n902_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n903_));
NOR2X1 NOR2X1_507 ( .A(u5__abc_78290_new_n905_), .B(u5__abc_78290_new_n456_), .Y(u5__abc_78290_new_n906_));
NOR2X1 NOR2X1_508 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n907_), .Y(u5__abc_78290_new_n908_));
NOR2X1 NOR2X1_509 ( .A(u5__abc_78290_new_n909_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n910_));
NOR2X1 NOR2X1_51 ( .A(u0__abc_74894_new_n3661_), .B(u0__abc_74894_new_n3770_), .Y(u0__abc_74894_new_n3950_));
NOR2X1 NOR2X1_510 ( .A(u5__abc_78290_new_n912_), .B(u5__abc_78290_new_n456_), .Y(u5__abc_78290_new_n913_));
NOR2X1 NOR2X1_511 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n914_), .Y(u5__abc_78290_new_n915_));
NOR2X1 NOR2X1_512 ( .A(u5__abc_78290_new_n904_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n917_));
NOR2X1 NOR2X1_513 ( .A(u5__abc_78290_new_n918_), .B(u5__abc_78290_new_n456_), .Y(u5__abc_78290_new_n919_));
NOR2X1 NOR2X1_514 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n920_), .Y(u5__abc_78290_new_n921_));
NOR2X1 NOR2X1_515 ( .A(u5__abc_78290_new_n911_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n924_));
NOR2X1 NOR2X1_516 ( .A(u5__abc_78290_new_n925_), .B(u5__abc_78290_new_n456_), .Y(u5__abc_78290_new_n926_));
NOR2X1 NOR2X1_517 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n927_), .Y(u5__abc_78290_new_n928_));
NOR2X1 NOR2X1_518 ( .A(u5__abc_78290_new_n932_), .B(u5__abc_78290_new_n933_), .Y(u5__abc_78290_new_n934_));
NOR2X1 NOR2X1_519 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n935_), .Y(u5__abc_78290_new_n936_));
NOR2X1 NOR2X1_52 ( .A(u0__abc_74894_new_n3961_), .B(u0__abc_74894_new_n3965_), .Y(u0__abc_74894_new_n3966_));
NOR2X1 NOR2X1_520 ( .A(u5__abc_78290_new_n941_), .B(u5__abc_78290_new_n942_), .Y(u5__abc_78290_new_n943_));
NOR2X1 NOR2X1_521 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n944_), .Y(u5__abc_78290_new_n945_));
NOR2X1 NOR2X1_522 ( .A(u5__abc_78290_new_n941_), .B(u5__abc_78290_new_n949_), .Y(u5__abc_78290_new_n950_));
NOR2X1 NOR2X1_523 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n951_), .Y(u5__abc_78290_new_n952_));
NOR2X1 NOR2X1_524 ( .A(u5__abc_78290_new_n954_), .B(u5__abc_78290_new_n923_), .Y(u5__abc_78290_new_n955_));
NOR2X1 NOR2X1_525 ( .A(u5__abc_78290_new_n956_), .B(u5__abc_78290_new_n886_), .Y(u5__abc_78290_new_n957_));
NOR2X1 NOR2X1_526 ( .A(u5_timer_1_), .B(u5_timer_2_), .Y(u5__abc_78290_new_n963_));
NOR2X1 NOR2X1_527 ( .A(u5_timer_3_), .B(u5__abc_78290_new_n964_), .Y(u5__abc_78290_new_n965_));
NOR2X1 NOR2X1_528 ( .A(u5_timer_5_), .B(u5_timer_4_), .Y(u5__abc_78290_new_n966_));
NOR2X1 NOR2X1_529 ( .A(u5_timer_7_), .B(u5__abc_78290_new_n967_), .Y(u5_timer_is_zero));
NOR2X1 NOR2X1_53 ( .A(u0__abc_74894_new_n3973_), .B(u0__abc_74894_new_n3969_), .Y(u0__abc_74894_new_n3974_));
NOR2X1 NOR2X1_530 ( .A(u5_ir_cnt_1_), .B(u5_ir_cnt_2_), .Y(u5__abc_78290_new_n970_));
NOR2X1 NOR2X1_531 ( .A(u5_ir_cnt_3_), .B(u5__abc_78290_new_n971_), .Y(u5__0ir_cnt_done_0_0_));
NOR2X1 NOR2X1_532 ( .A(u1_wb_write_go), .B(u3_wb_read_go), .Y(u5__0no_wb_cycle_0_0_));
NOR2X1 NOR2X1_533 ( .A(u5__abc_78290_new_n932_), .B(u5__abc_78290_new_n979_), .Y(u5__abc_78290_new_n980_));
NOR2X1 NOR2X1_534 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n981_), .Y(u5__abc_78290_new_n982_));
NOR2X1 NOR2X1_535 ( .A(u5__abc_78290_new_n954_), .B(u5__abc_78290_new_n984_), .Y(u5__abc_78290_new_n985_));
NOR2X1 NOR2X1_536 ( .A(u5__abc_78290_new_n988_), .B(u5__abc_78290_new_n989_), .Y(u5__abc_78290_new_n990_));
NOR2X1 NOR2X1_537 ( .A(u5__abc_78290_new_n697_), .B(u5__abc_78290_new_n991_), .Y(u5__abc_78290_new_n992_));
NOR2X1 NOR2X1_538 ( .A(u5__abc_78290_new_n994_), .B(u5__abc_78290_new_n993_), .Y(u5__abc_78290_new_n995_));
NOR2X1 NOR2X1_539 ( .A(u5__abc_78290_new_n986_), .B(u5__abc_78290_new_n996_), .Y(u5__abc_78290_new_n997_));
NOR2X1 NOR2X1_54 ( .A(u0__abc_74894_new_n3980_), .B(u0__abc_74894_new_n3984_), .Y(u0__abc_74894_new_n3985_));
NOR2X1 NOR2X1_540 ( .A(u5__abc_78290_new_n809_), .B(u5__abc_78290_new_n542_), .Y(u5__abc_78290_new_n1000_));
NOR2X1 NOR2X1_541 ( .A(u5__abc_78290_new_n1002_), .B(u5__abc_78290_new_n1003_), .Y(u5__abc_78290_new_n1004_));
NOR2X1 NOR2X1_542 ( .A(u5__abc_78290_new_n1005_), .B(u5__abc_78290_new_n1006_), .Y(u5__abc_78290_new_n1007_));
NOR2X1 NOR2X1_543 ( .A(u5__abc_78290_new_n1008_), .B(u5__abc_78290_new_n1009_), .Y(u5__abc_78290_new_n1010_));
NOR2X1 NOR2X1_544 ( .A(u5__abc_78290_new_n595_), .B(u5__abc_78290_new_n512_), .Y(u5__abc_78290_new_n1012_));
NOR2X1 NOR2X1_545 ( .A(u5__abc_78290_new_n1014_), .B(u5__abc_78290_new_n608_), .Y(u5__abc_78290_new_n1015_));
NOR2X1 NOR2X1_546 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1021_), .Y(u5__abc_78290_new_n1022_));
NOR2X1 NOR2X1_547 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1025_), .Y(u5__abc_78290_new_n1026_));
NOR2X1 NOR2X1_548 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1029_), .Y(u5__abc_78290_new_n1030_));
NOR2X1 NOR2X1_549 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n1032_), .Y(u5__abc_78290_new_n1033_));
NOR2X1 NOR2X1_55 ( .A(u0__abc_74894_new_n3992_), .B(u0__abc_74894_new_n3988_), .Y(u0__abc_74894_new_n3993_));
NOR2X1 NOR2X1_550 ( .A(u5__abc_78290_new_n457_), .B(u5__abc_78290_new_n1040_), .Y(u5__abc_78290_new_n1041_));
NOR2X1 NOR2X1_551 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1044_), .Y(u5__abc_78290_new_n1045_));
NOR2X1 NOR2X1_552 ( .A(u5_state_60_), .B(u5__abc_78290_new_n854_), .Y(u5__abc_78290_new_n1046_));
NOR2X1 NOR2X1_553 ( .A(u5__abc_78290_new_n457_), .B(u5__abc_78290_new_n1047_), .Y(u5__abc_78290_new_n1048_));
NOR2X1 NOR2X1_554 ( .A(u5_state_61_), .B(u5__abc_78290_new_n846_), .Y(u5__abc_78290_new_n1049_));
NOR2X1 NOR2X1_555 ( .A(u5__abc_78290_new_n457_), .B(u5__abc_78290_new_n1050_), .Y(u5__abc_78290_new_n1051_));
NOR2X1 NOR2X1_556 ( .A(u5__abc_78290_new_n445_), .B(u5__abc_78290_new_n1054_), .Y(u5__abc_78290_new_n1055_));
NOR2X1 NOR2X1_557 ( .A(u5_state_3_), .B(u5__abc_78290_new_n862_), .Y(u5__abc_78290_new_n1056_));
NOR2X1 NOR2X1_558 ( .A(u5__abc_78290_new_n1057_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1058_));
NOR2X1 NOR2X1_559 ( .A(u5_state_2_), .B(u5__abc_78290_new_n869_), .Y(u5__abc_78290_new_n1059_));
NOR2X1 NOR2X1_56 ( .A(u0__abc_74894_new_n3999_), .B(u0__abc_74894_new_n3998_), .Y(u0__abc_74894_new_n4000_));
NOR2X1 NOR2X1_560 ( .A(u5__abc_78290_new_n1060_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1061_));
NOR2X1 NOR2X1_561 ( .A(u5__abc_78290_new_n1058_), .B(u5__abc_78290_new_n1061_), .Y(u5__abc_78290_new_n1062_));
NOR2X1 NOR2X1_562 ( .A(u5__abc_78290_new_n1064_), .B(u5__abc_78290_new_n1066_), .Y(u5__abc_78290_new_n1067_));
NOR2X1 NOR2X1_563 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n1068_), .Y(u5__abc_78290_new_n1069_));
NOR2X1 NOR2X1_564 ( .A(u5__abc_78290_new_n1073_), .B(u5__abc_78290_new_n685_), .Y(u5__abc_78290_new_n1074_));
NOR2X1 NOR2X1_565 ( .A(u5_state_57_), .B(u5__abc_78290_new_n911_), .Y(u5__abc_78290_new_n1075_));
NOR2X1 NOR2X1_566 ( .A(u5__abc_78290_new_n1076_), .B(u5__abc_78290_new_n391_), .Y(u5__abc_78290_new_n1077_));
NOR2X1 NOR2X1_567 ( .A(u5__abc_78290_new_n384_), .B(u5__abc_78290_new_n477_), .Y(u5__abc_78290_new_n1079_));
NOR2X1 NOR2X1_568 ( .A(u5_state_54_), .B(u5__abc_78290_new_n976_), .Y(u5__abc_78290_new_n1080_));
NOR2X1 NOR2X1_569 ( .A(u5__abc_78290_new_n460_), .B(u5__abc_78290_new_n1081_), .Y(u5__abc_78290_new_n1082_));
NOR2X1 NOR2X1_57 ( .A(u0__abc_74894_new_n4010_), .B(u0__abc_74894_new_n4014_), .Y(u0__abc_74894_new_n4015_));
NOR2X1 NOR2X1_570 ( .A(u5_state_53_), .B(u5__abc_78290_new_n946_), .Y(u5__abc_78290_new_n1086_));
NOR2X1 NOR2X1_571 ( .A(u5__abc_78290_new_n460_), .B(u5__abc_78290_new_n1087_), .Y(u5__abc_78290_new_n1088_));
NOR2X1 NOR2X1_572 ( .A(u5_state_52_), .B(u5__abc_78290_new_n938_), .Y(u5__abc_78290_new_n1090_));
NOR2X1 NOR2X1_573 ( .A(u5__abc_78290_new_n460_), .B(u5__abc_78290_new_n1091_), .Y(u5__abc_78290_new_n1092_));
NOR2X1 NOR2X1_574 ( .A(u5__abc_78290_new_n1084_), .B(u5__abc_78290_new_n1094_), .Y(u5__abc_78290_new_n1095_));
NOR2X1 NOR2X1_575 ( .A(u5__abc_78290_new_n456_), .B(u5__abc_78290_new_n391_), .Y(u5__abc_78290_new_n1096_));
NOR2X1 NOR2X1_576 ( .A(u5__abc_78290_new_n1097_), .B(u5__abc_78290_new_n477_), .Y(u5__abc_78290_new_n1098_));
NOR2X1 NOR2X1_577 ( .A(u5_state_59_), .B(u5__abc_78290_new_n904_), .Y(u5__abc_78290_new_n1100_));
NOR2X1 NOR2X1_578 ( .A(u5__abc_78290_new_n1101_), .B(u5__abc_78290_new_n477_), .Y(u5__abc_78290_new_n1102_));
NOR2X1 NOR2X1_579 ( .A(u5_state_56_), .B(u5__abc_78290_new_n909_), .Y(u5__abc_78290_new_n1106_));
NOR2X1 NOR2X1_58 ( .A(u0__abc_74894_new_n4021_), .B(u0__abc_74894_new_n4020_), .Y(u0__abc_74894_new_n4022_));
NOR2X1 NOR2X1_580 ( .A(u5__abc_78290_new_n1107_), .B(u5__abc_78290_new_n391_), .Y(u5__abc_78290_new_n1108_));
NOR2X1 NOR2X1_581 ( .A(u5_state_55_), .B(u5__abc_78290_new_n929_), .Y(u5__abc_78290_new_n1110_));
NOR2X1 NOR2X1_582 ( .A(u5__abc_78290_new_n460_), .B(u5__abc_78290_new_n1111_), .Y(u5__abc_78290_new_n1112_));
NOR2X1 NOR2X1_583 ( .A(u5__abc_78290_new_n1105_), .B(u5__abc_78290_new_n1114_), .Y(u5__abc_78290_new_n1115_));
NOR2X1 NOR2X1_584 ( .A(u5__abc_78290_new_n475_), .B(u5__abc_78290_new_n1118_), .Y(u5__abc_78290_new_n1119_));
NOR2X1 NOR2X1_585 ( .A(u5__abc_78290_new_n475_), .B(u5__abc_78290_new_n1121_), .Y(u5__abc_78290_new_n1122_));
NOR2X1 NOR2X1_586 ( .A(u5__abc_78290_new_n463_), .B(u5__abc_78290_new_n1125_), .Y(u5__abc_78290_new_n1126_));
NOR2X1 NOR2X1_587 ( .A(u5__abc_78290_new_n464_), .B(u5__abc_78290_new_n1129_), .Y(u5__abc_78290_new_n1130_));
NOR2X1 NOR2X1_588 ( .A(u5__abc_78290_new_n1124_), .B(u5__abc_78290_new_n1132_), .Y(u5__abc_78290_new_n1133_));
NOR2X1 NOR2X1_589 ( .A(u5__abc_78290_new_n1138_), .B(u5__abc_78290_new_n685_), .Y(u5__abc_78290_new_n1139_));
NOR2X1 NOR2X1_59 ( .A(u0__abc_74894_new_n4032_), .B(u0__abc_74894_new_n4036_), .Y(u0__abc_74894_new_n4037_));
NOR2X1 NOR2X1_590 ( .A(u5_state_48_), .B(u5__abc_78290_new_n632_), .Y(u5__abc_78290_new_n1140_));
NOR2X1 NOR2X1_591 ( .A(u5__abc_78290_new_n1141_), .B(u5__abc_78290_new_n384_), .Y(u5__abc_78290_new_n1142_));
NOR2X1 NOR2X1_592 ( .A(u5_state_49_), .B(u5__abc_78290_new_n634_), .Y(u5__abc_78290_new_n1143_));
NOR2X1 NOR2X1_593 ( .A(u5__abc_78290_new_n1144_), .B(u5__abc_78290_new_n384_), .Y(u5__abc_78290_new_n1145_));
NOR2X1 NOR2X1_594 ( .A(u5__abc_78290_new_n464_), .B(u5__abc_78290_new_n1150_), .Y(u5__abc_78290_new_n1151_));
NOR2X1 NOR2X1_595 ( .A(u5__abc_78290_new_n463_), .B(u5__abc_78290_new_n1153_), .Y(u5__abc_78290_new_n1154_));
NOR2X1 NOR2X1_596 ( .A(u5__abc_78290_new_n464_), .B(u5__abc_78290_new_n1158_), .Y(u5__abc_78290_new_n1159_));
NOR2X1 NOR2X1_597 ( .A(u5__abc_78290_new_n1160_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1161_));
NOR2X1 NOR2X1_598 ( .A(u5__abc_78290_new_n464_), .B(u5__abc_78290_new_n1162_), .Y(u5__abc_78290_new_n1163_));
NOR2X1 NOR2X1_599 ( .A(u5__abc_78290_new_n1164_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1165_));
NOR2X1 NOR2X1_6 ( .A(1'h0), .B(u0_u0_wp_err), .Y(u0__abc_74894_new_n3473_));
NOR2X1 NOR2X1_60 ( .A(u0__abc_74894_new_n4042_), .B(u0__abc_74894_new_n4044_), .Y(u0__abc_74894_new_n4045_));
NOR2X1 NOR2X1_600 ( .A(u5__abc_78290_new_n1161_), .B(u5__abc_78290_new_n1165_), .Y(u5__abc_78290_new_n1166_));
NOR2X1 NOR2X1_601 ( .A(u5_state_43_), .B(u5__abc_78290_new_n711_), .Y(u5__abc_78290_new_n1168_));
NOR2X1 NOR2X1_602 ( .A(u5__abc_78290_new_n463_), .B(u5__abc_78290_new_n1169_), .Y(u5__abc_78290_new_n1170_));
NOR2X1 NOR2X1_603 ( .A(u5__abc_78290_new_n463_), .B(u5__abc_78290_new_n1172_), .Y(u5__abc_78290_new_n1173_));
NOR2X1 NOR2X1_604 ( .A(u5__abc_78290_new_n475_), .B(u5__abc_78290_new_n1176_), .Y(u5__abc_78290_new_n1177_));
NOR2X1 NOR2X1_605 ( .A(u5__abc_78290_new_n475_), .B(u5__abc_78290_new_n1179_), .Y(u5__abc_78290_new_n1180_));
NOR2X1 NOR2X1_606 ( .A(u5__abc_78290_new_n1175_), .B(u5__abc_78290_new_n1182_), .Y(u5__abc_78290_new_n1183_));
NOR2X1 NOR2X1_607 ( .A(u5__abc_78290_new_n1149_), .B(u5__abc_78290_new_n1184_), .Y(u5__abc_78290_new_n1185_));
NOR2X1 NOR2X1_608 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n408_), .Y(u5__abc_78290_new_n1188_));
NOR2X1 NOR2X1_609 ( .A(u5__abc_78290_new_n557_), .B(u5__abc_78290_new_n605_), .Y(u5__abc_78290_new_n1189_));
NOR2X1 NOR2X1_61 ( .A(u0__abc_74894_new_n4062_), .B(u0__abc_74894_new_n4066_), .Y(u0__abc_74894_new_n4067_));
NOR2X1 NOR2X1_610 ( .A(u5__abc_78290_new_n557_), .B(u5__abc_78290_new_n598_), .Y(u5__abc_78290_new_n1192_));
NOR2X1 NOR2X1_611 ( .A(u5__abc_78290_new_n501_), .B(u5__abc_78290_new_n581_), .Y(u5__abc_78290_new_n1194_));
NOR2X1 NOR2X1_612 ( .A(u5__abc_78290_new_n557_), .B(u5__abc_78290_new_n592_), .Y(u5__abc_78290_new_n1198_));
NOR2X1 NOR2X1_613 ( .A(u5__abc_78290_new_n1200_), .B(u5__abc_78290_new_n1197_), .Y(u5__abc_78290_new_n1201_));
NOR2X1 NOR2X1_614 ( .A(u5__abc_78290_new_n452_), .B(u5__abc_78290_new_n1202_), .Y(u5__abc_78290_new_n1203_));
NOR2X1 NOR2X1_615 ( .A(u5__abc_78290_new_n683_), .B(u5__abc_78290_new_n1205_), .Y(u5__abc_78290_new_n1206_));
NOR2X1 NOR2X1_616 ( .A(u5__abc_78290_new_n1191_), .B(u5__abc_78290_new_n1210_), .Y(u5__abc_78290_new_n1211_));
NOR2X1 NOR2X1_617 ( .A(u5__abc_78290_new_n436_), .B(u5__abc_78290_new_n1213_), .Y(u5__abc_78290_new_n1214_));
NOR2X1 NOR2X1_618 ( .A(u5__abc_78290_new_n474_), .B(u5__abc_78290_new_n1217_), .Y(u5__abc_78290_new_n1218_));
NOR2X1 NOR2X1_619 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n1220_), .Y(u5__abc_78290_new_n1221_));
NOR2X1 NOR2X1_62 ( .A(u0__abc_74894_new_n4074_), .B(u0__abc_74894_new_n4078_), .Y(u0__abc_74894_new_n4079_));
NOR2X1 NOR2X1_620 ( .A(u5__abc_78290_new_n1226_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n1227_));
NOR2X1 NOR2X1_621 ( .A(u5_state_14_), .B(u5__abc_78290_new_n763_), .Y(u5__abc_78290_new_n1230_));
NOR2X1 NOR2X1_622 ( .A(u5__abc_78290_new_n443_), .B(u5__abc_78290_new_n1231_), .Y(u5__abc_78290_new_n1232_));
NOR2X1 NOR2X1_623 ( .A(u5__abc_78290_new_n474_), .B(u5__abc_78290_new_n1236_), .Y(u5__abc_78290_new_n1237_));
NOR2X1 NOR2X1_624 ( .A(u5__abc_78290_new_n452_), .B(u5__abc_78290_new_n1241_), .Y(u5__abc_78290_new_n1242_));
NOR2X1 NOR2X1_625 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1243_), .Y(u5__abc_78290_new_n1244_));
NOR2X1 NOR2X1_626 ( .A(u5_state_34_), .B(u5__abc_78290_new_n513_), .Y(u5__abc_78290_new_n1245_));
NOR2X1 NOR2X1_627 ( .A(u5__abc_78290_new_n399_), .B(u5__abc_78290_new_n1246_), .Y(u5__abc_78290_new_n1247_));
NOR2X1 NOR2X1_628 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1248_), .Y(u5__abc_78290_new_n1249_));
NOR2X1 NOR2X1_629 ( .A(u5__abc_78290_new_n1216_), .B(u5__abc_78290_new_n1252_), .Y(u5__abc_78290_new_n1253_));
NOR2X1 NOR2X1_63 ( .A(u0__abc_74894_new_n4084_), .B(u0__abc_74894_new_n4086_), .Y(u0__abc_74894_new_n4087_));
NOR2X1 NOR2X1_630 ( .A(u5__abc_78290_new_n1254_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n1255_));
NOR2X1 NOR2X1_631 ( .A(u5__abc_78290_new_n1256_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1257_));
NOR2X1 NOR2X1_632 ( .A(u5_state_9_), .B(u5__abc_78290_new_n741_), .Y(u5__abc_78290_new_n1259_));
NOR2X1 NOR2X1_633 ( .A(u5__abc_78290_new_n1261_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1262_));
NOR2X1 NOR2X1_634 ( .A(u5__abc_78290_new_n1257_), .B(u5__abc_78290_new_n1262_), .Y(u5__abc_78290_new_n1263_));
NOR2X1 NOR2X1_635 ( .A(u5_state_8_), .B(u5__abc_78290_new_n726_), .Y(u5__abc_78290_new_n1264_));
NOR2X1 NOR2X1_636 ( .A(u5_state_15_), .B(u5__abc_78290_new_n829_), .Y(u5__abc_78290_new_n1269_));
NOR2X1 NOR2X1_637 ( .A(u5__abc_78290_new_n443_), .B(u5__abc_78290_new_n1270_), .Y(u5__abc_78290_new_n1271_));
NOR2X1 NOR2X1_638 ( .A(u5__abc_78290_new_n1272_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1273_));
NOR2X1 NOR2X1_639 ( .A(u5__abc_78290_new_n1273_), .B(u5__abc_78290_new_n1268_), .Y(u5__abc_78290_new_n1274_));
NOR2X1 NOR2X1_64 ( .A(u0__abc_74894_new_n4106_), .B(u0__abc_74894_new_n4108_), .Y(u0__abc_74894_new_n4109_));
NOR2X1 NOR2X1_640 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n408_), .Y(u5__abc_78290_new_n1278_));
NOR2X1 NOR2X1_641 ( .A(u5_state_11_), .B(u5__abc_78290_new_n757_), .Y(u5__abc_78290_new_n1279_));
NOR2X1 NOR2X1_642 ( .A(u5__abc_78290_new_n1280_), .B(u5__abc_78290_new_n1258_), .Y(u5__abc_78290_new_n1281_));
NOR2X1 NOR2X1_643 ( .A(u5_state_7_), .B(u5__abc_78290_new_n733_), .Y(u5__abc_78290_new_n1285_));
NOR2X1 NOR2X1_644 ( .A(u5_state_6_), .B(u5__abc_78290_new_n777_), .Y(u5__abc_78290_new_n1288_));
NOR2X1 NOR2X1_645 ( .A(u5__abc_78290_new_n1289_), .B(u5__abc_78290_new_n1284_), .Y(u5__abc_78290_new_n1290_));
NOR2X1 NOR2X1_646 ( .A(u5__abc_78290_new_n415_), .B(u5__abc_78290_new_n1295_), .Y(u5__abc_78290_new_n1296_));
NOR2X1 NOR2X1_647 ( .A(u5__abc_78290_new_n770_), .B(u5__abc_78290_new_n773_), .Y(u5__abc_78290_new_n1298_));
NOR2X1 NOR2X1_648 ( .A(u5__abc_78290_new_n1305_), .B(u5__abc_78290_new_n1303_), .Y(u5__abc_78290_new_n1306_));
NOR2X1 NOR2X1_649 ( .A(u5_state_1_), .B(u5__abc_78290_new_n787_), .Y(u5__abc_78290_new_n1308_));
NOR2X1 NOR2X1_65 ( .A(u0__abc_74894_new_n4129_), .B(u0__abc_74894_new_n4128_), .Y(u0__abc_74894_new_n4130_));
NOR2X1 NOR2X1_650 ( .A(u5__abc_78290_new_n1310_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1311_));
NOR2X1 NOR2X1_651 ( .A(u5__abc_78290_new_n574_), .B(u5__abc_78290_new_n1311_), .Y(u5__abc_78290_new_n1312_));
NOR2X1 NOR2X1_652 ( .A(u5__abc_78290_new_n1313_), .B(u5__abc_78290_new_n1294_), .Y(u5__abc_78290_new_n1314_));
NOR2X1 NOR2X1_653 ( .A(u5__abc_78290_new_n1212_), .B(u5__abc_78290_new_n1315_), .Y(u5__abc_78290_new_n1316_));
NOR2X1 NOR2X1_654 ( .A(csc_s_3_), .B(u5__abc_78290_new_n1320_), .Y(u5__abc_78290_new_n1321_));
NOR2X1 NOR2X1_655 ( .A(u5__abc_78290_new_n1319_), .B(u5__abc_78290_new_n1322_), .Y(u5__abc_78290_new_n1323_));
NOR2X1 NOR2X1_656 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1324_), .Y(u5__abc_78290_new_n1325_));
NOR2X1 NOR2X1_657 ( .A(obct_cs_2_), .B(obct_cs_3_), .Y(u5__abc_78290_new_n1327_));
NOR2X1 NOR2X1_658 ( .A(obct_cs_0_), .B(obct_cs_1_), .Y(u5__abc_78290_new_n1328_));
NOR2X1 NOR2X1_659 ( .A(obct_cs_6_), .B(obct_cs_7_), .Y(u5__abc_78290_new_n1330_));
NOR2X1 NOR2X1_66 ( .A(u0__abc_74894_new_n4140_), .B(u0__abc_74894_new_n4144_), .Y(u0__abc_74894_new_n4145_));
NOR2X1 NOR2X1_660 ( .A(obct_cs_4_), .B(obct_cs_5_), .Y(u5__abc_78290_new_n1331_));
NOR2X1 NOR2X1_661 ( .A(u5_wb_cycle), .B(u5__abc_78290_new_n1338_), .Y(u5__abc_78290_new_n1339_));
NOR2X1 NOR2X1_662 ( .A(init_req), .B(rfr_req), .Y(u5__abc_78290_new_n1343_));
NOR2X1 NOR2X1_663 ( .A(u5__abc_78290_new_n1335_), .B(u5__abc_78290_new_n1344_), .Y(u5__abc_78290_new_n1345_));
NOR2X1 NOR2X1_664 ( .A(u5__abc_78290_new_n1223_), .B(u5__abc_78290_new_n1353_), .Y(u5__abc_78290_new_n1354_));
NOR2X1 NOR2X1_665 ( .A(u5__abc_78290_new_n1127_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1358_));
NOR2X1 NOR2X1_666 ( .A(u5__abc_78290_new_n1246_), .B(u5__abc_78290_new_n670_), .Y(u5__abc_78290_new_n1362_));
NOR2X1 NOR2X1_667 ( .A(u5__abc_78290_new_n1365_), .B(u5__abc_78290_new_n1364_), .Y(u5__abc_78290_new_n1366_));
NOR2X1 NOR2X1_668 ( .A(u5__abc_78290_new_n1043_), .B(u5__abc_78290_new_n1369_), .Y(u5__abc_78290_new_n1370_));
NOR2X1 NOR2X1_669 ( .A(u5__abc_78290_new_n1355_), .B(u5__abc_78290_new_n1372_), .Y(u5__abc_78290_new_n1373_));
NOR2X1 NOR2X1_67 ( .A(u0__abc_74894_new_n4151_), .B(u0__abc_74894_new_n4155_), .Y(u0__abc_74894_new_n4156_));
NOR2X1 NOR2X1_670 ( .A(u5_kro), .B(u5__abc_78290_new_n1375_), .Y(u5__abc_78290_new_n1376_));
NOR2X1 NOR2X1_671 ( .A(u5__abc_78290_new_n1376_), .B(u5__abc_78290_new_n1374_), .Y(u5__abc_78290_new_n1377_));
NOR2X1 NOR2X1_672 ( .A(u5__abc_78290_new_n1268_), .B(u5__abc_78290_new_n1377_), .Y(u5__abc_78290_new_n1378_));
NOR2X1 NOR2X1_673 ( .A(u5__abc_78290_new_n1171_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1380_));
NOR2X1 NOR2X1_674 ( .A(u5__abc_78290_new_n1178_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1381_));
NOR2X1 NOR2X1_675 ( .A(u5__abc_78290_new_n1380_), .B(u5__abc_78290_new_n1381_), .Y(u5__abc_78290_new_n1382_));
NOR2X1 NOR2X1_676 ( .A(u5__abc_78290_new_n1152_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1383_));
NOR2X1 NOR2X1_677 ( .A(u5__abc_78290_new_n1161_), .B(u5__abc_78290_new_n1383_), .Y(u5__abc_78290_new_n1384_));
NOR2X1 NOR2X1_678 ( .A(u5__abc_78290_new_n1385_), .B(u5__abc_78290_new_n1389_), .Y(u5__abc_78290_new_n1390_));
NOR2X1 NOR2X1_679 ( .A(u5__abc_78290_new_n1181_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1394_));
NOR2X1 NOR2X1_68 ( .A(u0__abc_74894_new_n4163_), .B(u0__abc_74894_new_n4159_), .Y(u0__abc_74894_new_n4164_));
NOR2X1 NOR2X1_680 ( .A(u5__abc_78290_new_n1391_), .B(u5__abc_78290_new_n1396_), .Y(u5__abc_78290_new_n1397_));
NOR2X1 NOR2X1_681 ( .A(tms_s_0_), .B(tms_s_2_), .Y(u5__abc_78290_new_n1404_));
NOR2X1 NOR2X1_682 ( .A(tms_s_1_), .B(u5__abc_78290_new_n1405_), .Y(u5__abc_78290_new_n1406_));
NOR2X1 NOR2X1_683 ( .A(u5_wb_write_go_r), .B(u5__abc_78290_new_n1412_), .Y(u5__abc_78290_new_n1413_));
NOR2X1 NOR2X1_684 ( .A(u5__abc_78290_new_n1375_), .B(u5__abc_78290_new_n877_), .Y(u5__abc_78290_new_n1422_));
NOR2X1 NOR2X1_685 ( .A(u5__abc_78290_new_n1422_), .B(u5__abc_78290_new_n1423_), .Y(u5__abc_78290_new_n1424_));
NOR2X1 NOR2X1_686 ( .A(u5__abc_78290_new_n1398_), .B(u5__abc_78290_new_n1425_), .Y(u5__abc_78290_new_n1426_));
NOR2X1 NOR2X1_687 ( .A(u5__abc_78290_new_n1433_), .B(u5__abc_78290_new_n1398_), .Y(u5__abc_78290_new_n1434_));
NOR2X1 NOR2X1_688 ( .A(u5__abc_78290_new_n1439_), .B(u5__abc_78290_new_n1438_), .Y(u5__abc_78290_new_n1440_));
NOR2X1 NOR2X1_689 ( .A(u5__abc_78290_new_n1443_), .B(u5__abc_78290_new_n1442_), .Y(u5__abc_78290_new_n1444_));
NOR2X1 NOR2X1_69 ( .A(u0__abc_74894_new_n4171_), .B(u0__abc_74894_new_n4169_), .Y(u0__abc_74894_new_n4172_));
NOR2X1 NOR2X1_690 ( .A(u5__abc_78290_new_n1447_), .B(u5__abc_78290_new_n1403_), .Y(u5__abc_78290_new_n1448_));
NOR2X1 NOR2X1_691 ( .A(u5__abc_78290_new_n1287_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1456_));
NOR2X1 NOR2X1_692 ( .A(u5__abc_78290_new_n1454_), .B(u5__abc_78290_new_n1461_), .Y(u5__abc_78290_new_n1462_));
NOR2X1 NOR2X1_693 ( .A(rfr_ack), .B(susp_sel), .Y(u5__abc_78290_new_n1469_));
NOR2X1 NOR2X1_694 ( .A(tms_s_16_), .B(tms_s_17_), .Y(u5__abc_78290_new_n1474_));
NOR2X1 NOR2X1_695 ( .A(u5__abc_78290_new_n1475_), .B(u5__abc_78290_new_n1472_), .Y(u5__abc_78290_new_n1476_));
NOR2X1 NOR2X1_696 ( .A(u5__abc_78290_new_n1400_), .B(u5__abc_78290_new_n1476_), .Y(u5__abc_78290_new_n1477_));
NOR2X1 NOR2X1_697 ( .A(csc_s_3_), .B(u5__abc_78290_new_n1480_), .Y(u5__abc_78290_new_n1481_));
NOR2X1 NOR2X1_698 ( .A(u1_wb_write_go), .B(u5_wb_wait), .Y(u5__abc_78290_new_n1482_));
NOR2X1 NOR2X1_699 ( .A(u5__abc_78290_new_n1483_), .B(u5__abc_78290_new_n1479_), .Y(u5__abc_78290_new_n1484_));
NOR2X1 NOR2X1_7 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n3474_));
NOR2X1 NOR2X1_70 ( .A(u0__abc_74894_new_n4182_), .B(u0__abc_74894_new_n4186_), .Y(u0__abc_74894_new_n4187_));
NOR2X1 NOR2X1_700 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1486_), .Y(u5__abc_78290_new_n1487_));
NOR2X1 NOR2X1_701 ( .A(u5__abc_78290_new_n1423_), .B(u5__abc_78290_new_n1498_), .Y(u5__abc_78290_new_n1499_));
NOR2X1 NOR2X1_702 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n877_), .Y(u5__abc_78290_new_n1502_));
NOR2X1 NOR2X1_703 ( .A(u5__abc_78290_new_n1504_), .B(u5__abc_78290_new_n1505_), .Y(u5__abc_78290_new_n1506_));
NOR2X1 NOR2X1_704 ( .A(u5__abc_78290_new_n1507_), .B(u5__abc_78290_new_n1477_), .Y(u5__abc_78290_new_n1508_));
NOR2X1 NOR2X1_705 ( .A(u5__abc_78290_new_n1514_), .B(u5__abc_78290_new_n1512_), .Y(u5__abc_78290_new_n1515_));
NOR2X1 NOR2X1_706 ( .A(u5__abc_78290_new_n1433_), .B(u5__abc_78290_new_n1459_), .Y(u5__abc_78290_new_n1516_));
NOR2X1 NOR2X1_707 ( .A(csc_s_4_), .B(csc_s_5_), .Y(u5__abc_78290_new_n1526_));
NOR2X1 NOR2X1_708 ( .A(u5__abc_78290_new_n669_), .B(u5__abc_78290_new_n1529_), .Y(u5__abc_78290_new_n1530_));
NOR2X1 NOR2X1_709 ( .A(u5__abc_78290_new_n1534_), .B(u5__abc_78290_new_n1537_), .Y(u5__abc_78290_new_n1538_));
NOR2X1 NOR2X1_71 ( .A(u0__abc_74894_new_n4193_), .B(u0__abc_74894_new_n4197_), .Y(u0__abc_74894_new_n4198_));
NOR2X1 NOR2X1_710 ( .A(u5_state_0_), .B(u5__abc_78290_new_n793_), .Y(u5__abc_78290_new_n1539_));
NOR2X1 NOR2X1_711 ( .A(u5__abc_78290_new_n1545_), .B(u5__abc_78290_new_n1546_), .Y(u5__abc_78290_new_n1547_));
NOR2X1 NOR2X1_712 ( .A(u5__abc_78290_new_n1542_), .B(u5__abc_78290_new_n1548_), .Y(u5__abc_78290_new_n1549_));
NOR2X1 NOR2X1_713 ( .A(u5__abc_78290_new_n1273_), .B(u5__abc_78290_new_n1551_), .Y(u5__abc_78290_new_n1552_));
NOR2X1 NOR2X1_714 ( .A(u5__abc_78290_new_n1299_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1554_));
NOR2X1 NOR2X1_715 ( .A(u5__abc_78290_new_n1554_), .B(u5__abc_78290_new_n1456_), .Y(u5__abc_78290_new_n1555_));
NOR2X1 NOR2X1_716 ( .A(u5__abc_78290_new_n1238_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n1557_));
NOR2X1 NOR2X1_717 ( .A(u5__abc_78290_new_n1311_), .B(u5__abc_78290_new_n1557_), .Y(u5__abc_78290_new_n1558_));
NOR2X1 NOR2X1_718 ( .A(u5__abc_78290_new_n1560_), .B(u5__abc_78290_new_n1559_), .Y(u5__abc_78290_new_n1561_));
NOR2X1 NOR2X1_719 ( .A(u5__abc_78290_new_n1353_), .B(u5__abc_78290_new_n1562_), .Y(u5__abc_78290_new_n1563_));
NOR2X1 NOR2X1_72 ( .A(u0__abc_74894_new_n4205_), .B(u0__abc_74894_new_n4201_), .Y(u0__abc_74894_new_n4206_));
NOR2X1 NOR2X1_720 ( .A(u5__abc_78290_new_n1556_), .B(u5__abc_78290_new_n1564_), .Y(u5__abc_78290_new_n1565_));
NOR2X1 NOR2X1_721 ( .A(u5__abc_78290_new_n1532_), .B(u5__abc_78290_new_n1566_), .Y(u5__abc_78290_new_n1567_));
NOR2X1 NOR2X1_722 ( .A(u5__abc_78290_new_n1531_), .B(u5__abc_78290_new_n1568_), .Y(u5_pack_le2_d));
NOR2X1 NOR2X1_723 ( .A(u5__abc_78290_new_n1292_), .B(u5__abc_78290_new_n1300_), .Y(u5__abc_78290_new_n1570_));
NOR2X1 NOR2X1_724 ( .A(u5__abc_78290_new_n1572_), .B(u5__abc_78290_new_n1571_), .Y(u5__abc_78290_new_n1573_));
NOR2X1 NOR2X1_725 ( .A(u5_cnt), .B(u5__abc_78290_new_n1574_), .Y(u5__abc_78290_new_n1575_));
NOR2X1 NOR2X1_726 ( .A(u5__abc_78290_new_n1536_), .B(u5__abc_78290_new_n1548_), .Y(u5__abc_78290_new_n1578_));
NOR2X1 NOR2X1_727 ( .A(u5__abc_78290_new_n1580_), .B(u5__abc_78290_new_n1583_), .Y(u5__abc_78290_new_n1584_));
NOR2X1 NOR2X1_728 ( .A(u5__abc_78290_new_n1576_), .B(u5__abc_78290_new_n1585_), .Y(u5_cnt_next));
NOR2X1 NOR2X1_729 ( .A(u5__abc_78290_new_n1587_), .B(u5__abc_78290_new_n1008_), .Y(u5__abc_78290_new_n1588_));
NOR2X1 NOR2X1_73 ( .A(u0__abc_74894_new_n4209_), .B(u0__abc_74894_new_n4213_), .Y(u0__abc_74894_new_n4214_));
NOR2X1 NOR2X1_730 ( .A(u5__abc_78290_new_n731_), .B(u5__abc_78290_new_n1589_), .Y(u5__abc_78290_new_n1590_));
NOR2X1 NOR2X1_731 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n1591_), .Y(bank_set));
NOR2X1 NOR2X1_732 ( .A(u5_ack_cnt_1_), .B(u5_ack_cnt_0_), .Y(u5__abc_78290_new_n1593_));
NOR2X1 NOR2X1_733 ( .A(u5_ack_cnt_2_), .B(u5__abc_78290_new_n1594_), .Y(u5__abc_78290_new_n1595_));
NOR2X1 NOR2X1_734 ( .A(u5_ack_cnt_3_), .B(u5__abc_78290_new_n1596_), .Y(u5__abc_78290_new_n1597_));
NOR2X1 NOR2X1_735 ( .A(u5_wb_wait), .B(u5_mem_ack_r), .Y(u5__abc_78290_new_n1601_));
NOR2X1 NOR2X1_736 ( .A(u5__abc_78290_new_n1600_), .B(u5__abc_78290_new_n1602_), .Y(u5__abc_78290_new_n1603_));
NOR2X1 NOR2X1_737 ( .A(u5__abc_78290_new_n1606_), .B(u5__abc_78290_new_n1479_), .Y(u5__abc_78290_new_n1607_));
NOR2X1 NOR2X1_738 ( .A(u5__abc_78290_new_n1324_), .B(u5__abc_78290_new_n1602_), .Y(u5__abc_78290_new_n1610_));
NOR2X1 NOR2X1_739 ( .A(u5__abc_78290_new_n486_), .B(u5__abc_78290_new_n1612_), .Y(u5__abc_78290_new_n1613_));
NOR2X1 NOR2X1_74 ( .A(u0__abc_74894_new_n4221_), .B(u0__abc_74894_new_n4225_), .Y(u0__abc_74894_new_n4226_));
NOR2X1 NOR2X1_740 ( .A(u5_mem_ack_r), .B(u5__abc_78290_new_n1620_), .Y(u5__abc_78290_new_n1621_));
NOR2X1 NOR2X1_741 ( .A(u5__abc_78290_new_n1618_), .B(u5__abc_78290_new_n1623_), .Y(u5__abc_78290_new_n1624_));
NOR2X1 NOR2X1_742 ( .A(u5__abc_78290_new_n1607_), .B(u5__abc_78290_new_n1626_), .Y(u5__abc_78290_new_n1627_));
NOR2X1 NOR2X1_743 ( .A(u5__abc_78290_new_n1629_), .B(mem_ack), .Y(u5__0wb_stb_first_0_0_));
NOR2X1 NOR2X1_744 ( .A(u5_kro), .B(u5__abc_78290_new_n1019_), .Y(u5__abc_78290_new_n1633_));
NOR2X1 NOR2X1_745 ( .A(u5__abc_78290_new_n1636_), .B(u5__abc_78290_new_n1401_), .Y(u5__abc_78290_new_n1637_));
NOR2X1 NOR2X1_746 ( .A(u5__abc_78290_new_n1640_), .B(u5__abc_78290_new_n1638_), .Y(u5__abc_78290_new_n1641_));
NOR2X1 NOR2X1_747 ( .A(u5__abc_78290_new_n1351_), .B(u5__abc_78290_new_n1644_), .Y(u5__abc_78290_new_n1645_));
NOR2X1 NOR2X1_748 ( .A(u5__abc_78290_new_n1646_), .B(u5__abc_78290_new_n1642_), .Y(u5__abc_78290_new_n1647_));
NOR2X1 NOR2X1_749 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n1653_), .Y(u5__abc_78290_new_n1654_));
NOR2X1 NOR2X1_75 ( .A(u0__abc_74894_new_n4235_), .B(u0__abc_74894_new_n4231_), .Y(u0__abc_74894_new_n4236_));
NOR2X1 NOR2X1_750 ( .A(u5_burst_cnt_0_), .B(u5__abc_78290_new_n1666_), .Y(u5__abc_78290_new_n1667_));
NOR2X1 NOR2X1_751 ( .A(u5_burst_cnt_5_), .B(u5__abc_78290_new_n1694_), .Y(u5__abc_78290_new_n1699_));
NOR2X1 NOR2X1_752 ( .A(u5__abc_78290_new_n474_), .B(u5__abc_78290_new_n1713_), .Y(u5__abc_78290_new_n1714_));
NOR2X1 NOR2X1_753 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n1715_), .Y(u5__abc_78290_new_n1716_));
NOR2X1 NOR2X1_754 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1719_), .Y(u5__abc_78290_new_n1720_));
NOR2X1 NOR2X1_755 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1721_), .Y(u5__abc_78290_new_n1722_));
NOR2X1 NOR2X1_756 ( .A(u5__abc_78290_new_n1718_), .B(u5__abc_78290_new_n1724_), .Y(u5__abc_78290_new_n1725_));
NOR2X1 NOR2X1_757 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n1726_), .Y(u5__abc_78290_new_n1727_));
NOR2X1 NOR2X1_758 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1730_), .Y(u5__abc_78290_new_n1731_));
NOR2X1 NOR2X1_759 ( .A(u5__abc_78290_new_n452_), .B(u5__abc_78290_new_n1733_), .Y(u5__abc_78290_new_n1734_));
NOR2X1 NOR2X1_76 ( .A(u0__abc_74894_new_n4261_), .B(u0__abc_74894_new_n4257_), .Y(u0__abc_74894_new_n4262_));
NOR2X1 NOR2X1_760 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n1739_), .Y(u5__abc_78290_new_n1740_));
NOR2X1 NOR2X1_761 ( .A(u5__abc_78290_new_n426_), .B(u5__abc_78290_new_n1744_), .Y(u5__abc_78290_new_n1745_));
NOR2X1 NOR2X1_762 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1746_), .Y(u5__abc_78290_new_n1747_));
NOR2X1 NOR2X1_763 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n1749_), .Y(u5__abc_78290_new_n1750_));
NOR2X1 NOR2X1_764 ( .A(u5__abc_78290_new_n449_), .B(u5__abc_78290_new_n559_), .Y(u5__abc_78290_new_n1754_));
NOR2X1 NOR2X1_765 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1755_), .Y(u5__abc_78290_new_n1756_));
NOR2X1 NOR2X1_766 ( .A(u5__abc_78290_new_n449_), .B(u5__abc_78290_new_n576_), .Y(u5__abc_78290_new_n1757_));
NOR2X1 NOR2X1_767 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1758_), .Y(u5__abc_78290_new_n1759_));
NOR2X1 NOR2X1_768 ( .A(u5__abc_78290_new_n1761_), .B(u5__abc_78290_new_n1743_), .Y(u5__abc_78290_new_n1762_));
NOR2X1 NOR2X1_769 ( .A(u5__abc_78290_new_n436_), .B(u5__abc_78290_new_n482_), .Y(u5__abc_78290_new_n1763_));
NOR2X1 NOR2X1_77 ( .A(u0__abc_74894_new_n4287_), .B(u0__abc_74894_new_n4283_), .Y(u0__abc_74894_new_n4288_));
NOR2X1 NOR2X1_770 ( .A(u5__abc_78290_new_n426_), .B(u5__abc_78290_new_n1772_), .Y(u5__abc_78290_new_n1773_));
NOR2X1 NOR2X1_771 ( .A(u5__abc_78290_new_n443_), .B(u5__abc_78290_new_n1777_), .Y(u5__abc_78290_new_n1778_));
NOR2X1 NOR2X1_772 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1779_), .Y(u5__abc_78290_new_n1780_));
NOR2X1 NOR2X1_773 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1783_), .Y(u5__abc_78290_new_n1784_));
NOR2X1 NOR2X1_774 ( .A(u5__abc_78290_new_n449_), .B(u5__abc_78290_new_n572_), .Y(u5__abc_78290_new_n1788_));
NOR2X1 NOR2X1_775 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1789_), .Y(u5__abc_78290_new_n1790_));
NOR2X1 NOR2X1_776 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1792_), .Y(u5__abc_78290_new_n1793_));
NOR2X1 NOR2X1_777 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1798_), .Y(u5__abc_78290_new_n1799_));
NOR2X1 NOR2X1_778 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1804_), .Y(u5__abc_78290_new_n1805_));
NOR2X1 NOR2X1_779 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1808_), .Y(u5__abc_78290_new_n1809_));
NOR2X1 NOR2X1_78 ( .A(u0__abc_74894_new_n4313_), .B(u0__abc_74894_new_n4309_), .Y(u0__abc_74894_new_n4314_));
NOR2X1 NOR2X1_780 ( .A(u5__abc_78290_new_n443_), .B(u5__abc_78290_new_n1813_), .Y(u5__abc_78290_new_n1814_));
NOR2X1 NOR2X1_781 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1815_), .Y(u5__abc_78290_new_n1816_));
NOR2X1 NOR2X1_782 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1818_), .Y(u5__abc_78290_new_n1819_));
NOR2X1 NOR2X1_783 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1826_), .Y(u5__abc_78290_new_n1827_));
NOR2X1 NOR2X1_784 ( .A(u5__abc_78290_new_n1796_), .B(u5__abc_78290_new_n1831_), .Y(u5__abc_78290_new_n1832_));
NOR2X1 NOR2X1_785 ( .A(u5__abc_78290_new_n459_), .B(u5__abc_78290_new_n1834_), .Y(u5__abc_78290_new_n1835_));
NOR2X1 NOR2X1_786 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n1836_), .Y(u5__abc_78290_new_n1837_));
NOR2X1 NOR2X1_787 ( .A(u5__abc_78290_new_n459_), .B(u5__abc_78290_new_n1839_), .Y(u5__abc_78290_new_n1840_));
NOR2X1 NOR2X1_788 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1841_), .Y(u5__abc_78290_new_n1842_));
NOR2X1 NOR2X1_789 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n1845_), .Y(u5__abc_78290_new_n1846_));
NOR2X1 NOR2X1_79 ( .A(u0__abc_74894_new_n4340_), .B(u0__abc_74894_new_n4336_), .Y(u0__abc_74894_new_n4341_));
NOR2X1 NOR2X1_790 ( .A(u5__abc_78290_new_n459_), .B(u5__abc_78290_new_n1848_), .Y(u5__abc_78290_new_n1849_));
NOR2X1 NOR2X1_791 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1850_), .Y(u5__abc_78290_new_n1851_));
NOR2X1 NOR2X1_792 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n1854_), .Y(u5__abc_78290_new_n1855_));
NOR2X1 NOR2X1_793 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1857_), .Y(u5__abc_78290_new_n1858_));
NOR2X1 NOR2X1_794 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n1863_), .Y(u5__abc_78290_new_n1864_));
NOR2X1 NOR2X1_795 ( .A(u5__abc_78290_new_n1853_), .B(u5__abc_78290_new_n1866_), .Y(u5__abc_78290_new_n1867_));
NOR2X1 NOR2X1_796 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1871_), .Y(u5__abc_78290_new_n1872_));
NOR2X1 NOR2X1_797 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n1873_), .Y(u5__abc_78290_new_n1874_));
NOR2X1 NOR2X1_798 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1882_), .Y(u5__abc_78290_new_n1883_));
NOR2X1 NOR2X1_799 ( .A(u5__abc_78290_new_n462_), .B(u5__abc_78290_new_n1884_), .Y(u5__abc_78290_new_n1885_));
NOR2X1 NOR2X1_8 ( .A(cs_le), .B(cs_0_), .Y(u0__abc_74894_new_n3479_));
NOR2X1 NOR2X1_80 ( .A(u0__abc_74894_new_n4362_), .B(u0__abc_74894_new_n4365_), .Y(u0__abc_74894_new_n4366_));
NOR2X1 NOR2X1_800 ( .A(u5__abc_78290_new_n1888_), .B(u5__abc_78290_new_n1877_), .Y(u5__abc_78290_new_n1889_));
NOR2X1 NOR2X1_801 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1042_), .Y(u5__abc_78290_new_n1891_));
NOR2X1 NOR2X1_802 ( .A(u5__abc_78290_new_n457_), .B(u5__abc_78290_new_n1892_), .Y(u5__abc_78290_new_n1893_));
NOR2X1 NOR2X1_803 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1894_), .Y(u5__abc_78290_new_n1895_));
NOR2X1 NOR2X1_804 ( .A(u5__abc_78290_new_n457_), .B(u5__abc_78290_new_n1897_), .Y(u5__abc_78290_new_n1898_));
NOR2X1 NOR2X1_805 ( .A(u5__abc_78290_new_n457_), .B(u5__abc_78290_new_n1900_), .Y(u5__abc_78290_new_n1901_));
NOR2X1 NOR2X1_806 ( .A(u5__abc_78290_new_n445_), .B(u5__abc_78290_new_n1905_), .Y(u5__abc_78290_new_n1906_));
NOR2X1 NOR2X1_807 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1907_), .Y(u5__abc_78290_new_n1908_));
NOR2X1 NOR2X1_808 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n1910_), .Y(u5__abc_78290_new_n1911_));
NOR2X1 NOR2X1_809 ( .A(u5__abc_78290_new_n460_), .B(u5__abc_78290_new_n1916_), .Y(u5__abc_78290_new_n1917_));
NOR2X1 NOR2X1_81 ( .A(u0__abc_74894_new_n1737_), .B(u0__abc_74894_new_n3716_), .Y(u0__abc_74894_new_n4372_));
NOR2X1 NOR2X1_810 ( .A(u5__abc_78290_new_n460_), .B(u5__abc_78290_new_n1919_), .Y(u5__abc_78290_new_n1920_));
NOR2X1 NOR2X1_811 ( .A(u5__abc_78290_new_n456_), .B(u5__abc_78290_new_n1097_), .Y(u5__abc_78290_new_n1924_));
NOR2X1 NOR2X1_812 ( .A(u5__abc_78290_new_n456_), .B(u5__abc_78290_new_n1934_), .Y(u5__abc_78290_new_n1935_));
NOR2X1 NOR2X1_813 ( .A(u5__abc_78290_new_n460_), .B(u5__abc_78290_new_n1939_), .Y(u5__abc_78290_new_n1940_));
NOR2X1 NOR2X1_814 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1941_), .Y(u5__abc_78290_new_n1942_));
NOR2X1 NOR2X1_815 ( .A(u5__abc_78290_new_n477_), .B(u5__abc_78290_new_n1944_), .Y(u5__abc_78290_new_n1945_));
NOR2X1 NOR2X1_816 ( .A(u5__abc_78290_new_n1948_), .B(u5__abc_78290_new_n1915_), .Y(u5__abc_78290_new_n1949_));
NOR2X1 NOR2X1_817 ( .A(u5__abc_78290_new_n1833_), .B(u5__abc_78290_new_n1950_), .Y(u5__abc_78290_new_n1951_));
NOR2X1 NOR2X1_818 ( .A(u5__abc_78290_new_n372_), .B(u5__abc_78290_new_n1959_), .Y(u5__abc_78290_new_n1962_));
NOR2X1 NOR2X1_819 ( .A(u5__abc_78290_new_n372_), .B(u5__abc_78290_new_n1967_), .Y(u5__abc_78290_new_n1968_));
NOR2X1 NOR2X1_82 ( .A(u0__abc_74894_new_n4386_), .B(u0__abc_74894_new_n4389_), .Y(u0__abc_74894_new_n4390_));
NOR2X1 NOR2X1_820 ( .A(u5__abc_78290_new_n1541_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n1983_));
NOR2X1 NOR2X1_821 ( .A(u5__abc_78290_new_n1983_), .B(u5__abc_78290_new_n1311_), .Y(u5__abc_78290_new_n1984_));
NOR2X1 NOR2X1_822 ( .A(u5__abc_78290_new_n574_), .B(u5__abc_78290_new_n1305_), .Y(u5__abc_78290_new_n1985_));
NOR2X1 NOR2X1_823 ( .A(u5__abc_78290_new_n1982_), .B(u5__abc_78290_new_n1987_), .Y(u5__abc_78290_new_n1988_));
NOR2X1 NOR2X1_824 ( .A(u5__abc_78290_new_n1990_), .B(u5__abc_78290_new_n1991_), .Y(u5__abc_78290_new_n1992_));
NOR2X1 NOR2X1_825 ( .A(u5__abc_78290_new_n1993_), .B(u5__abc_78290_new_n1989_), .Y(u5__abc_78290_new_n1994_));
NOR2X1 NOR2X1_826 ( .A(u5__abc_78290_new_n2000_), .B(u5__abc_78290_new_n1995_), .Y(u5__abc_78290_new_n2001_));
NOR2X1 NOR2X1_827 ( .A(u5__abc_78290_new_n1532_), .B(u5__abc_78290_new_n1014_), .Y(u5__abc_78290_new_n2007_));
NOR2X1 NOR2X1_828 ( .A(u5__abc_78290_new_n2008_), .B(u5__abc_78290_new_n2000_), .Y(u5__abc_78290_new_n2009_));
NOR2X1 NOR2X1_829 ( .A(u5_ir_cnt_2_), .B(u5__abc_78290_new_n2015_), .Y(u5__abc_78290_new_n2017_));
NOR2X1 NOR2X1_83 ( .A(u0__abc_74894_new_n1757_), .B(u0__abc_74894_new_n3716_), .Y(u0__abc_74894_new_n4396_));
NOR2X1 NOR2X1_830 ( .A(u5__abc_78290_new_n1303_), .B(u5__abc_78290_new_n1216_), .Y(u5__abc_78290_new_n2024_));
NOR2X1 NOR2X1_831 ( .A(u5__abc_78290_new_n2027_), .B(u5__abc_78290_new_n2030_), .Y(u5__abc_78290_new_n2031_));
NOR2X1 NOR2X1_832 ( .A(u5_wb_wait_r), .B(u5__abc_78290_new_n1008_), .Y(u5__abc_78290_new_n2035_));
NOR2X1 NOR2X1_833 ( .A(u5__abc_78290_new_n1991_), .B(u5__abc_78290_new_n739_), .Y(u5__abc_78290_new_n2036_));
NOR2X1 NOR2X1_834 ( .A(u5__abc_78290_new_n2037_), .B(u5__abc_78290_new_n1564_), .Y(u5__abc_78290_new_n2038_));
NOR2X1 NOR2X1_835 ( .A(tms_s_4_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2041_));
NOR2X1 NOR2X1_836 ( .A(u5__abc_78290_new_n2042_), .B(u5__abc_78290_new_n1571_), .Y(u5__abc_78290_new_n2043_));
NOR2X1 NOR2X1_837 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n2044_), .Y(u5__abc_78290_new_n2045_));
NOR2X1 NOR2X1_838 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n804_), .Y(u5__abc_78290_new_n2052_));
NOR2X1 NOR2X1_839 ( .A(u5__abc_78290_new_n2048_), .B(u5__abc_78290_new_n2055_), .Y(u5__abc_78290_new_n2056_));
NOR2X1 NOR2X1_84 ( .A(u0__abc_74894_new_n4410_), .B(u0__abc_74894_new_n4413_), .Y(u0__abc_74894_new_n4414_));
NOR2X1 NOR2X1_840 ( .A(u5__abc_78290_new_n2057_), .B(u5__abc_78290_new_n2059_), .Y(u5__abc_78290_new_n2060_));
NOR2X1 NOR2X1_841 ( .A(u5__abc_78290_new_n2065_), .B(u5__abc_78290_new_n2064_), .Y(u5__abc_78290_new_n2066_));
NOR2X1 NOR2X1_842 ( .A(u5__abc_78290_new_n731_), .B(u5__abc_78290_new_n2069_), .Y(u5__abc_78290_new_n2070_));
NOR2X1 NOR2X1_843 ( .A(u5__abc_78290_new_n1991_), .B(u5__abc_78290_new_n2071_), .Y(u5__abc_78290_new_n2072_));
NOR2X1 NOR2X1_844 ( .A(u5__abc_78290_new_n2073_), .B(u5__abc_78290_new_n2067_), .Y(u5__abc_78290_new_n2074_));
NOR2X1 NOR2X1_845 ( .A(u5__abc_78290_new_n2077_), .B(u5__abc_78290_new_n1537_), .Y(u5__abc_78290_new_n2078_));
NOR2X1 NOR2X1_846 ( .A(u5__abc_78290_new_n1223_), .B(u5__abc_78290_new_n1234_), .Y(u5__abc_78290_new_n2079_));
NOR2X1 NOR2X1_847 ( .A(u5__abc_78290_new_n1999_), .B(u5__abc_78290_new_n2080_), .Y(u5__abc_78290_new_n2081_));
NOR2X1 NOR2X1_848 ( .A(u5__abc_78290_new_n2093_), .B(u5__abc_78290_new_n2092_), .Y(u5__abc_78290_new_n2094_));
NOR2X1 NOR2X1_849 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n2099_), .Y(u5__abc_78290_new_n2100_));
NOR2X1 NOR2X1_85 ( .A(\wb_addr_i[31] ), .B(u0__abc_74894_new_n4431_), .Y(u0__abc_74894_new_n4432_));
NOR2X1 NOR2X1_850 ( .A(u5__abc_78290_new_n1761_), .B(u5__abc_78290_new_n2104_), .Y(u5__abc_78290_new_n2105_));
NOR2X1 NOR2X1_851 ( .A(u5__abc_78290_new_n2108_), .B(u5__abc_78290_new_n1743_), .Y(u5__abc_78290_new_n2109_));
NOR2X1 NOR2X1_852 ( .A(u5__abc_78290_new_n2112_), .B(u5__abc_78290_new_n2114_), .Y(u5__abc_78290_new_n2115_));
NOR2X1 NOR2X1_853 ( .A(u5__abc_78290_new_n2103_), .B(u5__abc_78290_new_n2120_), .Y(u5__abc_78290_new_n2121_));
NOR2X1 NOR2X1_854 ( .A(u5__abc_78290_new_n1950_), .B(u5__abc_78290_new_n2123_), .Y(u5__abc_78290_new_n2124_));
NOR2X1 NOR2X1_855 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n2039_), .Y(u5__abc_78290_new_n2130_));
NOR2X1 NOR2X1_856 ( .A(tms_s_20_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2133_));
NOR2X1 NOR2X1_857 ( .A(u5__abc_78290_new_n1008_), .B(u5__abc_78290_new_n2136_), .Y(u5__abc_78290_new_n2137_));
NOR2X1 NOR2X1_858 ( .A(tms_s_15_), .B(u5__abc_78290_new_n2134_), .Y(u5__abc_78290_new_n2144_));
NOR2X1 NOR2X1_859 ( .A(tms_s_15_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2145_));
NOR2X1 NOR2X1_86 ( .A(u0_rf_we), .B(u0__abc_74894_new_n4433_), .Y(u0__0rf_we_0_0_));
NOR2X1 NOR2X1_860 ( .A(u5__abc_78290_new_n2147_), .B(u5__abc_78290_new_n2149_), .Y(u5__abc_78290_new_n2150_));
NOR2X1 NOR2X1_861 ( .A(u5__abc_78290_new_n2161_), .B(u5__abc_78290_new_n2159_), .Y(u5__abc_78290_new_n2162_));
NOR2X1 NOR2X1_862 ( .A(u5__abc_78290_new_n2163_), .B(u5__abc_78290_new_n2151_), .Y(u5__abc_78290_new_n2164_));
NOR2X1 NOR2X1_863 ( .A(u5__abc_78290_new_n1580_), .B(u5__abc_78290_new_n2174_), .Y(u5__abc_78290_new_n2175_));
NOR2X1 NOR2X1_864 ( .A(u5__abc_78290_new_n2176_), .B(u5__abc_78290_new_n2177_), .Y(u5__abc_78290_new_n2178_));
NOR2X1 NOR2X1_865 ( .A(u5__abc_78290_new_n1071_), .B(u5__abc_78290_new_n2180_), .Y(u5__abc_78290_new_n2181_));
NOR2X1 NOR2X1_866 ( .A(u5__abc_78290_new_n2183_), .B(u5__abc_78290_new_n2182_), .Y(u5__abc_78290_new_n2184_));
NOR2X1 NOR2X1_867 ( .A(u5__abc_78290_new_n2185_), .B(u5__abc_78290_new_n2179_), .Y(u5__abc_78290_new_n2186_));
NOR2X1 NOR2X1_868 ( .A(u5__abc_78290_new_n1042_), .B(u5__abc_78290_new_n1038_), .Y(u5__abc_78290_new_n2190_));
NOR2X1 NOR2X1_869 ( .A(u5__abc_78290_new_n1300_), .B(u5__abc_78290_new_n1132_), .Y(u5__abc_78290_new_n2191_));
NOR2X1 NOR2X1_87 ( .A(u0__abc_74894_new_n4438_), .B(u0__abc_74894_new_n4437_), .Y(cs_need_rfr_0_));
NOR2X1 NOR2X1_870 ( .A(u5__abc_78290_new_n1124_), .B(u5__abc_78290_new_n1175_), .Y(u5__abc_78290_new_n2193_));
NOR2X1 NOR2X1_871 ( .A(u5__abc_78290_new_n1114_), .B(u5__abc_78290_new_n2197_), .Y(u5__abc_78290_new_n2198_));
NOR2X1 NOR2X1_872 ( .A(u5__abc_78290_new_n1182_), .B(u5__abc_78290_new_n1105_), .Y(u5__abc_78290_new_n2199_));
NOR2X1 NOR2X1_873 ( .A(u5__abc_78290_new_n1375_), .B(u5__abc_78290_new_n2182_), .Y(u5__abc_78290_new_n2201_));
NOR2X1 NOR2X1_874 ( .A(u5__abc_78290_new_n2200_), .B(u5__abc_78290_new_n2202_), .Y(u5__abc_78290_new_n2203_));
NOR2X1 NOR2X1_875 ( .A(u5__abc_78290_new_n2194_), .B(u5__abc_78290_new_n2204_), .Y(u5__abc_78290_new_n2205_));
NOR2X1 NOR2X1_876 ( .A(u5__abc_78290_new_n2207_), .B(u5__abc_78290_new_n2176_), .Y(u5__abc_78290_new_n2208_));
NOR2X1 NOR2X1_877 ( .A(u5__abc_78290_new_n2190_), .B(u5__abc_78290_new_n2209_), .Y(u5__abc_78290_new_n2210_));
NOR2X1 NOR2X1_878 ( .A(u5__abc_78290_new_n1512_), .B(u5__abc_78290_new_n2149_), .Y(u5__abc_78290_new_n2214_));
NOR2X1 NOR2X1_879 ( .A(u5__abc_78290_new_n2214_), .B(u5__abc_78290_new_n1019_), .Y(u5__abc_78290_new_n2215_));
NOR2X1 NOR2X1_88 ( .A(u0__abc_74894_new_n4441_), .B(u0__abc_74894_new_n4440_), .Y(cs_need_rfr_1_));
NOR2X1 NOR2X1_880 ( .A(u5__abc_78290_new_n1433_), .B(u5__abc_78290_new_n2218_), .Y(u5__abc_78290_new_n2219_));
NOR2X1 NOR2X1_881 ( .A(u5__abc_78290_new_n2220_), .B(u5__abc_78290_new_n2179_), .Y(u5__abc_78290_new_n2221_));
NOR2X1 NOR2X1_882 ( .A(u5__abc_78290_new_n2215_), .B(u5__abc_78290_new_n2222_), .Y(u5__abc_78290_new_n2223_));
NOR2X1 NOR2X1_883 ( .A(tms_s_8_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2225_));
NOR2X1 NOR2X1_884 ( .A(tms_s_12_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2228_));
NOR2X1 NOR2X1_885 ( .A(tms_s_13_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2230_));
NOR2X1 NOR2X1_886 ( .A(tms_s_5_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2231_));
NOR2X1 NOR2X1_887 ( .A(u5_timer_1_), .B(u5__abc_78290_new_n2084_), .Y(u5__abc_78290_new_n2234_));
NOR2X1 NOR2X1_888 ( .A(tms_s_21_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2244_));
NOR2X1 NOR2X1_889 ( .A(u5__abc_78290_new_n2133_), .B(u5__abc_78290_new_n2145_), .Y(u5__abc_78290_new_n2248_));
NOR2X1 NOR2X1_89 ( .A(1'h0), .B(u0__abc_74894_new_n4443_), .Y(u0__abc_74894_new_n4444_));
NOR2X1 NOR2X1_890 ( .A(tms_s_9_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2259_));
NOR2X1 NOR2X1_891 ( .A(tms_s_22_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2264_));
NOR2X1 NOR2X1_892 ( .A(tms_s_21_), .B(u5__abc_78290_new_n2268_), .Y(u5__abc_78290_new_n2269_));
NOR2X1 NOR2X1_893 ( .A(u5__abc_78290_new_n2265_), .B(u5__abc_78290_new_n2270_), .Y(u5__abc_78290_new_n2271_));
NOR2X1 NOR2X1_894 ( .A(u5__abc_78290_new_n1998_), .B(u5__abc_78290_new_n2279_), .Y(u5__abc_78290_new_n2280_));
NOR2X1 NOR2X1_895 ( .A(u5__abc_78290_new_n1546_), .B(u5__abc_78290_new_n2285_), .Y(u5__abc_78290_new_n2286_));
NOR2X1 NOR2X1_896 ( .A(u5__abc_78290_new_n2287_), .B(u5__abc_78290_new_n2282_), .Y(u5__abc_78290_new_n2288_));
NOR2X1 NOR2X1_897 ( .A(u5__abc_78290_new_n2000_), .B(u5__abc_78290_new_n2289_), .Y(u5__abc_78290_new_n2290_));
NOR2X1 NOR2X1_898 ( .A(tms_s_10_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2303_));
NOR2X1 NOR2X1_899 ( .A(tms_s_14_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2306_));
NOR2X1 NOR2X1_9 ( .A(cs_le), .B(cs_1_), .Y(u0__abc_74894_new_n3481_));
NOR2X1 NOR2X1_90 ( .A(u0__abc_74894_new_n4447_), .B(u0__abc_74894_new_n4446_), .Y(cs_need_rfr_3_));
NOR2X1 NOR2X1_900 ( .A(tms_s_23_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2308_));
NOR2X1 NOR2X1_901 ( .A(u5__abc_78290_new_n2297_), .B(u5__abc_78290_new_n2033_), .Y(u5__abc_78290_new_n2320_));
NOR2X1 NOR2X1_902 ( .A(tms_s_3_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2323_));
NOR2X1 NOR2X1_903 ( .A(u5__abc_78290_new_n2330_), .B(u5__abc_78290_new_n2331_), .Y(u5__abc_78290_new_n2332_));
NOR2X1 NOR2X1_904 ( .A(u5__abc_78290_new_n2334_), .B(u5__abc_78290_new_n2332_), .Y(u5__abc_78290_new_n2335_));
NOR2X1 NOR2X1_905 ( .A(u5__abc_78290_new_n2314_), .B(u5__abc_78290_new_n2083_), .Y(u5__abc_78290_new_n2339_));
NOR2X1 NOR2X1_906 ( .A(u5_timer_4_), .B(u5__abc_78290_new_n2340_), .Y(u5__abc_78290_new_n2341_));
NOR2X1 NOR2X1_907 ( .A(u5_timer_5_), .B(u5__abc_78290_new_n2342_), .Y(u5__abc_78290_new_n2348_));
NOR2X1 NOR2X1_908 ( .A(u5_timer_5_), .B(u5_timer_6_), .Y(u5__abc_78290_new_n2356_));
NOR2X1 NOR2X1_909 ( .A(u5__abc_78290_new_n1486_), .B(u5__abc_78290_new_n1019_), .Y(u5__abc_78290_new_n2367_));
NOR2X1 NOR2X1_91 ( .A(1'h0), .B(u0__abc_74894_new_n4449_), .Y(u0__abc_74894_new_n4450_));
NOR2X1 NOR2X1_910 ( .A(u5__abc_78290_new_n2067_), .B(u5__abc_78290_new_n2370_), .Y(u5__abc_78290_new_n2371_));
NOR2X1 NOR2X1_911 ( .A(u5__abc_78290_new_n2376_), .B(u5__abc_78290_new_n2373_), .Y(u5__abc_78290_new_n2377_));
NOR2X1 NOR2X1_912 ( .A(u5__abc_78290_new_n2369_), .B(u5__abc_78290_new_n2378_), .Y(u5__abc_78290_new_n2379_));
NOR2X1 NOR2X1_913 ( .A(u5__abc_78290_new_n2383_), .B(u5__abc_78290_new_n2382_), .Y(u5__abc_78290_new_n2384_));
NOR2X1 NOR2X1_914 ( .A(u5__abc_78290_new_n2387_), .B(u5__abc_78290_new_n2382_), .Y(u5__abc_78290_new_n2388_));
NOR2X1 NOR2X1_915 ( .A(u5__abc_78290_new_n2389_), .B(u5__abc_78290_new_n2382_), .Y(u5__abc_78290_new_n2390_));
NOR2X1 NOR2X1_916 ( .A(u5_timer2_1_), .B(u5_timer2_0_), .Y(u5__abc_78290_new_n2396_));
NOR2X1 NOR2X1_917 ( .A(u5_timer2_2_), .B(u5__abc_78290_new_n2397_), .Y(u5__abc_78290_new_n2398_));
NOR2X1 NOR2X1_918 ( .A(u5_timer2_3_), .B(u5__abc_78290_new_n2399_), .Y(u5__abc_78290_new_n2400_));
NOR2X1 NOR2X1_919 ( .A(u5_timer2_6_), .B(u5__abc_78290_new_n2403_), .Y(u5__abc_78290_new_n2404_));
NOR2X1 NOR2X1_92 ( .A(u0__abc_74894_new_n4453_), .B(u0__abc_74894_new_n4452_), .Y(cs_need_rfr_5_));
NOR2X1 NOR2X1_920 ( .A(u5_timer2_7_), .B(u5__abc_78290_new_n2405_), .Y(u5__abc_78290_new_n2406_));
NOR2X1 NOR2X1_921 ( .A(u5__abc_78290_new_n1149_), .B(u5__abc_78290_new_n2410_), .Y(u5__abc_78290_new_n2411_));
NOR2X1 NOR2X1_922 ( .A(u5__abc_78290_new_n2412_), .B(u5__abc_78290_new_n2408_), .Y(u5__abc_78290_new_n2413_));
NOR2X1 NOR2X1_923 ( .A(u5__abc_78290_new_n1358_), .B(u5__abc_78290_new_n1124_), .Y(u5__abc_78290_new_n2418_));
NOR2X1 NOR2X1_924 ( .A(u5__abc_78290_new_n1300_), .B(u5__abc_78290_new_n1147_), .Y(u5__abc_78290_new_n2419_));
NOR2X1 NOR2X1_925 ( .A(u5__abc_78290_new_n2276_), .B(u5__abc_78290_new_n2420_), .Y(u5__abc_78290_new_n2421_));
NOR2X1 NOR2X1_926 ( .A(tms_s_17_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2433_));
NOR2X1 NOR2X1_927 ( .A(u5__abc_78290_new_n2434_), .B(u5__abc_78290_new_n2369_), .Y(u5__abc_78290_new_n2435_));
NOR2X1 NOR2X1_928 ( .A(u5__abc_78290_new_n682_), .B(u5__abc_78290_new_n2071_), .Y(u5__abc_78290_new_n2438_));
NOR2X1 NOR2X1_929 ( .A(u5__abc_78290_new_n2440_), .B(u5__abc_78290_new_n2439_), .Y(u5__abc_78290_new_n2441_));
NOR2X1 NOR2X1_93 ( .A(u0__abc_74894_new_n4455_), .B(u0__abc_74894_new_n4456_), .Y(cs_need_rfr_6_));
NOR2X1 NOR2X1_930 ( .A(u5__abc_78290_new_n986_), .B(u5__abc_78290_new_n2442_), .Y(u5__abc_78290_new_n2443_));
NOR2X1 NOR2X1_931 ( .A(u5__abc_78290_new_n1005_), .B(u5__abc_78290_new_n835_), .Y(u5__abc_78290_new_n2444_));
NOR2X1 NOR2X1_932 ( .A(u5__abc_78290_new_n2448_), .B(u5__abc_78290_new_n2447_), .Y(u5__abc_78290_new_n2449_));
NOR2X1 NOR2X1_933 ( .A(tms_s_18_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2464_));
NOR2X1 NOR2X1_934 ( .A(u5__abc_78290_new_n2265_), .B(u5__abc_78290_new_n2380_), .Y(u5__abc_78290_new_n2466_));
NOR2X1 NOR2X1_935 ( .A(u5__abc_78290_new_n2458_), .B(u5__abc_78290_new_n2429_), .Y(u5__abc_78290_new_n2479_));
NOR2X1 NOR2X1_936 ( .A(u5__abc_78290_new_n2395_), .B(u5__abc_78290_new_n2400_), .Y(u5__abc_78290_new_n2501_));
NOR2X1 NOR2X1_937 ( .A(tms_s_24_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2506_));
NOR2X1 NOR2X1_938 ( .A(u5__abc_78290_new_n2394_), .B(u5__abc_78290_new_n2402_), .Y(u5__abc_78290_new_n2512_));
NOR2X1 NOR2X1_939 ( .A(tms_s_25_), .B(u5__abc_78290_new_n1471_), .Y(u5__abc_78290_new_n2516_));
NOR2X1 NOR2X1_94 ( .A(1'h0), .B(u0__abc_74894_new_n4458_), .Y(u0__abc_74894_new_n4459_));
NOR2X1 NOR2X1_940 ( .A(u5__abc_78290_new_n1605_), .B(dv), .Y(u5__abc_78290_new_n2535_));
NOR2X1 NOR2X1_941 ( .A(u5__abc_78290_new_n1593_), .B(u5__abc_78290_new_n2542_), .Y(u5__abc_78290_new_n2543_));
NOR2X1 NOR2X1_942 ( .A(u5__abc_78290_new_n2218_), .B(u5__abc_78290_new_n2567_), .Y(u5__abc_78290_new_n2568_));
NOR2X1 NOR2X1_943 ( .A(u5__abc_78290_new_n2570_), .B(u5__abc_78290_new_n2194_), .Y(u5__abc_78290_new_n2571_));
NOR2X1 NOR2X1_944 ( .A(u5_cmd_asserted2), .B(u5__abc_78290_new_n2579_), .Y(u5__abc_78290_new_n2580_));
NOR2X1 NOR2X1_945 ( .A(u5__abc_78290_new_n2582_), .B(u5__abc_78290_new_n2577_), .Y(u5__abc_78290_new_n2583_));
NOR2X1 NOR2X1_946 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1335_), .Y(u5__abc_78290_new_n2591_));
NOR2X1 NOR2X1_947 ( .A(u5__abc_78290_new_n2598_), .B(u5__abc_78290_new_n1375_), .Y(u5__abc_78290_new_n2599_));
NOR2X1 NOR2X1_948 ( .A(u5__abc_78290_new_n1990_), .B(u5__abc_78290_new_n1490_), .Y(u5__abc_78290_new_n2601_));
NOR2X1 NOR2X1_949 ( .A(u5_ap_en), .B(u5__abc_78290_new_n2605_), .Y(u5__abc_78290_new_n2606_));
NOR2X1 NOR2X1_95 ( .A(u0_init_req0), .B(u0_init_req1), .Y(u0__abc_74894_new_n4467_));
NOR2X1 NOR2X1_950 ( .A(u5__abc_78290_new_n1418_), .B(u5__abc_78290_new_n2610_), .Y(u5__abc_78290_new_n2611_));
NOR2X1 NOR2X1_951 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n2615_), .Y(u5__abc_78290_new_n2616_));
NOR2X1 NOR2X1_952 ( .A(u5__abc_78290_new_n1422_), .B(u5__abc_78290_new_n2622_), .Y(u5__abc_78290_new_n2623_));
NOR2X1 NOR2X1_953 ( .A(u5_kro), .B(u5_ap_en), .Y(u5__abc_78290_new_n2626_));
NOR2X1 NOR2X1_954 ( .A(u5__abc_78290_new_n2628_), .B(u5__abc_78290_new_n1229_), .Y(u5__abc_78290_new_n2629_));
NOR2X1 NOR2X1_955 ( .A(u5__abc_78290_new_n2599_), .B(u5__abc_78290_new_n1374_), .Y(u5__abc_78290_new_n2631_));
NOR2X1 NOR2X1_956 ( .A(u5__abc_78290_new_n869_), .B(u5__abc_78290_new_n2589_), .Y(u5__abc_78290_new_n2644_));
NOR2X1 NOR2X1_957 ( .A(init_req), .B(u5__abc_78290_new_n1341_), .Y(u5__abc_78290_new_n2647_));
NOR2X1 NOR2X1_958 ( .A(u5__abc_78290_new_n2651_), .B(u5__abc_78290_new_n2650_), .Y(u5__abc_78290_new_n2652_));
NOR2X1 NOR2X1_959 ( .A(row_same), .B(u5__abc_78290_new_n2653_), .Y(u5__abc_78290_new_n2654_));
NOR2X1 NOR2X1_96 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n4468_));
NOR2X1 NOR2X1_960 ( .A(u5_state_5_), .B(u5_cmd_asserted), .Y(u5__abc_78290_new_n2661_));
NOR2X1 NOR2X1_961 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1514_), .Y(u5__abc_78290_new_n2664_));
NOR2X1 NOR2X1_962 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1336_), .Y(u5__abc_78290_new_n2666_));
NOR2X1 NOR2X1_963 ( .A(u5__abc_78290_new_n491_), .B(u5__abc_78290_new_n1828_), .Y(u5__abc_78290_new_n2671_));
NOR2X1 NOR2X1_964 ( .A(u5__abc_78290_new_n1375_), .B(u5__abc_78290_new_n2672_), .Y(u5__abc_78290_new_n2673_));
NOR2X1 NOR2X1_965 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n733_), .Y(u5__abc_78290_new_n2675_));
NOR2X1 NOR2X1_966 ( .A(u5__abc_78290_new_n2581_), .B(u5__abc_78290_new_n2578_), .Y(u5__abc_78290_new_n2678_));
NOR2X1 NOR2X1_967 ( .A(u5__abc_78290_new_n2679_), .B(u5__abc_78290_new_n2678_), .Y(u5__abc_78290_new_n2680_));
NOR2X1 NOR2X1_968 ( .A(u5__abc_78290_new_n777_), .B(u5__abc_78290_new_n2683_), .Y(u5__abc_78290_new_n2684_));
NOR2X1 NOR2X1_969 ( .A(u5__abc_78290_new_n741_), .B(u5__abc_78290_new_n1414_), .Y(u5__abc_78290_new_n2689_));
NOR2X1 NOR2X1_97 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n4470_));
NOR2X1 NOR2X1_970 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n1267_), .Y(u5__abc_78290_new_n2701_));
NOR2X1 NOR2X1_971 ( .A(u5__abc_78290_new_n1277_), .B(u5__abc_78290_new_n1053_), .Y(u5__abc_78290_new_n2713_));
NOR2X1 NOR2X1_972 ( .A(u5__abc_78290_new_n492_), .B(u5__abc_78290_new_n2591_), .Y(u5__abc_78290_new_n2717_));
NOR2X1 NOR2X1_973 ( .A(u5_state_12_), .B(u5__abc_78290_new_n1609_), .Y(u5__abc_78290_new_n2721_));
NOR2X1 NOR2X1_974 ( .A(u5__abc_78290_new_n747_), .B(u5__abc_78290_new_n2591_), .Y(u5__abc_78290_new_n2722_));
NOR2X1 NOR2X1_975 ( .A(u5__abc_78290_new_n747_), .B(u5__abc_78290_new_n2625_), .Y(u5__abc_78290_new_n2723_));
NOR2X1 NOR2X1_976 ( .A(u1_wb_write_go), .B(u5__abc_78290_new_n1990_), .Y(u5__abc_78290_new_n2732_));
NOR2X1 NOR2X1_977 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n834_), .Y(u5__abc_78290_new_n2740_));
NOR2X1 NOR2X1_978 ( .A(u5__abc_78290_new_n564_), .B(u5__abc_78290_new_n2601_), .Y(u5__abc_78290_new_n2759_));
NOR2X1 NOR2X1_979 ( .A(u5_state_16_), .B(u5_cmd_asserted), .Y(u5__abc_78290_new_n2760_));
NOR2X1 NOR2X1_98 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n4471_));
NOR2X1 NOR2X1_980 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n571_), .Y(u5__abc_78290_new_n2774_));
NOR2X1 NOR2X1_981 ( .A(u5__abc_78290_new_n1336_), .B(u5__abc_78290_new_n1337_), .Y(u5__abc_78290_new_n2782_));
NOR2X1 NOR2X1_982 ( .A(u5__abc_78290_new_n2784_), .B(u5__abc_78290_new_n2593_), .Y(u5__abc_78290_new_n2785_));
NOR2X1 NOR2X1_983 ( .A(u5__abc_78290_new_n2789_), .B(u5__abc_78290_new_n2577_), .Y(u5__abc_78290_new_n2790_));
NOR2X1 NOR2X1_984 ( .A(rfr_req), .B(u5__abc_78290_new_n1019_), .Y(u5__abc_78290_new_n2795_));
NOR2X1 NOR2X1_985 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n603_), .Y(u5__abc_78290_new_n2799_));
NOR2X1 NOR2X1_986 ( .A(u5__abc_78290_new_n2802_), .B(u5__abc_78290_new_n2796_), .Y(u5_next_state_21_));
NOR2X1 NOR2X1_987 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n596_), .Y(u5__abc_78290_new_n2805_));
NOR2X1 NOR2X1_988 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n590_), .Y(u5__abc_78290_new_n2810_));
NOR2X1 NOR2X1_989 ( .A(u5__abc_78290_new_n2813_), .B(u5__abc_78290_new_n2577_), .Y(u5__abc_78290_new_n2814_));
NOR2X1 NOR2X1_99 ( .A(1'h0), .B(u0__abc_74894_new_n4473_), .Y(u0__abc_74894_new_n4474_));
NOR2X1 NOR2X1_990 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n582_), .Y(u5__abc_78290_new_n2822_));
NOR2X1 NOR2X1_991 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n548_), .Y(u5__abc_78290_new_n2827_));
NOR2X1 NOR2X1_992 ( .A(u5__abc_78290_new_n2833_), .B(u5__abc_78290_new_n2577_), .Y(u5__abc_78290_new_n2834_));
NOR2X1 NOR2X1_993 ( .A(u5_state_31_), .B(u5_resume_req_r), .Y(u5__abc_78290_new_n2850_));
NOR2X1 NOR2X1_994 ( .A(u5__abc_78290_new_n2679_), .B(u5__abc_78290_new_n2856_), .Y(u5_next_state_33_));
NOR2X1 NOR2X1_995 ( .A(csc_s_1_), .B(u5__abc_78290_new_n1322_), .Y(u5__abc_78290_new_n2863_));
NOR2X1 NOR2X1_996 ( .A(u5__abc_78290_new_n2866_), .B(u5__abc_78290_new_n2867_), .Y(u5_next_state_36_));
NOR2X1 NOR2X1_997 ( .A(u5__abc_78290_new_n2869_), .B(u5__abc_78290_new_n1382_), .Y(u5__abc_78290_new_n2870_));
NOR2X1 NOR2X1_998 ( .A(u5__abc_78290_new_n1394_), .B(u5__abc_78290_new_n2870_), .Y(u5__abc_78290_new_n2871_));
NOR2X1 NOR2X1_999 ( .A(csc_s_5_), .B(u5__abc_78290_new_n2565_), .Y(u5__abc_78290_new_n2873_));
NOR3X1 NOR3X1_1 ( .A(init_ack), .B(lmr_ack), .C(cs_0_), .Y(_abc_81086_new_n238_));
NOR3X1 NOR3X1_10 ( .A(u0__abc_74894_new_n3790_), .B(u0__abc_74894_new_n3792_), .C(u0__abc_74894_new_n3794_), .Y(u0__abc_74894_new_n3795_));
NOR3X1 NOR3X1_11 ( .A(u0__abc_74894_new_n3833_), .B(u0__abc_74894_new_n3835_), .C(u0__abc_74894_new_n3837_), .Y(u0__abc_74894_new_n3838_));
NOR3X1 NOR3X1_12 ( .A(u0__abc_74894_new_n3842_), .B(u0__abc_74894_new_n3844_), .C(u0__abc_74894_new_n3847_), .Y(u0__abc_74894_new_n3848_));
NOR3X1 NOR3X1_13 ( .A(u0__abc_74894_new_n3874_), .B(u0__abc_74894_new_n3876_), .C(u0__abc_74894_new_n3878_), .Y(u0__abc_74894_new_n3879_));
NOR3X1 NOR3X1_14 ( .A(u0__abc_74894_new_n3950_), .B(u0__abc_74894_new_n3952_), .C(u0__abc_74894_new_n3954_), .Y(u0__abc_74894_new_n3955_));
NOR3X1 NOR3X1_15 ( .A(u0__abc_74894_new_n4251_), .B(u0__abc_74894_new_n4249_), .C(u0__abc_74894_new_n4245_), .Y(u0__abc_74894_new_n4252_));
NOR3X1 NOR3X1_16 ( .A(u0__abc_74894_new_n4277_), .B(u0__abc_74894_new_n4271_), .C(u0__abc_74894_new_n4275_), .Y(u0__abc_74894_new_n4278_));
NOR3X1 NOR3X1_17 ( .A(u0__abc_74894_new_n4303_), .B(u0__abc_74894_new_n4301_), .C(u0__abc_74894_new_n4297_), .Y(u0__abc_74894_new_n4304_));
NOR3X1 NOR3X1_18 ( .A(u0__abc_74894_new_n4330_), .B(u0__abc_74894_new_n4327_), .C(u0__abc_74894_new_n4323_), .Y(u0__abc_74894_new_n4331_));
NOR3X1 NOR3X1_19 ( .A(u0__abc_74894_new_n4356_), .B(u0__abc_74894_new_n4354_), .C(u0__abc_74894_new_n4350_), .Y(u0__abc_74894_new_n4357_));
NOR3X1 NOR3X1_2 ( .A(init_ack), .B(lmr_ack), .C(cs_1_), .Y(_abc_81086_new_n243_));
NOR3X1 NOR3X1_20 ( .A(u0__abc_74894_new_n4372_), .B(u0__abc_74894_new_n4376_), .C(u0__abc_74894_new_n4380_), .Y(u0__abc_74894_new_n4381_));
NOR3X1 NOR3X1_21 ( .A(u0__abc_74894_new_n4396_), .B(u0__abc_74894_new_n4400_), .C(u0__abc_74894_new_n4404_), .Y(u0__abc_74894_new_n4405_));
NOR3X1 NOR3X1_22 ( .A(u0__abc_74894_new_n4420_), .B(u0__abc_74894_new_n4424_), .C(u0__abc_74894_new_n4428_), .Y(u0__abc_74894_new_n4429_));
NOR3X1 NOR3X1_23 ( .A(u0_u0_addr_r_6_), .B(u0_u0_addr_r_5_), .C(u0_u0__abc_72207_new_n320_), .Y(u0_u0__abc_72207_new_n321_));
NOR3X1 NOR3X1_24 ( .A(u1__abc_72801_new_n332_), .B(u1__abc_72801_new_n334_), .C(u1__abc_72801_new_n338_), .Y(u1__abc_72801_new_n339_));
NOR3X1 NOR3X1_25 ( .A(u1_bas), .B(u1__abc_72801_new_n342_), .C(u1__abc_72801_new_n339_), .Y(u1__abc_72801_new_n343_));
NOR3X1 NOR3X1_26 ( .A(u1__abc_72801_new_n340_), .B(u1__abc_72801_new_n264_), .C(u1__abc_72801_new_n350_), .Y(u1__abc_72801_new_n351_));
NOR3X1 NOR3X1_27 ( .A(u1__abc_72801_new_n399_), .B(u1__abc_72801_new_n334_), .C(u1__abc_72801_new_n338_), .Y(u1__abc_72801_new_n400_));
NOR3X1 NOR3X1_28 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n401_), .C(u1__abc_72801_new_n400_), .Y(u1__abc_72801_new_n402_));
NOR3X1 NOR3X1_29 ( .A(u1__abc_72801_new_n408_), .B(u1__abc_72801_new_n334_), .C(u1__abc_72801_new_n338_), .Y(u1__abc_72801_new_n409_));
NOR3X1 NOR3X1_3 ( .A(init_ack), .B(lmr_ack), .C(cs_2_), .Y(_abc_81086_new_n247_));
NOR3X1 NOR3X1_30 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n410_), .C(u1__abc_72801_new_n409_), .Y(u1__abc_72801_new_n411_));
NOR3X1 NOR3X1_31 ( .A(u1__abc_72801_new_n432_), .B(u1__abc_72801_new_n334_), .C(u1__abc_72801_new_n338_), .Y(u1__abc_72801_new_n433_));
NOR3X1 NOR3X1_32 ( .A(u1__abc_72801_new_n423_), .B(u1__abc_72801_new_n334_), .C(u1__abc_72801_new_n338_), .Y(u1__abc_72801_new_n442_));
NOR3X1 NOR3X1_33 ( .A(u1__abc_72801_new_n444_), .B(u1__abc_72801_new_n445_), .C(u1__abc_72801_new_n442_), .Y(u1__abc_72801_new_n446_));
NOR3X1 NOR3X1_34 ( .A(u1_u0__abc_72719_new_n99_), .B(u1_u0__abc_72719_new_n103_), .C(u1_u0__abc_72719_new_n91_), .Y(u1_u0__abc_72719_new_n104_));
NOR3X1 NOR3X1_35 ( .A(u1_u0__abc_72719_new_n119_), .B(u1_u0__abc_72719_new_n115_), .C(u1_u0__abc_72719_new_n97_), .Y(u1_u0__abc_72719_new_n126_));
NOR3X1 NOR3X1_36 ( .A(u2_u0__abc_73914_new_n292_), .B(u2_u0__abc_73914_new_n287_), .C(u2_u0__abc_73914_new_n296_), .Y(u2_u0__abc_73914_new_n297_));
NOR3X1 NOR3X1_37 ( .A(u2_u0__abc_73914_new_n327_), .B(u2_u0__abc_73914_new_n318_), .C(u2_u0__abc_73914_new_n322_), .Y(u2_u0__abc_73914_new_n328_));
NOR3X1 NOR3X1_38 ( .A(u2_u0__abc_73914_new_n344_), .B(u2_u0__abc_73914_new_n338_), .C(u2_u0__abc_73914_new_n333_), .Y(u2_u0__abc_73914_new_n345_));
NOR3X1 NOR3X1_39 ( .A(u2_u0__abc_73914_new_n391_), .B(u2_u0__abc_73914_new_n387_), .C(u2_u0__abc_73914_new_n394_), .Y(u2_u0__abc_73914_new_n395_));
NOR3X1 NOR3X1_4 ( .A(init_ack), .B(lmr_ack), .C(cs_3_), .Y(_abc_81086_new_n251_));
NOR3X1 NOR3X1_40 ( .A(u2_u1__abc_73914_new_n292_), .B(u2_u1__abc_73914_new_n287_), .C(u2_u1__abc_73914_new_n296_), .Y(u2_u1__abc_73914_new_n297_));
NOR3X1 NOR3X1_41 ( .A(u2_u1__abc_73914_new_n327_), .B(u2_u1__abc_73914_new_n318_), .C(u2_u1__abc_73914_new_n322_), .Y(u2_u1__abc_73914_new_n328_));
NOR3X1 NOR3X1_42 ( .A(u2_u1__abc_73914_new_n344_), .B(u2_u1__abc_73914_new_n338_), .C(u2_u1__abc_73914_new_n333_), .Y(u2_u1__abc_73914_new_n345_));
NOR3X1 NOR3X1_43 ( .A(u2_u1__abc_73914_new_n391_), .B(u2_u1__abc_73914_new_n387_), .C(u2_u1__abc_73914_new_n394_), .Y(u2_u1__abc_73914_new_n395_));
NOR3X1 NOR3X1_44 ( .A(u4__abc_74770_new_n101_), .B(u4__abc_74770_new_n111_), .C(u4__abc_74770_new_n102_), .Y(u4__abc_74770_new_n112_));
NOR3X1 NOR3X1_45 ( .A(u4__abc_74770_new_n147_), .B(u4__abc_74770_new_n139_), .C(u4__abc_74770_new_n154_), .Y(u4__abc_74770_new_n165_));
NOR3X1 NOR3X1_46 ( .A(u5__abc_78290_new_n384_), .B(u5__abc_78290_new_n622_), .C(u5__abc_78290_new_n477_), .Y(u5__abc_78290_new_n623_));
NOR3X1 NOR3X1_47 ( .A(u5__abc_78290_new_n770_), .B(u5__abc_78290_new_n773_), .C(u5__abc_78290_new_n415_), .Y(u5__abc_78290_new_n774_));
NOR3X1 NOR3X1_48 ( .A(u5__abc_78290_new_n601_), .B(u5__abc_78290_new_n415_), .C(u5__abc_78290_new_n422_), .Y(u5__abc_78290_new_n820_));
NOR3X1 NOR3X1_49 ( .A(u5_state_62_), .B(u5__abc_78290_new_n878_), .C(u5__abc_78290_new_n457_), .Y(u5__abc_78290_new_n879_));
NOR3X1 NOR3X1_5 ( .A(init_ack), .B(lmr_ack), .C(cs_4_), .Y(_abc_81086_new_n255_));
NOR3X1 NOR3X1_50 ( .A(u5__abc_78290_new_n998_), .B(u5__abc_78290_new_n835_), .C(u5__abc_78290_new_n822_), .Y(u5__abc_78290_new_n999_));
NOR3X1 NOR3X1_51 ( .A(u5__abc_78290_new_n1011_), .B(u5__abc_78290_new_n1001_), .C(u5__abc_78290_new_n1017_), .Y(u5__abc_78290_new_n1018_));
NOR3X1 NOR3X1_52 ( .A(u5__abc_78290_new_n1043_), .B(u5__abc_78290_new_n1071_), .C(u5__abc_78290_new_n1063_), .Y(u5__abc_78290_new_n1072_));
NOR3X1 NOR3X1_53 ( .A(u5__abc_78290_new_n1718_), .B(u5__abc_78290_new_n1950_), .C(u5__abc_78290_new_n2110_), .Y(u5__abc_78290_new_n2111_));
NOR3X1 NOR3X1_6 ( .A(init_ack), .B(lmr_ack), .C(cs_5_), .Y(_abc_81086_new_n259_));
NOR3X1 NOR3X1_7 ( .A(init_ack), .B(lmr_ack), .C(cs_6_), .Y(_abc_81086_new_n263_));
NOR3X1 NOR3X1_8 ( .A(init_ack), .B(lmr_ack), .C(cs_7_), .Y(_abc_81086_new_n267_));
NOR3X1 NOR3X1_9 ( .A(u0__abc_74894_new_n3771_), .B(u0__abc_74894_new_n3773_), .C(u0__abc_74894_new_n3775_), .Y(u0__abc_74894_new_n3776_));
OAI21X1 OAI21X1_1 ( .A(susp_sel), .B(rfr_ack), .C(cs_need_rfr_0_), .Y(_abc_81086_new_n239_));
OAI21X1 OAI21X1_10 ( .A(susp_sel), .B(rfr_ack), .C(cs_need_rfr_3_), .Y(_abc_81086_new_n252_));
OAI21X1 OAI21X1_100 ( .A(u0__abc_74894_new_n1101_), .B(u0_init_req1), .C(u0__abc_74894_new_n1109_), .Y(u0__abc_74894_new_n1110_));
OAI21X1 OAI21X1_1000 ( .A(csc_5_), .B(u3_byte0_5_), .C(u3__abc_73372_new_n518_), .Y(u3__abc_73372_new_n519_));
OAI21X1 OAI21X1_1001 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n519_), .C(u3__abc_73372_new_n520_), .Y(mem_dout_5_));
OAI21X1 OAI21X1_1002 ( .A(csc_5_), .B(u3_byte0_6_), .C(u3__abc_73372_new_n522_), .Y(u3__abc_73372_new_n523_));
OAI21X1 OAI21X1_1003 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n523_), .C(u3__abc_73372_new_n524_), .Y(mem_dout_6_));
OAI21X1 OAI21X1_1004 ( .A(csc_5_), .B(u3_byte0_7_), .C(u3__abc_73372_new_n526_), .Y(u3__abc_73372_new_n527_));
OAI21X1 OAI21X1_1005 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n527_), .C(u3__abc_73372_new_n528_), .Y(mem_dout_7_));
OAI21X1 OAI21X1_1006 ( .A(csc_5_), .B(u3_byte1_0_), .C(u3__abc_73372_new_n530_), .Y(u3__abc_73372_new_n531_));
OAI21X1 OAI21X1_1007 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n531_), .C(u3__abc_73372_new_n532_), .Y(mem_dout_8_));
OAI21X1 OAI21X1_1008 ( .A(csc_5_), .B(u3_byte1_1_), .C(u3__abc_73372_new_n534_), .Y(u3__abc_73372_new_n535_));
OAI21X1 OAI21X1_1009 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n535_), .C(u3__abc_73372_new_n536_), .Y(mem_dout_9_));
OAI21X1 OAI21X1_101 ( .A(u0__abc_74894_new_n1101_), .B(1'h0), .C(u0__abc_74894_new_n1114_), .Y(u0__abc_74894_new_n1115_));
OAI21X1 OAI21X1_1010 ( .A(csc_5_), .B(u3_byte1_2_), .C(u3__abc_73372_new_n538_), .Y(u3__abc_73372_new_n539_));
OAI21X1 OAI21X1_1011 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n539_), .C(u3__abc_73372_new_n540_), .Y(mem_dout_10_));
OAI21X1 OAI21X1_1012 ( .A(csc_5_), .B(u3_byte1_3_), .C(u3__abc_73372_new_n542_), .Y(u3__abc_73372_new_n543_));
OAI21X1 OAI21X1_1013 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n543_), .C(u3__abc_73372_new_n544_), .Y(mem_dout_11_));
OAI21X1 OAI21X1_1014 ( .A(csc_5_), .B(u3_byte1_4_), .C(u3__abc_73372_new_n546_), .Y(u3__abc_73372_new_n547_));
OAI21X1 OAI21X1_1015 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n547_), .C(u3__abc_73372_new_n548_), .Y(mem_dout_12_));
OAI21X1 OAI21X1_1016 ( .A(csc_5_), .B(u3_byte1_5_), .C(u3__abc_73372_new_n550_), .Y(u3__abc_73372_new_n551_));
OAI21X1 OAI21X1_1017 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n551_), .C(u3__abc_73372_new_n552_), .Y(mem_dout_13_));
OAI21X1 OAI21X1_1018 ( .A(csc_5_), .B(u3_byte1_6_), .C(u3__abc_73372_new_n554_), .Y(u3__abc_73372_new_n555_));
OAI21X1 OAI21X1_1019 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n555_), .C(u3__abc_73372_new_n556_), .Y(mem_dout_14_));
OAI21X1 OAI21X1_102 ( .A(init_req), .B(u0__abc_74894_new_n1120_), .C(u0__abc_74894_new_n1121_), .Y(u0__abc_74894_new_n1122_));
OAI21X1 OAI21X1_1020 ( .A(csc_5_), .B(u3_byte1_7_), .C(u3__abc_73372_new_n558_), .Y(u3__abc_73372_new_n559_));
OAI21X1 OAI21X1_1021 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n559_), .C(u3__abc_73372_new_n560_), .Y(mem_dout_15_));
OAI21X1 OAI21X1_1022 ( .A(u3__abc_73372_new_n626_), .B(u3__abc_73372_new_n627_), .C(wb_cyc_i), .Y(u3_rd_fifo_clr));
OAI21X1 OAI21X1_1023 ( .A(u3__abc_73372_new_n635_), .B(u3__abc_73372_new_n636_), .C(u3__abc_73372_new_n634_), .Y(u3__abc_73372_new_n637_));
OAI21X1 OAI21X1_1024 ( .A(u3__abc_73372_new_n635_), .B(u3__abc_73372_new_n636_), .C(u3_rd_fifo_out_33_), .Y(u3__abc_73372_new_n640_));
OAI21X1 OAI21X1_1025 ( .A(u3__abc_73372_new_n655_), .B(u3__abc_73372_new_n658_), .C(u3__abc_73372_new_n651_), .Y(u3__abc_73372_new_n659_));
OAI21X1 OAI21X1_1026 ( .A(u3__abc_73372_new_n680_), .B(u3__abc_73372_new_n685_), .C(u3__abc_73372_new_n684_), .Y(u3__abc_73372_new_n686_));
OAI21X1 OAI21X1_1027 ( .A(u3__abc_73372_new_n680_), .B(u3__abc_73372_new_n685_), .C(u3_rd_fifo_out_32_), .Y(u3__abc_73372_new_n689_));
OAI21X1 OAI21X1_1028 ( .A(u3__abc_73372_new_n705_), .B(u3__abc_73372_new_n708_), .C(u3__abc_73372_new_n701_), .Y(u3__abc_73372_new_n709_));
OAI21X1 OAI21X1_1029 ( .A(u3_u0__abc_74260_new_n382_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n384_), .Y(u3_u0__0r1_35_0__0_));
OAI21X1 OAI21X1_103 ( .A(init_req), .B(u0__abc_74894_new_n1126_), .C(u0__abc_74894_new_n1127_), .Y(u0__abc_74894_new_n1128_));
OAI21X1 OAI21X1_1030 ( .A(u3_u0__abc_74260_new_n386_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n387_), .Y(u3_u0__0r1_35_0__1_));
OAI21X1 OAI21X1_1031 ( .A(u3_u0__abc_74260_new_n389_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n390_), .Y(u3_u0__0r1_35_0__2_));
OAI21X1 OAI21X1_1032 ( .A(u3_u0__abc_74260_new_n392_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n393_), .Y(u3_u0__0r1_35_0__3_));
OAI21X1 OAI21X1_1033 ( .A(u3_u0__abc_74260_new_n395_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n396_), .Y(u3_u0__0r1_35_0__4_));
OAI21X1 OAI21X1_1034 ( .A(u3_u0__abc_74260_new_n398_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n399_), .Y(u3_u0__0r1_35_0__5_));
OAI21X1 OAI21X1_1035 ( .A(u3_u0__abc_74260_new_n401_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n402_), .Y(u3_u0__0r1_35_0__6_));
OAI21X1 OAI21X1_1036 ( .A(u3_u0__abc_74260_new_n404_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n405_), .Y(u3_u0__0r1_35_0__7_));
OAI21X1 OAI21X1_1037 ( .A(u3_u0__abc_74260_new_n407_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n408_), .Y(u3_u0__0r1_35_0__8_));
OAI21X1 OAI21X1_1038 ( .A(u3_u0__abc_74260_new_n410_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n411_), .Y(u3_u0__0r1_35_0__9_));
OAI21X1 OAI21X1_1039 ( .A(u3_u0__abc_74260_new_n413_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n414_), .Y(u3_u0__0r1_35_0__10_));
OAI21X1 OAI21X1_104 ( .A(init_req), .B(u0__abc_74894_new_n1135_), .C(u0__abc_74894_new_n1136_), .Y(u0__abc_74894_new_n1137_));
OAI21X1 OAI21X1_1040 ( .A(u3_u0__abc_74260_new_n416_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n417_), .Y(u3_u0__0r1_35_0__11_));
OAI21X1 OAI21X1_1041 ( .A(u3_u0__abc_74260_new_n419_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n420_), .Y(u3_u0__0r1_35_0__12_));
OAI21X1 OAI21X1_1042 ( .A(u3_u0__abc_74260_new_n422_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n423_), .Y(u3_u0__0r1_35_0__13_));
OAI21X1 OAI21X1_1043 ( .A(u3_u0__abc_74260_new_n425_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n426_), .Y(u3_u0__0r1_35_0__14_));
OAI21X1 OAI21X1_1044 ( .A(u3_u0__abc_74260_new_n428_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n429_), .Y(u3_u0__0r1_35_0__15_));
OAI21X1 OAI21X1_1045 ( .A(u3_u0__abc_74260_new_n431_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n432_), .Y(u3_u0__0r1_35_0__16_));
OAI21X1 OAI21X1_1046 ( .A(u3_u0__abc_74260_new_n434_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n435_), .Y(u3_u0__0r1_35_0__17_));
OAI21X1 OAI21X1_1047 ( .A(u3_u0__abc_74260_new_n437_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n438_), .Y(u3_u0__0r1_35_0__18_));
OAI21X1 OAI21X1_1048 ( .A(u3_u0__abc_74260_new_n440_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n441_), .Y(u3_u0__0r1_35_0__19_));
OAI21X1 OAI21X1_1049 ( .A(u3_u0__abc_74260_new_n443_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n444_), .Y(u3_u0__0r1_35_0__20_));
OAI21X1 OAI21X1_105 ( .A(init_req), .B(u0__abc_74894_new_n1141_), .C(u0__abc_74894_new_n1142_), .Y(u0__abc_74894_new_n1143_));
OAI21X1 OAI21X1_1050 ( .A(u3_u0__abc_74260_new_n446_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n447_), .Y(u3_u0__0r1_35_0__21_));
OAI21X1 OAI21X1_1051 ( .A(u3_u0__abc_74260_new_n449_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n450_), .Y(u3_u0__0r1_35_0__22_));
OAI21X1 OAI21X1_1052 ( .A(u3_u0__abc_74260_new_n452_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n453_), .Y(u3_u0__0r1_35_0__23_));
OAI21X1 OAI21X1_1053 ( .A(u3_u0__abc_74260_new_n455_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n456_), .Y(u3_u0__0r1_35_0__24_));
OAI21X1 OAI21X1_1054 ( .A(u3_u0__abc_74260_new_n458_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n459_), .Y(u3_u0__0r1_35_0__25_));
OAI21X1 OAI21X1_1055 ( .A(u3_u0__abc_74260_new_n461_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n462_), .Y(u3_u0__0r1_35_0__26_));
OAI21X1 OAI21X1_1056 ( .A(u3_u0__abc_74260_new_n464_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n465_), .Y(u3_u0__0r1_35_0__27_));
OAI21X1 OAI21X1_1057 ( .A(u3_u0__abc_74260_new_n467_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n468_), .Y(u3_u0__0r1_35_0__28_));
OAI21X1 OAI21X1_1058 ( .A(u3_u0__abc_74260_new_n470_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n471_), .Y(u3_u0__0r1_35_0__29_));
OAI21X1 OAI21X1_1059 ( .A(u3_u0__abc_74260_new_n473_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n474_), .Y(u3_u0__0r1_35_0__30_));
OAI21X1 OAI21X1_106 ( .A(init_req), .B(u0__abc_74894_new_n1149_), .C(u0__abc_74894_new_n1150_), .Y(u0__abc_74894_new_n1151_));
OAI21X1 OAI21X1_1060 ( .A(u3_u0__abc_74260_new_n476_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n477_), .Y(u3_u0__0r1_35_0__31_));
OAI21X1 OAI21X1_1061 ( .A(u3_u0__abc_74260_new_n479_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n480_), .Y(u3_u0__0r1_35_0__32_));
OAI21X1 OAI21X1_1062 ( .A(u3_u0__abc_74260_new_n482_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n483_), .Y(u3_u0__0r1_35_0__33_));
OAI21X1 OAI21X1_1063 ( .A(u3_u0__abc_74260_new_n485_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n486_), .Y(u3_u0__0r1_35_0__34_));
OAI21X1 OAI21X1_1064 ( .A(u3_u0__abc_74260_new_n488_), .B(u3_u0__abc_74260_new_n383_), .C(u3_u0__abc_74260_new_n489_), .Y(u3_u0__0r1_35_0__35_));
OAI21X1 OAI21X1_1065 ( .A(u3_u0__abc_74260_new_n382_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n492_), .Y(u3_u0__0r3_35_0__0_));
OAI21X1 OAI21X1_1066 ( .A(u3_u0__abc_74260_new_n386_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n494_), .Y(u3_u0__0r3_35_0__1_));
OAI21X1 OAI21X1_1067 ( .A(u3_u0__abc_74260_new_n389_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n496_), .Y(u3_u0__0r3_35_0__2_));
OAI21X1 OAI21X1_1068 ( .A(u3_u0__abc_74260_new_n392_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n498_), .Y(u3_u0__0r3_35_0__3_));
OAI21X1 OAI21X1_1069 ( .A(u3_u0__abc_74260_new_n395_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n500_), .Y(u3_u0__0r3_35_0__4_));
OAI21X1 OAI21X1_107 ( .A(cs_le_d), .B(u0_rf_we), .C(u0__abc_74894_new_n1154_), .Y(u0__abc_74894_new_n1155_));
OAI21X1 OAI21X1_1070 ( .A(u3_u0__abc_74260_new_n398_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n502_), .Y(u3_u0__0r3_35_0__5_));
OAI21X1 OAI21X1_1071 ( .A(u3_u0__abc_74260_new_n401_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n504_), .Y(u3_u0__0r3_35_0__6_));
OAI21X1 OAI21X1_1072 ( .A(u3_u0__abc_74260_new_n404_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n506_), .Y(u3_u0__0r3_35_0__7_));
OAI21X1 OAI21X1_1073 ( .A(u3_u0__abc_74260_new_n407_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n508_), .Y(u3_u0__0r3_35_0__8_));
OAI21X1 OAI21X1_1074 ( .A(u3_u0__abc_74260_new_n410_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n510_), .Y(u3_u0__0r3_35_0__9_));
OAI21X1 OAI21X1_1075 ( .A(u3_u0__abc_74260_new_n413_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n512_), .Y(u3_u0__0r3_35_0__10_));
OAI21X1 OAI21X1_1076 ( .A(u3_u0__abc_74260_new_n416_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n514_), .Y(u3_u0__0r3_35_0__11_));
OAI21X1 OAI21X1_1077 ( .A(u3_u0__abc_74260_new_n419_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n516_), .Y(u3_u0__0r3_35_0__12_));
OAI21X1 OAI21X1_1078 ( .A(u3_u0__abc_74260_new_n422_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n518_), .Y(u3_u0__0r3_35_0__13_));
OAI21X1 OAI21X1_1079 ( .A(u3_u0__abc_74260_new_n425_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n520_), .Y(u3_u0__0r3_35_0__14_));
OAI21X1 OAI21X1_108 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1170_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1171_));
OAI21X1 OAI21X1_1080 ( .A(u3_u0__abc_74260_new_n428_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n522_), .Y(u3_u0__0r3_35_0__15_));
OAI21X1 OAI21X1_1081 ( .A(u3_u0__abc_74260_new_n431_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n524_), .Y(u3_u0__0r3_35_0__16_));
OAI21X1 OAI21X1_1082 ( .A(u3_u0__abc_74260_new_n434_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n526_), .Y(u3_u0__0r3_35_0__17_));
OAI21X1 OAI21X1_1083 ( .A(u3_u0__abc_74260_new_n437_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n528_), .Y(u3_u0__0r3_35_0__18_));
OAI21X1 OAI21X1_1084 ( .A(u3_u0__abc_74260_new_n440_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n530_), .Y(u3_u0__0r3_35_0__19_));
OAI21X1 OAI21X1_1085 ( .A(u3_u0__abc_74260_new_n443_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n532_), .Y(u3_u0__0r3_35_0__20_));
OAI21X1 OAI21X1_1086 ( .A(u3_u0__abc_74260_new_n446_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n534_), .Y(u3_u0__0r3_35_0__21_));
OAI21X1 OAI21X1_1087 ( .A(u3_u0__abc_74260_new_n449_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n536_), .Y(u3_u0__0r3_35_0__22_));
OAI21X1 OAI21X1_1088 ( .A(u3_u0__abc_74260_new_n452_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n538_), .Y(u3_u0__0r3_35_0__23_));
OAI21X1 OAI21X1_1089 ( .A(u3_u0__abc_74260_new_n455_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n540_), .Y(u3_u0__0r3_35_0__24_));
OAI21X1 OAI21X1_109 ( .A(u0__abc_74894_new_n1171_), .B(u0__abc_74894_new_n1169_), .C(u0__abc_74894_new_n1173_), .Y(u0__abc_74894_new_n1174_));
OAI21X1 OAI21X1_1090 ( .A(u3_u0__abc_74260_new_n458_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n542_), .Y(u3_u0__0r3_35_0__25_));
OAI21X1 OAI21X1_1091 ( .A(u3_u0__abc_74260_new_n461_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n544_), .Y(u3_u0__0r3_35_0__26_));
OAI21X1 OAI21X1_1092 ( .A(u3_u0__abc_74260_new_n464_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n546_), .Y(u3_u0__0r3_35_0__27_));
OAI21X1 OAI21X1_1093 ( .A(u3_u0__abc_74260_new_n467_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n548_), .Y(u3_u0__0r3_35_0__28_));
OAI21X1 OAI21X1_1094 ( .A(u3_u0__abc_74260_new_n470_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n550_), .Y(u3_u0__0r3_35_0__29_));
OAI21X1 OAI21X1_1095 ( .A(u3_u0__abc_74260_new_n473_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n552_), .Y(u3_u0__0r3_35_0__30_));
OAI21X1 OAI21X1_1096 ( .A(u3_u0__abc_74260_new_n476_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n554_), .Y(u3_u0__0r3_35_0__31_));
OAI21X1 OAI21X1_1097 ( .A(u3_u0__abc_74260_new_n479_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n556_), .Y(u3_u0__0r3_35_0__32_));
OAI21X1 OAI21X1_1098 ( .A(u3_u0__abc_74260_new_n482_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n558_), .Y(u3_u0__0r3_35_0__33_));
OAI21X1 OAI21X1_1099 ( .A(u3_u0__abc_74260_new_n485_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n560_), .Y(u3_u0__0r3_35_0__34_));
OAI21X1 OAI21X1_11 ( .A(spec_req_cs_3_), .B(_abc_81086_new_n236_), .C(_abc_81086_new_n240_), .Y(_abc_81086_new_n253_));
OAI21X1 OAI21X1_110 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1190_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1191_));
OAI21X1 OAI21X1_1100 ( .A(u3_u0__abc_74260_new_n488_), .B(u3_u0__abc_74260_new_n491_), .C(u3_u0__abc_74260_new_n562_), .Y(u3_u0__0r3_35_0__35_));
OAI21X1 OAI21X1_1101 ( .A(u3_u0__abc_74260_new_n382_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n565_), .Y(u3_u0__0r2_35_0__0_));
OAI21X1 OAI21X1_1102 ( .A(u3_u0__abc_74260_new_n386_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n567_), .Y(u3_u0__0r2_35_0__1_));
OAI21X1 OAI21X1_1103 ( .A(u3_u0__abc_74260_new_n389_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n569_), .Y(u3_u0__0r2_35_0__2_));
OAI21X1 OAI21X1_1104 ( .A(u3_u0__abc_74260_new_n392_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n571_), .Y(u3_u0__0r2_35_0__3_));
OAI21X1 OAI21X1_1105 ( .A(u3_u0__abc_74260_new_n395_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n573_), .Y(u3_u0__0r2_35_0__4_));
OAI21X1 OAI21X1_1106 ( .A(u3_u0__abc_74260_new_n398_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n575_), .Y(u3_u0__0r2_35_0__5_));
OAI21X1 OAI21X1_1107 ( .A(u3_u0__abc_74260_new_n401_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n577_), .Y(u3_u0__0r2_35_0__6_));
OAI21X1 OAI21X1_1108 ( .A(u3_u0__abc_74260_new_n404_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n579_), .Y(u3_u0__0r2_35_0__7_));
OAI21X1 OAI21X1_1109 ( .A(u3_u0__abc_74260_new_n407_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n581_), .Y(u3_u0__0r2_35_0__8_));
OAI21X1 OAI21X1_111 ( .A(u0__abc_74894_new_n1191_), .B(u0__abc_74894_new_n1189_), .C(u0__abc_74894_new_n1193_), .Y(u0__abc_74894_new_n1194_));
OAI21X1 OAI21X1_1110 ( .A(u3_u0__abc_74260_new_n410_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n583_), .Y(u3_u0__0r2_35_0__9_));
OAI21X1 OAI21X1_1111 ( .A(u3_u0__abc_74260_new_n413_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n585_), .Y(u3_u0__0r2_35_0__10_));
OAI21X1 OAI21X1_1112 ( .A(u3_u0__abc_74260_new_n416_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n587_), .Y(u3_u0__0r2_35_0__11_));
OAI21X1 OAI21X1_1113 ( .A(u3_u0__abc_74260_new_n419_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n589_), .Y(u3_u0__0r2_35_0__12_));
OAI21X1 OAI21X1_1114 ( .A(u3_u0__abc_74260_new_n422_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n591_), .Y(u3_u0__0r2_35_0__13_));
OAI21X1 OAI21X1_1115 ( .A(u3_u0__abc_74260_new_n425_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n593_), .Y(u3_u0__0r2_35_0__14_));
OAI21X1 OAI21X1_1116 ( .A(u3_u0__abc_74260_new_n428_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n595_), .Y(u3_u0__0r2_35_0__15_));
OAI21X1 OAI21X1_1117 ( .A(u3_u0__abc_74260_new_n431_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n597_), .Y(u3_u0__0r2_35_0__16_));
OAI21X1 OAI21X1_1118 ( .A(u3_u0__abc_74260_new_n434_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n599_), .Y(u3_u0__0r2_35_0__17_));
OAI21X1 OAI21X1_1119 ( .A(u3_u0__abc_74260_new_n437_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n601_), .Y(u3_u0__0r2_35_0__18_));
OAI21X1 OAI21X1_112 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1210_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1211_));
OAI21X1 OAI21X1_1120 ( .A(u3_u0__abc_74260_new_n440_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n603_), .Y(u3_u0__0r2_35_0__19_));
OAI21X1 OAI21X1_1121 ( .A(u3_u0__abc_74260_new_n443_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n605_), .Y(u3_u0__0r2_35_0__20_));
OAI21X1 OAI21X1_1122 ( .A(u3_u0__abc_74260_new_n446_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n607_), .Y(u3_u0__0r2_35_0__21_));
OAI21X1 OAI21X1_1123 ( .A(u3_u0__abc_74260_new_n449_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n609_), .Y(u3_u0__0r2_35_0__22_));
OAI21X1 OAI21X1_1124 ( .A(u3_u0__abc_74260_new_n452_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n611_), .Y(u3_u0__0r2_35_0__23_));
OAI21X1 OAI21X1_1125 ( .A(u3_u0__abc_74260_new_n455_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n613_), .Y(u3_u0__0r2_35_0__24_));
OAI21X1 OAI21X1_1126 ( .A(u3_u0__abc_74260_new_n458_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n615_), .Y(u3_u0__0r2_35_0__25_));
OAI21X1 OAI21X1_1127 ( .A(u3_u0__abc_74260_new_n461_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n617_), .Y(u3_u0__0r2_35_0__26_));
OAI21X1 OAI21X1_1128 ( .A(u3_u0__abc_74260_new_n464_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n619_), .Y(u3_u0__0r2_35_0__27_));
OAI21X1 OAI21X1_1129 ( .A(u3_u0__abc_74260_new_n467_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n621_), .Y(u3_u0__0r2_35_0__28_));
OAI21X1 OAI21X1_113 ( .A(u0__abc_74894_new_n1211_), .B(u0__abc_74894_new_n1209_), .C(u0__abc_74894_new_n1213_), .Y(u0__abc_74894_new_n1214_));
OAI21X1 OAI21X1_1130 ( .A(u3_u0__abc_74260_new_n470_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n623_), .Y(u3_u0__0r2_35_0__29_));
OAI21X1 OAI21X1_1131 ( .A(u3_u0__abc_74260_new_n473_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n625_), .Y(u3_u0__0r2_35_0__30_));
OAI21X1 OAI21X1_1132 ( .A(u3_u0__abc_74260_new_n476_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n627_), .Y(u3_u0__0r2_35_0__31_));
OAI21X1 OAI21X1_1133 ( .A(u3_u0__abc_74260_new_n479_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n629_), .Y(u3_u0__0r2_35_0__32_));
OAI21X1 OAI21X1_1134 ( .A(u3_u0__abc_74260_new_n482_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n631_), .Y(u3_u0__0r2_35_0__33_));
OAI21X1 OAI21X1_1135 ( .A(u3_u0__abc_74260_new_n485_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n633_), .Y(u3_u0__0r2_35_0__34_));
OAI21X1 OAI21X1_1136 ( .A(u3_u0__abc_74260_new_n488_), .B(u3_u0__abc_74260_new_n564_), .C(u3_u0__abc_74260_new_n635_), .Y(u3_u0__0r2_35_0__35_));
OAI21X1 OAI21X1_1137 ( .A(u3_u0__abc_74260_new_n637_), .B(u3_re), .C(u3_u0__abc_74260_new_n638_), .Y(u3_u0__0rd_adr_3_0__0_));
OAI21X1 OAI21X1_1138 ( .A(u3_u0_rd_adr_0_), .B(u3_u0__abc_74260_new_n640_), .C(u3_u0__abc_74260_new_n642_), .Y(u3_u0__abc_74260_new_n643_));
OAI21X1 OAI21X1_1139 ( .A(u3_u0_rd_adr_1_), .B(u3_u0__abc_74260_new_n640_), .C(u3_u0__abc_74260_new_n642_), .Y(u3_u0__abc_74260_new_n646_));
OAI21X1 OAI21X1_114 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1230_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1231_));
OAI21X1 OAI21X1_1140 ( .A(u3_u0_rd_adr_2_), .B(u3_u0__abc_74260_new_n640_), .C(u3_u0__abc_74260_new_n642_), .Y(u3_u0__abc_74260_new_n649_));
OAI21X1 OAI21X1_1141 ( .A(dv), .B(u3_u0__abc_74260_new_n651_), .C(u3_u0__abc_74260_new_n652_), .Y(u3_u0__0wr_adr_3_0__0_));
OAI21X1 OAI21X1_1142 ( .A(u3_u0__abc_74260_new_n738_), .B(u3_u0__abc_74260_new_n739_), .C(u3_u0__abc_74260_new_n737_), .Y(u3_u0__abc_74260_new_n740_));
OAI21X1 OAI21X1_1143 ( .A(u4_rfr_ce), .B(u4_rfr_cnt_0_), .C(u4__abc_74770_new_n94_), .Y(u4__abc_74770_new_n95_));
OAI21X1 OAI21X1_1144 ( .A(u4_rfr_cnt_1_), .B(u4__abc_74770_new_n93_), .C(u4__abc_74770_new_n94_), .Y(u4__abc_74770_new_n99_));
OAI21X1 OAI21X1_1145 ( .A(u4_rfr_cnt_2_), .B(u4__abc_74770_new_n98_), .C(u4__abc_74770_new_n94_), .Y(u4__abc_74770_new_n104_));
OAI21X1 OAI21X1_1146 ( .A(u4_rfr_cnt_3_), .B(u4__abc_74770_new_n103_), .C(u4__abc_74770_new_n94_), .Y(u4__abc_74770_new_n108_));
OAI21X1 OAI21X1_1147 ( .A(u4_rfr_cnt_5_), .B(u4__abc_74770_new_n112_), .C(u4__abc_74770_new_n94_), .Y(u4__abc_74770_new_n115_));
OAI21X1 OAI21X1_1148 ( .A(u4__abc_74770_new_n117_), .B(u4__abc_74770_new_n118_), .C(u4__abc_74770_new_n94_), .Y(u4__abc_74770_new_n119_));
OAI21X1 OAI21X1_1149 ( .A(u4__abc_74770_new_n117_), .B(u4__abc_74770_new_n118_), .C(u4_rfr_cnt_7_), .Y(u4__abc_74770_new_n121_));
OAI21X1 OAI21X1_115 ( .A(u0__abc_74894_new_n1231_), .B(u0__abc_74894_new_n1229_), .C(u0__abc_74894_new_n1233_), .Y(u0__abc_74894_new_n1234_));
OAI21X1 OAI21X1_1150 ( .A(u4__abc_74770_new_n136_), .B(u4__abc_74770_new_n134_), .C(u4__abc_74770_new_n140_), .Y(u4__abc_74770_new_n141_));
OAI21X1 OAI21X1_1151 ( .A(u4__abc_74770_new_n157_), .B(u4__abc_74770_new_n158_), .C(u4_ps_cnt_6_), .Y(u4__abc_74770_new_n163_));
OAI21X1 OAI21X1_1152 ( .A(u4_rfr_cnt_3_), .B(u4__abc_74770_new_n174_), .C(ref_int_1_), .Y(u4__abc_74770_new_n175_));
OAI21X1 OAI21X1_1153 ( .A(u4_rfr_cnt_5_), .B(u4__abc_74770_new_n174_), .C(u4__abc_74770_new_n177_), .Y(u4__abc_74770_new_n182_));
OAI21X1 OAI21X1_1154 ( .A(u4__abc_74770_new_n123_), .B(u4__abc_74770_new_n183_), .C(u4__abc_74770_new_n182_), .Y(u4__abc_74770_new_n184_));
OAI21X1 OAI21X1_1155 ( .A(u5__abc_78290_new_n618_), .B(u5__abc_78290_new_n623_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n624_));
OAI21X1 OAI21X1_1156 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n631_), .C(u5__abc_78290_new_n639_), .Y(u5__abc_78290_new_n640_));
OAI21X1 OAI21X1_1157 ( .A(u5__abc_78290_new_n671_), .B(u5__abc_78290_new_n707_), .C(u5__abc_78290_new_n702_), .Y(u5__abc_78290_new_n708_));
OAI21X1 OAI21X1_1158 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n738_), .C(u5__abc_78290_new_n732_), .Y(u5__abc_78290_new_n739_));
OAI21X1 OAI21X1_1159 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n745_), .C(u5__abc_78290_new_n752_), .Y(u5__abc_78290_new_n753_));
OAI21X1 OAI21X1_116 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1250_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1251_));
OAI21X1 OAI21X1_1160 ( .A(u5__abc_78290_new_n756_), .B(u5__abc_78290_new_n759_), .C(u5__abc_78290_new_n767_), .Y(u5__abc_78290_new_n768_));
OAI21X1 OAI21X1_1161 ( .A(u5__abc_78290_new_n819_), .B(u5__abc_78290_new_n821_), .C(u5__abc_78290_new_n816_), .Y(u5__abc_78290_new_n822_));
OAI21X1 OAI21X1_1162 ( .A(u5__abc_78290_new_n853_), .B(u5__abc_78290_new_n860_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n861_));
OAI21X1 OAI21X1_1163 ( .A(u5__abc_78290_new_n908_), .B(u5__abc_78290_new_n915_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n916_));
OAI21X1 OAI21X1_1164 ( .A(u5__abc_78290_new_n936_), .B(u5__abc_78290_new_n928_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n937_));
OAI21X1 OAI21X1_1165 ( .A(u5__abc_78290_new_n945_), .B(u5__abc_78290_new_n952_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n953_));
OAI21X1 OAI21X1_1166 ( .A(u5__abc_78290_new_n488_), .B(u5__abc_78290_new_n498_), .C(u5__abc_78290_new_n958_), .Y(dv));
OAI21X1 OAI21X1_1167 ( .A(u5__abc_78290_new_n908_), .B(u5__abc_78290_new_n921_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n975_));
OAI21X1 OAI21X1_1168 ( .A(u5__abc_78290_new_n982_), .B(u5__abc_78290_new_n915_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n983_));
OAI21X1 OAI21X1_1169 ( .A(u5__abc_78290_new_n638_), .B(u5__abc_78290_new_n653_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n987_));
OAI21X1 OAI21X1_117 ( .A(u0__abc_74894_new_n1251_), .B(u0__abc_74894_new_n1249_), .C(u0__abc_74894_new_n1253_), .Y(u0__abc_74894_new_n1254_));
OAI21X1 OAI21X1_1170 ( .A(u5__abc_78290_new_n670_), .B(u5__abc_78290_new_n681_), .C(u5__abc_78290_new_n901_), .Y(u5__abc_78290_new_n994_));
OAI21X1 OAI21X1_1171 ( .A(u5__abc_78290_new_n974_), .B(u5__abc_78290_new_n1019_), .C(u5__abc_78290_new_n1036_), .Y(u5_rfr_ack_d));
OAI21X1 OAI21X1_1172 ( .A(u5__abc_78290_new_n1042_), .B(u5__abc_78290_new_n1038_), .C(u5__abc_78290_new_n1039_), .Y(u5__abc_78290_new_n1043_));
OAI21X1 OAI21X1_1173 ( .A(u5__abc_78290_new_n1048_), .B(u5__abc_78290_new_n1051_), .C(u5__abc_78290_new_n1045_), .Y(u5__abc_78290_new_n1052_));
OAI21X1 OAI21X1_1174 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1099_), .C(u5__abc_78290_new_n1104_), .Y(u5__abc_78290_new_n1105_));
OAI21X1 OAI21X1_1175 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1131_), .C(u5__abc_78290_new_n1128_), .Y(u5__abc_78290_new_n1132_));
OAI21X1 OAI21X1_1176 ( .A(u5__abc_78290_new_n1134_), .B(u5__abc_78290_new_n1136_), .C(u5__abc_78290_new_n1085_), .Y(u5__abc_78290_new_n1137_));
OAI21X1 OAI21X1_1177 ( .A(u5__abc_78290_new_n1142_), .B(u5__abc_78290_new_n1145_), .C(u5__abc_78290_new_n1139_), .Y(u5__abc_78290_new_n1146_));
OAI21X1 OAI21X1_1178 ( .A(u5__abc_78290_new_n440_), .B(u5__abc_78290_new_n1214_), .C(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n1215_));
OAI21X1 OAI21X1_1179 ( .A(u5__abc_78290_new_n1219_), .B(u5__abc_78290_new_n1038_), .C(u5__abc_78290_new_n1222_), .Y(u5__abc_78290_new_n1223_));
OAI21X1 OAI21X1_118 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1270_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1271_));
OAI21X1 OAI21X1_1180 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1233_), .C(u5__abc_78290_new_n1229_), .Y(u5__abc_78290_new_n1234_));
OAI21X1 OAI21X1_1181 ( .A(u5__abc_78290_new_n1249_), .B(u5__abc_78290_new_n1244_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1250_));
OAI21X1 OAI21X1_1182 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1277_), .C(u5__abc_78290_new_n1282_), .Y(u5__abc_78290_new_n1283_));
OAI21X1 OAI21X1_1183 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1287_), .C(u5__abc_78290_new_n1291_), .Y(u5__abc_78290_new_n1292_));
OAI21X1 OAI21X1_1184 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1299_), .C(u5__abc_78290_new_n1297_), .Y(u5__abc_78290_new_n1300_));
OAI21X1 OAI21X1_1185 ( .A(u1_wb_write_go), .B(u3_wb_read_go), .C(u5_lookup_ready2), .Y(u5__abc_78290_new_n1333_));
OAI21X1 OAI21X1_1186 ( .A(u5__abc_78290_new_n1336_), .B(u5__abc_78290_new_n1337_), .C(u5__abc_78290_new_n1340_), .Y(u5__abc_78290_new_n1341_));
OAI21X1 OAI21X1_1187 ( .A(u5__abc_78290_new_n1326_), .B(u5__abc_78290_new_n1346_), .C(u5__abc_78290_new_n1318_), .Y(u5__abc_78290_new_n1347_));
OAI21X1 OAI21X1_1188 ( .A(u5__abc_78290_new_n1092_), .B(u5__abc_78290_new_n1112_), .C(u5__abc_78290_new_n1085_), .Y(u5__abc_78290_new_n1350_));
OAI21X1 OAI21X1_1189 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1277_), .C(u5__abc_78290_new_n1229_), .Y(u5__abc_78290_new_n1353_));
OAI21X1 OAI21X1_119 ( .A(u0__abc_74894_new_n1271_), .B(u0__abc_74894_new_n1269_), .C(u0__abc_74894_new_n1273_), .Y(u0__abc_74894_new_n1274_));
OAI21X1 OAI21X1_1190 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1261_), .C(u5__abc_78290_new_n1291_), .Y(u5__abc_78290_new_n1356_));
OAI21X1 OAI21X1_1191 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1310_), .C(u5__abc_78290_new_n1363_), .Y(u5__abc_78290_new_n1364_));
OAI21X1 OAI21X1_1192 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1299_), .C(u5__abc_78290_new_n561_), .Y(u5__abc_78290_new_n1365_));
OAI21X1 OAI21X1_1193 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1164_), .C(u5__abc_78290_new_n1386_), .Y(u5__abc_78290_new_n1387_));
OAI21X1 OAI21X1_1194 ( .A(u5__abc_78290_new_n622_), .B(u5__abc_78290_new_n1399_), .C(u5__abc_78290_new_n1400_), .Y(u5__abc_78290_new_n1401_));
OAI21X1 OAI21X1_1195 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1287_), .C(u5__abc_78290_new_n1402_), .Y(u5__abc_78290_new_n1403_));
OAI21X1 OAI21X1_1196 ( .A(tms_s_9_), .B(u5__abc_78290_new_n1406_), .C(u5_wb_cycle), .Y(u5__abc_78290_new_n1407_));
OAI21X1 OAI21X1_1197 ( .A(tms_s_1_), .B(u5__abc_78290_new_n1405_), .C(u5__abc_78290_new_n1409_), .Y(u5__abc_78290_new_n1410_));
OAI21X1 OAI21X1_1198 ( .A(u5_cnt), .B(u5__abc_78290_new_n1410_), .C(u5__abc_78290_new_n1416_), .Y(u5__abc_78290_new_n1417_));
OAI21X1 OAI21X1_1199 ( .A(u5__abc_78290_new_n1414_), .B(u5__abc_78290_new_n1415_), .C(u5__abc_78290_new_n1417_), .Y(u5__abc_78290_new_n1418_));
OAI21X1 OAI21X1_12 ( .A(_abc_81086_new_n251_), .B(_abc_81086_new_n253_), .C(_abc_81086_new_n252_), .Y(obct_cs_3_));
OAI21X1 OAI21X1_120 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1290_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1291_));
OAI21X1 OAI21X1_1200 ( .A(u5__abc_78290_new_n1428_), .B(u5__abc_78290_new_n1429_), .C(u5__abc_78290_new_n1430_), .Y(u5_we_));
OAI21X1 OAI21X1_1201 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n1432_), .C(u5__abc_78290_new_n1434_), .Y(u5__abc_78290_new_n1435_));
OAI21X1 OAI21X1_1202 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1233_), .C(u5__abc_78290_new_n1297_), .Y(u5__abc_78290_new_n1439_));
OAI21X1 OAI21X1_1203 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1131_), .C(u5__abc_78290_new_n1441_), .Y(u5__abc_78290_new_n1442_));
OAI21X1 OAI21X1_1204 ( .A(u5__abc_78290_new_n1446_), .B(u5__abc_78290_new_n1408_), .C(u5__abc_78290_new_n1374_), .Y(u5__abc_78290_new_n1447_));
OAI21X1 OAI21X1_1205 ( .A(u5__abc_78290_new_n1449_), .B(u5__abc_78290_new_n1435_), .C(u5__abc_78290_new_n1429_), .Y(u5__abc_78290_new_n1452_));
OAI21X1 OAI21X1_1206 ( .A(u5__abc_78290_new_n1429_), .B(u5__abc_78290_new_n1451_), .C(u5__abc_78290_new_n1452_), .Y(cas_));
OAI21X1 OAI21X1_1207 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1233_), .C(u5__abc_78290_new_n1402_), .Y(u5__abc_78290_new_n1454_));
OAI21X1 OAI21X1_1208 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1272_), .C(u5__abc_78290_new_n1458_), .Y(u5__abc_78290_new_n1459_));
OAI21X1 OAI21X1_1209 ( .A(u5__abc_78290_new_n1455_), .B(u5__abc_78290_new_n1457_), .C(u5__abc_78290_new_n1460_), .Y(u5__abc_78290_new_n1461_));
OAI21X1 OAI21X1_121 ( .A(u0__abc_74894_new_n1291_), .B(u0__abc_74894_new_n1289_), .C(u0__abc_74894_new_n1293_), .Y(u0__abc_74894_new_n1294_));
OAI21X1 OAI21X1_1210 ( .A(u5__abc_78290_new_n1463_), .B(u5__abc_78290_new_n1435_), .C(u5__abc_78290_new_n1429_), .Y(u5__abc_78290_new_n1466_));
OAI21X1 OAI21X1_1211 ( .A(u5__abc_78290_new_n1429_), .B(u5__abc_78290_new_n1465_), .C(u5__abc_78290_new_n1466_), .Y(ras_));
OAI21X1 OAI21X1_1212 ( .A(u5__abc_78290_new_n1481_), .B(u5__abc_78290_new_n1323_), .C(u5__abc_78290_new_n1482_), .Y(u5__abc_78290_new_n1483_));
OAI21X1 OAI21X1_1213 ( .A(u5__abc_78290_new_n1374_), .B(u5__abc_78290_new_n1490_), .C(u5__abc_78290_new_n1492_), .Y(u5__abc_78290_new_n1493_));
OAI21X1 OAI21X1_1214 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1256_), .C(u5__abc_78290_new_n1267_), .Y(u5__abc_78290_new_n1496_));
OAI21X1 OAI21X1_1215 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n1495_), .C(u5__abc_78290_new_n1497_), .Y(u5__abc_78290_new_n1498_));
OAI21X1 OAI21X1_1216 ( .A(u5__abc_78290_new_n1418_), .B(u5__abc_78290_new_n1500_), .C(u5__abc_78290_new_n1407_), .Y(u5__abc_78290_new_n1501_));
OAI21X1 OAI21X1_1217 ( .A(u1_wr_cycle), .B(u5__abc_78290_new_n1508_), .C(u5__abc_78290_new_n1510_), .Y(cs_en));
OAI21X1 OAI21X1_1218 ( .A(csc_s_2_), .B(csc_s_1_), .C(u5__abc_78290_new_n1513_), .Y(u5__abc_78290_new_n1514_));
OAI21X1 OAI21X1_1219 ( .A(u5__abc_78290_new_n1262_), .B(u5__abc_78290_new_n1517_), .C(u5__abc_78290_new_n1325_), .Y(u5__abc_78290_new_n1518_));
OAI21X1 OAI21X1_122 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1310_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1311_));
OAI21X1 OAI21X1_1220 ( .A(u5__abc_78290_new_n1400_), .B(u5__abc_78290_new_n1476_), .C(u5__abc_78290_new_n1520_), .Y(u5_data_oe_d));
OAI21X1 OAI21X1_1221 ( .A(u5__abc_78290_new_n1429_), .B(u5__abc_78290_new_n1522_), .C(u5__abc_78290_new_n1523_), .Y(u5__0data_oe_0_0_));
OAI21X1 OAI21X1_1222 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1160_), .C(u5__abc_78290_new_n1386_), .Y(u5__abc_78290_new_n1527_));
OAI21X1 OAI21X1_1223 ( .A(u5__abc_78290_new_n1242_), .B(u5__abc_78290_new_n545_), .C(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n1533_));
OAI21X1 OAI21X1_1224 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1541_), .C(u5__abc_78290_new_n1374_), .Y(u5__abc_78290_new_n1542_));
OAI21X1 OAI21X1_1225 ( .A(u5__abc_78290_new_n1198_), .B(u5__abc_78290_new_n1189_), .C(u5__abc_78290_new_n1188_), .Y(u5__abc_78290_new_n1544_));
OAI21X1 OAI21X1_1226 ( .A(u5__abc_78290_new_n570_), .B(u5__abc_78290_new_n1013_), .C(u5__abc_78290_new_n1193_), .Y(u5__abc_78290_new_n1546_));
OAI21X1 OAI21X1_1227 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1219_), .C(u5__abc_78290_new_n484_), .Y(u5__abc_78290_new_n1559_));
OAI21X1 OAI21X1_1228 ( .A(u5__abc_78290_new_n1233_), .B(u5__abc_78290_new_n1053_), .C(u5__abc_78290_new_n1222_), .Y(u5__abc_78290_new_n1560_));
OAI21X1 OAI21X1_1229 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1261_), .C(u5__abc_78290_new_n1267_), .Y(u5__abc_78290_new_n1572_));
OAI21X1 OAI21X1_123 ( .A(u0__abc_74894_new_n1311_), .B(u0__abc_74894_new_n1309_), .C(u0__abc_74894_new_n1313_), .Y(u0__abc_74894_new_n1314_));
OAI21X1 OAI21X1_1230 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1228_), .C(u5__abc_78290_new_n1282_), .Y(u5__abc_78290_new_n1574_));
OAI21X1 OAI21X1_1231 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n782_), .C(u5_kro), .Y(u5__abc_78290_new_n1587_));
OAI21X1 OAI21X1_1232 ( .A(u5__abc_78290_new_n1598_), .B(u5__abc_78290_new_n1599_), .C(u5__abc_78290_new_n1603_), .Y(u5__abc_78290_new_n1604_));
OAI21X1 OAI21X1_1233 ( .A(u5__abc_78290_new_n1608_), .B(u5__abc_78290_new_n1471_), .C(u5__0burst_act_rd_0_0_), .Y(u5__abc_78290_new_n1609_));
OAI21X1 OAI21X1_1234 ( .A(u5__abc_78290_new_n1433_), .B(u5__abc_78290_new_n1616_), .C(u5_tmr_done), .Y(u5__abc_78290_new_n1617_));
OAI21X1 OAI21X1_1235 ( .A(u5__abc_78290_new_n1104_), .B(u5__abc_78290_new_n1612_), .C(u5__abc_78290_new_n1622_), .Y(u5__abc_78290_new_n1623_));
OAI21X1 OAI21X1_1236 ( .A(u5__abc_78290_new_n1614_), .B(u5__abc_78290_new_n1609_), .C(u5__abc_78290_new_n1625_), .Y(u5__abc_78290_new_n1626_));
OAI21X1 OAI21X1_1237 ( .A(u5__abc_78290_new_n1631_), .B(u5__abc_78290_new_n1478_), .C(u5__abc_78290_new_n1634_), .Y(u5__0ap_en_0_0_));
OAI21X1 OAI21X1_1238 ( .A(u5__abc_78290_new_n1135_), .B(u5__abc_78290_new_n1399_), .C(u5__abc_78290_new_n1297_), .Y(u5__abc_78290_new_n1636_));
OAI21X1 OAI21X1_1239 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1127_), .C(u5__abc_78290_new_n1639_), .Y(u5__abc_78290_new_n1640_));
OAI21X1 OAI21X1_124 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1330_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1331_));
OAI21X1 OAI21X1_1240 ( .A(u5__abc_78290_new_n1650_), .B(u5__abc_78290_new_n1651_), .C(u5__abc_78290_new_n1632_), .Y(u5__abc_78290_new_n1652_));
OAI21X1 OAI21X1_1241 ( .A(tms_s_2_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n1652_), .Y(u5__abc_78290_new_n1653_));
OAI21X1 OAI21X1_1242 ( .A(u5__abc_78290_new_n1657_), .B(u5__abc_78290_new_n1655_), .C(u5__abc_78290_new_n1478_), .Y(u5__abc_78290_new_n1658_));
OAI21X1 OAI21X1_1243 ( .A(u5__abc_78290_new_n1607_), .B(u5__abc_78290_new_n1626_), .C(u1_wr_cycle), .Y(u5__abc_78290_new_n1665_));
OAI21X1 OAI21X1_1244 ( .A(u5__abc_78290_new_n1667_), .B(u5__abc_78290_new_n1669_), .C(u5__abc_78290_new_n1317_), .Y(u5__abc_78290_new_n1670_));
OAI21X1 OAI21X1_1245 ( .A(u5_burst_cnt_0_), .B(u5__abc_78290_new_n1666_), .C(u5_burst_cnt_1_), .Y(u5__abc_78290_new_n1672_));
OAI21X1 OAI21X1_1246 ( .A(u5__abc_78290_new_n1658_), .B(u5__abc_78290_new_n1676_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1677_));
OAI21X1 OAI21X1_1247 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n1661_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1682_));
OAI21X1 OAI21X1_1248 ( .A(u5__abc_78290_new_n1318_), .B(u5__abc_78290_new_n1681_), .C(u5__abc_78290_new_n1683_), .Y(u5__0burst_cnt_10_0__2_));
OAI21X1 OAI21X1_1249 ( .A(u5__abc_78290_new_n368_), .B(u5__abc_78290_new_n1666_), .C(u5_burst_cnt_3_), .Y(u5__abc_78290_new_n1685_));
OAI21X1 OAI21X1_125 ( .A(u0__abc_74894_new_n1331_), .B(u0__abc_74894_new_n1329_), .C(u0__abc_74894_new_n1333_), .Y(u0__abc_74894_new_n1334_));
OAI21X1 OAI21X1_1250 ( .A(u5__abc_78290_new_n1687_), .B(u5__abc_78290_new_n1660_), .C(u5__abc_78290_new_n1688_), .Y(u5__abc_78290_new_n1689_));
OAI21X1 OAI21X1_1251 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n1689_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1690_));
OAI21X1 OAI21X1_1252 ( .A(u5__abc_78290_new_n1693_), .B(u5__abc_78290_new_n1695_), .C(u5__abc_78290_new_n1317_), .Y(u5__abc_78290_new_n1696_));
OAI21X1 OAI21X1_1253 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n1702_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1703_));
OAI21X1 OAI21X1_1254 ( .A(u5_burst_cnt_5_), .B(u5__abc_78290_new_n1694_), .C(u5_burst_cnt_6_), .Y(u5__abc_78290_new_n1705_));
OAI21X1 OAI21X1_1255 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n1708_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1709_));
OAI21X1 OAI21X1_1256 ( .A(u5__abc_78290_new_n1720_), .B(u5__abc_78290_new_n1722_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1723_));
OAI21X1 OAI21X1_1257 ( .A(u5__abc_78290_new_n1731_), .B(u5__abc_78290_new_n1729_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1732_));
OAI21X1 OAI21X1_1258 ( .A(u5__abc_78290_new_n1741_), .B(u5__abc_78290_new_n1737_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1742_));
OAI21X1 OAI21X1_1259 ( .A(u5__abc_78290_new_n1747_), .B(u5__abc_78290_new_n1752_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1753_));
OAI21X1 OAI21X1_126 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1350_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1351_));
OAI21X1 OAI21X1_1260 ( .A(u5__abc_78290_new_n1756_), .B(u5__abc_78290_new_n1759_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1760_));
OAI21X1 OAI21X1_1261 ( .A(u5__abc_78290_new_n1786_), .B(u5__abc_78290_new_n1776_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1787_));
OAI21X1 OAI21X1_1262 ( .A(u5__abc_78290_new_n1794_), .B(u5__abc_78290_new_n1790_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1795_));
OAI21X1 OAI21X1_1263 ( .A(u5__abc_78290_new_n1816_), .B(u5__abc_78290_new_n1819_), .C(u5__abc_78290_new_n478_), .Y(u5__abc_78290_new_n1820_));
OAI21X1 OAI21X1_1264 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n1824_), .C(u5__abc_78290_new_n1828_), .Y(u5__abc_78290_new_n1829_));
OAI21X1 OAI21X1_1265 ( .A(u5__abc_78290_new_n1829_), .B(u5__abc_78290_new_n1821_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1830_));
OAI21X1 OAI21X1_1266 ( .A(u5__abc_78290_new_n1838_), .B(u5__abc_78290_new_n1842_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1843_));
OAI21X1 OAI21X1_1267 ( .A(u5__abc_78290_new_n1847_), .B(u5__abc_78290_new_n1851_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1852_));
OAI21X1 OAI21X1_1268 ( .A(u5__abc_78290_new_n1856_), .B(u5__abc_78290_new_n1858_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1859_));
OAI21X1 OAI21X1_1269 ( .A(u5__abc_78290_new_n491_), .B(u5__abc_78290_new_n1865_), .C(u5__abc_78290_new_n1859_), .Y(u5__abc_78290_new_n1866_));
OAI21X1 OAI21X1_127 ( .A(u0__abc_74894_new_n1351_), .B(u0__abc_74894_new_n1349_), .C(u0__abc_74894_new_n1353_), .Y(u0__abc_74894_new_n1354_));
OAI21X1 OAI21X1_1270 ( .A(u5__abc_78290_new_n1875_), .B(u5__abc_78290_new_n1872_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1876_));
OAI21X1 OAI21X1_1271 ( .A(u5__abc_78290_new_n1886_), .B(u5__abc_78290_new_n1883_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1887_));
OAI21X1 OAI21X1_1272 ( .A(u5__abc_78290_new_n839_), .B(u5__abc_78290_new_n876_), .C(u5__abc_78290_new_n838_), .Y(u5__abc_78290_new_n1890_));
OAI21X1 OAI21X1_1273 ( .A(u5__abc_78290_new_n1895_), .B(u5__abc_78290_new_n1891_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1896_));
OAI21X1 OAI21X1_1274 ( .A(u5__abc_78290_new_n1912_), .B(u5__abc_78290_new_n1908_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1913_));
OAI21X1 OAI21X1_1275 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n1929_), .C(u5__abc_78290_new_n1926_), .Y(u5__abc_78290_new_n1930_));
OAI21X1 OAI21X1_1276 ( .A(u5__abc_78290_new_n1937_), .B(u5__abc_78290_new_n1930_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1938_));
OAI21X1 OAI21X1_1277 ( .A(u5__abc_78290_new_n1946_), .B(u5__abc_78290_new_n1942_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n1947_));
OAI21X1 OAI21X1_1278 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n1956_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1957_));
OAI21X1 OAI21X1_1279 ( .A(u5__abc_78290_new_n372_), .B(u5__abc_78290_new_n1959_), .C(u5_burst_cnt_8_), .Y(u5__abc_78290_new_n1960_));
OAI21X1 OAI21X1_128 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1370_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1371_));
OAI21X1 OAI21X1_1280 ( .A(u5__abc_78290_new_n1952_), .B(u5__abc_78290_new_n1964_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1965_));
OAI21X1 OAI21X1_1281 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n1972_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1973_));
OAI21X1 OAI21X1_1282 ( .A(u5__abc_78290_new_n1666_), .B(u5__abc_78290_new_n1976_), .C(u5__abc_78290_new_n1977_), .Y(u5__abc_78290_new_n1978_));
OAI21X1 OAI21X1_1283 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n1979_), .C(u5__abc_78290_new_n1648_), .Y(u5__abc_78290_new_n1980_));
OAI21X1 OAI21X1_1284 ( .A(u5_ir_cnt_1_), .B(u5__abc_78290_new_n2003_), .C(u5__abc_78290_new_n2013_), .Y(u5__0ir_cnt_3_0__1_));
OAI21X1 OAI21X1_1285 ( .A(u5__abc_78290_new_n2017_), .B(u5__abc_78290_new_n2016_), .C(u5__abc_78290_new_n2010_), .Y(u5__abc_78290_new_n2018_));
OAI21X1 OAI21X1_1286 ( .A(u5__abc_78290_new_n560_), .B(u5__abc_78290_new_n1304_), .C(u5__abc_78290_new_n480_), .Y(u5__abc_78290_new_n2025_));
OAI21X1 OAI21X1_1287 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n834_), .C(u5__abc_78290_new_n2047_), .Y(u5__abc_78290_new_n2048_));
OAI21X1 OAI21X1_1288 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n828_), .C(u5__abc_78290_new_n895_), .Y(u5__abc_78290_new_n2049_));
OAI21X1 OAI21X1_1289 ( .A(u5__abc_78290_new_n1013_), .B(u5__abc_78290_new_n570_), .C(u5__abc_78290_new_n600_), .Y(u5__abc_78290_new_n2063_));
OAI21X1 OAI21X1_129 ( .A(u0__abc_74894_new_n1371_), .B(u0__abc_74894_new_n1369_), .C(u0__abc_74894_new_n1373_), .Y(u0__abc_74894_new_n1374_));
OAI21X1 OAI21X1_1290 ( .A(u5__abc_78290_new_n578_), .B(u5__abc_78290_new_n570_), .C(u5__abc_78290_new_n569_), .Y(u5__abc_78290_new_n2065_));
OAI21X1 OAI21X1_1291 ( .A(u5_timer_7_), .B(u5__abc_78290_new_n967_), .C(u5__0mc_le_0_0_), .Y(u5__abc_78290_new_n2083_));
OAI21X1 OAI21X1_1292 ( .A(u5__abc_78290_new_n1950_), .B(u5__abc_78290_new_n2082_), .C(u5__abc_78290_new_n2086_), .Y(u5__abc_78290_new_n2087_));
OAI21X1 OAI21X1_1293 ( .A(u5__abc_78290_new_n1768_), .B(u5__abc_78290_new_n1776_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n2088_));
OAI21X1 OAI21X1_1294 ( .A(u5__abc_78290_new_n1786_), .B(u5__abc_78290_new_n1801_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n2089_));
OAI21X1 OAI21X1_1295 ( .A(u5__abc_78290_new_n491_), .B(u5__abc_78290_new_n1820_), .C(u5__abc_78290_new_n1812_), .Y(u5__abc_78290_new_n2093_));
OAI21X1 OAI21X1_1296 ( .A(u5__abc_78290_new_n1722_), .B(u5__abc_78290_new_n1244_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n2107_));
OAI21X1 OAI21X1_1297 ( .A(u5__abc_78290_new_n1741_), .B(u5__abc_78290_new_n1731_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n2116_));
OAI21X1 OAI21X1_1298 ( .A(u5__abc_78290_new_n1747_), .B(u5__abc_78290_new_n1756_), .C(u5__abc_78290_new_n428_), .Y(u5__abc_78290_new_n2117_));
OAI21X1 OAI21X1_1299 ( .A(u5__abc_78290_new_n491_), .B(u5__abc_78290_new_n2119_), .C(u5__abc_78290_new_n2096_), .Y(u5__abc_78290_new_n2120_));
OAI21X1 OAI21X1_13 ( .A(susp_sel), .B(rfr_ack), .C(cs_need_rfr_4_), .Y(_abc_81086_new_n256_));
OAI21X1 OAI21X1_130 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1390_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1391_));
OAI21X1 OAI21X1_1300 ( .A(u5__abc_78290_new_n2111_), .B(u5__abc_78290_new_n2087_), .C(u5__abc_78290_new_n2125_), .Y(u5__abc_78290_new_n2126_));
OAI21X1 OAI21X1_1301 ( .A(tms_s_24_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2124_), .Y(u5__abc_78290_new_n2127_));
OAI21X1 OAI21X1_1302 ( .A(tms_s_17_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2130_), .Y(u5__abc_78290_new_n2131_));
OAI21X1 OAI21X1_1303 ( .A(u5__abc_78290_new_n2134_), .B(u5__abc_78290_new_n2034_), .C(u5__abc_78290_new_n2141_), .Y(u5__abc_78290_new_n2142_));
OAI21X1 OAI21X1_1304 ( .A(u5__abc_78290_new_n2133_), .B(u5__abc_78290_new_n2145_), .C(u5__abc_78290_new_n2140_), .Y(u5__abc_78290_new_n2146_));
OAI21X1 OAI21X1_1305 ( .A(u5__abc_78290_new_n1320_), .B(u5__abc_78290_new_n1319_), .C(u5__abc_78290_new_n1513_), .Y(u5__abc_78290_new_n2148_));
OAI21X1 OAI21X1_1306 ( .A(u5__abc_78290_new_n853_), .B(u5__abc_78290_new_n844_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n2153_));
OAI21X1 OAI21X1_1307 ( .A(u5__abc_78290_new_n1019_), .B(u5__abc_78290_new_n2150_), .C(u5__abc_78290_new_n2164_), .Y(u5__abc_78290_new_n2165_));
OAI21X1 OAI21X1_1308 ( .A(u5__abc_78290_new_n2146_), .B(u5__abc_78290_new_n2144_), .C(u5__abc_78290_new_n2165_), .Y(u5__abc_78290_new_n2166_));
OAI21X1 OAI21X1_1309 ( .A(u5__abc_78290_new_n1206_), .B(u5__abc_78290_new_n1198_), .C(u5__abc_78290_new_n1188_), .Y(u5__abc_78290_new_n2170_));
OAI21X1 OAI21X1_131 ( .A(u0__abc_74894_new_n1391_), .B(u0__abc_74894_new_n1389_), .C(u0__abc_74894_new_n1393_), .Y(u0__abc_74894_new_n1394_));
OAI21X1 OAI21X1_1310 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1042_), .C(u5__abc_78290_new_n1615_), .Y(u5__abc_78290_new_n2183_));
OAI21X1 OAI21X1_1311 ( .A(u5__abc_78290_new_n1317_), .B(u5__abc_78290_new_n2150_), .C(u5__abc_78290_new_n2187_), .Y(u5__abc_78290_new_n2188_));
OAI21X1 OAI21X1_1312 ( .A(u5__abc_78290_new_n839_), .B(u5__abc_78290_new_n876_), .C(u5__abc_78290_new_n838_), .Y(u5__abc_78290_new_n2195_));
OAI21X1 OAI21X1_1313 ( .A(u5__abc_78290_new_n2166_), .B(u5__abc_78290_new_n2143_), .C(u5__abc_78290_new_n2212_), .Y(u5__abc_78290_new_n2213_));
OAI21X1 OAI21X1_1314 ( .A(u5__abc_78290_new_n2215_), .B(u5__abc_78290_new_n2222_), .C(u5__abc_78290_new_n2210_), .Y(u5__abc_78290_new_n2224_));
OAI21X1 OAI21X1_1315 ( .A(u5__abc_78290_new_n2226_), .B(u5__abc_78290_new_n2223_), .C(u5__abc_78290_new_n2224_), .Y(u5__abc_78290_new_n2227_));
OAI21X1 OAI21X1_1316 ( .A(u5_timer_0_), .B(u5__abc_78290_new_n2083_), .C(u5_timer_1_), .Y(u5__abc_78290_new_n2233_));
OAI21X1 OAI21X1_1317 ( .A(u5__abc_78290_new_n1950_), .B(u5__abc_78290_new_n2082_), .C(u5__abc_78290_new_n2236_), .Y(u5__abc_78290_new_n2237_));
OAI21X1 OAI21X1_1318 ( .A(u5__abc_78290_new_n2111_), .B(u5__abc_78290_new_n2237_), .C(u5__abc_78290_new_n2125_), .Y(u5__abc_78290_new_n2238_));
OAI21X1 OAI21X1_1319 ( .A(tms_s_25_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2124_), .Y(u5__abc_78290_new_n2239_));
OAI21X1 OAI21X1_132 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1410_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1411_));
OAI21X1 OAI21X1_1320 ( .A(tms_s_18_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2130_), .Y(u5__abc_78290_new_n2242_));
OAI21X1 OAI21X1_1321 ( .A(u5__abc_78290_new_n2245_), .B(u5__abc_78290_new_n2034_), .C(u5__abc_78290_new_n2141_), .Y(u5__abc_78290_new_n2246_));
OAI21X1 OAI21X1_1322 ( .A(u5__abc_78290_new_n2249_), .B(u5__abc_78290_new_n2250_), .C(u5__abc_78290_new_n1632_), .Y(u5__abc_78290_new_n2251_));
OAI21X1 OAI21X1_1323 ( .A(u5__abc_78290_new_n2248_), .B(u5__abc_78290_new_n2252_), .C(u5__abc_78290_new_n2253_), .Y(u5__abc_78290_new_n2254_));
OAI21X1 OAI21X1_1324 ( .A(u5__abc_78290_new_n2255_), .B(u5__abc_78290_new_n2247_), .C(u5__abc_78290_new_n2257_), .Y(u5__abc_78290_new_n2258_));
OAI21X1 OAI21X1_1325 ( .A(u5__abc_78290_new_n2260_), .B(u5__abc_78290_new_n2223_), .C(u5__abc_78290_new_n2224_), .Y(u5__abc_78290_new_n2261_));
OAI21X1 OAI21X1_1326 ( .A(u5__abc_78290_new_n2269_), .B(u5__abc_78290_new_n2266_), .C(u5__abc_78290_new_n2267_), .Y(u5__abc_78290_new_n2270_));
OAI21X1 OAI21X1_1327 ( .A(u5__abc_78290_new_n2264_), .B(u5__abc_78290_new_n2272_), .C(u5__abc_78290_new_n2140_), .Y(u5__abc_78290_new_n2273_));
OAI21X1 OAI21X1_1328 ( .A(u5__abc_78290_new_n2147_), .B(u5__abc_78290_new_n2149_), .C(u5__abc_78290_new_n1478_), .Y(u5__abc_78290_new_n2274_));
OAI21X1 OAI21X1_1329 ( .A(tms_s_26_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2124_), .Y(u5__abc_78290_new_n2292_));
OAI21X1 OAI21X1_133 ( .A(u0__abc_74894_new_n1411_), .B(u0__abc_74894_new_n1409_), .C(u0__abc_74894_new_n1413_), .Y(u0__abc_74894_new_n1414_));
OAI21X1 OAI21X1_1330 ( .A(u5__abc_78290_new_n1950_), .B(u5__abc_78290_new_n2082_), .C(u5__abc_78290_new_n2294_), .Y(u5__abc_78290_new_n2295_));
OAI21X1 OAI21X1_1331 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n2039_), .C(u5__abc_78290_new_n2075_), .Y(u5__abc_78290_new_n2297_));
OAI21X1 OAI21X1_1332 ( .A(u5__abc_78290_new_n2297_), .B(u5__abc_78290_new_n2296_), .C(u5__abc_78290_new_n2275_), .Y(u5__abc_78290_new_n2298_));
OAI21X1 OAI21X1_1333 ( .A(u5__abc_78290_new_n2271_), .B(u5__abc_78290_new_n2273_), .C(u5__abc_78290_new_n2300_), .Y(u5__abc_78290_new_n2301_));
OAI21X1 OAI21X1_1334 ( .A(u5__abc_78290_new_n2264_), .B(u5__abc_78290_new_n2272_), .C(u5__abc_78290_new_n2310_), .Y(u5__abc_78290_new_n2311_));
OAI21X1 OAI21X1_1335 ( .A(tms_s_27_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2124_), .Y(u5__abc_78290_new_n2313_));
OAI21X1 OAI21X1_1336 ( .A(u5_timer_2_), .B(u5__abc_78290_new_n2235_), .C(u5_timer_3_), .Y(u5__abc_78290_new_n2315_));
OAI21X1 OAI21X1_1337 ( .A(u5__abc_78290_new_n2314_), .B(u5__abc_78290_new_n2083_), .C(u5__abc_78290_new_n2315_), .Y(u5__abc_78290_new_n2316_));
OAI21X1 OAI21X1_1338 ( .A(u5__abc_78290_new_n1950_), .B(u5__abc_78290_new_n2082_), .C(u5__abc_78290_new_n2316_), .Y(u5__abc_78290_new_n2317_));
OAI21X1 OAI21X1_1339 ( .A(u5__abc_78290_new_n2124_), .B(u5__abc_78290_new_n2318_), .C(u5__abc_78290_new_n2313_), .Y(u5__abc_78290_new_n2319_));
OAI21X1 OAI21X1_134 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1430_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1431_));
OAI21X1 OAI21X1_1340 ( .A(u5__abc_78290_new_n2140_), .B(u5__abc_78290_new_n2321_), .C(u5__abc_78290_new_n2165_), .Y(u5__abc_78290_new_n2322_));
OAI21X1 OAI21X1_1341 ( .A(u5__abc_78290_new_n2322_), .B(u5__abc_78290_new_n2312_), .C(u5__abc_78290_new_n2324_), .Y(u5__abc_78290_new_n2325_));
OAI21X1 OAI21X1_1342 ( .A(u5__abc_78290_new_n1950_), .B(u5__abc_78290_new_n2082_), .C(u5__abc_78290_new_n2333_), .Y(u5__abc_78290_new_n2334_));
OAI21X1 OAI21X1_1343 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n2044_), .C(u5__abc_78290_new_n2040_), .Y(u5__abc_78290_new_n2337_));
OAI21X1 OAI21X1_1344 ( .A(u5__abc_78290_new_n2314_), .B(u5__abc_78290_new_n2083_), .C(u5_timer_4_), .Y(u5__abc_78290_new_n2343_));
OAI21X1 OAI21X1_1345 ( .A(tms_s_4_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2189_), .Y(u5__abc_78290_new_n2346_));
OAI21X1 OAI21X1_1346 ( .A(u5__abc_78290_new_n2348_), .B(u5__abc_78290_new_n2349_), .C(u5__abc_78290_new_n2350_), .Y(u5__abc_78290_new_n2351_));
OAI21X1 OAI21X1_1347 ( .A(u5__abc_78290_new_n2188_), .B(u5__abc_78290_new_n2353_), .C(u5__abc_78290_new_n2352_), .Y(u5__abc_78290_new_n2354_));
OAI21X1 OAI21X1_1348 ( .A(u5__abc_78290_new_n961_), .B(u5__abc_78290_new_n2348_), .C(u5__abc_78290_new_n2357_), .Y(u5__abc_78290_new_n2358_));
OAI21X1 OAI21X1_1349 ( .A(u5__abc_78290_new_n2188_), .B(u5__abc_78290_new_n2360_), .C(u5__abc_78290_new_n2352_), .Y(u5__abc_78290_new_n2361_));
OAI21X1 OAI21X1_135 ( .A(u0__abc_74894_new_n1431_), .B(u0__abc_74894_new_n1429_), .C(u0__abc_74894_new_n1433_), .Y(u0__abc_74894_new_n1434_));
OAI21X1 OAI21X1_1350 ( .A(u5__abc_78290_new_n2188_), .B(u5__abc_78290_new_n2364_), .C(u5__abc_78290_new_n2352_), .Y(u5__abc_78290_new_n2365_));
OAI21X1 OAI21X1_1351 ( .A(tms_s_16_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2367_), .Y(u5__abc_78290_new_n2368_));
OAI21X1 OAI21X1_1352 ( .A(u5__abc_78290_new_n535_), .B(u5__abc_78290_new_n623_), .C(u5__abc_78290_new_n455_), .Y(u5__abc_78290_new_n2375_));
OAI21X1 OAI21X1_1353 ( .A(u5__abc_78290_new_n2388_), .B(u5__abc_78290_new_n2390_), .C(u5__abc_78290_new_n1567_), .Y(u5__abc_78290_new_n2391_));
OAI21X1 OAI21X1_1354 ( .A(u5__abc_78290_new_n2134_), .B(u5__abc_78290_new_n2380_), .C(u5__abc_78290_new_n2415_), .Y(u5__abc_78290_new_n2416_));
OAI21X1 OAI21X1_1355 ( .A(csc_s_3_), .B(u5__abc_78290_new_n1480_), .C(u5__abc_78290_new_n1478_), .Y(u5__abc_78290_new_n2426_));
OAI21X1 OAI21X1_1356 ( .A(u5__abc_78290_new_n2427_), .B(u5__abc_78290_new_n2428_), .C(u5__abc_78290_new_n2425_), .Y(u5__abc_78290_new_n2429_));
OAI21X1 OAI21X1_1357 ( .A(u5__abc_78290_new_n2424_), .B(u5__abc_78290_new_n2422_), .C(u5__abc_78290_new_n2430_), .Y(u5__abc_78290_new_n2431_));
OAI21X1 OAI21X1_1358 ( .A(u5__abc_78290_new_n2431_), .B(u5__abc_78290_new_n2423_), .C(u5__abc_78290_new_n2368_), .Y(u5__0timer2_8_0__0_));
OAI21X1 OAI21X1_1359 ( .A(tms_s_0_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2450_), .Y(u5__abc_78290_new_n2451_));
OAI21X1 OAI21X1_136 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1450_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1451_));
OAI21X1 OAI21X1_1360 ( .A(u5__abc_78290_new_n2379_), .B(u5__abc_78290_new_n2455_), .C(u5__abc_78290_new_n2456_), .Y(u5__abc_78290_new_n2457_));
OAI21X1 OAI21X1_1361 ( .A(u5__abc_78290_new_n2461_), .B(u5__abc_78290_new_n2422_), .C(u5__abc_78290_new_n2430_), .Y(u5__abc_78290_new_n2462_));
OAI21X1 OAI21X1_1362 ( .A(tms_s_1_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2450_), .Y(u5__abc_78290_new_n2469_));
OAI21X1 OAI21X1_1363 ( .A(u5_timer2_1_), .B(u5_timer2_0_), .C(u5_timer2_2_), .Y(u5__abc_78290_new_n2470_));
OAI21X1 OAI21X1_1364 ( .A(u5__abc_78290_new_n2466_), .B(u5__abc_78290_new_n2474_), .C(u5__abc_78290_new_n2465_), .Y(u5__abc_78290_new_n2475_));
OAI21X1 OAI21X1_1365 ( .A(u5__abc_78290_new_n2478_), .B(u5__abc_78290_new_n2429_), .C(u5__abc_78290_new_n2480_), .Y(u5__abc_78290_new_n2481_));
OAI21X1 OAI21X1_1366 ( .A(tms_s_19_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2367_), .Y(u5__abc_78290_new_n2483_));
OAI21X1 OAI21X1_1367 ( .A(u5__abc_78290_new_n2484_), .B(u5__abc_78290_new_n2422_), .C(u5__abc_78290_new_n2430_), .Y(u5__abc_78290_new_n2485_));
OAI21X1 OAI21X1_1368 ( .A(tms_s_2_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2450_), .Y(u5__abc_78290_new_n2486_));
OAI21X1 OAI21X1_1369 ( .A(u5_timer2_2_), .B(u5__abc_78290_new_n2397_), .C(u5_timer2_3_), .Y(u5__abc_78290_new_n2488_));
OAI21X1 OAI21X1_137 ( .A(u0__abc_74894_new_n1451_), .B(u0__abc_74894_new_n1449_), .C(u0__abc_74894_new_n1453_), .Y(u0__abc_74894_new_n1454_));
OAI21X1 OAI21X1_1370 ( .A(u5__abc_78290_new_n2464_), .B(u5__abc_78290_new_n2465_), .C(u5__abc_78290_new_n2422_), .Y(u5__abc_78290_new_n2494_));
OAI21X1 OAI21X1_1371 ( .A(u5__abc_78290_new_n2485_), .B(u5__abc_78290_new_n2495_), .C(u5__abc_78290_new_n2483_), .Y(u5__0timer2_8_0__3_));
OAI21X1 OAI21X1_1372 ( .A(tms_s_11_), .B(u5__abc_78290_new_n1471_), .C(u5__abc_78290_new_n2497_), .Y(u5__abc_78290_new_n2498_));
OAI21X1 OAI21X1_1373 ( .A(u5__abc_78290_new_n2402_), .B(u5__abc_78290_new_n2501_), .C(u5__abc_78290_new_n2407_), .Y(u5__abc_78290_new_n2502_));
OAI21X1 OAI21X1_1374 ( .A(u5__abc_78290_new_n2499_), .B(u5__abc_78290_new_n2500_), .C(u5__abc_78290_new_n2503_), .Y(u5__abc_78290_new_n2504_));
OAI21X1 OAI21X1_1375 ( .A(u5__abc_78290_new_n2511_), .B(u5__abc_78290_new_n2512_), .C(u5__abc_78290_new_n2407_), .Y(u5__abc_78290_new_n2513_));
OAI21X1 OAI21X1_1376 ( .A(u5_timer2_5_), .B(u5__abc_78290_new_n2401_), .C(u5_timer2_6_), .Y(u5__abc_78290_new_n2520_));
OAI21X1 OAI21X1_1377 ( .A(u5__abc_78290_new_n2413_), .B(u5__abc_78290_new_n2521_), .C(u5__abc_78290_new_n2522_), .Y(u5__abc_78290_new_n2523_));
OAI21X1 OAI21X1_1378 ( .A(u5_timer2_6_), .B(u5__abc_78290_new_n2403_), .C(u5_timer2_7_), .Y(u5__abc_78290_new_n2527_));
OAI21X1 OAI21X1_1379 ( .A(u5__abc_78290_new_n2393_), .B(u5__abc_78290_new_n2526_), .C(u5__abc_78290_new_n2527_), .Y(u5__abc_78290_new_n2528_));
OAI21X1 OAI21X1_138 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1470_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1471_));
OAI21X1 OAI21X1_1380 ( .A(u5__abc_78290_new_n2393_), .B(u5__abc_78290_new_n2406_), .C(u5__abc_78290_new_n2500_), .Y(u5__abc_78290_new_n2531_));
OAI21X1 OAI21X1_1381 ( .A(u5__abc_78290_new_n2364_), .B(u5__abc_78290_new_n2500_), .C(u5__abc_78290_new_n2531_), .Y(u5__abc_78290_new_n2532_));
OAI21X1 OAI21X1_1382 ( .A(u5__abc_78290_new_n1597_), .B(u5__abc_78290_new_n1604_), .C(dv), .Y(u5__abc_78290_new_n2534_));
OAI21X1 OAI21X1_1383 ( .A(u5_ack_cnt_0_), .B(u5__abc_78290_new_n2537_), .C(u5__abc_78290_new_n2538_), .Y(u5__abc_78290_new_n2539_));
OAI21X1 OAI21X1_1384 ( .A(u5_ack_cnt_1_), .B(u5__abc_78290_new_n2535_), .C(u5__abc_78290_new_n2544_), .Y(u5__abc_78290_new_n2545_));
OAI21X1 OAI21X1_1385 ( .A(u5__abc_78290_new_n2543_), .B(u5__abc_78290_new_n2534_), .C(u5__abc_78290_new_n2538_), .Y(u5__abc_78290_new_n2546_));
OAI21X1 OAI21X1_1386 ( .A(u5_ack_cnt_1_), .B(u5_ack_cnt_0_), .C(u5__abc_78290_new_n2534_), .Y(u5__abc_78290_new_n2549_));
OAI21X1 OAI21X1_1387 ( .A(u5__abc_78290_new_n2535_), .B(u5__abc_78290_new_n2542_), .C(u5__abc_78290_new_n2549_), .Y(u5__abc_78290_new_n2550_));
OAI21X1 OAI21X1_1388 ( .A(u5__abc_78290_new_n2548_), .B(u5__abc_78290_new_n2550_), .C(u5__abc_78290_new_n2538_), .Y(u5__abc_78290_new_n2551_));
OAI21X1 OAI21X1_1389 ( .A(u5__abc_78290_new_n1596_), .B(u5__abc_78290_new_n2536_), .C(u5_ack_cnt_3_), .Y(u5__abc_78290_new_n2553_));
OAI21X1 OAI21X1_139 ( .A(u0__abc_74894_new_n1471_), .B(u0__abc_74894_new_n1469_), .C(u0__abc_74894_new_n1473_), .Y(u0__abc_74894_new_n1474_));
OAI21X1 OAI21X1_1390 ( .A(u5__abc_78290_new_n2555_), .B(u5__abc_78290_new_n2534_), .C(u5__abc_78290_new_n2538_), .Y(u5__abc_78290_new_n2556_));
OAI21X1 OAI21X1_1391 ( .A(u5_mc_le), .B(u5__abc_78290_new_n1990_), .C(u5__abc_78290_new_n2558_), .Y(u5__0cmd_asserted2_0_0_));
OAI21X1 OAI21X1_1392 ( .A(u5__abc_78290_new_n1507_), .B(u5__abc_78290_new_n1477_), .C(u5__0mc_le_0_0_), .Y(u5__abc_78290_new_n2560_));
OAI21X1 OAI21X1_1393 ( .A(u5__0mc_le_0_0_), .B(u5__abc_78290_new_n1990_), .C(u5__abc_78290_new_n2560_), .Y(u5__0cmd_asserted_0_0_));
OAI21X1 OAI21X1_1394 ( .A(u5_mc_le), .B(u5__abc_78290_new_n2562_), .C(u5__abc_78290_new_n2563_), .Y(u5__0mc_adv_r_0_0_));
OAI21X1 OAI21X1_1395 ( .A(u5__0mc_le_0_0_), .B(u5__abc_78290_new_n2562_), .C(u5__abc_78290_new_n2574_), .Y(u5__0mc_adv_r1_0_0_));
OAI21X1 OAI21X1_1396 ( .A(u5__abc_78290_new_n1058_), .B(u5__abc_78290_new_n1311_), .C(u5__abc_78290_new_n1375_), .Y(u5__abc_78290_new_n2576_));
OAI21X1 OAI21X1_1397 ( .A(u5__abc_78290_new_n2581_), .B(u5__abc_78290_new_n2578_), .C(u5__abc_78290_new_n1342_), .Y(u5__abc_78290_new_n2582_));
OAI21X1 OAI21X1_1398 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1335_), .C(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2584_));
OAI21X1 OAI21X1_1399 ( .A(u5__abc_78290_new_n486_), .B(u5__abc_78290_new_n1414_), .C(u5_tmr2_done), .Y(u5__abc_78290_new_n2586_));
OAI21X1 OAI21X1_14 ( .A(spec_req_cs_4_), .B(_abc_81086_new_n236_), .C(_abc_81086_new_n240_), .Y(_abc_81086_new_n257_));
OAI21X1 OAI21X1_140 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1490_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1491_));
OAI21X1 OAI21X1_1400 ( .A(u5__abc_78290_new_n486_), .B(u5_cs_le_r), .C(u5__abc_78290_new_n2587_), .Y(u5__abc_78290_new_n2588_));
OAI21X1 OAI21X1_1401 ( .A(u5__abc_78290_new_n2578_), .B(u5__abc_78290_new_n2581_), .C(u5__abc_78290_new_n2592_), .Y(u5__abc_78290_new_n2593_));
OAI21X1 OAI21X1_1402 ( .A(u5__abc_78290_new_n793_), .B(u5__abc_78290_new_n2594_), .C(u5__abc_78290_new_n2590_), .Y(u5__abc_78290_new_n2595_));
OAI21X1 OAI21X1_1403 ( .A(u5_state_1_), .B(u5__abc_78290_new_n2589_), .C(u5__abc_78290_new_n2595_), .Y(u5__abc_78290_new_n2596_));
OAI21X1 OAI21X1_1404 ( .A(u5__abc_78290_new_n793_), .B(u5__abc_78290_new_n2601_), .C(u5__abc_78290_new_n2600_), .Y(u5__abc_78290_new_n2602_));
OAI21X1 OAI21X1_1405 ( .A(u5_wb_write_go_r), .B(u5__abc_78290_new_n1600_), .C(u5__abc_78290_new_n862_), .Y(u5__abc_78290_new_n2607_));
OAI21X1 OAI21X1_1406 ( .A(u5__abc_78290_new_n2607_), .B(u5__abc_78290_new_n1609_), .C(u5__abc_78290_new_n1500_), .Y(u5__abc_78290_new_n2608_));
OAI21X1 OAI21X1_1407 ( .A(tms_s_9_), .B(u5__abc_78290_new_n1406_), .C(u5__abc_78290_new_n486_), .Y(u5__abc_78290_new_n2609_));
OAI21X1 OAI21X1_1408 ( .A(u5__abc_78290_new_n2608_), .B(u5__abc_78290_new_n2606_), .C(u5__abc_78290_new_n2609_), .Y(u5__abc_78290_new_n2610_));
OAI21X1 OAI21X1_1409 ( .A(u5_state_2_), .B(u5__abc_78290_new_n1419_), .C(u5__abc_78290_new_n1273_), .Y(u5__abc_78290_new_n2612_));
OAI21X1 OAI21X1_141 ( .A(u0__abc_74894_new_n1491_), .B(u0__abc_74894_new_n1489_), .C(u0__abc_74894_new_n1493_), .Y(u0__abc_74894_new_n1494_));
OAI21X1 OAI21X1_1410 ( .A(u5__abc_78290_new_n2591_), .B(u5__abc_78290_new_n2613_), .C(u5__abc_78290_new_n2576_), .Y(u5__abc_78290_new_n2614_));
OAI21X1 OAI21X1_1411 ( .A(u5__abc_78290_new_n2616_), .B(u5__abc_78290_new_n2614_), .C(u5_state_2_), .Y(u5__abc_78290_new_n2617_));
OAI21X1 OAI21X1_1412 ( .A(u5_state_2_), .B(u5_cmd_asserted), .C(u5__abc_78290_new_n2618_), .Y(u5__abc_78290_new_n2619_));
OAI21X1 OAI21X1_1413 ( .A(u5_state_2_), .B(u5__abc_78290_new_n2579_), .C(u5__abc_78290_new_n2620_), .Y(u5__abc_78290_new_n2621_));
OAI21X1 OAI21X1_1414 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1042_), .C(u5__abc_78290_new_n2621_), .Y(u5__abc_78290_new_n2622_));
OAI21X1 OAI21X1_1415 ( .A(u1_wb_write_go), .B(u5__abc_78290_new_n1597_), .C(u5__abc_78290_new_n1601_), .Y(u5__abc_78290_new_n2624_));
OAI21X1 OAI21X1_1416 ( .A(u1_wb_write_go), .B(u5__abc_78290_new_n1597_), .C(u5__abc_78290_new_n2626_), .Y(u5__abc_78290_new_n2627_));
OAI21X1 OAI21X1_1417 ( .A(u5_state_2_), .B(u5__abc_78290_new_n2625_), .C(u5__abc_78290_new_n2629_), .Y(u5__abc_78290_new_n2630_));
OAI21X1 OAI21X1_1418 ( .A(u5_state_2_), .B(u5__abc_78290_new_n2601_), .C(u5__abc_78290_new_n2631_), .Y(u5__abc_78290_new_n2632_));
OAI21X1 OAI21X1_1419 ( .A(u5_state_2_), .B(u5_cmd_asserted), .C(u5__abc_78290_new_n1257_), .Y(u5__abc_78290_new_n2639_));
OAI21X1 OAI21X1_142 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1510_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1511_));
OAI21X1 OAI21X1_1420 ( .A(u5__abc_78290_new_n2612_), .B(u5__abc_78290_new_n2611_), .C(u5__abc_78290_new_n2641_), .Y(u5_next_state_2_));
OAI21X1 OAI21X1_1421 ( .A(u5__abc_78290_new_n2643_), .B(u5__abc_78290_new_n1019_), .C(u5__abc_78290_new_n2645_), .Y(u5_next_state_3_));
OAI21X1 OAI21X1_1422 ( .A(u5__abc_78290_new_n627_), .B(u5__abc_78290_new_n2580_), .C(u5__abc_78290_new_n1335_), .Y(u5__abc_78290_new_n2648_));
OAI21X1 OAI21X1_1423 ( .A(u5__abc_78290_new_n2649_), .B(u5__abc_78290_new_n2655_), .C(u5__abc_78290_new_n974_), .Y(u5__abc_78290_new_n2656_));
OAI21X1 OAI21X1_1424 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n2374_), .C(u5__abc_78290_new_n2657_), .Y(u5_next_state_4_));
OAI21X1 OAI21X1_1425 ( .A(u5__abc_78290_new_n2664_), .B(u5__abc_78290_new_n2652_), .C(u5__abc_78290_new_n2578_), .Y(u5__abc_78290_new_n2665_));
OAI21X1 OAI21X1_1426 ( .A(u5__abc_78290_new_n2667_), .B(u5__abc_78290_new_n1335_), .C(u5__abc_78290_new_n733_), .Y(u5__abc_78290_new_n2668_));
OAI21X1 OAI21X1_1427 ( .A(u5__abc_78290_new_n2669_), .B(u5__abc_78290_new_n2577_), .C(u5__abc_78290_new_n2676_), .Y(u5_next_state_6_));
OAI21X1 OAI21X1_1428 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1335_), .C(u5__abc_78290_new_n1342_), .Y(u5__abc_78290_new_n2679_));
OAI21X1 OAI21X1_1429 ( .A(u5_wb_wait_r), .B(u5__abc_78290_new_n1375_), .C(u5__abc_78290_new_n1620_), .Y(u5__abc_78290_new_n2683_));
OAI21X1 OAI21X1_143 ( .A(u0__abc_74894_new_n1511_), .B(u0__abc_74894_new_n1509_), .C(u0__abc_74894_new_n1513_), .Y(u0__abc_74894_new_n1514_));
OAI21X1 OAI21X1_1430 ( .A(u5__abc_78290_new_n2681_), .B(u5__abc_78290_new_n2577_), .C(u5__abc_78290_new_n2685_), .Y(u5_next_state_7_));
OAI21X1 OAI21X1_1431 ( .A(u5__abc_78290_new_n2653_), .B(u5__abc_78290_new_n2688_), .C(u5__abc_78290_new_n2690_), .Y(u5__abc_78290_new_n2691_));
OAI21X1 OAI21X1_1432 ( .A(u5_state_8_), .B(u5__abc_78290_new_n2578_), .C(u5__abc_78290_new_n2691_), .Y(u5__abc_78290_new_n2692_));
OAI21X1 OAI21X1_1433 ( .A(u5__abc_78290_new_n2598_), .B(u5__abc_78290_new_n1455_), .C(u5__abc_78290_new_n1414_), .Y(u5__abc_78290_new_n2693_));
OAI21X1 OAI21X1_1434 ( .A(u5__abc_78290_new_n1324_), .B(u5_wb_wait), .C(u5__abc_78290_new_n2693_), .Y(u5__abc_78290_new_n2694_));
OAI21X1 OAI21X1_1435 ( .A(u5__abc_78290_new_n1514_), .B(u5__abc_78290_new_n1335_), .C(u5__abc_78290_new_n726_), .Y(u5__abc_78290_new_n2696_));
OAI21X1 OAI21X1_1436 ( .A(u5__abc_78290_new_n726_), .B(u5__abc_78290_new_n1414_), .C(u5__abc_78290_new_n2697_), .Y(u5__abc_78290_new_n2698_));
OAI21X1 OAI21X1_1437 ( .A(u5_wb_wait_r), .B(u5__abc_78290_new_n1375_), .C(u5__abc_78290_new_n726_), .Y(u5__abc_78290_new_n2702_));
OAI21X1 OAI21X1_1438 ( .A(u5__abc_78290_new_n1324_), .B(u5__abc_78290_new_n1375_), .C(u5__abc_78290_new_n2702_), .Y(u5__abc_78290_new_n2703_));
OAI21X1 OAI21X1_1439 ( .A(u5__abc_78290_new_n726_), .B(u5__abc_78290_new_n1414_), .C(u5__abc_78290_new_n2147_), .Y(u5__abc_78290_new_n2704_));
OAI21X1 OAI21X1_144 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1530_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1531_));
OAI21X1 OAI21X1_1440 ( .A(u5__abc_78290_new_n1291_), .B(u5__abc_78290_new_n2703_), .C(u5__abc_78290_new_n2705_), .Y(u5__abc_78290_new_n2706_));
OAI21X1 OAI21X1_1441 ( .A(u5__abc_78290_new_n2701_), .B(u5__abc_78290_new_n2706_), .C(u5__abc_78290_new_n2700_), .Y(u5__abc_78290_new_n2707_));
OAI21X1 OAI21X1_1442 ( .A(u5__abc_78290_new_n2699_), .B(u5__abc_78290_new_n2613_), .C(u5__abc_78290_new_n2707_), .Y(u5_next_state_9_));
OAI21X1 OAI21X1_1443 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1335_), .C(u5_state_10_), .Y(u5__abc_78290_new_n2709_));
OAI21X1 OAI21X1_1444 ( .A(u5__abc_78290_new_n2709_), .B(u5__abc_78290_new_n2613_), .C(u5__abc_78290_new_n2710_), .Y(u5_next_state_10_));
OAI21X1 OAI21X1_1445 ( .A(u5_wb_cycle), .B(u5__abc_78290_new_n1609_), .C(u5__abc_78290_new_n2715_), .Y(u5__abc_78290_new_n2716_));
OAI21X1 OAI21X1_1446 ( .A(u5__abc_78290_new_n2716_), .B(u5__abc_78290_new_n2712_), .C(u5__abc_78290_new_n2719_), .Y(u5_next_state_11_));
OAI21X1 OAI21X1_1447 ( .A(u5__abc_78290_new_n2721_), .B(u5__abc_78290_new_n2716_), .C(u5__abc_78290_new_n2724_), .Y(u5_next_state_12_));
OAI21X1 OAI21X1_1448 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1335_), .C(u5_state_13_), .Y(u5__abc_78290_new_n2726_));
OAI21X1 OAI21X1_1449 ( .A(u5__abc_78290_new_n1291_), .B(u5__abc_78290_new_n1620_), .C(u5__abc_78290_new_n2727_), .Y(u5__abc_78290_new_n2728_));
OAI21X1 OAI21X1_145 ( .A(u0__abc_74894_new_n1531_), .B(u0__abc_74894_new_n1529_), .C(u0__abc_74894_new_n1533_), .Y(u0__abc_74894_new_n1534_));
OAI21X1 OAI21X1_1450 ( .A(u5__abc_78290_new_n2726_), .B(u5__abc_78290_new_n2613_), .C(u5__abc_78290_new_n2729_), .Y(u5_next_state_13_));
OAI21X1 OAI21X1_1451 ( .A(u5__abc_78290_new_n1600_), .B(u5_wb_write_go_r), .C(u5__abc_78290_new_n2609_), .Y(u5__abc_78290_new_n2736_));
OAI21X1 OAI21X1_1452 ( .A(u5__abc_78290_new_n2736_), .B(u5__abc_78290_new_n1609_), .C(u5__abc_78290_new_n1419_), .Y(u5__abc_78290_new_n2737_));
OAI21X1 OAI21X1_1453 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n2741_), .C(u5__abc_78290_new_n2747_), .Y(u5__abc_78290_new_n2748_));
OAI21X1 OAI21X1_1454 ( .A(u5_state_15_), .B(u5__abc_78290_new_n486_), .C(u5__abc_78290_new_n2605_), .Y(u5__abc_78290_new_n2749_));
OAI21X1 OAI21X1_1455 ( .A(u5__abc_78290_new_n486_), .B(u5__abc_78290_new_n1324_), .C(u5__abc_78290_new_n2749_), .Y(u5__abc_78290_new_n2750_));
OAI21X1 OAI21X1_1456 ( .A(u5_wb_write_go_r), .B(u5__abc_78290_new_n1600_), .C(u5_state_15_), .Y(u5__abc_78290_new_n2752_));
OAI21X1 OAI21X1_1457 ( .A(u5__abc_78290_new_n2752_), .B(u5__abc_78290_new_n1609_), .C(u5__abc_78290_new_n1500_), .Y(u5__abc_78290_new_n2753_));
OAI21X1 OAI21X1_1458 ( .A(u5__abc_78290_new_n2612_), .B(u5__abc_78290_new_n2754_), .C(u5__abc_78290_new_n2751_), .Y(u5_next_state_15_));
OAI21X1 OAI21X1_1459 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n1335_), .C(u5_state_16_), .Y(u5__abc_78290_new_n2758_));
OAI21X1 OAI21X1_146 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1550_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1551_));
OAI21X1 OAI21X1_1460 ( .A(u5__abc_78290_new_n2758_), .B(u5__abc_78290_new_n2613_), .C(u5__abc_78290_new_n2763_), .Y(u5__abc_78290_new_n2764_));
OAI21X1 OAI21X1_1461 ( .A(u5_wb_write_go_r), .B(u5__abc_78290_new_n1600_), .C(u5_state_16_), .Y(u5__abc_78290_new_n2767_));
OAI21X1 OAI21X1_1462 ( .A(u5__abc_78290_new_n1609_), .B(u5__abc_78290_new_n2767_), .C(u5__abc_78290_new_n2766_), .Y(u5__abc_78290_new_n2768_));
OAI21X1 OAI21X1_1463 ( .A(u5__abc_78290_new_n2612_), .B(u5__abc_78290_new_n2770_), .C(u5__abc_78290_new_n2765_), .Y(u5_next_state_16_));
OAI21X1 OAI21X1_1464 ( .A(u5__abc_78290_new_n2773_), .B(u5__abc_78290_new_n2618_), .C(u5__abc_78290_new_n2774_), .Y(u5__abc_78290_new_n2775_));
OAI21X1 OAI21X1_1465 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n2076_), .C(u5__abc_78290_new_n472_), .Y(u5__abc_78290_new_n2777_));
OAI21X1 OAI21X1_1466 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n571_), .C(u5__abc_78290_new_n2778_), .Y(u5__abc_78290_new_n2779_));
OAI21X1 OAI21X1_1467 ( .A(u5_wb_cycle), .B(u5__abc_78290_new_n1338_), .C(u5_state_18_), .Y(u5__abc_78290_new_n2784_));
OAI21X1 OAI21X1_1468 ( .A(u5__abc_78290_new_n2782_), .B(u5__abc_78290_new_n2785_), .C(u5__abc_78290_new_n2783_), .Y(u5__abc_78290_new_n2786_));
OAI21X1 OAI21X1_1469 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n1437_), .C(u5__abc_78290_new_n2786_), .Y(u5_next_state_18_));
OAI21X1 OAI21X1_147 ( .A(u0__abc_74894_new_n1551_), .B(u0__abc_74894_new_n1549_), .C(u0__abc_74894_new_n1553_), .Y(u0__abc_74894_new_n1554_));
OAI21X1 OAI21X1_1470 ( .A(u5_state_19_), .B(u5_cmd_asserted), .C(u5__abc_78290_new_n579_), .Y(u5__abc_78290_new_n2792_));
OAI21X1 OAI21X1_1471 ( .A(u5__abc_78290_new_n561_), .B(u5__abc_78290_new_n2791_), .C(u5__abc_78290_new_n2792_), .Y(u5__abc_78290_new_n2793_));
OAI21X1 OAI21X1_1472 ( .A(u5__abc_78290_new_n2797_), .B(u5__abc_78290_new_n2796_), .C(u5__abc_78290_new_n2800_), .Y(u5_next_state_20_));
OAI21X1 OAI21X1_1473 ( .A(u5__abc_78290_new_n2804_), .B(u5__abc_78290_new_n2577_), .C(u5__abc_78290_new_n2806_), .Y(u5_next_state_22_));
OAI21X1 OAI21X1_1474 ( .A(u5__abc_78290_new_n2808_), .B(u5__abc_78290_new_n2577_), .C(u5__abc_78290_new_n2811_), .Y(u5_next_state_23_));
OAI21X1 OAI21X1_1475 ( .A(u5__abc_78290_new_n2815_), .B(u5__abc_78290_new_n1200_), .C(u5__abc_78290_new_n2816_), .Y(u5__abc_78290_new_n2817_));
OAI21X1 OAI21X1_1476 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n587_), .C(u5__abc_78290_new_n2817_), .Y(u5__abc_78290_new_n2818_));
OAI21X1 OAI21X1_1477 ( .A(u5__abc_78290_new_n2820_), .B(u5__abc_78290_new_n2577_), .C(u5__abc_78290_new_n2823_), .Y(u5_next_state_25_));
OAI21X1 OAI21X1_1478 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n548_), .C(u5__abc_78290_new_n2815_), .Y(u5__abc_78290_new_n2826_));
OAI21X1 OAI21X1_1479 ( .A(u5__abc_78290_new_n2825_), .B(u5__abc_78290_new_n2577_), .C(u5__abc_78290_new_n2828_), .Y(u5_next_state_26_));
OAI21X1 OAI21X1_148 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1570_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1571_));
OAI21X1 OAI21X1_1480 ( .A(u5__abc_78290_new_n1336_), .B(u5__abc_78290_new_n1337_), .C(u5__abc_78290_new_n2783_), .Y(u5__abc_78290_new_n2830_));
OAI21X1 OAI21X1_1481 ( .A(u5_state_28_), .B(u5_cmd_asserted), .C(u5__abc_78290_new_n2835_), .Y(u5__abc_78290_new_n2836_));
OAI21X1 OAI21X1_1482 ( .A(u5_tmr_done), .B(u5__abc_78290_new_n2076_), .C(u5__abc_78290_new_n2836_), .Y(u5__abc_78290_new_n2837_));
OAI21X1 OAI21X1_1483 ( .A(u5__abc_78290_new_n1375_), .B(u5__abc_78290_new_n2076_), .C(u5__abc_78290_new_n522_), .Y(u5__abc_78290_new_n2840_));
OAI21X1 OAI21X1_1484 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n1302_), .C(u5__abc_78290_new_n2076_), .Y(u5__abc_78290_new_n2841_));
OAI21X1 OAI21X1_1485 ( .A(u5__abc_78290_new_n2839_), .B(u5__abc_78290_new_n2577_), .C(u5__abc_78290_new_n2842_), .Y(u5_next_state_29_));
OAI21X1 OAI21X1_1486 ( .A(u5__abc_78290_new_n1990_), .B(u5__abc_78290_new_n1302_), .C(u5__abc_78290_new_n481_), .Y(u5__abc_78290_new_n2845_));
OAI21X1 OAI21X1_1487 ( .A(u5_resume_req_r), .B(u5__abc_78290_new_n441_), .C(u5__abc_78290_new_n1302_), .Y(u5__abc_78290_new_n2846_));
OAI21X1 OAI21X1_1488 ( .A(u5__abc_78290_new_n2844_), .B(u5__abc_78290_new_n2577_), .C(u5__abc_78290_new_n2847_), .Y(u5_next_state_30_));
OAI21X1 OAI21X1_1489 ( .A(u5__abc_78290_new_n441_), .B(u5__abc_78290_new_n2850_), .C(u5__abc_78290_new_n2849_), .Y(u5_next_state_31_));
OAI21X1 OAI21X1_149 ( .A(u0__abc_74894_new_n1571_), .B(u0__abc_74894_new_n1569_), .C(u0__abc_74894_new_n1573_), .Y(u0__abc_74894_new_n1574_));
OAI21X1 OAI21X1_1490 ( .A(u5__abc_78290_new_n536_), .B(u5__abc_78290_new_n2852_), .C(u5__abc_78290_new_n2854_), .Y(u5_next_state_32_));
OAI21X1 OAI21X1_1491 ( .A(u5_state_33_), .B(u5__abc_78290_new_n2678_), .C(u5__abc_78290_new_n2783_), .Y(u5__abc_78290_new_n2856_));
OAI21X1 OAI21X1_1492 ( .A(u5__abc_78290_new_n515_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n816_), .Y(u5_next_state_34_));
OAI21X1 OAI21X1_1493 ( .A(u5__abc_78290_new_n513_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2859_), .Y(u5_next_state_35_));
OAI21X1 OAI21X1_1494 ( .A(u5_lookup_ready2), .B(u5__abc_78290_new_n2653_), .C(u5__abc_78290_new_n1414_), .Y(u5__abc_78290_new_n2861_));
OAI21X1 OAI21X1_1495 ( .A(u5__abc_78290_new_n2147_), .B(u5__abc_78290_new_n2864_), .C(u5__abc_78290_new_n2578_), .Y(u5__abc_78290_new_n2865_));
OAI21X1 OAI21X1_1496 ( .A(u5__abc_78290_new_n2862_), .B(u5__abc_78290_new_n2865_), .C(u5__abc_78290_new_n2663_), .Y(u5__abc_78290_new_n2866_));
OAI21X1 OAI21X1_1497 ( .A(u5_state_36_), .B(u5__abc_78290_new_n2578_), .C(u5__abc_78290_new_n2783_), .Y(u5__abc_78290_new_n2867_));
OAI21X1 OAI21X1_1498 ( .A(u5__abc_78290_new_n898_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2871_), .Y(u5_next_state_37_));
OAI21X1 OAI21X1_1499 ( .A(u5_state_38_), .B(u5_tmr2_done), .C(u5__abc_78290_new_n2874_), .Y(u5__abc_78290_new_n2875_));
OAI21X1 OAI21X1_15 ( .A(_abc_81086_new_n255_), .B(_abc_81086_new_n257_), .C(_abc_81086_new_n256_), .Y(obct_cs_4_));
OAI21X1 OAI21X1_150 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1590_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1591_));
OAI21X1 OAI21X1_1500 ( .A(u5__abc_78290_new_n2878_), .B(u5__abc_78290_new_n2877_), .C(u5__abc_78290_new_n1527_), .Y(u5__abc_78290_new_n2879_));
OAI21X1 OAI21X1_1501 ( .A(u5__abc_78290_new_n698_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2879_), .Y(u5_next_state_39_));
OAI21X1 OAI21X1_1502 ( .A(u5__abc_78290_new_n644_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n1393_), .Y(u5_next_state_40_));
OAI21X1 OAI21X1_1503 ( .A(u5__abc_78290_new_n2882_), .B(u5__abc_78290_new_n2883_), .C(u5__abc_78290_new_n1381_), .Y(u5__abc_78290_new_n2884_));
OAI21X1 OAI21X1_1504 ( .A(u5__abc_78290_new_n643_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2884_), .Y(u5_next_state_41_));
OAI21X1 OAI21X1_1505 ( .A(u5__abc_78290_new_n711_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2888_), .Y(u5_next_state_42_));
OAI21X1 OAI21X1_1506 ( .A(u5__abc_78290_new_n671_), .B(u5__abc_78290_new_n714_), .C(u5__abc_78290_new_n2894_), .Y(u5_next_state_44_));
OAI21X1 OAI21X1_1507 ( .A(csc_s_5_), .B(u5__abc_78290_new_n2896_), .C(u5_tmr2_done), .Y(u5__abc_78290_new_n2897_));
OAI21X1 OAI21X1_1508 ( .A(u5__abc_78290_new_n671_), .B(u5__abc_78290_new_n707_), .C(u5__abc_78290_new_n2898_), .Y(u5__abc_78290_new_n2899_));
OAI21X1 OAI21X1_1509 ( .A(u5_state_45_), .B(u5_tmr2_done), .C(u5__abc_78290_new_n2899_), .Y(u5__abc_78290_new_n2900_));
OAI21X1 OAI21X1_151 ( .A(u0__abc_74894_new_n1591_), .B(u0__abc_74894_new_n1589_), .C(u0__abc_74894_new_n1593_), .Y(u0__abc_74894_new_n1594_));
OAI21X1 OAI21X1_1510 ( .A(u5__abc_78290_new_n703_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2900_), .Y(u5_next_state_45_));
OAI21X1 OAI21X1_1511 ( .A(u5__abc_78290_new_n655_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2903_), .Y(u5_next_state_46_));
OAI21X1 OAI21X1_1512 ( .A(u5__abc_78290_new_n2908_), .B(u5__abc_78290_new_n2909_), .C(u5__abc_78290_new_n1442_), .Y(u5__abc_78290_new_n2910_));
OAI21X1 OAI21X1_1513 ( .A(u5__abc_78290_new_n634_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2910_), .Y(u5_next_state_48_));
OAI21X1 OAI21X1_1514 ( .A(u5__abc_78290_new_n614_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2915_), .Y(u5_next_state_50_));
OAI21X1 OAI21X1_1515 ( .A(u5_state_52_), .B(u5__abc_78290_new_n1414_), .C(u5__abc_78290_new_n2922_), .Y(u5__abc_78290_new_n2923_));
OAI21X1 OAI21X1_1516 ( .A(u5__abc_78290_new_n938_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2928_), .Y(u5_next_state_53_));
OAI21X1 OAI21X1_1517 ( .A(u5__abc_78290_new_n2565_), .B(u5__abc_78290_new_n1093_), .C(u5__abc_78290_new_n929_), .Y(u5__abc_78290_new_n2931_));
OAI21X1 OAI21X1_1518 ( .A(u5__abc_78290_new_n2926_), .B(u5__abc_78290_new_n2659_), .C(u5__abc_78290_new_n2931_), .Y(u5__abc_78290_new_n2932_));
OAI21X1 OAI21X1_1519 ( .A(u5__abc_78290_new_n1113_), .B(u5__abc_78290_new_n2930_), .C(u5__abc_78290_new_n2932_), .Y(u5_next_state_54_));
OAI21X1 OAI21X1_152 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1610_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1611_));
OAI21X1 OAI21X1_1520 ( .A(u5__abc_78290_new_n1113_), .B(u5__abc_78290_new_n2934_), .C(u5__abc_78290_new_n2938_), .Y(u5_next_state_55_));
OAI21X1 OAI21X1_1521 ( .A(u5__abc_78290_new_n2940_), .B(u5__abc_78290_new_n2941_), .C(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2942_));
OAI21X1 OAI21X1_1522 ( .A(u5_state_56_), .B(u5__abc_78290_new_n1597_), .C(u3_wb_read_go), .Y(u5__abc_78290_new_n2943_));
OAI21X1 OAI21X1_1523 ( .A(u5__abc_78290_new_n909_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2954_), .Y(u5_next_state_57_));
OAI21X1 OAI21X1_1524 ( .A(u5__abc_78290_new_n2956_), .B(u5__abc_78290_new_n2957_), .C(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2958_));
OAI21X1 OAI21X1_1525 ( .A(u1_wb_write_go), .B(u5__abc_78290_new_n1990_), .C(u5_state_58_), .Y(u5__abc_78290_new_n2959_));
OAI21X1 OAI21X1_1526 ( .A(u5__abc_78290_new_n902_), .B(u5__abc_78290_new_n2732_), .C(u5__abc_78290_new_n2963_), .Y(u5__abc_78290_new_n2964_));
OAI21X1 OAI21X1_1527 ( .A(u5__abc_78290_new_n902_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2965_), .Y(u5_next_state_59_));
OAI21X1 OAI21X1_1528 ( .A(u5__abc_78290_new_n2196_), .B(u5__abc_78290_new_n2971_), .C(u5__abc_78290_new_n2969_), .Y(u5_next_state_60_));
OAI21X1 OAI21X1_1529 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n854_), .C(u5__abc_78290_new_n2975_), .Y(u5__abc_78290_new_n2976_));
OAI21X1 OAI21X1_153 ( .A(u0__abc_74894_new_n1611_), .B(u0__abc_74894_new_n1609_), .C(u0__abc_74894_new_n1613_), .Y(u0__abc_74894_new_n1614_));
OAI21X1 OAI21X1_1530 ( .A(u5__abc_78290_new_n854_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2977_), .Y(u5_next_state_61_));
OAI21X1 OAI21X1_1531 ( .A(u5__abc_78290_new_n2982_), .B(u5__abc_78290_new_n2983_), .C(u5__abc_78290_new_n2583_), .Y(u5__abc_78290_new_n2984_));
OAI21X1 OAI21X1_1532 ( .A(u5__abc_78290_new_n2981_), .B(u5__abc_78290_new_n2985_), .C(u5__abc_78290_new_n2984_), .Y(u5_next_state_63_));
OAI21X1 OAI21X1_1533 ( .A(u5_tmr2_done), .B(u5__abc_78290_new_n490_), .C(u5__abc_78290_new_n2975_), .Y(u5__abc_78290_new_n2988_));
OAI21X1 OAI21X1_1534 ( .A(u5__abc_78290_new_n490_), .B(u5__abc_78290_new_n2584_), .C(u5__abc_78290_new_n2989_), .Y(u5_next_state_64_));
OAI21X1 OAI21X1_1535 ( .A(u5__abc_78290_new_n2896_), .B(csc_s_5_), .C(u5__abc_78290_new_n1165_), .Y(u5__abc_78290_new_n2993_));
OAI21X1 OAI21X1_1536 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1155_), .C(u5__abc_78290_new_n2890_), .Y(u5__abc_78290_new_n2996_));
OAI21X1 OAI21X1_1537 ( .A(u5__abc_78290_new_n3005_), .B(u5__abc_78290_new_n1609_), .C(u5__abc_78290_new_n1416_), .Y(u5__abc_78290_new_n3006_));
OAI21X1 OAI21X1_1538 ( .A(u5__abc_78290_new_n3007_), .B(u5__abc_78290_new_n3004_), .C(u5__abc_78290_new_n3014_), .Y(u5_cke_d));
OAI21X1 OAI21X1_1539 ( .A(u5__abc_78290_new_n1186_), .B(u5__abc_78290_new_n3021_), .C(u5__abc_78290_new_n1190_), .Y(u5_lmr_ack_d));
OAI21X1 OAI21X1_154 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1630_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1631_));
OAI21X1 OAI21X1_1540 ( .A(u5_wb_wait), .B(u5__abc_78290_new_n2742_), .C(u5__abc_78290_new_n2647_), .Y(u5__abc_78290_new_n3035_));
OAI21X1 OAI21X1_1541 ( .A(u5__abc_78290_new_n3038_), .B(u5__abc_78290_new_n3039_), .C(u5__abc_78290_new_n3040_), .Y(u5__abc_78290_new_n3041_));
OAI21X1 OAI21X1_1542 ( .A(u5__abc_78290_new_n1238_), .B(u5__abc_78290_new_n1038_), .C(u5__abc_78290_new_n1222_), .Y(u5__abc_78290_new_n3044_));
OAI21X1 OAI21X1_1543 ( .A(u5__abc_78290_new_n1344_), .B(u5__abc_78290_new_n3050_), .C(u5__abc_78290_new_n1478_), .Y(u5__abc_78290_new_n3051_));
OAI21X1 OAI21X1_1544 ( .A(u5__abc_78290_new_n1203_), .B(u5__abc_78290_new_n1242_), .C(u5__abc_78290_new_n433_), .Y(u5__abc_78290_new_n3052_));
OAI21X1 OAI21X1_1545 ( .A(u5__abc_78290_new_n2579_), .B(u5__abc_78290_new_n1363_), .C(u5__abc_78290_new_n3028_), .Y(u5__abc_78290_new_n3054_));
OAI21X1 OAI21X1_1546 ( .A(u5__abc_78290_new_n1374_), .B(u5__abc_78290_new_n1490_), .C(u5__abc_78290_new_n3070_), .Y(bank_clr));
OAI21X1 OAI21X1_1547 ( .A(u5__abc_78290_new_n1164_), .B(u5__abc_78290_new_n1038_), .C(u5__abc_78290_new_n2873_), .Y(u5__abc_78290_new_n3073_));
OAI21X1 OAI21X1_1548 ( .A(u5__abc_78290_new_n1380_), .B(u5__abc_78290_new_n1383_), .C(u5_tmr2_done), .Y(u5__abc_78290_new_n3082_));
OAI21X1 OAI21X1_1549 ( .A(u5__abc_78290_new_n1585_), .B(u5__abc_78290_new_n3081_), .C(u5__abc_78290_new_n3082_), .Y(next_adr));
OAI21X1 OAI21X1_155 ( .A(u0__abc_74894_new_n1631_), .B(u0__abc_74894_new_n1629_), .C(u0__abc_74894_new_n1633_), .Y(u0__abc_74894_new_n1634_));
OAI21X1 OAI21X1_1550 ( .A(u5__abc_78290_new_n3085_), .B(u5__abc_78290_new_n2331_), .C(u5__abc_78290_new_n1291_), .Y(row_sel));
OAI21X1 OAI21X1_1551 ( .A(u5__abc_78290_new_n1135_), .B(u5__abc_78290_new_n1399_), .C(u5__abc_78290_new_n2196_), .Y(u5__abc_78290_new_n3089_));
OAI21X1 OAI21X1_1552 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1060_), .C(u5__abc_78290_new_n1267_), .Y(u5__abc_78290_new_n3090_));
OAI21X1 OAI21X1_1553 ( .A(u5__abc_78290_new_n454_), .B(u5__abc_78290_new_n631_), .C(u5_cmd_a10_r), .Y(u5__abc_78290_new_n3099_));
OAI21X1 OAI21X1_1554 ( .A(u5__abc_78290_new_n3088_), .B(u5__abc_78290_new_n3097_), .C(u5_ap_en), .Y(u5__abc_78290_new_n3103_));
OAI21X1 OAI21X1_1555 ( .A(tms_s_9_), .B(u5__abc_78290_new_n1406_), .C(u5__abc_78290_new_n2598_), .Y(u5__abc_78290_new_n3104_));
OAI21X1 OAI21X1_1556 ( .A(u5__abc_78290_new_n1324_), .B(u5__abc_78290_new_n1375_), .C(u5__abc_78290_new_n1460_), .Y(u5__abc_78290_new_n3105_));
OAI21X1 OAI21X1_1557 ( .A(u5__abc_78290_new_n3104_), .B(u5__abc_78290_new_n3106_), .C(u5__abc_78290_new_n1631_), .Y(u5__abc_78290_new_n3107_));
OAI21X1 OAI21X1_1558 ( .A(u5_ap_en), .B(u5__abc_78290_new_n1325_), .C(u5__abc_78290_new_n1262_), .Y(u5__abc_78290_new_n3108_));
OAI21X1 OAI21X1_1559 ( .A(u5__abc_78290_new_n2672_), .B(u5__abc_78290_new_n1297_), .C(u5__abc_78290_new_n3060_), .Y(u5__abc_78290_new_n3111_));
OAI21X1 OAI21X1_156 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1650_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1651_));
OAI21X1 OAI21X1_1560 ( .A(u5__abc_78290_new_n3098_), .B(u5__abc_78290_new_n3102_), .C(u5__abc_78290_new_n3114_), .Y(cmd_a10));
OAI21X1 OAI21X1_1561 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1123_), .C(u5__abc_78290_new_n1052_), .Y(u5__abc_78290_new_n3116_));
OAI21X1 OAI21X1_1562 ( .A(u5__abc_78290_new_n1113_), .B(u5__abc_78290_new_n2930_), .C(u5__abc_78290_new_n3118_), .Y(u5__abc_78290_new_n3119_));
OAI21X1 OAI21X1_1563 ( .A(u5_wb_cycle), .B(u5__abc_78290_new_n1609_), .C(u5_cnt), .Y(u5__abc_78290_new_n3132_));
OAI21X1 OAI21X1_1564 ( .A(mc_cke_pad_o_), .B(u5__abc_78290_new_n3133_), .C(u5__abc_78290_new_n3134_), .Y(u5__abc_78290_new_n3135_));
OAI21X1 OAI21X1_1565 ( .A(u5__abc_78290_new_n3150_), .B(u5__abc_78290_new_n2005_), .C(susp_sel), .Y(u5__abc_78290_new_n3151_));
OAI21X1 OAI21X1_1566 ( .A(u5__abc_78290_new_n1340_), .B(u5__abc_78290_new_n2830_), .C(u5__abc_78290_new_n3151_), .Y(u5__0susp_sel_r_0_0_));
OAI21X1 OAI21X1_1567 ( .A(not_mem_cyc), .B(u5__abc_78290_new_n3153_), .C(u5__abc_78290_new_n1479_), .Y(u5__0wb_cycle_0_0_));
OAI21X1 OAI21X1_1568 ( .A(u5__abc_78290_new_n1598_), .B(u5__abc_78290_new_n1599_), .C(u5__abc_78290_new_n1324_), .Y(u5__abc_78290_new_n3155_));
OAI21X1 OAI21X1_1569 ( .A(u5__abc_78290_new_n2667_), .B(u5__abc_78290_new_n1479_), .C(u5__abc_78290_new_n1357_), .Y(u5__abc_78290_new_n3156_));
OAI21X1 OAI21X1_157 ( .A(u0__abc_74894_new_n1651_), .B(u0__abc_74894_new_n1649_), .C(u0__abc_74894_new_n1653_), .Y(u0__abc_74894_new_n1654_));
OAI21X1 OAI21X1_1570 ( .A(u5__abc_78290_new_n1429_), .B(u5__abc_78290_new_n1318_), .C(u5__abc_78290_new_n3157_), .Y(u5__0wr_cycle_0_0_));
OAI21X1 OAI21X1_1571 ( .A(err), .B(u6__abc_81318_new_n139_), .C(u6__abc_81318_new_n138_), .Y(u6__abc_81318_new_n140_));
OAI21X1 OAI21X1_1572 ( .A(u6__abc_81318_new_n146_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n147_), .Y(u6__0wb_data_o_31_0__0_));
OAI21X1 OAI21X1_1573 ( .A(u6__abc_81318_new_n149_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n150_), .Y(u6__0wb_data_o_31_0__1_));
OAI21X1 OAI21X1_1574 ( .A(u6__abc_81318_new_n152_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n153_), .Y(u6__0wb_data_o_31_0__2_));
OAI21X1 OAI21X1_1575 ( .A(u6__abc_81318_new_n155_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n156_), .Y(u6__0wb_data_o_31_0__3_));
OAI21X1 OAI21X1_1576 ( .A(u6__abc_81318_new_n158_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n159_), .Y(u6__0wb_data_o_31_0__4_));
OAI21X1 OAI21X1_1577 ( .A(u6__abc_81318_new_n161_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n162_), .Y(u6__0wb_data_o_31_0__5_));
OAI21X1 OAI21X1_1578 ( .A(u6__abc_81318_new_n164_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n165_), .Y(u6__0wb_data_o_31_0__6_));
OAI21X1 OAI21X1_1579 ( .A(u6__abc_81318_new_n167_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n168_), .Y(u6__0wb_data_o_31_0__7_));
OAI21X1 OAI21X1_158 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1670_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1671_));
OAI21X1 OAI21X1_1580 ( .A(u6__abc_81318_new_n170_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n171_), .Y(u6__0wb_data_o_31_0__8_));
OAI21X1 OAI21X1_1581 ( .A(u6__abc_81318_new_n173_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n174_), .Y(u6__0wb_data_o_31_0__9_));
OAI21X1 OAI21X1_1582 ( .A(u6__abc_81318_new_n176_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n177_), .Y(u6__0wb_data_o_31_0__10_));
OAI21X1 OAI21X1_1583 ( .A(u6__abc_81318_new_n179_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n180_), .Y(u6__0wb_data_o_31_0__11_));
OAI21X1 OAI21X1_1584 ( .A(u6__abc_81318_new_n182_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n183_), .Y(u6__0wb_data_o_31_0__12_));
OAI21X1 OAI21X1_1585 ( .A(u6__abc_81318_new_n185_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n186_), .Y(u6__0wb_data_o_31_0__13_));
OAI21X1 OAI21X1_1586 ( .A(u6__abc_81318_new_n188_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n189_), .Y(u6__0wb_data_o_31_0__14_));
OAI21X1 OAI21X1_1587 ( .A(u6__abc_81318_new_n191_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n192_), .Y(u6__0wb_data_o_31_0__15_));
OAI21X1 OAI21X1_1588 ( .A(u6__abc_81318_new_n194_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n195_), .Y(u6__0wb_data_o_31_0__16_));
OAI21X1 OAI21X1_1589 ( .A(u6__abc_81318_new_n197_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n198_), .Y(u6__0wb_data_o_31_0__17_));
OAI21X1 OAI21X1_159 ( .A(u0__abc_74894_new_n1671_), .B(u0__abc_74894_new_n1669_), .C(u0__abc_74894_new_n1673_), .Y(u0__abc_74894_new_n1674_));
OAI21X1 OAI21X1_1590 ( .A(u6__abc_81318_new_n200_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n201_), .Y(u6__0wb_data_o_31_0__18_));
OAI21X1 OAI21X1_1591 ( .A(u6__abc_81318_new_n203_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n204_), .Y(u6__0wb_data_o_31_0__19_));
OAI21X1 OAI21X1_1592 ( .A(u6__abc_81318_new_n206_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n207_), .Y(u6__0wb_data_o_31_0__20_));
OAI21X1 OAI21X1_1593 ( .A(u6__abc_81318_new_n209_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n210_), .Y(u6__0wb_data_o_31_0__21_));
OAI21X1 OAI21X1_1594 ( .A(u6__abc_81318_new_n212_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n213_), .Y(u6__0wb_data_o_31_0__22_));
OAI21X1 OAI21X1_1595 ( .A(u6__abc_81318_new_n215_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n216_), .Y(u6__0wb_data_o_31_0__23_));
OAI21X1 OAI21X1_1596 ( .A(u6__abc_81318_new_n218_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n219_), .Y(u6__0wb_data_o_31_0__24_));
OAI21X1 OAI21X1_1597 ( .A(u6__abc_81318_new_n221_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n222_), .Y(u6__0wb_data_o_31_0__25_));
OAI21X1 OAI21X1_1598 ( .A(u6__abc_81318_new_n224_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n225_), .Y(u6__0wb_data_o_31_0__26_));
OAI21X1 OAI21X1_1599 ( .A(u6__abc_81318_new_n227_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n228_), .Y(u6__0wb_data_o_31_0__27_));
OAI21X1 OAI21X1_16 ( .A(susp_sel), .B(rfr_ack), .C(cs_need_rfr_5_), .Y(_abc_81086_new_n260_));
OAI21X1 OAI21X1_160 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1690_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1691_));
OAI21X1 OAI21X1_1600 ( .A(u6__abc_81318_new_n230_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n231_), .Y(u6__0wb_data_o_31_0__28_));
OAI21X1 OAI21X1_1601 ( .A(u6__abc_81318_new_n233_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n234_), .Y(u6__0wb_data_o_31_0__29_));
OAI21X1 OAI21X1_1602 ( .A(u6__abc_81318_new_n236_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n237_), .Y(u6__0wb_data_o_31_0__30_));
OAI21X1 OAI21X1_1603 ( .A(u6__abc_81318_new_n239_), .B(u6__abc_81318_new_n135_), .C(u6__abc_81318_new_n240_), .Y(u6__0wb_data_o_31_0__31_));
OAI21X1 OAI21X1_1604 ( .A(u6__abc_81318_new_n242_), .B(u6__abc_81318_new_n138_), .C(u6__abc_81318_new_n243_), .Y(u6__0wr_hold_0_0_));
OAI21X1 OAI21X1_1605 ( .A(u6__abc_81318_new_n135_), .B(u6__abc_81318_new_n269_), .C(u6__abc_81318_new_n271_), .Y(u5_wb_first));
OAI21X1 OAI21X1_1606 ( .A(u6__abc_81318_new_n136_), .B(u6__abc_81318_new_n253_), .C(u6__abc_81318_new_n143_), .Y(u6__0rmw_en_0_0_));
OAI21X1 OAI21X1_1607 ( .A(u6__abc_81318_new_n135_), .B(u6__abc_81318_new_n269_), .C(u6__abc_81318_new_n271_), .Y(u6__0wb_first_r_0_0_));
OAI21X1 OAI21X1_1608 ( .A(u1_wr_cycle), .B(u7__abc_73829_new_n78_), .C(u7__abc_73829_new_n76_), .Y(u7__abc_73829_new_n79_));
OAI21X1 OAI21X1_1609 ( .A(u7__abc_73829_new_n87_), .B(u7__abc_73829_new_n88_), .C(u7__abc_73829_new_n89_), .Y(u7__0mc_dqm_r_3_0__0_));
OAI21X1 OAI21X1_161 ( .A(u0__abc_74894_new_n1691_), .B(u0__abc_74894_new_n1689_), .C(u0__abc_74894_new_n1693_), .Y(u0__abc_74894_new_n1694_));
OAI21X1 OAI21X1_1610 ( .A(u7__abc_73829_new_n91_), .B(u7__abc_73829_new_n88_), .C(u7__abc_73829_new_n92_), .Y(u7__0mc_dqm_r_3_0__1_));
OAI21X1 OAI21X1_1611 ( .A(u7__abc_73829_new_n94_), .B(u7__abc_73829_new_n88_), .C(u7__abc_73829_new_n95_), .Y(u7__0mc_dqm_r_3_0__2_));
OAI21X1 OAI21X1_1612 ( .A(u7__abc_73829_new_n97_), .B(u7__abc_73829_new_n88_), .C(u7__abc_73829_new_n98_), .Y(u7__0mc_dqm_r_3_0__3_));
OAI21X1 OAI21X1_162 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1710_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1711_));
OAI21X1 OAI21X1_163 ( .A(u0__abc_74894_new_n1711_), .B(u0__abc_74894_new_n1709_), .C(u0__abc_74894_new_n1713_), .Y(u0__abc_74894_new_n1714_));
OAI21X1 OAI21X1_164 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1831_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1832_));
OAI21X1 OAI21X1_165 ( .A(u0__abc_74894_new_n1832_), .B(u0__abc_74894_new_n1830_), .C(u0__abc_74894_new_n1834_), .Y(u0__abc_74894_new_n1835_));
OAI21X1 OAI21X1_166 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1851_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1852_));
OAI21X1 OAI21X1_167 ( .A(u0__abc_74894_new_n1852_), .B(u0__abc_74894_new_n1850_), .C(u0__abc_74894_new_n1854_), .Y(u0__abc_74894_new_n1855_));
OAI21X1 OAI21X1_168 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1871_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1872_));
OAI21X1 OAI21X1_169 ( .A(u0__abc_74894_new_n1872_), .B(u0__abc_74894_new_n1870_), .C(u0__abc_74894_new_n1874_), .Y(u0__abc_74894_new_n1875_));
OAI21X1 OAI21X1_17 ( .A(spec_req_cs_5_), .B(_abc_81086_new_n236_), .C(_abc_81086_new_n240_), .Y(_abc_81086_new_n261_));
OAI21X1 OAI21X1_170 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1891_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1892_));
OAI21X1 OAI21X1_171 ( .A(u0__abc_74894_new_n1892_), .B(u0__abc_74894_new_n1890_), .C(u0__abc_74894_new_n1894_), .Y(u0__abc_74894_new_n1895_));
OAI21X1 OAI21X1_172 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1911_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1912_));
OAI21X1 OAI21X1_173 ( .A(u0__abc_74894_new_n1912_), .B(u0__abc_74894_new_n1910_), .C(u0__abc_74894_new_n1914_), .Y(u0__abc_74894_new_n1915_));
OAI21X1 OAI21X1_174 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1931_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1932_));
OAI21X1 OAI21X1_175 ( .A(u0__abc_74894_new_n1932_), .B(u0__abc_74894_new_n1930_), .C(u0__abc_74894_new_n1934_), .Y(u0__abc_74894_new_n1935_));
OAI21X1 OAI21X1_176 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1951_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1952_));
OAI21X1 OAI21X1_177 ( .A(u0__abc_74894_new_n1952_), .B(u0__abc_74894_new_n1950_), .C(u0__abc_74894_new_n1954_), .Y(u0__abc_74894_new_n1955_));
OAI21X1 OAI21X1_178 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n1991_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n1992_));
OAI21X1 OAI21X1_179 ( .A(u0__abc_74894_new_n1992_), .B(u0__abc_74894_new_n1990_), .C(u0__abc_74894_new_n1994_), .Y(u0__abc_74894_new_n1995_));
OAI21X1 OAI21X1_18 ( .A(_abc_81086_new_n259_), .B(_abc_81086_new_n261_), .C(_abc_81086_new_n260_), .Y(obct_cs_5_));
OAI21X1 OAI21X1_180 ( .A(u0__abc_74894_new_n1106_), .B(u0__abc_74894_new_n2011_), .C(u0__abc_74894_new_n1100_), .Y(u0__abc_74894_new_n2012_));
OAI21X1 OAI21X1_181 ( .A(u0__abc_74894_new_n2012_), .B(u0__abc_74894_new_n2010_), .C(u0__abc_74894_new_n2014_), .Y(u0__abc_74894_new_n2015_));
OAI21X1 OAI21X1_182 ( .A(u0__abc_74894_new_n1170_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2456_));
OAI21X1 OAI21X1_183 ( .A(u0__abc_74894_new_n2456_), .B(u0__abc_74894_new_n2453_), .C(u0__abc_74894_new_n2457_), .Y(u0__abc_74894_new_n2458_));
OAI21X1 OAI21X1_184 ( .A(u0__abc_74894_new_n1190_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2472_));
OAI21X1 OAI21X1_185 ( .A(u0__abc_74894_new_n2472_), .B(u0__abc_74894_new_n2471_), .C(u0__abc_74894_new_n2473_), .Y(u0__abc_74894_new_n2474_));
OAI21X1 OAI21X1_186 ( .A(u0__abc_74894_new_n1210_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2488_));
OAI21X1 OAI21X1_187 ( .A(u0__abc_74894_new_n2488_), .B(u0__abc_74894_new_n2487_), .C(u0__abc_74894_new_n2489_), .Y(u0__abc_74894_new_n2490_));
OAI21X1 OAI21X1_188 ( .A(u0__abc_74894_new_n1230_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2504_));
OAI21X1 OAI21X1_189 ( .A(u0__abc_74894_new_n2504_), .B(u0__abc_74894_new_n2503_), .C(u0__abc_74894_new_n2505_), .Y(u0__abc_74894_new_n2506_));
OAI21X1 OAI21X1_19 ( .A(susp_sel), .B(rfr_ack), .C(cs_need_rfr_6_), .Y(_abc_81086_new_n264_));
OAI21X1 OAI21X1_190 ( .A(u0__abc_74894_new_n1250_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2520_));
OAI21X1 OAI21X1_191 ( .A(u0__abc_74894_new_n2520_), .B(u0__abc_74894_new_n2519_), .C(u0__abc_74894_new_n2521_), .Y(u0__abc_74894_new_n2522_));
OAI21X1 OAI21X1_192 ( .A(u0__abc_74894_new_n1270_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2536_));
OAI21X1 OAI21X1_193 ( .A(u0__abc_74894_new_n2536_), .B(u0__abc_74894_new_n2535_), .C(u0__abc_74894_new_n2537_), .Y(u0__abc_74894_new_n2538_));
OAI21X1 OAI21X1_194 ( .A(u0__abc_74894_new_n1290_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2552_));
OAI21X1 OAI21X1_195 ( .A(u0__abc_74894_new_n2552_), .B(u0__abc_74894_new_n2551_), .C(u0__abc_74894_new_n2553_), .Y(u0__abc_74894_new_n2554_));
OAI21X1 OAI21X1_196 ( .A(u0__abc_74894_new_n1310_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2568_));
OAI21X1 OAI21X1_197 ( .A(u0__abc_74894_new_n2568_), .B(u0__abc_74894_new_n2567_), .C(u0__abc_74894_new_n2569_), .Y(u0__abc_74894_new_n2570_));
OAI21X1 OAI21X1_198 ( .A(u0__abc_74894_new_n1330_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2584_));
OAI21X1 OAI21X1_199 ( .A(u0__abc_74894_new_n2584_), .B(u0__abc_74894_new_n2583_), .C(u0__abc_74894_new_n2585_), .Y(u0__abc_74894_new_n2586_));
OAI21X1 OAI21X1_2 ( .A(spec_req_cs_0_), .B(_abc_81086_new_n236_), .C(_abc_81086_new_n240_), .Y(_abc_81086_new_n241_));
OAI21X1 OAI21X1_20 ( .A(spec_req_cs_6_), .B(_abc_81086_new_n236_), .C(_abc_81086_new_n240_), .Y(_abc_81086_new_n265_));
OAI21X1 OAI21X1_200 ( .A(u0__abc_74894_new_n1350_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2600_));
OAI21X1 OAI21X1_201 ( .A(u0__abc_74894_new_n2600_), .B(u0__abc_74894_new_n2599_), .C(u0__abc_74894_new_n2601_), .Y(u0__abc_74894_new_n2602_));
OAI21X1 OAI21X1_202 ( .A(u0__abc_74894_new_n1370_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2616_));
OAI21X1 OAI21X1_203 ( .A(u0__abc_74894_new_n2616_), .B(u0__abc_74894_new_n2615_), .C(u0__abc_74894_new_n2617_), .Y(u0__abc_74894_new_n2618_));
OAI21X1 OAI21X1_204 ( .A(u0__abc_74894_new_n1390_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2632_));
OAI21X1 OAI21X1_205 ( .A(u0__abc_74894_new_n2632_), .B(u0__abc_74894_new_n2631_), .C(u0__abc_74894_new_n2633_), .Y(u0__abc_74894_new_n2634_));
OAI21X1 OAI21X1_206 ( .A(u0__abc_74894_new_n1410_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2648_));
OAI21X1 OAI21X1_207 ( .A(u0__abc_74894_new_n2648_), .B(u0__abc_74894_new_n2647_), .C(u0__abc_74894_new_n2649_), .Y(u0__abc_74894_new_n2650_));
OAI21X1 OAI21X1_208 ( .A(u0__abc_74894_new_n1430_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2664_));
OAI21X1 OAI21X1_209 ( .A(u0__abc_74894_new_n2664_), .B(u0__abc_74894_new_n2663_), .C(u0__abc_74894_new_n2665_), .Y(u0__abc_74894_new_n2666_));
OAI21X1 OAI21X1_21 ( .A(_abc_81086_new_n263_), .B(_abc_81086_new_n265_), .C(_abc_81086_new_n264_), .Y(obct_cs_6_));
OAI21X1 OAI21X1_210 ( .A(u0__abc_74894_new_n1450_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2680_));
OAI21X1 OAI21X1_211 ( .A(u0__abc_74894_new_n2680_), .B(u0__abc_74894_new_n2679_), .C(u0__abc_74894_new_n2681_), .Y(u0__abc_74894_new_n2682_));
OAI21X1 OAI21X1_212 ( .A(u0__abc_74894_new_n1470_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2696_));
OAI21X1 OAI21X1_213 ( .A(u0__abc_74894_new_n2696_), .B(u0__abc_74894_new_n2695_), .C(u0__abc_74894_new_n2697_), .Y(u0__abc_74894_new_n2698_));
OAI21X1 OAI21X1_214 ( .A(u0__abc_74894_new_n1490_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2712_));
OAI21X1 OAI21X1_215 ( .A(u0__abc_74894_new_n2712_), .B(u0__abc_74894_new_n2711_), .C(u0__abc_74894_new_n2713_), .Y(u0__abc_74894_new_n2714_));
OAI21X1 OAI21X1_216 ( .A(u0__abc_74894_new_n1510_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2728_));
OAI21X1 OAI21X1_217 ( .A(u0__abc_74894_new_n2728_), .B(u0__abc_74894_new_n2727_), .C(u0__abc_74894_new_n2729_), .Y(u0__abc_74894_new_n2730_));
OAI21X1 OAI21X1_218 ( .A(u0__abc_74894_new_n1530_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2744_));
OAI21X1 OAI21X1_219 ( .A(u0__abc_74894_new_n2744_), .B(u0__abc_74894_new_n2743_), .C(u0__abc_74894_new_n2745_), .Y(u0__abc_74894_new_n2746_));
OAI21X1 OAI21X1_22 ( .A(susp_sel), .B(rfr_ack), .C(cs_need_rfr_7_), .Y(_abc_81086_new_n268_));
OAI21X1 OAI21X1_220 ( .A(u0__abc_74894_new_n1550_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2760_));
OAI21X1 OAI21X1_221 ( .A(u0__abc_74894_new_n2760_), .B(u0__abc_74894_new_n2759_), .C(u0__abc_74894_new_n2761_), .Y(u0__abc_74894_new_n2762_));
OAI21X1 OAI21X1_222 ( .A(u0__abc_74894_new_n1570_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2776_));
OAI21X1 OAI21X1_223 ( .A(u0__abc_74894_new_n2776_), .B(u0__abc_74894_new_n2775_), .C(u0__abc_74894_new_n2777_), .Y(u0__abc_74894_new_n2778_));
OAI21X1 OAI21X1_224 ( .A(u0__abc_74894_new_n1590_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2792_));
OAI21X1 OAI21X1_225 ( .A(u0__abc_74894_new_n2792_), .B(u0__abc_74894_new_n2791_), .C(u0__abc_74894_new_n2793_), .Y(u0__abc_74894_new_n2794_));
OAI21X1 OAI21X1_226 ( .A(u0__abc_74894_new_n1610_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2808_));
OAI21X1 OAI21X1_227 ( .A(u0__abc_74894_new_n2808_), .B(u0__abc_74894_new_n2807_), .C(u0__abc_74894_new_n2809_), .Y(u0__abc_74894_new_n2810_));
OAI21X1 OAI21X1_228 ( .A(u0__abc_74894_new_n1630_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2824_));
OAI21X1 OAI21X1_229 ( .A(u0__abc_74894_new_n2824_), .B(u0__abc_74894_new_n2823_), .C(u0__abc_74894_new_n2825_), .Y(u0__abc_74894_new_n2826_));
OAI21X1 OAI21X1_23 ( .A(spec_req_cs_7_), .B(_abc_81086_new_n236_), .C(_abc_81086_new_n240_), .Y(_abc_81086_new_n269_));
OAI21X1 OAI21X1_230 ( .A(u0__abc_74894_new_n1650_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2840_));
OAI21X1 OAI21X1_231 ( .A(u0__abc_74894_new_n2840_), .B(u0__abc_74894_new_n2839_), .C(u0__abc_74894_new_n2841_), .Y(u0__abc_74894_new_n2842_));
OAI21X1 OAI21X1_232 ( .A(u0__abc_74894_new_n1670_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2856_));
OAI21X1 OAI21X1_233 ( .A(u0__abc_74894_new_n2856_), .B(u0__abc_74894_new_n2855_), .C(u0__abc_74894_new_n2857_), .Y(u0__abc_74894_new_n2858_));
OAI21X1 OAI21X1_234 ( .A(u0__abc_74894_new_n1690_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2872_));
OAI21X1 OAI21X1_235 ( .A(u0__abc_74894_new_n2872_), .B(u0__abc_74894_new_n2871_), .C(u0__abc_74894_new_n2873_), .Y(u0__abc_74894_new_n2874_));
OAI21X1 OAI21X1_236 ( .A(u0__abc_74894_new_n1710_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2888_));
OAI21X1 OAI21X1_237 ( .A(u0__abc_74894_new_n2888_), .B(u0__abc_74894_new_n2887_), .C(u0__abc_74894_new_n2889_), .Y(u0__abc_74894_new_n2890_));
OAI21X1 OAI21X1_238 ( .A(u0__abc_74894_new_n1831_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n2985_));
OAI21X1 OAI21X1_239 ( .A(u0_csc0_1_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n2987_));
OAI21X1 OAI21X1_24 ( .A(_abc_81086_new_n267_), .B(_abc_81086_new_n269_), .C(_abc_81086_new_n268_), .Y(obct_cs_7_));
OAI21X1 OAI21X1_240 ( .A(u0__abc_74894_new_n2987_), .B(u0__abc_74894_new_n2986_), .C(u0__abc_74894_new_n2973_), .Y(u0__0csc_31_0__1_));
OAI21X1 OAI21X1_241 ( .A(u0__abc_74894_new_n1851_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3001_));
OAI21X1 OAI21X1_242 ( .A(u0_csc0_2_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3003_));
OAI21X1 OAI21X1_243 ( .A(u0__abc_74894_new_n3003_), .B(u0__abc_74894_new_n3002_), .C(u0__abc_74894_new_n2989_), .Y(u0__0csc_31_0__2_));
OAI21X1 OAI21X1_244 ( .A(u0__abc_74894_new_n1871_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3017_));
OAI21X1 OAI21X1_245 ( .A(u0_csc0_3_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3019_));
OAI21X1 OAI21X1_246 ( .A(u0__abc_74894_new_n3019_), .B(u0__abc_74894_new_n3018_), .C(u0__abc_74894_new_n3005_), .Y(u0__0csc_31_0__3_));
OAI21X1 OAI21X1_247 ( .A(u0__abc_74894_new_n1891_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3033_));
OAI21X1 OAI21X1_248 ( .A(u0_csc0_4_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3035_));
OAI21X1 OAI21X1_249 ( .A(u0__abc_74894_new_n3035_), .B(u0__abc_74894_new_n3034_), .C(u0__abc_74894_new_n3021_), .Y(u0__0csc_31_0__4_));
OAI21X1 OAI21X1_25 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_0_), .Y(_abc_81086_new_n272_));
OAI21X1 OAI21X1_250 ( .A(u0__abc_74894_new_n1911_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3049_));
OAI21X1 OAI21X1_251 ( .A(u0_csc0_5_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3051_));
OAI21X1 OAI21X1_252 ( .A(u0__abc_74894_new_n3051_), .B(u0__abc_74894_new_n3050_), .C(u0__abc_74894_new_n3037_), .Y(u0__0csc_31_0__5_));
OAI21X1 OAI21X1_253 ( .A(u0__abc_74894_new_n1931_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3065_));
OAI21X1 OAI21X1_254 ( .A(u0_csc0_6_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3067_));
OAI21X1 OAI21X1_255 ( .A(u0__abc_74894_new_n3067_), .B(u0__abc_74894_new_n3066_), .C(u0__abc_74894_new_n3053_), .Y(u0__0csc_31_0__6_));
OAI21X1 OAI21X1_256 ( .A(u0__abc_74894_new_n1951_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3081_));
OAI21X1 OAI21X1_257 ( .A(u0_csc0_7_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3083_));
OAI21X1 OAI21X1_258 ( .A(u0__abc_74894_new_n3083_), .B(u0__abc_74894_new_n3082_), .C(u0__abc_74894_new_n3069_), .Y(u0__0csc_31_0__7_));
OAI21X1 OAI21X1_259 ( .A(u0__abc_74894_new_n1991_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3113_));
OAI21X1 OAI21X1_26 ( .A(_abc_81086_new_n271_), .B(lmr_sel), .C(_abc_81086_new_n272_), .Y(tms_s_0_));
OAI21X1 OAI21X1_260 ( .A(u0_csc0_9_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3115_));
OAI21X1 OAI21X1_261 ( .A(u0__abc_74894_new_n3115_), .B(u0__abc_74894_new_n3114_), .C(u0__abc_74894_new_n3101_), .Y(u0__0csc_31_0__9_));
OAI21X1 OAI21X1_262 ( .A(u0__abc_74894_new_n2011_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3129_));
OAI21X1 OAI21X1_263 ( .A(u0_csc0_10_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3131_));
OAI21X1 OAI21X1_264 ( .A(u0__abc_74894_new_n3131_), .B(u0__abc_74894_new_n3130_), .C(u0__abc_74894_new_n3117_), .Y(u0__0csc_31_0__10_));
OAI21X1 OAI21X1_265 ( .A(u0__abc_74894_new_n2031_), .B(u0__abc_74894_new_n2454_), .C(u0__abc_74894_new_n2455_), .Y(u0__abc_74894_new_n3145_));
OAI21X1 OAI21X1_266 ( .A(u0_csc0_11_), .B(u0__abc_74894_new_n2455_), .C(u0__abc_74894_new_n2970_), .Y(u0__abc_74894_new_n3147_));
OAI21X1 OAI21X1_267 ( .A(u0__abc_74894_new_n3147_), .B(u0__abc_74894_new_n3146_), .C(u0__abc_74894_new_n3133_), .Y(u0__0csc_31_0__11_));
OAI21X1 OAI21X1_268 ( .A(u0__abc_74894_new_n3471_), .B(u0__abc_74894_new_n3475_), .C(u0__abc_74894_new_n3470_), .Y(u0__abc_74894_new_n3476_));
OAI21X1 OAI21X1_269 ( .A(u0__abc_74894_new_n3470_), .B(u0__abc_74894_new_n3477_), .C(u0__abc_74894_new_n3476_), .Y(u0__0wp_err_0_0_));
OAI21X1 OAI21X1_27 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_1_), .Y(_abc_81086_new_n275_));
OAI21X1 OAI21X1_270 ( .A(cs_le), .B(u0__abc_74894_new_n3493_), .C(u0__abc_74894_new_n3494_), .Y(u0__0cs_7_0__7_));
OAI21X1 OAI21X1_271 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3496_), .C(u0__abc_74894_new_n3497_), .Y(u0__0poc_31_0__0_));
OAI21X1 OAI21X1_272 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3499_), .C(u0__abc_74894_new_n3500_), .Y(u0__0poc_31_0__1_));
OAI21X1 OAI21X1_273 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3502_), .C(u0__abc_74894_new_n3503_), .Y(u0__0poc_31_0__2_));
OAI21X1 OAI21X1_274 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3505_), .C(u0__abc_74894_new_n3506_), .Y(u0__0poc_31_0__3_));
OAI21X1 OAI21X1_275 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3508_), .C(u0__abc_74894_new_n3509_), .Y(u0__0poc_31_0__4_));
OAI21X1 OAI21X1_276 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3511_), .C(u0__abc_74894_new_n3512_), .Y(u0__0poc_31_0__5_));
OAI21X1 OAI21X1_277 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3514_), .C(u0__abc_74894_new_n3515_), .Y(u0__0poc_31_0__6_));
OAI21X1 OAI21X1_278 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3517_), .C(u0__abc_74894_new_n3518_), .Y(u0__0poc_31_0__7_));
OAI21X1 OAI21X1_279 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3520_), .C(u0__abc_74894_new_n3521_), .Y(u0__0poc_31_0__8_));
OAI21X1 OAI21X1_28 ( .A(_abc_81086_new_n274_), .B(lmr_sel), .C(_abc_81086_new_n275_), .Y(tms_s_1_));
OAI21X1 OAI21X1_280 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3523_), .C(u0__abc_74894_new_n3524_), .Y(u0__0poc_31_0__9_));
OAI21X1 OAI21X1_281 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3526_), .C(u0__abc_74894_new_n3527_), .Y(u0__0poc_31_0__10_));
OAI21X1 OAI21X1_282 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3529_), .C(u0__abc_74894_new_n3530_), .Y(u0__0poc_31_0__11_));
OAI21X1 OAI21X1_283 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3532_), .C(u0__abc_74894_new_n3533_), .Y(u0__0poc_31_0__12_));
OAI21X1 OAI21X1_284 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3535_), .C(u0__abc_74894_new_n3536_), .Y(u0__0poc_31_0__13_));
OAI21X1 OAI21X1_285 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3538_), .C(u0__abc_74894_new_n3539_), .Y(u0__0poc_31_0__14_));
OAI21X1 OAI21X1_286 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3541_), .C(u0__abc_74894_new_n3542_), .Y(u0__0poc_31_0__15_));
OAI21X1 OAI21X1_287 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3544_), .C(u0__abc_74894_new_n3545_), .Y(u0__0poc_31_0__16_));
OAI21X1 OAI21X1_288 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3547_), .C(u0__abc_74894_new_n3548_), .Y(u0__0poc_31_0__17_));
OAI21X1 OAI21X1_289 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3550_), .C(u0__abc_74894_new_n3551_), .Y(u0__0poc_31_0__18_));
OAI21X1 OAI21X1_29 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_2_), .Y(_abc_81086_new_n278_));
OAI21X1 OAI21X1_290 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3553_), .C(u0__abc_74894_new_n3554_), .Y(u0__0poc_31_0__19_));
OAI21X1 OAI21X1_291 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3556_), .C(u0__abc_74894_new_n3557_), .Y(u0__0poc_31_0__20_));
OAI21X1 OAI21X1_292 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3559_), .C(u0__abc_74894_new_n3560_), .Y(u0__0poc_31_0__21_));
OAI21X1 OAI21X1_293 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3562_), .C(u0__abc_74894_new_n3563_), .Y(u0__0poc_31_0__22_));
OAI21X1 OAI21X1_294 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3565_), .C(u0__abc_74894_new_n3566_), .Y(u0__0poc_31_0__23_));
OAI21X1 OAI21X1_295 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3568_), .C(u0__abc_74894_new_n3569_), .Y(u0__0poc_31_0__24_));
OAI21X1 OAI21X1_296 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3571_), .C(u0__abc_74894_new_n3572_), .Y(u0__0poc_31_0__25_));
OAI21X1 OAI21X1_297 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3574_), .C(u0__abc_74894_new_n3575_), .Y(u0__0poc_31_0__26_));
OAI21X1 OAI21X1_298 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3577_), .C(u0__abc_74894_new_n3578_), .Y(u0__0poc_31_0__27_));
OAI21X1 OAI21X1_299 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3580_), .C(u0__abc_74894_new_n3581_), .Y(u0__0poc_31_0__28_));
OAI21X1 OAI21X1_3 ( .A(_abc_81086_new_n238_), .B(_abc_81086_new_n241_), .C(_abc_81086_new_n239_), .Y(obct_cs_0_));
OAI21X1 OAI21X1_30 ( .A(_abc_81086_new_n277_), .B(lmr_sel), .C(_abc_81086_new_n278_), .Y(tms_s_2_));
OAI21X1 OAI21X1_300 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3583_), .C(u0__abc_74894_new_n3584_), .Y(u0__0poc_31_0__29_));
OAI21X1 OAI21X1_301 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3586_), .C(u0__abc_74894_new_n3587_), .Y(u0__0poc_31_0__30_));
OAI21X1 OAI21X1_302 ( .A(u0_rst_r3), .B(u0__abc_74894_new_n3589_), .C(u0__abc_74894_new_n3590_), .Y(u0__0poc_31_0__31_));
OAI21X1 OAI21X1_303 ( .A(u0__abc_74894_new_n3592_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3599_), .Y(u0__0csc_mask_r_10_0__0_));
OAI21X1 OAI21X1_304 ( .A(u0__abc_74894_new_n3601_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3602_), .Y(u0__0csc_mask_r_10_0__1_));
OAI21X1 OAI21X1_305 ( .A(u0__abc_74894_new_n3604_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3605_), .Y(u0__0csc_mask_r_10_0__2_));
OAI21X1 OAI21X1_306 ( .A(u0__abc_74894_new_n3607_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3608_), .Y(u0__0csc_mask_r_10_0__3_));
OAI21X1 OAI21X1_307 ( .A(u0__abc_74894_new_n3610_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3611_), .Y(u0__0csc_mask_r_10_0__4_));
OAI21X1 OAI21X1_308 ( .A(u0__abc_74894_new_n3613_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3614_), .Y(u0__0csc_mask_r_10_0__5_));
OAI21X1 OAI21X1_309 ( .A(u0__abc_74894_new_n3616_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3617_), .Y(u0__0csc_mask_r_10_0__6_));
OAI21X1 OAI21X1_31 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_3_), .Y(_abc_81086_new_n281_));
OAI21X1 OAI21X1_310 ( .A(u0__abc_74894_new_n3619_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3620_), .Y(u0__0csc_mask_r_10_0__7_));
OAI21X1 OAI21X1_311 ( .A(u0__abc_74894_new_n3622_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3623_), .Y(u0__0csc_mask_r_10_0__8_));
OAI21X1 OAI21X1_312 ( .A(u0__abc_74894_new_n3625_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3626_), .Y(u0__0csc_mask_r_10_0__9_));
OAI21X1 OAI21X1_313 ( .A(u0__abc_74894_new_n3628_), .B(u0__abc_74894_new_n3598_), .C(u0__abc_74894_new_n3629_), .Y(u0__0csc_mask_r_10_0__10_));
OAI21X1 OAI21X1_314 ( .A(u0__abc_74894_new_n3631_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3635_), .Y(u0__0csr_r_10_1__0_));
OAI21X1 OAI21X1_315 ( .A(u0__abc_74894_new_n3637_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3638_), .Y(u0__0csr_r_10_1__1_));
OAI21X1 OAI21X1_316 ( .A(u0__abc_74894_new_n3640_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3641_), .Y(u0__0csr_r_10_1__2_));
OAI21X1 OAI21X1_317 ( .A(u0__abc_74894_new_n3643_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3644_), .Y(u0__0csr_r_10_1__3_));
OAI21X1 OAI21X1_318 ( .A(u0__abc_74894_new_n3646_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3647_), .Y(u0__0csr_r_10_1__4_));
OAI21X1 OAI21X1_319 ( .A(u0__abc_74894_new_n3649_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3650_), .Y(u0__0csr_r_10_1__5_));
OAI21X1 OAI21X1_32 ( .A(_abc_81086_new_n280_), .B(lmr_sel), .C(_abc_81086_new_n281_), .Y(tms_s_3_));
OAI21X1 OAI21X1_320 ( .A(u0__abc_74894_new_n3652_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3653_), .Y(u0__0csr_r_10_1__6_));
OAI21X1 OAI21X1_321 ( .A(u0__abc_74894_new_n3655_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3656_), .Y(u0__0csr_r_10_1__7_));
OAI21X1 OAI21X1_322 ( .A(u0__abc_74894_new_n3658_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3659_), .Y(u0__0csr_r_10_1__8_));
OAI21X1 OAI21X1_323 ( .A(u0__abc_74894_new_n3661_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3662_), .Y(u0__0csr_r_10_1__9_));
OAI21X1 OAI21X1_324 ( .A(u0__abc_74894_new_n3664_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3665_), .Y(u0__0csr_r2_7_0__0_));
OAI21X1 OAI21X1_325 ( .A(u0__abc_74894_new_n3667_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3668_), .Y(u0__0csr_r2_7_0__1_));
OAI21X1 OAI21X1_326 ( .A(u0__abc_74894_new_n3670_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3671_), .Y(u0__0csr_r2_7_0__2_));
OAI21X1 OAI21X1_327 ( .A(u0__abc_74894_new_n3673_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3674_), .Y(u0__0csr_r2_7_0__3_));
OAI21X1 OAI21X1_328 ( .A(u0__abc_74894_new_n3676_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3677_), .Y(u0__0csr_r2_7_0__4_));
OAI21X1 OAI21X1_329 ( .A(u0__abc_74894_new_n3679_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3680_), .Y(u0__0csr_r2_7_0__5_));
OAI21X1 OAI21X1_33 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_4_), .Y(_abc_81086_new_n284_));
OAI21X1 OAI21X1_330 ( .A(u0__abc_74894_new_n3682_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3683_), .Y(u0__0csr_r2_7_0__6_));
OAI21X1 OAI21X1_331 ( .A(u0__abc_74894_new_n3685_), .B(u0__abc_74894_new_n3634_), .C(u0__abc_74894_new_n3686_), .Y(u0__0csr_r2_7_0__7_));
OAI21X1 OAI21X1_332 ( .A(u0__abc_74894_new_n3725_), .B(u0__abc_74894_new_n3726_), .C(u0__abc_74894_new_n3727_), .Y(u0__abc_74894_new_n3728_));
OAI21X1 OAI21X1_333 ( .A(u0__abc_74894_new_n3724_), .B(u0__abc_74894_new_n3688_), .C(u0__abc_74894_new_n3728_), .Y(u0__abc_74894_new_n3729_));
OAI21X1 OAI21X1_334 ( .A(u0__abc_74894_new_n1811_), .B(u0__abc_74894_new_n3732_), .C(u0__abc_74894_new_n3738_), .Y(u0__abc_74894_new_n3739_));
OAI21X1 OAI21X1_335 ( .A(u0__abc_74894_new_n1170_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n3752_), .Y(u0__abc_74894_new_n3753_));
OAI21X1 OAI21X1_336 ( .A(u0__abc_74894_new_n3764_), .B(u0__abc_74894_new_n3765_), .C(u0__abc_74894_new_n3766_), .Y(u0__abc_74894_new_n3767_));
OAI21X1 OAI21X1_337 ( .A(\wb_addr_i[5] ), .B(\wb_addr_i[4] ), .C(\wb_addr_i[6] ), .Y(u0__abc_74894_new_n3769_));
OAI21X1 OAI21X1_338 ( .A(u0__abc_74894_new_n1190_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n3772_), .Y(u0__abc_74894_new_n3773_));
OAI21X1 OAI21X1_339 ( .A(u0__abc_74894_new_n1831_), .B(u0__abc_74894_new_n3732_), .C(u0__abc_74894_new_n3774_), .Y(u0__abc_74894_new_n3775_));
OAI21X1 OAI21X1_34 ( .A(_abc_81086_new_n283_), .B(lmr_sel), .C(_abc_81086_new_n284_), .Y(tms_s_4_));
OAI21X1 OAI21X1_340 ( .A(u0__abc_74894_new_n3785_), .B(u0__abc_74894_new_n3765_), .C(u0__abc_74894_new_n3786_), .Y(u0__abc_74894_new_n3787_));
OAI21X1 OAI21X1_341 ( .A(u0__abc_74894_new_n1210_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n3791_), .Y(u0__abc_74894_new_n3792_));
OAI21X1 OAI21X1_342 ( .A(u0__abc_74894_new_n1851_), .B(u0__abc_74894_new_n3732_), .C(u0__abc_74894_new_n3793_), .Y(u0__abc_74894_new_n3794_));
OAI21X1 OAI21X1_343 ( .A(u0__abc_74894_new_n3797_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n3799_), .Y(u0__abc_74894_new_n3800_));
OAI21X1 OAI21X1_344 ( .A(u0__abc_74894_new_n1878_), .B(u0__abc_74894_new_n3707_), .C(u0__abc_74894_new_n3830_), .Y(u0__abc_74894_new_n3831_));
OAI21X1 OAI21X1_345 ( .A(u0__abc_74894_new_n1250_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n3834_), .Y(u0__abc_74894_new_n3835_));
OAI21X1 OAI21X1_346 ( .A(u0__abc_74894_new_n1891_), .B(u0__abc_74894_new_n3732_), .C(u0__abc_74894_new_n3836_), .Y(u0__abc_74894_new_n3837_));
OAI21X1 OAI21X1_347 ( .A(u0__abc_74894_new_n3840_), .B(u0__abc_74894_new_n3765_), .C(u0__abc_74894_new_n3841_), .Y(u0__abc_74894_new_n3842_));
OAI21X1 OAI21X1_348 ( .A(u0__abc_74894_new_n1259_), .B(u0__abc_74894_new_n3719_), .C(u0__abc_74894_new_n3843_), .Y(u0__abc_74894_new_n3844_));
OAI21X1 OAI21X1_349 ( .A(u0__abc_74894_new_n3613_), .B(u0__abc_74894_new_n3845_), .C(u0__abc_74894_new_n3846_), .Y(u0__abc_74894_new_n3847_));
OAI21X1 OAI21X1_35 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_5_), .Y(_abc_81086_new_n287_));
OAI21X1 OAI21X1_350 ( .A(u0__abc_74894_new_n1918_), .B(u0__abc_74894_new_n3707_), .C(u0__abc_74894_new_n3871_), .Y(u0__abc_74894_new_n3872_));
OAI21X1 OAI21X1_351 ( .A(u0__abc_74894_new_n1290_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n3875_), .Y(u0__abc_74894_new_n3876_));
OAI21X1 OAI21X1_352 ( .A(u0__abc_74894_new_n1931_), .B(u0__abc_74894_new_n3732_), .C(u0__abc_74894_new_n3877_), .Y(u0__abc_74894_new_n3878_));
OAI21X1 OAI21X1_353 ( .A(u0__abc_74894_new_n3652_), .B(u0__abc_74894_new_n3770_), .C(u0__abc_74894_new_n3891_), .Y(u0__abc_74894_new_n3892_));
OAI21X1 OAI21X1_354 ( .A(u0__abc_74894_new_n1958_), .B(u0__abc_74894_new_n3707_), .C(u0__abc_74894_new_n3908_), .Y(u0__abc_74894_new_n3909_));
OAI21X1 OAI21X1_355 ( .A(u0__abc_74894_new_n3918_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n3919_), .Y(u0__abc_74894_new_n3920_));
OAI21X1 OAI21X1_356 ( .A(u0__abc_74894_new_n1998_), .B(u0__abc_74894_new_n3707_), .C(u0__abc_74894_new_n3947_), .Y(u0__abc_74894_new_n3948_));
OAI21X1 OAI21X1_357 ( .A(u0__abc_74894_new_n1370_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n3951_), .Y(u0__abc_74894_new_n3952_));
OAI21X1 OAI21X1_358 ( .A(u0__abc_74894_new_n2011_), .B(u0__abc_74894_new_n3732_), .C(u0__abc_74894_new_n3953_), .Y(u0__abc_74894_new_n3954_));
OAI21X1 OAI21X1_359 ( .A(u0__abc_74894_new_n4001_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n4002_), .Y(u0__abc_74894_new_n4003_));
OAI21X1 OAI21X1_36 ( .A(_abc_81086_new_n286_), .B(lmr_sel), .C(_abc_81086_new_n287_), .Y(tms_s_5_));
OAI21X1 OAI21X1_360 ( .A(u0__abc_74894_new_n3535_), .B(u0__abc_74894_new_n3750_), .C(u0__abc_74894_new_n4005_), .Y(u0__abc_74894_new_n4006_));
OAI21X1 OAI21X1_361 ( .A(u0__abc_74894_new_n2058_), .B(u0__abc_74894_new_n3707_), .C(u0__abc_74894_new_n4009_), .Y(u0__abc_74894_new_n4010_));
OAI21X1 OAI21X1_362 ( .A(u0__abc_74894_new_n4023_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n4024_), .Y(u0__abc_74894_new_n4025_));
OAI21X1 OAI21X1_363 ( .A(u0__abc_74894_new_n3538_), .B(u0__abc_74894_new_n3750_), .C(u0__abc_74894_new_n4027_), .Y(u0__abc_74894_new_n4028_));
OAI21X1 OAI21X1_364 ( .A(u0__abc_74894_new_n2078_), .B(u0__abc_74894_new_n3707_), .C(u0__abc_74894_new_n4031_), .Y(u0__abc_74894_new_n4032_));
OAI21X1 OAI21X1_365 ( .A(u0__abc_74894_new_n1457_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n4039_), .Y(u0__abc_74894_new_n4040_));
OAI21X1 OAI21X1_366 ( .A(u0__abc_74894_new_n1470_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n4043_), .Y(u0__abc_74894_new_n4044_));
OAI21X1 OAI21X1_367 ( .A(u0__abc_74894_new_n4052_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n4053_), .Y(u0__abc_74894_new_n4054_));
OAI21X1 OAI21X1_368 ( .A(u0__abc_74894_new_n3541_), .B(u0__abc_74894_new_n3750_), .C(u0__abc_74894_new_n4056_), .Y(u0__abc_74894_new_n4057_));
OAI21X1 OAI21X1_369 ( .A(u0__abc_74894_new_n2133_), .B(u0__abc_74894_new_n3733_), .C(u0__abc_74894_new_n4061_), .Y(u0__abc_74894_new_n4062_));
OAI21X1 OAI21X1_37 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_6_), .Y(_abc_81086_new_n290_));
OAI21X1 OAI21X1_370 ( .A(u0__abc_74894_new_n1492_), .B(u0__abc_74894_new_n3736_), .C(u0__abc_74894_new_n4068_), .Y(u0__abc_74894_new_n4069_));
OAI21X1 OAI21X1_371 ( .A(u0__abc_74894_new_n1497_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n4081_), .Y(u0__abc_74894_new_n4082_));
OAI21X1 OAI21X1_372 ( .A(u0__abc_74894_new_n1510_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n4085_), .Y(u0__abc_74894_new_n4086_));
OAI21X1 OAI21X1_373 ( .A(u0__abc_74894_new_n4094_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n4095_), .Y(u0__abc_74894_new_n4096_));
OAI21X1 OAI21X1_374 ( .A(u0__abc_74894_new_n3547_), .B(u0__abc_74894_new_n3750_), .C(u0__abc_74894_new_n4098_), .Y(u0__abc_74894_new_n4099_));
OAI21X1 OAI21X1_375 ( .A(u0__abc_74894_new_n1517_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n4103_), .Y(u0__abc_74894_new_n4104_));
OAI21X1 OAI21X1_376 ( .A(u0__abc_74894_new_n1530_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n4107_), .Y(u0__abc_74894_new_n4108_));
OAI21X1 OAI21X1_377 ( .A(u0__abc_74894_new_n4116_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n4117_), .Y(u0__abc_74894_new_n4118_));
OAI21X1 OAI21X1_378 ( .A(u0__abc_74894_new_n3550_), .B(u0__abc_74894_new_n3750_), .C(u0__abc_74894_new_n4120_), .Y(u0__abc_74894_new_n4121_));
OAI21X1 OAI21X1_379 ( .A(u0__abc_74894_new_n4131_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n4132_), .Y(u0__abc_74894_new_n4133_));
OAI21X1 OAI21X1_38 ( .A(_abc_81086_new_n289_), .B(lmr_sel), .C(_abc_81086_new_n290_), .Y(tms_s_6_));
OAI21X1 OAI21X1_380 ( .A(u0__abc_74894_new_n3553_), .B(u0__abc_74894_new_n3750_), .C(u0__abc_74894_new_n4135_), .Y(u0__abc_74894_new_n4136_));
OAI21X1 OAI21X1_381 ( .A(u0__abc_74894_new_n2178_), .B(u0__abc_74894_new_n3707_), .C(u0__abc_74894_new_n4139_), .Y(u0__abc_74894_new_n4140_));
OAI21X1 OAI21X1_382 ( .A(u0__abc_74894_new_n1579_), .B(u0__abc_74894_new_n3719_), .C(u0__abc_74894_new_n4170_), .Y(u0__abc_74894_new_n4171_));
OAI21X1 OAI21X1_383 ( .A(u0__abc_74894_new_n4173_), .B(u0__abc_74894_new_n3798_), .C(u0__abc_74894_new_n4174_), .Y(u0__abc_74894_new_n4175_));
OAI21X1 OAI21X1_384 ( .A(u0__abc_74894_new_n3559_), .B(u0__abc_74894_new_n3750_), .C(u0__abc_74894_new_n4177_), .Y(u0__abc_74894_new_n4178_));
OAI21X1 OAI21X1_385 ( .A(u0__abc_74894_new_n2218_), .B(u0__abc_74894_new_n3707_), .C(u0__abc_74894_new_n4181_), .Y(u0__abc_74894_new_n4182_));
OAI21X1 OAI21X1_386 ( .A(u0__abc_74894_new_n2273_), .B(u0__abc_74894_new_n3733_), .C(u0__abc_74894_new_n4208_), .Y(u0__abc_74894_new_n4209_));
OAI21X1 OAI21X1_387 ( .A(u0__abc_74894_new_n1632_), .B(u0__abc_74894_new_n3736_), .C(u0__abc_74894_new_n4215_), .Y(u0__abc_74894_new_n4216_));
OAI21X1 OAI21X1_388 ( .A(u0__abc_74894_new_n1637_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n4250_), .Y(u0__abc_74894_new_n4251_));
OAI21X1 OAI21X1_389 ( .A(u0__abc_74894_new_n4272_), .B(u0__abc_74894_new_n4273_), .C(u0__abc_74894_new_n4274_), .Y(u0__abc_74894_new_n4275_));
OAI21X1 OAI21X1_39 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_7_), .Y(_abc_81086_new_n293_));
OAI21X1 OAI21X1_390 ( .A(u0__abc_74894_new_n1657_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n4276_), .Y(u0__abc_74894_new_n4277_));
OAI21X1 OAI21X1_391 ( .A(u0__abc_74894_new_n1677_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n4302_), .Y(u0__abc_74894_new_n4303_));
OAI21X1 OAI21X1_392 ( .A(u0__abc_74894_new_n4328_), .B(u0__abc_74894_new_n4273_), .C(u0__abc_74894_new_n4329_), .Y(u0__abc_74894_new_n4330_));
OAI21X1 OAI21X1_393 ( .A(u0__abc_74894_new_n1717_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n4355_), .Y(u0__abc_74894_new_n4356_));
OAI21X1 OAI21X1_394 ( .A(u0_u0__abc_72207_new_n209_), .B(u0_u0__abc_72207_new_n212_), .C(u0_u0__abc_72207_new_n210_), .Y(u0_u0__0lmr_req_0_0_));
OAI21X1 OAI21X1_395 ( .A(\poc_o[3] ), .B(\poc_o[2] ), .C(u0_u0_rst_r2), .Y(u0_u0__abc_72207_new_n330_));
OAI21X1 OAI21X1_396 ( .A(\wb_data_i[1] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n334_));
OAI21X1 OAI21X1_397 ( .A(u0_u0__abc_72207_new_n333_), .B(u0_u0__abc_72207_new_n334_), .C(u0_u0__abc_72207_new_n332_), .Y(u0_u0__0csc_31_0__1_));
OAI21X1 OAI21X1_398 ( .A(\wb_data_i[2] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n338_));
OAI21X1 OAI21X1_399 ( .A(u0_u0__abc_72207_new_n337_), .B(u0_u0__abc_72207_new_n338_), .C(u0_u0__abc_72207_new_n336_), .Y(u0_u0__0csc_31_0__2_));
OAI21X1 OAI21X1_4 ( .A(susp_sel), .B(rfr_ack), .C(cs_need_rfr_1_), .Y(_abc_81086_new_n244_));
OAI21X1 OAI21X1_40 ( .A(_abc_81086_new_n292_), .B(lmr_sel), .C(_abc_81086_new_n293_), .Y(tms_s_7_));
OAI21X1 OAI21X1_400 ( .A(\wb_data_i[3] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n340_));
OAI21X1 OAI21X1_401 ( .A(\wb_data_i[6] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n357_));
OAI21X1 OAI21X1_402 ( .A(\wb_data_i[7] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n360_));
OAI21X1 OAI21X1_403 ( .A(\wb_data_i[8] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n363_));
OAI21X1 OAI21X1_404 ( .A(\wb_data_i[9] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n366_));
OAI21X1 OAI21X1_405 ( .A(\wb_data_i[10] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n369_));
OAI21X1 OAI21X1_406 ( .A(\wb_data_i[11] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n372_));
OAI21X1 OAI21X1_407 ( .A(\wb_data_i[12] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n375_));
OAI21X1 OAI21X1_408 ( .A(\wb_data_i[13] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n378_));
OAI21X1 OAI21X1_409 ( .A(\wb_data_i[14] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n381_));
OAI21X1 OAI21X1_41 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_8_), .Y(_abc_81086_new_n296_));
OAI21X1 OAI21X1_410 ( .A(\wb_data_i[15] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n384_));
OAI21X1 OAI21X1_411 ( .A(\wb_data_i[16] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n387_));
OAI21X1 OAI21X1_412 ( .A(\wb_data_i[17] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n390_));
OAI21X1 OAI21X1_413 ( .A(\wb_data_i[18] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n393_));
OAI21X1 OAI21X1_414 ( .A(\wb_data_i[19] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n396_));
OAI21X1 OAI21X1_415 ( .A(\wb_data_i[20] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n399_));
OAI21X1 OAI21X1_416 ( .A(\wb_data_i[21] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n402_));
OAI21X1 OAI21X1_417 ( .A(\wb_data_i[22] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n405_));
OAI21X1 OAI21X1_418 ( .A(\wb_data_i[23] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n408_));
OAI21X1 OAI21X1_419 ( .A(\wb_data_i[24] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n411_));
OAI21X1 OAI21X1_42 ( .A(_abc_81086_new_n295_), .B(lmr_sel), .C(_abc_81086_new_n296_), .Y(tms_s_8_));
OAI21X1 OAI21X1_420 ( .A(\wb_data_i[25] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n414_));
OAI21X1 OAI21X1_421 ( .A(\wb_data_i[26] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n417_));
OAI21X1 OAI21X1_422 ( .A(\wb_data_i[27] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n420_));
OAI21X1 OAI21X1_423 ( .A(\wb_data_i[28] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n423_));
OAI21X1 OAI21X1_424 ( .A(\wb_data_i[29] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n426_));
OAI21X1 OAI21X1_425 ( .A(\wb_data_i[30] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n429_));
OAI21X1 OAI21X1_426 ( .A(\wb_data_i[31] ), .B(u0_u0__abc_72207_new_n322_), .C(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n432_));
OAI21X1 OAI21X1_427 ( .A(u0_csc0_21_), .B(\wb_addr_i[26] ), .C(u0_csc_mask_5_), .Y(u0_u0__abc_72207_new_n436_));
OAI21X1 OAI21X1_428 ( .A(u0_csc0_19_), .B(\wb_addr_i[24] ), .C(u0_csc_mask_3_), .Y(u0_u0__abc_72207_new_n438_));
OAI21X1 OAI21X1_429 ( .A(u0_csc0_17_), .B(\wb_addr_i[22] ), .C(u0_csc_mask_1_), .Y(u0_u0__abc_72207_new_n441_));
OAI21X1 OAI21X1_43 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_9_), .Y(_abc_81086_new_n299_));
OAI21X1 OAI21X1_430 ( .A(u0_csc0_16_), .B(\wb_addr_i[21] ), .C(u0_csc_mask_0_), .Y(u0_u0__abc_72207_new_n444_));
OAI21X1 OAI21X1_431 ( .A(u0_csc0_18_), .B(\wb_addr_i[23] ), .C(u0_csc_mask_2_), .Y(u0_u0__abc_72207_new_n446_));
OAI21X1 OAI21X1_432 ( .A(u0_csc0_23_), .B(\wb_addr_i[28] ), .C(u0_csc_mask_7_), .Y(u0_u0__abc_72207_new_n450_));
OAI21X1 OAI21X1_433 ( .A(u0_u0__abc_72207_new_n449_), .B(u0_u0__abc_72207_new_n450_), .C(u0_csc0_0_), .Y(u0_u0__abc_72207_new_n451_));
OAI21X1 OAI21X1_434 ( .A(u0_csc0_22_), .B(\wb_addr_i[27] ), .C(u0_csc_mask_6_), .Y(u0_u0__abc_72207_new_n453_));
OAI21X1 OAI21X1_435 ( .A(u0_csc0_20_), .B(\wb_addr_i[25] ), .C(u0_csc_mask_4_), .Y(u0_u0__abc_72207_new_n455_));
OAI21X1 OAI21X1_436 ( .A(u0_u1__abc_72470_new_n205_), .B(u0_u1__abc_72470_new_n208_), .C(u0_u1__abc_72470_new_n206_), .Y(u0_u1__0lmr_req_0_0_));
OAI21X1 OAI21X1_437 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_0_), .Y(u0_u1__abc_72470_new_n219_));
OAI21X1 OAI21X1_438 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_1_), .Y(u0_u1__abc_72470_new_n222_));
OAI21X1 OAI21X1_439 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_2_), .Y(u0_u1__abc_72470_new_n225_));
OAI21X1 OAI21X1_44 ( .A(_abc_81086_new_n298_), .B(lmr_sel), .C(_abc_81086_new_n299_), .Y(tms_s_9_));
OAI21X1 OAI21X1_440 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_3_), .Y(u0_u1__abc_72470_new_n228_));
OAI21X1 OAI21X1_441 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_4_), .Y(u0_u1__abc_72470_new_n231_));
OAI21X1 OAI21X1_442 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_5_), .Y(u0_u1__abc_72470_new_n234_));
OAI21X1 OAI21X1_443 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_6_), .Y(u0_u1__abc_72470_new_n237_));
OAI21X1 OAI21X1_444 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_7_), .Y(u0_u1__abc_72470_new_n240_));
OAI21X1 OAI21X1_445 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_8_), .Y(u0_u1__abc_72470_new_n243_));
OAI21X1 OAI21X1_446 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_9_), .Y(u0_u1__abc_72470_new_n246_));
OAI21X1 OAI21X1_447 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_10_), .Y(u0_u1__abc_72470_new_n249_));
OAI21X1 OAI21X1_448 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_11_), .Y(u0_u1__abc_72470_new_n252_));
OAI21X1 OAI21X1_449 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_12_), .Y(u0_u1__abc_72470_new_n255_));
OAI21X1 OAI21X1_45 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_10_), .Y(_abc_81086_new_n302_));
OAI21X1 OAI21X1_450 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_13_), .Y(u0_u1__abc_72470_new_n258_));
OAI21X1 OAI21X1_451 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_14_), .Y(u0_u1__abc_72470_new_n261_));
OAI21X1 OAI21X1_452 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_15_), .Y(u0_u1__abc_72470_new_n264_));
OAI21X1 OAI21X1_453 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_16_), .Y(u0_u1__abc_72470_new_n267_));
OAI21X1 OAI21X1_454 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_17_), .Y(u0_u1__abc_72470_new_n270_));
OAI21X1 OAI21X1_455 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_18_), .Y(u0_u1__abc_72470_new_n273_));
OAI21X1 OAI21X1_456 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_19_), .Y(u0_u1__abc_72470_new_n276_));
OAI21X1 OAI21X1_457 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_20_), .Y(u0_u1__abc_72470_new_n279_));
OAI21X1 OAI21X1_458 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_21_), .Y(u0_u1__abc_72470_new_n282_));
OAI21X1 OAI21X1_459 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_22_), .Y(u0_u1__abc_72470_new_n285_));
OAI21X1 OAI21X1_46 ( .A(_abc_81086_new_n301_), .B(lmr_sel), .C(_abc_81086_new_n302_), .Y(tms_s_10_));
OAI21X1 OAI21X1_460 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_23_), .Y(u0_u1__abc_72470_new_n288_));
OAI21X1 OAI21X1_461 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_24_), .Y(u0_u1__abc_72470_new_n291_));
OAI21X1 OAI21X1_462 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_25_), .Y(u0_u1__abc_72470_new_n294_));
OAI21X1 OAI21X1_463 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_26_), .Y(u0_u1__abc_72470_new_n297_));
OAI21X1 OAI21X1_464 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_27_), .Y(u0_u1__abc_72470_new_n300_));
OAI21X1 OAI21X1_465 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_28_), .Y(u0_u1__abc_72470_new_n303_));
OAI21X1 OAI21X1_466 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_29_), .Y(u0_u1__abc_72470_new_n306_));
OAI21X1 OAI21X1_467 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_30_), .Y(u0_u1__abc_72470_new_n309_));
OAI21X1 OAI21X1_468 ( .A(u0_u1__abc_72470_new_n210_), .B(u0_u1__abc_72470_new_n215_), .C(u0_tms1_31_), .Y(u0_u1__abc_72470_new_n312_));
OAI21X1 OAI21X1_469 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_0_), .Y(u0_u1__abc_72470_new_n316_));
OAI21X1 OAI21X1_47 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_11_), .Y(_abc_81086_new_n305_));
OAI21X1 OAI21X1_470 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_1_), .Y(u0_u1__abc_72470_new_n319_));
OAI21X1 OAI21X1_471 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_2_), .Y(u0_u1__abc_72470_new_n322_));
OAI21X1 OAI21X1_472 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_3_), .Y(u0_u1__abc_72470_new_n325_));
OAI21X1 OAI21X1_473 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_4_), .Y(u0_u1__abc_72470_new_n328_));
OAI21X1 OAI21X1_474 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_5_), .Y(u0_u1__abc_72470_new_n331_));
OAI21X1 OAI21X1_475 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_6_), .Y(u0_u1__abc_72470_new_n334_));
OAI21X1 OAI21X1_476 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_7_), .Y(u0_u1__abc_72470_new_n337_));
OAI21X1 OAI21X1_477 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_8_), .Y(u0_u1__abc_72470_new_n340_));
OAI21X1 OAI21X1_478 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_9_), .Y(u0_u1__abc_72470_new_n343_));
OAI21X1 OAI21X1_479 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_10_), .Y(u0_u1__abc_72470_new_n346_));
OAI21X1 OAI21X1_48 ( .A(_abc_81086_new_n304_), .B(lmr_sel), .C(_abc_81086_new_n305_), .Y(tms_s_11_));
OAI21X1 OAI21X1_480 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_11_), .Y(u0_u1__abc_72470_new_n349_));
OAI21X1 OAI21X1_481 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_12_), .Y(u0_u1__abc_72470_new_n352_));
OAI21X1 OAI21X1_482 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_13_), .Y(u0_u1__abc_72470_new_n355_));
OAI21X1 OAI21X1_483 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_14_), .Y(u0_u1__abc_72470_new_n358_));
OAI21X1 OAI21X1_484 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_15_), .Y(u0_u1__abc_72470_new_n361_));
OAI21X1 OAI21X1_485 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_16_), .Y(u0_u1__abc_72470_new_n364_));
OAI21X1 OAI21X1_486 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_17_), .Y(u0_u1__abc_72470_new_n367_));
OAI21X1 OAI21X1_487 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_18_), .Y(u0_u1__abc_72470_new_n370_));
OAI21X1 OAI21X1_488 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_19_), .Y(u0_u1__abc_72470_new_n373_));
OAI21X1 OAI21X1_489 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_20_), .Y(u0_u1__abc_72470_new_n376_));
OAI21X1 OAI21X1_49 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_12_), .Y(_abc_81086_new_n308_));
OAI21X1 OAI21X1_490 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_21_), .Y(u0_u1__abc_72470_new_n379_));
OAI21X1 OAI21X1_491 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_22_), .Y(u0_u1__abc_72470_new_n382_));
OAI21X1 OAI21X1_492 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_23_), .Y(u0_u1__abc_72470_new_n385_));
OAI21X1 OAI21X1_493 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_24_), .Y(u0_u1__abc_72470_new_n388_));
OAI21X1 OAI21X1_494 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_25_), .Y(u0_u1__abc_72470_new_n391_));
OAI21X1 OAI21X1_495 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_26_), .Y(u0_u1__abc_72470_new_n394_));
OAI21X1 OAI21X1_496 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_27_), .Y(u0_u1__abc_72470_new_n397_));
OAI21X1 OAI21X1_497 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_28_), .Y(u0_u1__abc_72470_new_n400_));
OAI21X1 OAI21X1_498 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_29_), .Y(u0_u1__abc_72470_new_n403_));
OAI21X1 OAI21X1_499 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_30_), .Y(u0_u1__abc_72470_new_n406_));
OAI21X1 OAI21X1_5 ( .A(spec_req_cs_1_), .B(_abc_81086_new_n236_), .C(_abc_81086_new_n240_), .Y(_abc_81086_new_n245_));
OAI21X1 OAI21X1_50 ( .A(_abc_81086_new_n307_), .B(lmr_sel), .C(_abc_81086_new_n308_), .Y(tms_s_12_));
OAI21X1 OAI21X1_500 ( .A(u0_u1_addr_r_2_), .B(u0_u1__abc_72470_new_n215_), .C(u0_csc1_31_), .Y(u0_u1__abc_72470_new_n409_));
OAI21X1 OAI21X1_501 ( .A(u0_csc1_21_), .B(\wb_addr_i[26] ), .C(u0_csc_mask_5_), .Y(u0_u1__abc_72470_new_n413_));
OAI21X1 OAI21X1_502 ( .A(u0_csc1_19_), .B(\wb_addr_i[24] ), .C(u0_csc_mask_3_), .Y(u0_u1__abc_72470_new_n415_));
OAI21X1 OAI21X1_503 ( .A(u0_csc1_16_), .B(\wb_addr_i[21] ), .C(u0_csc_mask_0_), .Y(u0_u1__abc_72470_new_n420_));
OAI21X1 OAI21X1_504 ( .A(u0_csc1_18_), .B(\wb_addr_i[23] ), .C(u0_csc_mask_2_), .Y(u0_u1__abc_72470_new_n422_));
OAI21X1 OAI21X1_505 ( .A(u0_csc1_23_), .B(\wb_addr_i[28] ), .C(u0_csc_mask_7_), .Y(u0_u1__abc_72470_new_n426_));
OAI21X1 OAI21X1_506 ( .A(u0_u1__abc_72470_new_n425_), .B(u0_u1__abc_72470_new_n426_), .C(u0_csc1_0_), .Y(u0_u1__abc_72470_new_n427_));
OAI21X1 OAI21X1_507 ( .A(u0_csc1_22_), .B(\wb_addr_i[27] ), .C(u0_csc_mask_6_), .Y(u0_u1__abc_72470_new_n429_));
OAI21X1 OAI21X1_508 ( .A(u0_csc1_20_), .B(\wb_addr_i[25] ), .C(u0_csc_mask_4_), .Y(u0_u1__abc_72470_new_n431_));
OAI21X1 OAI21X1_509 ( .A(u1__abc_72801_new_n259_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n271_), .Y(page_size_8_));
OAI21X1 OAI21X1_51 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_13_), .Y(_abc_81086_new_n311_));
OAI21X1 OAI21X1_510 ( .A(u1__abc_72801_new_n261_), .B(u1__abc_72801_new_n266_), .C(u1__abc_72801_new_n282_), .Y(page_size_9_));
OAI21X1 OAI21X1_511 ( .A(u1__abc_72801_new_n277_), .B(u1__abc_72801_new_n274_), .C(u1__abc_72801_new_n284_), .Y(u1__abc_72801_new_n285_));
OAI21X1 OAI21X1_512 ( .A(u1__abc_72801_new_n289_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[23] ), .Y(u1__abc_72801_new_n296_));
OAI21X1 OAI21X1_513 ( .A(u1__abc_72801_new_n261_), .B(u1__abc_72801_new_n266_), .C(u1__abc_72801_new_n291_), .Y(u1__abc_72801_new_n297_));
OAI21X1 OAI21X1_514 ( .A(u1__abc_72801_new_n300_), .B(u1__abc_72801_new_n301_), .C(u1_bas), .Y(u1__abc_72801_new_n302_));
OAI21X1 OAI21X1_515 ( .A(u1__abc_72801_new_n304_), .B(u1__abc_72801_new_n295_), .C(cs_le), .Y(u1__abc_72801_new_n305_));
OAI21X1 OAI21X1_516 ( .A(u1__abc_72801_new_n308_), .B(u1__abc_72801_new_n274_), .C(u1__abc_72801_new_n309_), .Y(u1__abc_72801_new_n310_));
OAI21X1 OAI21X1_517 ( .A(u1__abc_72801_new_n289_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[24] ), .Y(u1__abc_72801_new_n314_));
OAI21X1 OAI21X1_518 ( .A(u1__abc_72801_new_n259_), .B(u1__abc_72801_new_n316_), .C(u1_bas), .Y(u1__abc_72801_new_n317_));
OAI21X1 OAI21X1_519 ( .A(u1__abc_72801_new_n319_), .B(u1__abc_72801_new_n313_), .C(cs_le), .Y(u1__abc_72801_new_n320_));
OAI21X1 OAI21X1_52 ( .A(_abc_81086_new_n310_), .B(lmr_sel), .C(_abc_81086_new_n311_), .Y(tms_s_13_));
OAI21X1 OAI21X1_520 ( .A(u1__abc_72801_new_n324_), .B(u1__abc_72801_new_n274_), .C(u1__abc_72801_new_n325_), .Y(u1__abc_72801_new_n326_));
OAI21X1 OAI21X1_521 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n285_), .C(cs_le), .Y(u1__abc_72801_new_n329_));
OAI21X1 OAI21X1_522 ( .A(u1__abc_72801_new_n327_), .B(u1__abc_72801_new_n329_), .C(u1__abc_72801_new_n323_), .Y(u1__0row_adr_12_0__0_));
OAI21X1 OAI21X1_523 ( .A(u1__abc_72801_new_n266_), .B(u1__abc_72801_new_n288_), .C(u1__abc_72801_new_n333_), .Y(u1__abc_72801_new_n334_));
OAI21X1 OAI21X1_524 ( .A(u1__abc_72801_new_n324_), .B(u1__abc_72801_new_n268_), .C(u1__abc_72801_new_n341_), .Y(u1__abc_72801_new_n342_));
OAI21X1 OAI21X1_525 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n310_), .C(cs_le), .Y(u1__abc_72801_new_n344_));
OAI21X1 OAI21X1_526 ( .A(u1__abc_72801_new_n343_), .B(u1__abc_72801_new_n344_), .C(u1__abc_72801_new_n331_), .Y(u1__0row_adr_12_0__1_));
OAI21X1 OAI21X1_527 ( .A(u1__abc_72801_new_n267_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[15] ), .Y(u1__abc_72801_new_n353_));
OAI21X1 OAI21X1_528 ( .A(cs_le), .B(u1__abc_72801_new_n346_), .C(u1__abc_72801_new_n357_), .Y(u1__0row_adr_12_0__2_));
OAI21X1 OAI21X1_529 ( .A(u1__abc_72801_new_n267_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[14] ), .Y(u1__abc_72801_new_n361_));
OAI21X1 OAI21X1_53 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_14_), .Y(_abc_81086_new_n314_));
OAI21X1 OAI21X1_530 ( .A(u1__abc_72801_new_n267_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[16] ), .Y(u1__abc_72801_new_n365_));
OAI21X1 OAI21X1_531 ( .A(u1__abc_72801_new_n267_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[17] ), .Y(u1__abc_72801_new_n373_));
OAI21X1 OAI21X1_532 ( .A(u1__abc_72801_new_n267_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[18] ), .Y(u1__abc_72801_new_n383_));
OAI21X1 OAI21X1_533 ( .A(u1__abc_72801_new_n267_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[19] ), .Y(u1__abc_72801_new_n392_));
OAI21X1 OAI21X1_534 ( .A(u1__abc_72801_new_n300_), .B(u1__abc_72801_new_n274_), .C(u1__abc_72801_new_n403_), .Y(u1__abc_72801_new_n404_));
OAI21X1 OAI21X1_535 ( .A(u1_bas), .B(u1__abc_72801_new_n404_), .C(cs_le), .Y(u1__abc_72801_new_n405_));
OAI21X1 OAI21X1_536 ( .A(u1__abc_72801_new_n402_), .B(u1__abc_72801_new_n405_), .C(u1__abc_72801_new_n398_), .Y(u1__0row_adr_12_0__7_));
OAI21X1 OAI21X1_537 ( .A(u1__abc_72801_new_n399_), .B(u1__abc_72801_new_n268_), .C(u1__abc_72801_new_n393_), .Y(u1__abc_72801_new_n410_));
OAI21X1 OAI21X1_538 ( .A(u1_bas), .B(u1__abc_72801_new_n414_), .C(cs_le), .Y(u1__abc_72801_new_n415_));
OAI21X1 OAI21X1_539 ( .A(u1__abc_72801_new_n411_), .B(u1__abc_72801_new_n415_), .C(u1__abc_72801_new_n407_), .Y(u1__0row_adr_12_0__8_));
OAI21X1 OAI21X1_54 ( .A(_abc_81086_new_n313_), .B(lmr_sel), .C(_abc_81086_new_n314_), .Y(tms_s_14_));
OAI21X1 OAI21X1_540 ( .A(u1__abc_72801_new_n300_), .B(u1__abc_72801_new_n301_), .C(u1__abc_72801_new_n328_), .Y(u1__abc_72801_new_n425_));
OAI21X1 OAI21X1_541 ( .A(cs_le), .B(u1__abc_72801_new_n417_), .C(u1__abc_72801_new_n428_), .Y(u1__0row_adr_12_0__9_));
OAI21X1 OAI21X1_542 ( .A(u1__abc_72801_new_n259_), .B(u1__abc_72801_new_n316_), .C(u1__abc_72801_new_n328_), .Y(u1__abc_72801_new_n434_));
OAI21X1 OAI21X1_543 ( .A(u1__abc_72801_new_n438_), .B(u1__abc_72801_new_n433_), .C(cs_le), .Y(u1__abc_72801_new_n439_));
OAI21X1 OAI21X1_544 ( .A(u1__abc_72801_new_n439_), .B(u1__abc_72801_new_n431_), .C(u1__abc_72801_new_n430_), .Y(u1__0row_adr_12_0__10_));
OAI21X1 OAI21X1_545 ( .A(u1__abc_72801_new_n300_), .B(u1__abc_72801_new_n349_), .C(u1__abc_72801_new_n443_), .Y(u1__abc_72801_new_n444_));
OAI21X1 OAI21X1_546 ( .A(u1__abc_72801_new_n267_), .B(u1__abc_72801_new_n264_), .C(\wb_addr_i[24] ), .Y(u1__abc_72801_new_n448_));
OAI21X1 OAI21X1_547 ( .A(u1__abc_72801_new_n289_), .B(u1__abc_72801_new_n299_), .C(\wb_addr_i[23] ), .Y(u1__abc_72801_new_n449_));
OAI21X1 OAI21X1_548 ( .A(u1__abc_72801_new_n450_), .B(u1__abc_72801_new_n447_), .C(cs_le), .Y(u1__abc_72801_new_n451_));
OAI21X1 OAI21X1_549 ( .A(u1__abc_72801_new_n266_), .B(u1__abc_72801_new_n316_), .C(u1__abc_72801_new_n436_), .Y(u1__abc_72801_new_n456_));
OAI21X1 OAI21X1_55 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_15_), .Y(_abc_81086_new_n317_));
OAI21X1 OAI21X1_550 ( .A(u1__abc_72801_new_n328_), .B(u1__abc_72801_new_n456_), .C(u1__abc_72801_new_n455_), .Y(u1__abc_72801_new_n457_));
OAI21X1 OAI21X1_551 ( .A(u1__abc_72801_new_n322_), .B(u1__abc_72801_new_n457_), .C(u1__abc_72801_new_n458_), .Y(u1__0row_adr_12_0__12_));
OAI21X1 OAI21X1_552 ( .A(u1__abc_72801_new_n460_), .B(u1__abc_72801_new_n461_), .C(u1__abc_72801_new_n462_), .Y(u1__0col_adr_9_0__0_));
OAI21X1 OAI21X1_553 ( .A(u1__abc_72801_new_n464_), .B(u1__abc_72801_new_n461_), .C(u1__abc_72801_new_n465_), .Y(u1__0col_adr_9_0__1_));
OAI21X1 OAI21X1_554 ( .A(u1__abc_72801_new_n467_), .B(u1__abc_72801_new_n461_), .C(u1__abc_72801_new_n468_), .Y(u1__0col_adr_9_0__2_));
OAI21X1 OAI21X1_555 ( .A(u1__abc_72801_new_n470_), .B(u1__abc_72801_new_n461_), .C(u1__abc_72801_new_n471_), .Y(u1__0col_adr_9_0__3_));
OAI21X1 OAI21X1_556 ( .A(u1__abc_72801_new_n473_), .B(u1__abc_72801_new_n461_), .C(u1__abc_72801_new_n474_), .Y(u1__0col_adr_9_0__4_));
OAI21X1 OAI21X1_557 ( .A(u1__abc_72801_new_n476_), .B(u1__abc_72801_new_n461_), .C(u1__abc_72801_new_n477_), .Y(u1__0col_adr_9_0__5_));
OAI21X1 OAI21X1_558 ( .A(u1__abc_72801_new_n479_), .B(u1__abc_72801_new_n461_), .C(u1__abc_72801_new_n480_), .Y(u1__0col_adr_9_0__6_));
OAI21X1 OAI21X1_559 ( .A(u1__abc_72801_new_n482_), .B(u1__abc_72801_new_n461_), .C(u1__abc_72801_new_n483_), .Y(u1__0col_adr_9_0__7_));
OAI21X1 OAI21X1_56 ( .A(_abc_81086_new_n316_), .B(lmr_sel), .C(_abc_81086_new_n317_), .Y(tms_s_15_));
OAI21X1 OAI21X1_560 ( .A(u1__abc_72801_new_n461_), .B(u1__abc_72801_new_n485_), .C(u1__abc_72801_new_n486_), .Y(u1__0col_adr_9_0__8_));
OAI21X1 OAI21X1_561 ( .A(u1__abc_72801_new_n461_), .B(u1__abc_72801_new_n488_), .C(u1__abc_72801_new_n489_), .Y(u1__0col_adr_9_0__9_));
OAI21X1 OAI21X1_562 ( .A(u1__abc_72801_new_n460_), .B(u1__abc_72801_new_n288_), .C(u1__abc_72801_new_n494_), .Y(u1__abc_72801_new_n495_));
OAI21X1 OAI21X1_563 ( .A(u1__abc_72801_new_n464_), .B(u1__abc_72801_new_n288_), .C(u1__abc_72801_new_n501_), .Y(u1__abc_72801_new_n502_));
OAI21X1 OAI21X1_564 ( .A(u1__abc_72801_new_n500_), .B(u1__abc_72801_new_n502_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n503_));
OAI21X1 OAI21X1_565 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n499_), .C(u1__abc_72801_new_n503_), .Y(u1__0acs_addr_23_0__1_));
OAI21X1 OAI21X1_566 ( .A(u1__abc_72801_new_n507_), .B(u1__abc_72801_new_n506_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n508_));
OAI21X1 OAI21X1_567 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n505_), .C(u1__abc_72801_new_n508_), .Y(u1__0acs_addr_23_0__2_));
OAI21X1 OAI21X1_568 ( .A(u1__abc_72801_new_n512_), .B(u1__abc_72801_new_n511_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n513_));
OAI21X1 OAI21X1_569 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n510_), .C(u1__abc_72801_new_n513_), .Y(u1__0acs_addr_23_0__3_));
OAI21X1 OAI21X1_57 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_16_), .Y(_abc_81086_new_n320_));
OAI21X1 OAI21X1_570 ( .A(u1__abc_72801_new_n517_), .B(u1__abc_72801_new_n516_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n518_));
OAI21X1 OAI21X1_571 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n515_), .C(u1__abc_72801_new_n518_), .Y(u1__0acs_addr_23_0__4_));
OAI21X1 OAI21X1_572 ( .A(u1__abc_72801_new_n522_), .B(u1__abc_72801_new_n521_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n523_));
OAI21X1 OAI21X1_573 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n520_), .C(u1__abc_72801_new_n523_), .Y(u1__0acs_addr_23_0__5_));
OAI21X1 OAI21X1_574 ( .A(u1__abc_72801_new_n527_), .B(u1__abc_72801_new_n526_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n528_));
OAI21X1 OAI21X1_575 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n525_), .C(u1__abc_72801_new_n528_), .Y(u1__0acs_addr_23_0__6_));
OAI21X1 OAI21X1_576 ( .A(u1__abc_72801_new_n532_), .B(u1__abc_72801_new_n531_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n533_));
OAI21X1 OAI21X1_577 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n530_), .C(u1__abc_72801_new_n533_), .Y(u1__0acs_addr_23_0__7_));
OAI21X1 OAI21X1_578 ( .A(u1__abc_72801_new_n538_), .B(u1__abc_72801_new_n536_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n539_));
OAI21X1 OAI21X1_579 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n535_), .C(u1__abc_72801_new_n539_), .Y(u1__0acs_addr_23_0__8_));
OAI21X1 OAI21X1_58 ( .A(_abc_81086_new_n319_), .B(lmr_sel), .C(_abc_81086_new_n320_), .Y(tms_s_16_));
OAI21X1 OAI21X1_580 ( .A(u1__abc_72801_new_n543_), .B(u1__abc_72801_new_n288_), .C(u1__abc_72801_new_n544_), .Y(u1__abc_72801_new_n545_));
OAI21X1 OAI21X1_581 ( .A(u1__abc_72801_new_n542_), .B(u1__abc_72801_new_n545_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n546_));
OAI21X1 OAI21X1_582 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n541_), .C(u1__abc_72801_new_n546_), .Y(u1__0acs_addr_23_0__9_));
OAI21X1 OAI21X1_583 ( .A(u1__abc_72801_new_n550_), .B(u1__abc_72801_new_n549_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n551_));
OAI21X1 OAI21X1_584 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n548_), .C(u1__abc_72801_new_n551_), .Y(u1__0acs_addr_23_0__10_));
OAI21X1 OAI21X1_585 ( .A(u1__abc_72801_new_n555_), .B(u1__abc_72801_new_n554_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n556_));
OAI21X1 OAI21X1_586 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n553_), .C(u1__abc_72801_new_n556_), .Y(u1__0acs_addr_23_0__11_));
OAI21X1 OAI21X1_587 ( .A(u1__abc_72801_new_n560_), .B(u1__abc_72801_new_n559_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n561_));
OAI21X1 OAI21X1_588 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n558_), .C(u1__abc_72801_new_n561_), .Y(u1__0acs_addr_23_0__12_));
OAI21X1 OAI21X1_589 ( .A(u1__abc_72801_new_n565_), .B(u1__abc_72801_new_n564_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n566_));
OAI21X1 OAI21X1_59 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_17_), .Y(_abc_81086_new_n323_));
OAI21X1 OAI21X1_590 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n563_), .C(u1__abc_72801_new_n566_), .Y(u1__0acs_addr_23_0__13_));
OAI21X1 OAI21X1_591 ( .A(u1__abc_72801_new_n332_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n569_), .Y(u1__abc_72801_new_n570_));
OAI21X1 OAI21X1_592 ( .A(u1__abc_72801_new_n332_), .B(u1__abc_72801_new_n574_), .C(u1__abc_72801_new_n575_), .Y(u1__abc_72801_new_n576_));
OAI21X1 OAI21X1_593 ( .A(cs_le), .B(wb_we_i), .C(u1__abc_72801_new_n576_), .Y(u1__abc_72801_new_n577_));
OAI21X1 OAI21X1_594 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n573_), .C(u1__abc_72801_new_n577_), .Y(u1__0acs_addr_23_0__15_));
OAI21X1 OAI21X1_595 ( .A(u1__abc_72801_new_n580_), .B(u1__abc_72801_new_n574_), .C(u1__abc_72801_new_n581_), .Y(u1__abc_72801_new_n582_));
OAI21X1 OAI21X1_596 ( .A(cs_le), .B(wb_we_i), .C(u1__abc_72801_new_n582_), .Y(u1__abc_72801_new_n583_));
OAI21X1 OAI21X1_597 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n579_), .C(u1__abc_72801_new_n583_), .Y(u1__0acs_addr_23_0__16_));
OAI21X1 OAI21X1_598 ( .A(u1__abc_72801_new_n399_), .B(u1__abc_72801_new_n288_), .C(u1__abc_72801_new_n587_), .Y(u1__abc_72801_new_n588_));
OAI21X1 OAI21X1_599 ( .A(u1__abc_72801_new_n586_), .B(u1__abc_72801_new_n588_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n589_));
OAI21X1 OAI21X1_6 ( .A(_abc_81086_new_n243_), .B(_abc_81086_new_n245_), .C(_abc_81086_new_n244_), .Y(obct_cs_1_));
OAI21X1 OAI21X1_60 ( .A(_abc_81086_new_n322_), .B(lmr_sel), .C(_abc_81086_new_n323_), .Y(tms_s_17_));
OAI21X1 OAI21X1_600 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n585_), .C(u1__abc_72801_new_n589_), .Y(u1__0acs_addr_23_0__17_));
OAI21X1 OAI21X1_601 ( .A(u1__abc_72801_new_n593_), .B(u1__abc_72801_new_n592_), .C(u1__abc_72801_new_n498_), .Y(u1__abc_72801_new_n594_));
OAI21X1 OAI21X1_602 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n591_), .C(u1__abc_72801_new_n594_), .Y(u1__0acs_addr_23_0__18_));
OAI21X1 OAI21X1_603 ( .A(u1__abc_72801_new_n399_), .B(u1__abc_72801_new_n574_), .C(u1__abc_72801_new_n597_), .Y(u1__abc_72801_new_n598_));
OAI21X1 OAI21X1_604 ( .A(cs_le), .B(wb_we_i), .C(u1__abc_72801_new_n598_), .Y(u1__abc_72801_new_n599_));
OAI21X1 OAI21X1_605 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n596_), .C(u1__abc_72801_new_n599_), .Y(u1__0acs_addr_23_0__19_));
OAI21X1 OAI21X1_606 ( .A(u1__abc_72801_new_n300_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n316_), .Y(u1__abc_72801_new_n602_));
OAI21X1 OAI21X1_607 ( .A(u1__abc_72801_new_n300_), .B(u1__abc_72801_new_n574_), .C(u1__abc_72801_new_n606_), .Y(u1__abc_72801_new_n607_));
OAI21X1 OAI21X1_608 ( .A(cs_le), .B(wb_we_i), .C(u1__abc_72801_new_n607_), .Y(u1__abc_72801_new_n608_));
OAI21X1 OAI21X1_609 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n605_), .C(u1__abc_72801_new_n608_), .Y(u1__0acs_addr_23_0__21_));
OAI21X1 OAI21X1_61 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_18_), .Y(_abc_81086_new_n326_));
OAI21X1 OAI21X1_610 ( .A(u1__abc_72801_new_n422_), .B(u1__abc_72801_new_n574_), .C(u1__abc_72801_new_n611_), .Y(u1__abc_72801_new_n612_));
OAI21X1 OAI21X1_611 ( .A(cs_le), .B(wb_we_i), .C(u1__abc_72801_new_n612_), .Y(u1__abc_72801_new_n613_));
OAI21X1 OAI21X1_612 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n610_), .C(u1__abc_72801_new_n613_), .Y(u1__0acs_addr_23_0__22_));
OAI21X1 OAI21X1_613 ( .A(u1__abc_72801_new_n423_), .B(u1__abc_72801_new_n574_), .C(u1__abc_72801_new_n616_), .Y(u1__abc_72801_new_n617_));
OAI21X1 OAI21X1_614 ( .A(cs_le), .B(wb_we_i), .C(u1__abc_72801_new_n617_), .Y(u1__abc_72801_new_n618_));
OAI21X1 OAI21X1_615 ( .A(u1__abc_72801_new_n498_), .B(u1__abc_72801_new_n615_), .C(u1__abc_72801_new_n618_), .Y(u1__0acs_addr_23_0__23_));
OAI21X1 OAI21X1_616 ( .A(wb_stb_i), .B(u1__abc_72801_new_n648_), .C(u1__abc_72801_new_n649_), .Y(u1__0sram_addr_23_0__14_));
OAI21X1 OAI21X1_617 ( .A(wb_stb_i), .B(u1__abc_72801_new_n651_), .C(u1__abc_72801_new_n652_), .Y(u1__0sram_addr_23_0__15_));
OAI21X1 OAI21X1_618 ( .A(wb_stb_i), .B(u1__abc_72801_new_n654_), .C(u1__abc_72801_new_n655_), .Y(u1__0sram_addr_23_0__16_));
OAI21X1 OAI21X1_619 ( .A(u1__abc_72801_new_n460_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n679_), .Y(u1__abc_72801_new_n680_));
OAI21X1 OAI21X1_62 ( .A(_abc_81086_new_n325_), .B(lmr_sel), .C(_abc_81086_new_n326_), .Y(tms_s_18_));
OAI21X1 OAI21X1_620 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n685_), .Y(u1__abc_72801_new_n686_));
OAI21X1 OAI21X1_621 ( .A(tms_s_0_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n686_), .Y(u1__abc_72801_new_n687_));
OAI21X1 OAI21X1_622 ( .A(u1_acs_addr_0_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n688_));
OAI21X1 OAI21X1_623 ( .A(u1__abc_72801_new_n464_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n690_), .Y(u1__abc_72801_new_n691_));
OAI21X1 OAI21X1_624 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n693_), .Y(u1__abc_72801_new_n694_));
OAI21X1 OAI21X1_625 ( .A(tms_s_1_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n694_), .Y(u1__abc_72801_new_n695_));
OAI21X1 OAI21X1_626 ( .A(u1_acs_addr_1_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n696_));
OAI21X1 OAI21X1_627 ( .A(u1__abc_72801_new_n467_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n698_), .Y(u1__abc_72801_new_n699_));
OAI21X1 OAI21X1_628 ( .A(u1_col_adr_2_), .B(row_sel), .C(u1__abc_72801_new_n701_), .Y(u1__abc_72801_new_n702_));
OAI21X1 OAI21X1_629 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n702_), .Y(u1__abc_72801_new_n703_));
OAI21X1 OAI21X1_63 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_19_), .Y(_abc_81086_new_n329_));
OAI21X1 OAI21X1_630 ( .A(tms_s_2_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n703_), .Y(u1__abc_72801_new_n704_));
OAI21X1 OAI21X1_631 ( .A(u1_acs_addr_2_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n705_));
OAI21X1 OAI21X1_632 ( .A(u1__abc_72801_new_n470_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n707_), .Y(u1__abc_72801_new_n708_));
OAI21X1 OAI21X1_633 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n710_), .Y(u1__abc_72801_new_n711_));
OAI21X1 OAI21X1_634 ( .A(tms_s_3_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n711_), .Y(u1__abc_72801_new_n712_));
OAI21X1 OAI21X1_635 ( .A(u1_acs_addr_3_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n713_));
OAI21X1 OAI21X1_636 ( .A(u1__abc_72801_new_n473_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n715_), .Y(u1__abc_72801_new_n716_));
OAI21X1 OAI21X1_637 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n718_), .Y(u1__abc_72801_new_n719_));
OAI21X1 OAI21X1_638 ( .A(tms_s_4_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n719_), .Y(u1__abc_72801_new_n720_));
OAI21X1 OAI21X1_639 ( .A(u1_acs_addr_4_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n721_));
OAI21X1 OAI21X1_64 ( .A(_abc_81086_new_n328_), .B(lmr_sel), .C(_abc_81086_new_n329_), .Y(tms_s_19_));
OAI21X1 OAI21X1_640 ( .A(u1__abc_72801_new_n476_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n723_), .Y(u1__abc_72801_new_n724_));
OAI21X1 OAI21X1_641 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n726_), .Y(u1__abc_72801_new_n727_));
OAI21X1 OAI21X1_642 ( .A(tms_s_5_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n727_), .Y(u1__abc_72801_new_n728_));
OAI21X1 OAI21X1_643 ( .A(u1_acs_addr_5_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n729_));
OAI21X1 OAI21X1_644 ( .A(u1__abc_72801_new_n479_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n731_), .Y(u1__abc_72801_new_n732_));
OAI21X1 OAI21X1_645 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n734_), .Y(u1__abc_72801_new_n735_));
OAI21X1 OAI21X1_646 ( .A(tms_s_6_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n735_), .Y(u1__abc_72801_new_n736_));
OAI21X1 OAI21X1_647 ( .A(u1_acs_addr_6_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n737_));
OAI21X1 OAI21X1_648 ( .A(u1__abc_72801_new_n482_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n739_), .Y(u1__abc_72801_new_n740_));
OAI21X1 OAI21X1_649 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n742_), .Y(u1__abc_72801_new_n743_));
OAI21X1 OAI21X1_65 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_20_), .Y(_abc_81086_new_n332_));
OAI21X1 OAI21X1_650 ( .A(tms_s_7_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n743_), .Y(u1__abc_72801_new_n744_));
OAI21X1 OAI21X1_651 ( .A(u1_acs_addr_7_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n745_));
OAI21X1 OAI21X1_652 ( .A(u1__abc_72801_new_n537_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n747_), .Y(u1__abc_72801_new_n748_));
OAI21X1 OAI21X1_653 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n750_), .Y(u1__abc_72801_new_n751_));
OAI21X1 OAI21X1_654 ( .A(tms_s_8_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n751_), .Y(u1__abc_72801_new_n752_));
OAI21X1 OAI21X1_655 ( .A(u1_acs_addr_8_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n753_));
OAI21X1 OAI21X1_656 ( .A(u1__abc_72801_new_n543_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n755_), .Y(u1__abc_72801_new_n756_));
OAI21X1 OAI21X1_657 ( .A(u1_col_adr_9_), .B(row_sel), .C(u1__abc_72801_new_n758_), .Y(u1__abc_72801_new_n759_));
OAI21X1 OAI21X1_658 ( .A(u1__abc_72801_new_n682_), .B(cas_), .C(u1__abc_72801_new_n759_), .Y(u1__abc_72801_new_n760_));
OAI21X1 OAI21X1_659 ( .A(tms_s_9_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n760_), .Y(u1__abc_72801_new_n761_));
OAI21X1 OAI21X1_66 ( .A(_abc_81086_new_n331_), .B(lmr_sel), .C(_abc_81086_new_n332_), .Y(tms_s_20_));
OAI21X1 OAI21X1_660 ( .A(u1_acs_addr_9_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n762_));
OAI21X1 OAI21X1_661 ( .A(u1__abc_72801_new_n308_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n764_), .Y(u1__abc_72801_new_n765_));
OAI21X1 OAI21X1_662 ( .A(u1__abc_72801_new_n441_), .B(u1__abc_72801_new_n767_), .C(u1__abc_72801_new_n684_), .Y(u1__abc_72801_new_n768_));
OAI21X1 OAI21X1_663 ( .A(tms_s_11_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n768_), .Y(u1__abc_72801_new_n769_));
OAI21X1 OAI21X1_664 ( .A(u1_acs_addr_11_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n770_));
OAI21X1 OAI21X1_665 ( .A(u1__abc_72801_new_n324_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n772_), .Y(u1__abc_72801_new_n773_));
OAI21X1 OAI21X1_666 ( .A(u1__abc_72801_new_n775_), .B(u1__abc_72801_new_n767_), .C(u1__abc_72801_new_n684_), .Y(u1__abc_72801_new_n776_));
OAI21X1 OAI21X1_667 ( .A(tms_s_12_), .B(u1__abc_72801_new_n684_), .C(u1__abc_72801_new_n776_), .Y(u1__abc_72801_new_n777_));
OAI21X1 OAI21X1_668 ( .A(u1_acs_addr_12_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n778_));
OAI21X1 OAI21X1_669 ( .A(u1__abc_72801_new_n332_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n780_), .Y(u1__abc_72801_new_n781_));
OAI21X1 OAI21X1_67 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_21_), .Y(_abc_81086_new_n335_));
OAI21X1 OAI21X1_670 ( .A(u1_acs_addr_13_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n783_));
OAI21X1 OAI21X1_671 ( .A(u1__abc_72801_new_n580_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n785_), .Y(u1__abc_72801_new_n786_));
OAI21X1 OAI21X1_672 ( .A(u1_acs_addr_14_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n788_));
OAI21X1 OAI21X1_673 ( .A(\wb_addr_i[17] ), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n790_), .Y(u1__abc_72801_new_n791_));
OAI21X1 OAI21X1_674 ( .A(u1_acs_addr_15_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n792_));
OAI21X1 OAI21X1_675 ( .A(\wb_addr_i[18] ), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n794_), .Y(u1__abc_72801_new_n795_));
OAI21X1 OAI21X1_676 ( .A(u1_acs_addr_16_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n796_));
OAI21X1 OAI21X1_677 ( .A(u1_acs_addr_17_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n799_));
OAI21X1 OAI21X1_678 ( .A(u1_acs_addr_18_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n802_));
OAI21X1 OAI21X1_679 ( .A(u1_acs_addr_19_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n805_));
OAI21X1 OAI21X1_68 ( .A(_abc_81086_new_n334_), .B(lmr_sel), .C(_abc_81086_new_n335_), .Y(tms_s_21_));
OAI21X1 OAI21X1_680 ( .A(u1_acs_addr_20_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n808_));
OAI21X1 OAI21X1_681 ( .A(u1_acs_addr_21_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n811_));
OAI21X1 OAI21X1_682 ( .A(u1_acs_addr_22_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n814_));
OAI21X1 OAI21X1_683 ( .A(u1_acs_addr_23_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n817_));
OAI21X1 OAI21X1_684 ( .A(u1__abc_72801_new_n277_), .B(u1__abc_72801_new_n678_), .C(u1__abc_72801_new_n819_), .Y(u1__abc_72801_new_n820_));
OAI21X1 OAI21X1_685 ( .A(u1_acs_addr_10_), .B(u1__abc_72801_new_n675_), .C(u1__abc_72801_new_n673_), .Y(u1__abc_72801_new_n822_));
OAI21X1 OAI21X1_686 ( .A(u1__abc_72801_new_n683_), .B(u1__abc_72801_new_n823_), .C(u1__abc_72801_new_n824_), .Y(u1__abc_72801_new_n825_));
OAI21X1 OAI21X1_687 ( .A(u1__abc_72801_new_n822_), .B(u1__abc_72801_new_n821_), .C(u1__abc_72801_new_n826_), .Y(mc_addr_d_10_));
OAI21X1 OAI21X1_688 ( .A(u1_u0__abc_72719_new_n65_), .B(u1_u0__abc_72719_new_n61_), .C(u1_u0__abc_72719_new_n66_), .Y(u1_u0__abc_72719_new_n67_));
OAI21X1 OAI21X1_689 ( .A(u1_u0__abc_72719_new_n74_), .B(u1_u0__abc_72719_new_n71_), .C(u1_u0__abc_72719_new_n75_), .Y(u1_u0__abc_72719_new_n76_));
OAI21X1 OAI21X1_69 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_22_), .Y(_abc_81086_new_n338_));
OAI21X1 OAI21X1_690 ( .A(u1_u0__abc_72719_new_n81_), .B(u1_u0__abc_72719_new_n78_), .C(u1_u0__abc_72719_new_n82_), .Y(u1_u0__abc_72719_new_n86_));
OAI21X1 OAI21X1_691 ( .A(u1_u0__abc_72719_new_n93_), .B(u1_u0__abc_72719_new_n91_), .C(u1_u0__abc_72719_new_n94_), .Y(u1_u0__abc_72719_new_n95_));
OAI21X1 OAI21X1_692 ( .A(u1_u0__abc_72719_new_n115_), .B(u1_u0__abc_72719_new_n97_), .C(u1_u0__abc_72719_new_n112_), .Y(u1_u0__abc_72719_new_n116_));
OAI21X1 OAI21X1_693 ( .A(u1_u0__abc_72719_new_n123_), .B(u1_u0__abc_72719_new_n121_), .C(u1_acs_addr_23_), .Y(u1_u0__abc_72719_new_n124_));
OAI21X1 OAI21X1_694 ( .A(u2__abc_74202_new_n65_), .B(u2__abc_74202_new_n90_), .C(u2__abc_74202_new_n91_), .Y(u2_bank_clr_all_0));
OAI21X1 OAI21X1_695 ( .A(u2__abc_74202_new_n67_), .B(u2__abc_74202_new_n90_), .C(u2__abc_74202_new_n91_), .Y(u2_bank_clr_all_1));
OAI21X1 OAI21X1_696 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_0_), .Y(u2_u0__abc_73914_new_n141_));
OAI21X1 OAI21X1_697 ( .A(u2_u0__abc_73914_new_n136_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n141_), .Y(u2_u0__0b3_last_row_12_0__0_));
OAI21X1 OAI21X1_698 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_1_), .Y(u2_u0__abc_73914_new_n144_));
OAI21X1 OAI21X1_699 ( .A(u2_u0__abc_73914_new_n143_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n144_), .Y(u2_u0__0b3_last_row_12_0__1_));
OAI21X1 OAI21X1_7 ( .A(susp_sel), .B(rfr_ack), .C(cs_need_rfr_2_), .Y(_abc_81086_new_n248_));
OAI21X1 OAI21X1_70 ( .A(_abc_81086_new_n337_), .B(lmr_sel), .C(_abc_81086_new_n338_), .Y(tms_s_22_));
OAI21X1 OAI21X1_700 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_2_), .Y(u2_u0__abc_73914_new_n147_));
OAI21X1 OAI21X1_701 ( .A(u2_u0__abc_73914_new_n146_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n147_), .Y(u2_u0__0b3_last_row_12_0__2_));
OAI21X1 OAI21X1_702 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_3_), .Y(u2_u0__abc_73914_new_n150_));
OAI21X1 OAI21X1_703 ( .A(u2_u0__abc_73914_new_n149_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n150_), .Y(u2_u0__0b3_last_row_12_0__3_));
OAI21X1 OAI21X1_704 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_4_), .Y(u2_u0__abc_73914_new_n153_));
OAI21X1 OAI21X1_705 ( .A(u2_u0__abc_73914_new_n152_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n153_), .Y(u2_u0__0b3_last_row_12_0__4_));
OAI21X1 OAI21X1_706 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_5_), .Y(u2_u0__abc_73914_new_n156_));
OAI21X1 OAI21X1_707 ( .A(u2_u0__abc_73914_new_n155_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n156_), .Y(u2_u0__0b3_last_row_12_0__5_));
OAI21X1 OAI21X1_708 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_6_), .Y(u2_u0__abc_73914_new_n159_));
OAI21X1 OAI21X1_709 ( .A(u2_u0__abc_73914_new_n158_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n159_), .Y(u2_u0__0b3_last_row_12_0__6_));
OAI21X1 OAI21X1_71 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_23_), .Y(_abc_81086_new_n341_));
OAI21X1 OAI21X1_710 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_7_), .Y(u2_u0__abc_73914_new_n162_));
OAI21X1 OAI21X1_711 ( .A(u2_u0__abc_73914_new_n161_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n162_), .Y(u2_u0__0b3_last_row_12_0__7_));
OAI21X1 OAI21X1_712 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_8_), .Y(u2_u0__abc_73914_new_n165_));
OAI21X1 OAI21X1_713 ( .A(u2_u0__abc_73914_new_n164_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n165_), .Y(u2_u0__0b3_last_row_12_0__8_));
OAI21X1 OAI21X1_714 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_9_), .Y(u2_u0__abc_73914_new_n168_));
OAI21X1 OAI21X1_715 ( .A(u2_u0__abc_73914_new_n167_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n168_), .Y(u2_u0__0b3_last_row_12_0__9_));
OAI21X1 OAI21X1_716 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_10_), .Y(u2_u0__abc_73914_new_n171_));
OAI21X1 OAI21X1_717 ( .A(u2_u0__abc_73914_new_n170_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n171_), .Y(u2_u0__0b3_last_row_12_0__10_));
OAI21X1 OAI21X1_718 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_11_), .Y(u2_u0__abc_73914_new_n174_));
OAI21X1 OAI21X1_719 ( .A(u2_u0__abc_73914_new_n173_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n174_), .Y(u2_u0__0b3_last_row_12_0__11_));
OAI21X1 OAI21X1_72 ( .A(_abc_81086_new_n340_), .B(lmr_sel), .C(_abc_81086_new_n341_), .Y(tms_s_23_));
OAI21X1 OAI21X1_720 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0_b3_last_row_12_), .Y(u2_u0__abc_73914_new_n177_));
OAI21X1 OAI21X1_721 ( .A(u2_u0__abc_73914_new_n176_), .B(u2_u0__abc_73914_new_n139_), .C(u2_u0__abc_73914_new_n177_), .Y(u2_u0__0b3_last_row_12_0__12_));
OAI21X1 OAI21X1_722 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_73914_new_n182_));
OAI21X1 OAI21X1_723 ( .A(u2_u0__abc_73914_new_n136_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n182_), .Y(u2_u0__0b0_last_row_12_0__0_));
OAI21X1 OAI21X1_724 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_73914_new_n184_));
OAI21X1 OAI21X1_725 ( .A(u2_u0__abc_73914_new_n143_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n184_), .Y(u2_u0__0b0_last_row_12_0__1_));
OAI21X1 OAI21X1_726 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_2_), .Y(u2_u0__abc_73914_new_n186_));
OAI21X1 OAI21X1_727 ( .A(u2_u0__abc_73914_new_n146_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n186_), .Y(u2_u0__0b0_last_row_12_0__2_));
OAI21X1 OAI21X1_728 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_3_), .Y(u2_u0__abc_73914_new_n188_));
OAI21X1 OAI21X1_729 ( .A(u2_u0__abc_73914_new_n149_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n188_), .Y(u2_u0__0b0_last_row_12_0__3_));
OAI21X1 OAI21X1_73 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_24_), .Y(_abc_81086_new_n344_));
OAI21X1 OAI21X1_730 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_4_), .Y(u2_u0__abc_73914_new_n190_));
OAI21X1 OAI21X1_731 ( .A(u2_u0__abc_73914_new_n152_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n190_), .Y(u2_u0__0b0_last_row_12_0__4_));
OAI21X1 OAI21X1_732 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_5_), .Y(u2_u0__abc_73914_new_n192_));
OAI21X1 OAI21X1_733 ( .A(u2_u0__abc_73914_new_n155_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n192_), .Y(u2_u0__0b0_last_row_12_0__5_));
OAI21X1 OAI21X1_734 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_6_), .Y(u2_u0__abc_73914_new_n194_));
OAI21X1 OAI21X1_735 ( .A(u2_u0__abc_73914_new_n158_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n194_), .Y(u2_u0__0b0_last_row_12_0__6_));
OAI21X1 OAI21X1_736 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_73914_new_n196_));
OAI21X1 OAI21X1_737 ( .A(u2_u0__abc_73914_new_n161_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n196_), .Y(u2_u0__0b0_last_row_12_0__7_));
OAI21X1 OAI21X1_738 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_8_), .Y(u2_u0__abc_73914_new_n198_));
OAI21X1 OAI21X1_739 ( .A(u2_u0__abc_73914_new_n164_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n198_), .Y(u2_u0__0b0_last_row_12_0__8_));
OAI21X1 OAI21X1_74 ( .A(_abc_81086_new_n343_), .B(lmr_sel), .C(_abc_81086_new_n344_), .Y(tms_s_24_));
OAI21X1 OAI21X1_740 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_9_), .Y(u2_u0__abc_73914_new_n200_));
OAI21X1 OAI21X1_741 ( .A(u2_u0__abc_73914_new_n167_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n200_), .Y(u2_u0__0b0_last_row_12_0__9_));
OAI21X1 OAI21X1_742 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_73914_new_n202_));
OAI21X1 OAI21X1_743 ( .A(u2_u0__abc_73914_new_n170_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n202_), .Y(u2_u0__0b0_last_row_12_0__10_));
OAI21X1 OAI21X1_744 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_73914_new_n204_));
OAI21X1 OAI21X1_745 ( .A(u2_u0__abc_73914_new_n173_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n204_), .Y(u2_u0__0b0_last_row_12_0__11_));
OAI21X1 OAI21X1_746 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0_b0_last_row_12_), .Y(u2_u0__abc_73914_new_n206_));
OAI21X1 OAI21X1_747 ( .A(u2_u0__abc_73914_new_n176_), .B(u2_u0__abc_73914_new_n181_), .C(u2_u0__abc_73914_new_n206_), .Y(u2_u0__0b0_last_row_12_0__12_));
OAI21X1 OAI21X1_748 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_0_), .Y(u2_u0__abc_73914_new_n211_));
OAI21X1 OAI21X1_749 ( .A(u2_u0__abc_73914_new_n136_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n211_), .Y(u2_u0__0b1_last_row_12_0__0_));
OAI21X1 OAI21X1_75 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_25_), .Y(_abc_81086_new_n347_));
OAI21X1 OAI21X1_750 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_1_), .Y(u2_u0__abc_73914_new_n213_));
OAI21X1 OAI21X1_751 ( .A(u2_u0__abc_73914_new_n143_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n213_), .Y(u2_u0__0b1_last_row_12_0__1_));
OAI21X1 OAI21X1_752 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_2_), .Y(u2_u0__abc_73914_new_n215_));
OAI21X1 OAI21X1_753 ( .A(u2_u0__abc_73914_new_n146_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n215_), .Y(u2_u0__0b1_last_row_12_0__2_));
OAI21X1 OAI21X1_754 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_3_), .Y(u2_u0__abc_73914_new_n217_));
OAI21X1 OAI21X1_755 ( .A(u2_u0__abc_73914_new_n149_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n217_), .Y(u2_u0__0b1_last_row_12_0__3_));
OAI21X1 OAI21X1_756 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_73914_new_n219_));
OAI21X1 OAI21X1_757 ( .A(u2_u0__abc_73914_new_n152_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n219_), .Y(u2_u0__0b1_last_row_12_0__4_));
OAI21X1 OAI21X1_758 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_5_), .Y(u2_u0__abc_73914_new_n221_));
OAI21X1 OAI21X1_759 ( .A(u2_u0__abc_73914_new_n155_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n221_), .Y(u2_u0__0b1_last_row_12_0__5_));
OAI21X1 OAI21X1_76 ( .A(_abc_81086_new_n346_), .B(lmr_sel), .C(_abc_81086_new_n347_), .Y(tms_s_25_));
OAI21X1 OAI21X1_760 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_73914_new_n223_));
OAI21X1 OAI21X1_761 ( .A(u2_u0__abc_73914_new_n158_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n223_), .Y(u2_u0__0b1_last_row_12_0__6_));
OAI21X1 OAI21X1_762 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_7_), .Y(u2_u0__abc_73914_new_n225_));
OAI21X1 OAI21X1_763 ( .A(u2_u0__abc_73914_new_n161_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n225_), .Y(u2_u0__0b1_last_row_12_0__7_));
OAI21X1 OAI21X1_764 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_73914_new_n227_));
OAI21X1 OAI21X1_765 ( .A(u2_u0__abc_73914_new_n164_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n227_), .Y(u2_u0__0b1_last_row_12_0__8_));
OAI21X1 OAI21X1_766 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_9_), .Y(u2_u0__abc_73914_new_n229_));
OAI21X1 OAI21X1_767 ( .A(u2_u0__abc_73914_new_n167_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n229_), .Y(u2_u0__0b1_last_row_12_0__9_));
OAI21X1 OAI21X1_768 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_10_), .Y(u2_u0__abc_73914_new_n231_));
OAI21X1 OAI21X1_769 ( .A(u2_u0__abc_73914_new_n170_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n231_), .Y(u2_u0__0b1_last_row_12_0__10_));
OAI21X1 OAI21X1_77 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_26_), .Y(_abc_81086_new_n350_));
OAI21X1 OAI21X1_770 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_11_), .Y(u2_u0__abc_73914_new_n233_));
OAI21X1 OAI21X1_771 ( .A(u2_u0__abc_73914_new_n173_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n233_), .Y(u2_u0__0b1_last_row_12_0__11_));
OAI21X1 OAI21X1_772 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0_b1_last_row_12_), .Y(u2_u0__abc_73914_new_n235_));
OAI21X1 OAI21X1_773 ( .A(u2_u0__abc_73914_new_n176_), .B(u2_u0__abc_73914_new_n210_), .C(u2_u0__abc_73914_new_n235_), .Y(u2_u0__0b1_last_row_12_0__12_));
OAI21X1 OAI21X1_774 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_0_), .Y(u2_u0__abc_73914_new_n240_));
OAI21X1 OAI21X1_775 ( .A(u2_u0__abc_73914_new_n136_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n240_), .Y(u2_u0__0b2_last_row_12_0__0_));
OAI21X1 OAI21X1_776 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_1_), .Y(u2_u0__abc_73914_new_n242_));
OAI21X1 OAI21X1_777 ( .A(u2_u0__abc_73914_new_n143_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n242_), .Y(u2_u0__0b2_last_row_12_0__1_));
OAI21X1 OAI21X1_778 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_73914_new_n244_));
OAI21X1 OAI21X1_779 ( .A(u2_u0__abc_73914_new_n146_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n244_), .Y(u2_u0__0b2_last_row_12_0__2_));
OAI21X1 OAI21X1_78 ( .A(_abc_81086_new_n349_), .B(lmr_sel), .C(_abc_81086_new_n350_), .Y(tms_s_26_));
OAI21X1 OAI21X1_780 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_73914_new_n246_));
OAI21X1 OAI21X1_781 ( .A(u2_u0__abc_73914_new_n149_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n246_), .Y(u2_u0__0b2_last_row_12_0__3_));
OAI21X1 OAI21X1_782 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_4_), .Y(u2_u0__abc_73914_new_n248_));
OAI21X1 OAI21X1_783 ( .A(u2_u0__abc_73914_new_n152_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n248_), .Y(u2_u0__0b2_last_row_12_0__4_));
OAI21X1 OAI21X1_784 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_73914_new_n250_));
OAI21X1 OAI21X1_785 ( .A(u2_u0__abc_73914_new_n155_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n250_), .Y(u2_u0__0b2_last_row_12_0__5_));
OAI21X1 OAI21X1_786 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_6_), .Y(u2_u0__abc_73914_new_n252_));
OAI21X1 OAI21X1_787 ( .A(u2_u0__abc_73914_new_n158_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n252_), .Y(u2_u0__0b2_last_row_12_0__6_));
OAI21X1 OAI21X1_788 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_73914_new_n254_));
OAI21X1 OAI21X1_789 ( .A(u2_u0__abc_73914_new_n161_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n254_), .Y(u2_u0__0b2_last_row_12_0__7_));
OAI21X1 OAI21X1_79 ( .A(init_ack), .B(lmr_ack), .C(sp_tms_27_), .Y(_abc_81086_new_n353_));
OAI21X1 OAI21X1_790 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_8_), .Y(u2_u0__abc_73914_new_n256_));
OAI21X1 OAI21X1_791 ( .A(u2_u0__abc_73914_new_n164_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n256_), .Y(u2_u0__0b2_last_row_12_0__8_));
OAI21X1 OAI21X1_792 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_9_), .Y(u2_u0__abc_73914_new_n258_));
OAI21X1 OAI21X1_793 ( .A(u2_u0__abc_73914_new_n167_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n258_), .Y(u2_u0__0b2_last_row_12_0__9_));
OAI21X1 OAI21X1_794 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_73914_new_n260_));
OAI21X1 OAI21X1_795 ( .A(u2_u0__abc_73914_new_n170_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n260_), .Y(u2_u0__0b2_last_row_12_0__10_));
OAI21X1 OAI21X1_796 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_11_), .Y(u2_u0__abc_73914_new_n262_));
OAI21X1 OAI21X1_797 ( .A(u2_u0__abc_73914_new_n173_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n262_), .Y(u2_u0__0b2_last_row_12_0__11_));
OAI21X1 OAI21X1_798 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0_b2_last_row_12_), .Y(u2_u0__abc_73914_new_n264_));
OAI21X1 OAI21X1_799 ( .A(u2_u0__abc_73914_new_n176_), .B(u2_u0__abc_73914_new_n238_), .C(u2_u0__abc_73914_new_n264_), .Y(u2_u0__0b2_last_row_12_0__12_));
OAI21X1 OAI21X1_8 ( .A(spec_req_cs_2_), .B(_abc_81086_new_n236_), .C(_abc_81086_new_n240_), .Y(_abc_81086_new_n249_));
OAI21X1 OAI21X1_80 ( .A(_abc_81086_new_n352_), .B(lmr_sel), .C(_abc_81086_new_n353_), .Y(tms_s_27_));
OAI21X1 OAI21X1_800 ( .A(u2_u0__abc_73914_new_n285_), .B(u2_u0__abc_73914_new_n286_), .C(u2_u0__abc_73914_new_n284_), .Y(u2_u0__abc_73914_new_n287_));
OAI21X1 OAI21X1_801 ( .A(u2_u0__abc_73914_new_n289_), .B(u2_u0__abc_73914_new_n288_), .C(u2_u0__abc_73914_new_n291_), .Y(u2_u0__abc_73914_new_n292_));
OAI21X1 OAI21X1_802 ( .A(u2_u0__abc_73914_new_n385_), .B(u2_u0__abc_73914_new_n386_), .C(u2_u0__abc_73914_new_n384_), .Y(u2_u0__abc_73914_new_n387_));
OAI21X1 OAI21X1_803 ( .A(u2_u0__abc_73914_new_n390_), .B(u2_u0__abc_73914_new_n389_), .C(u2_u0__abc_73914_new_n388_), .Y(u2_u0__abc_73914_new_n391_));
OAI21X1 OAI21X1_804 ( .A(u2_u0__abc_73914_new_n399_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0__abc_73914_new_n400_), .Y(u2_u0__abc_73914_new_n401_));
OAI21X1 OAI21X1_805 ( .A(u2_u0__abc_73914_new_n398_), .B(u2_u0__abc_73914_new_n179_), .C(u2_u0__abc_73914_new_n402_), .Y(u2_bank_open_0));
OAI21X1 OAI21X1_806 ( .A(u2_u0__abc_73914_new_n404_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0__abc_73914_new_n406_), .Y(u2_u0__abc_73914_new_n407_));
OAI21X1 OAI21X1_807 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n239_), .C(u2_u0__abc_73914_new_n407_), .Y(u2_u0__0bank2_open_0_0_));
OAI21X1 OAI21X1_808 ( .A(u2_u0__abc_73914_new_n404_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0__abc_73914_new_n410_), .Y(u2_u0__abc_73914_new_n411_));
OAI21X1 OAI21X1_809 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n137_), .C(u2_u0__abc_73914_new_n411_), .Y(u2_u0__0bank3_open_0_0_));
OAI21X1 OAI21X1_81 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_1_), .Y(_abc_81086_new_n371_));
OAI21X1 OAI21X1_810 ( .A(u2_u0__abc_73914_new_n404_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0__abc_73914_new_n415_), .Y(u2_u0__abc_73914_new_n416_));
OAI21X1 OAI21X1_811 ( .A(u2_u0__abc_73914_new_n140_), .B(u2_u0__abc_73914_new_n209_), .C(u2_u0__abc_73914_new_n416_), .Y(u2_u0__0bank1_open_0_0_));
OAI21X1 OAI21X1_812 ( .A(u2_u0__abc_73914_new_n419_), .B(u2_u0__abc_73914_new_n418_), .C(u2_u0__abc_73914_new_n181_), .Y(u2_u0__0bank0_open_0_0_));
OAI21X1 OAI21X1_813 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_0_), .Y(u2_u1__abc_73914_new_n141_));
OAI21X1 OAI21X1_814 ( .A(u2_u1__abc_73914_new_n136_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n141_), .Y(u2_u1__0b3_last_row_12_0__0_));
OAI21X1 OAI21X1_815 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_1_), .Y(u2_u1__abc_73914_new_n144_));
OAI21X1 OAI21X1_816 ( .A(u2_u1__abc_73914_new_n143_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n144_), .Y(u2_u1__0b3_last_row_12_0__1_));
OAI21X1 OAI21X1_817 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_2_), .Y(u2_u1__abc_73914_new_n147_));
OAI21X1 OAI21X1_818 ( .A(u2_u1__abc_73914_new_n146_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n147_), .Y(u2_u1__0b3_last_row_12_0__2_));
OAI21X1 OAI21X1_819 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_3_), .Y(u2_u1__abc_73914_new_n150_));
OAI21X1 OAI21X1_82 ( .A(_abc_81086_new_n370_), .B(lmr_sel), .C(_abc_81086_new_n371_), .Y(csc_s_1_));
OAI21X1 OAI21X1_820 ( .A(u2_u1__abc_73914_new_n149_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n150_), .Y(u2_u1__0b3_last_row_12_0__3_));
OAI21X1 OAI21X1_821 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_4_), .Y(u2_u1__abc_73914_new_n153_));
OAI21X1 OAI21X1_822 ( .A(u2_u1__abc_73914_new_n152_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n153_), .Y(u2_u1__0b3_last_row_12_0__4_));
OAI21X1 OAI21X1_823 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_5_), .Y(u2_u1__abc_73914_new_n156_));
OAI21X1 OAI21X1_824 ( .A(u2_u1__abc_73914_new_n155_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n156_), .Y(u2_u1__0b3_last_row_12_0__5_));
OAI21X1 OAI21X1_825 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_6_), .Y(u2_u1__abc_73914_new_n159_));
OAI21X1 OAI21X1_826 ( .A(u2_u1__abc_73914_new_n158_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n159_), .Y(u2_u1__0b3_last_row_12_0__6_));
OAI21X1 OAI21X1_827 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_7_), .Y(u2_u1__abc_73914_new_n162_));
OAI21X1 OAI21X1_828 ( .A(u2_u1__abc_73914_new_n161_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n162_), .Y(u2_u1__0b3_last_row_12_0__7_));
OAI21X1 OAI21X1_829 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_8_), .Y(u2_u1__abc_73914_new_n165_));
OAI21X1 OAI21X1_83 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_2_), .Y(_abc_81086_new_n374_));
OAI21X1 OAI21X1_830 ( .A(u2_u1__abc_73914_new_n164_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n165_), .Y(u2_u1__0b3_last_row_12_0__8_));
OAI21X1 OAI21X1_831 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_9_), .Y(u2_u1__abc_73914_new_n168_));
OAI21X1 OAI21X1_832 ( .A(u2_u1__abc_73914_new_n167_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n168_), .Y(u2_u1__0b3_last_row_12_0__9_));
OAI21X1 OAI21X1_833 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_10_), .Y(u2_u1__abc_73914_new_n171_));
OAI21X1 OAI21X1_834 ( .A(u2_u1__abc_73914_new_n170_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n171_), .Y(u2_u1__0b3_last_row_12_0__10_));
OAI21X1 OAI21X1_835 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_11_), .Y(u2_u1__abc_73914_new_n174_));
OAI21X1 OAI21X1_836 ( .A(u2_u1__abc_73914_new_n173_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n174_), .Y(u2_u1__0b3_last_row_12_0__11_));
OAI21X1 OAI21X1_837 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1_b3_last_row_12_), .Y(u2_u1__abc_73914_new_n177_));
OAI21X1 OAI21X1_838 ( .A(u2_u1__abc_73914_new_n176_), .B(u2_u1__abc_73914_new_n139_), .C(u2_u1__abc_73914_new_n177_), .Y(u2_u1__0b3_last_row_12_0__12_));
OAI21X1 OAI21X1_839 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_73914_new_n182_));
OAI21X1 OAI21X1_84 ( .A(_abc_81086_new_n373_), .B(lmr_sel), .C(_abc_81086_new_n374_), .Y(csc_s_2_));
OAI21X1 OAI21X1_840 ( .A(u2_u1__abc_73914_new_n136_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n182_), .Y(u2_u1__0b0_last_row_12_0__0_));
OAI21X1 OAI21X1_841 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_73914_new_n184_));
OAI21X1 OAI21X1_842 ( .A(u2_u1__abc_73914_new_n143_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n184_), .Y(u2_u1__0b0_last_row_12_0__1_));
OAI21X1 OAI21X1_843 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_2_), .Y(u2_u1__abc_73914_new_n186_));
OAI21X1 OAI21X1_844 ( .A(u2_u1__abc_73914_new_n146_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n186_), .Y(u2_u1__0b0_last_row_12_0__2_));
OAI21X1 OAI21X1_845 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_3_), .Y(u2_u1__abc_73914_new_n188_));
OAI21X1 OAI21X1_846 ( .A(u2_u1__abc_73914_new_n149_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n188_), .Y(u2_u1__0b0_last_row_12_0__3_));
OAI21X1 OAI21X1_847 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_4_), .Y(u2_u1__abc_73914_new_n190_));
OAI21X1 OAI21X1_848 ( .A(u2_u1__abc_73914_new_n152_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n190_), .Y(u2_u1__0b0_last_row_12_0__4_));
OAI21X1 OAI21X1_849 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_5_), .Y(u2_u1__abc_73914_new_n192_));
OAI21X1 OAI21X1_85 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_3_), .Y(_abc_81086_new_n377_));
OAI21X1 OAI21X1_850 ( .A(u2_u1__abc_73914_new_n155_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n192_), .Y(u2_u1__0b0_last_row_12_0__5_));
OAI21X1 OAI21X1_851 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_6_), .Y(u2_u1__abc_73914_new_n194_));
OAI21X1 OAI21X1_852 ( .A(u2_u1__abc_73914_new_n158_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n194_), .Y(u2_u1__0b0_last_row_12_0__6_));
OAI21X1 OAI21X1_853 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_73914_new_n196_));
OAI21X1 OAI21X1_854 ( .A(u2_u1__abc_73914_new_n161_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n196_), .Y(u2_u1__0b0_last_row_12_0__7_));
OAI21X1 OAI21X1_855 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_8_), .Y(u2_u1__abc_73914_new_n198_));
OAI21X1 OAI21X1_856 ( .A(u2_u1__abc_73914_new_n164_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n198_), .Y(u2_u1__0b0_last_row_12_0__8_));
OAI21X1 OAI21X1_857 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_9_), .Y(u2_u1__abc_73914_new_n200_));
OAI21X1 OAI21X1_858 ( .A(u2_u1__abc_73914_new_n167_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n200_), .Y(u2_u1__0b0_last_row_12_0__9_));
OAI21X1 OAI21X1_859 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_73914_new_n202_));
OAI21X1 OAI21X1_86 ( .A(_abc_81086_new_n376_), .B(lmr_sel), .C(_abc_81086_new_n377_), .Y(csc_s_3_));
OAI21X1 OAI21X1_860 ( .A(u2_u1__abc_73914_new_n170_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n202_), .Y(u2_u1__0b0_last_row_12_0__10_));
OAI21X1 OAI21X1_861 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_73914_new_n204_));
OAI21X1 OAI21X1_862 ( .A(u2_u1__abc_73914_new_n173_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n204_), .Y(u2_u1__0b0_last_row_12_0__11_));
OAI21X1 OAI21X1_863 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1_b0_last_row_12_), .Y(u2_u1__abc_73914_new_n206_));
OAI21X1 OAI21X1_864 ( .A(u2_u1__abc_73914_new_n176_), .B(u2_u1__abc_73914_new_n181_), .C(u2_u1__abc_73914_new_n206_), .Y(u2_u1__0b0_last_row_12_0__12_));
OAI21X1 OAI21X1_865 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_0_), .Y(u2_u1__abc_73914_new_n211_));
OAI21X1 OAI21X1_866 ( .A(u2_u1__abc_73914_new_n136_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n211_), .Y(u2_u1__0b1_last_row_12_0__0_));
OAI21X1 OAI21X1_867 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_1_), .Y(u2_u1__abc_73914_new_n213_));
OAI21X1 OAI21X1_868 ( .A(u2_u1__abc_73914_new_n143_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n213_), .Y(u2_u1__0b1_last_row_12_0__1_));
OAI21X1 OAI21X1_869 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_2_), .Y(u2_u1__abc_73914_new_n215_));
OAI21X1 OAI21X1_87 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_4_), .Y(_abc_81086_new_n380_));
OAI21X1 OAI21X1_870 ( .A(u2_u1__abc_73914_new_n146_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n215_), .Y(u2_u1__0b1_last_row_12_0__2_));
OAI21X1 OAI21X1_871 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_3_), .Y(u2_u1__abc_73914_new_n217_));
OAI21X1 OAI21X1_872 ( .A(u2_u1__abc_73914_new_n149_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n217_), .Y(u2_u1__0b1_last_row_12_0__3_));
OAI21X1 OAI21X1_873 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_73914_new_n219_));
OAI21X1 OAI21X1_874 ( .A(u2_u1__abc_73914_new_n152_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n219_), .Y(u2_u1__0b1_last_row_12_0__4_));
OAI21X1 OAI21X1_875 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_5_), .Y(u2_u1__abc_73914_new_n221_));
OAI21X1 OAI21X1_876 ( .A(u2_u1__abc_73914_new_n155_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n221_), .Y(u2_u1__0b1_last_row_12_0__5_));
OAI21X1 OAI21X1_877 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_73914_new_n223_));
OAI21X1 OAI21X1_878 ( .A(u2_u1__abc_73914_new_n158_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n223_), .Y(u2_u1__0b1_last_row_12_0__6_));
OAI21X1 OAI21X1_879 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_7_), .Y(u2_u1__abc_73914_new_n225_));
OAI21X1 OAI21X1_88 ( .A(_abc_81086_new_n379_), .B(lmr_sel), .C(_abc_81086_new_n380_), .Y(csc_s_4_));
OAI21X1 OAI21X1_880 ( .A(u2_u1__abc_73914_new_n161_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n225_), .Y(u2_u1__0b1_last_row_12_0__7_));
OAI21X1 OAI21X1_881 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_73914_new_n227_));
OAI21X1 OAI21X1_882 ( .A(u2_u1__abc_73914_new_n164_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n227_), .Y(u2_u1__0b1_last_row_12_0__8_));
OAI21X1 OAI21X1_883 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_9_), .Y(u2_u1__abc_73914_new_n229_));
OAI21X1 OAI21X1_884 ( .A(u2_u1__abc_73914_new_n167_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n229_), .Y(u2_u1__0b1_last_row_12_0__9_));
OAI21X1 OAI21X1_885 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_10_), .Y(u2_u1__abc_73914_new_n231_));
OAI21X1 OAI21X1_886 ( .A(u2_u1__abc_73914_new_n170_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n231_), .Y(u2_u1__0b1_last_row_12_0__10_));
OAI21X1 OAI21X1_887 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_11_), .Y(u2_u1__abc_73914_new_n233_));
OAI21X1 OAI21X1_888 ( .A(u2_u1__abc_73914_new_n173_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n233_), .Y(u2_u1__0b1_last_row_12_0__11_));
OAI21X1 OAI21X1_889 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1_b1_last_row_12_), .Y(u2_u1__abc_73914_new_n235_));
OAI21X1 OAI21X1_89 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_5_), .Y(_abc_81086_new_n383_));
OAI21X1 OAI21X1_890 ( .A(u2_u1__abc_73914_new_n176_), .B(u2_u1__abc_73914_new_n210_), .C(u2_u1__abc_73914_new_n235_), .Y(u2_u1__0b1_last_row_12_0__12_));
OAI21X1 OAI21X1_891 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_0_), .Y(u2_u1__abc_73914_new_n240_));
OAI21X1 OAI21X1_892 ( .A(u2_u1__abc_73914_new_n136_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n240_), .Y(u2_u1__0b2_last_row_12_0__0_));
OAI21X1 OAI21X1_893 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_1_), .Y(u2_u1__abc_73914_new_n242_));
OAI21X1 OAI21X1_894 ( .A(u2_u1__abc_73914_new_n143_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n242_), .Y(u2_u1__0b2_last_row_12_0__1_));
OAI21X1 OAI21X1_895 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_73914_new_n244_));
OAI21X1 OAI21X1_896 ( .A(u2_u1__abc_73914_new_n146_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n244_), .Y(u2_u1__0b2_last_row_12_0__2_));
OAI21X1 OAI21X1_897 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_73914_new_n246_));
OAI21X1 OAI21X1_898 ( .A(u2_u1__abc_73914_new_n149_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n246_), .Y(u2_u1__0b2_last_row_12_0__3_));
OAI21X1 OAI21X1_899 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_4_), .Y(u2_u1__abc_73914_new_n248_));
OAI21X1 OAI21X1_9 ( .A(_abc_81086_new_n247_), .B(_abc_81086_new_n249_), .C(_abc_81086_new_n248_), .Y(obct_cs_2_));
OAI21X1 OAI21X1_90 ( .A(_abc_81086_new_n382_), .B(lmr_sel), .C(_abc_81086_new_n383_), .Y(csc_s_5_));
OAI21X1 OAI21X1_900 ( .A(u2_u1__abc_73914_new_n152_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n248_), .Y(u2_u1__0b2_last_row_12_0__4_));
OAI21X1 OAI21X1_901 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_73914_new_n250_));
OAI21X1 OAI21X1_902 ( .A(u2_u1__abc_73914_new_n155_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n250_), .Y(u2_u1__0b2_last_row_12_0__5_));
OAI21X1 OAI21X1_903 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_6_), .Y(u2_u1__abc_73914_new_n252_));
OAI21X1 OAI21X1_904 ( .A(u2_u1__abc_73914_new_n158_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n252_), .Y(u2_u1__0b2_last_row_12_0__6_));
OAI21X1 OAI21X1_905 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_73914_new_n254_));
OAI21X1 OAI21X1_906 ( .A(u2_u1__abc_73914_new_n161_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n254_), .Y(u2_u1__0b2_last_row_12_0__7_));
OAI21X1 OAI21X1_907 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_8_), .Y(u2_u1__abc_73914_new_n256_));
OAI21X1 OAI21X1_908 ( .A(u2_u1__abc_73914_new_n164_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n256_), .Y(u2_u1__0b2_last_row_12_0__8_));
OAI21X1 OAI21X1_909 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_9_), .Y(u2_u1__abc_73914_new_n258_));
OAI21X1 OAI21X1_91 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_6_), .Y(_abc_81086_new_n386_));
OAI21X1 OAI21X1_910 ( .A(u2_u1__abc_73914_new_n167_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n258_), .Y(u2_u1__0b2_last_row_12_0__9_));
OAI21X1 OAI21X1_911 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_73914_new_n260_));
OAI21X1 OAI21X1_912 ( .A(u2_u1__abc_73914_new_n170_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n260_), .Y(u2_u1__0b2_last_row_12_0__10_));
OAI21X1 OAI21X1_913 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_11_), .Y(u2_u1__abc_73914_new_n262_));
OAI21X1 OAI21X1_914 ( .A(u2_u1__abc_73914_new_n173_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n262_), .Y(u2_u1__0b2_last_row_12_0__11_));
OAI21X1 OAI21X1_915 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1_b2_last_row_12_), .Y(u2_u1__abc_73914_new_n264_));
OAI21X1 OAI21X1_916 ( .A(u2_u1__abc_73914_new_n176_), .B(u2_u1__abc_73914_new_n238_), .C(u2_u1__abc_73914_new_n264_), .Y(u2_u1__0b2_last_row_12_0__12_));
OAI21X1 OAI21X1_917 ( .A(u2_u1__abc_73914_new_n285_), .B(u2_u1__abc_73914_new_n286_), .C(u2_u1__abc_73914_new_n284_), .Y(u2_u1__abc_73914_new_n287_));
OAI21X1 OAI21X1_918 ( .A(u2_u1__abc_73914_new_n289_), .B(u2_u1__abc_73914_new_n288_), .C(u2_u1__abc_73914_new_n291_), .Y(u2_u1__abc_73914_new_n292_));
OAI21X1 OAI21X1_919 ( .A(u2_u1__abc_73914_new_n385_), .B(u2_u1__abc_73914_new_n386_), .C(u2_u1__abc_73914_new_n384_), .Y(u2_u1__abc_73914_new_n387_));
OAI21X1 OAI21X1_92 ( .A(_abc_81086_new_n385_), .B(lmr_sel), .C(_abc_81086_new_n386_), .Y(csc_s_6_));
OAI21X1 OAI21X1_920 ( .A(u2_u1__abc_73914_new_n390_), .B(u2_u1__abc_73914_new_n389_), .C(u2_u1__abc_73914_new_n388_), .Y(u2_u1__abc_73914_new_n391_));
OAI21X1 OAI21X1_921 ( .A(u2_u1__abc_73914_new_n399_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1__abc_73914_new_n400_), .Y(u2_u1__abc_73914_new_n401_));
OAI21X1 OAI21X1_922 ( .A(u2_u1__abc_73914_new_n398_), .B(u2_u1__abc_73914_new_n179_), .C(u2_u1__abc_73914_new_n402_), .Y(u2_bank_open_1));
OAI21X1 OAI21X1_923 ( .A(u2_u1__abc_73914_new_n404_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1__abc_73914_new_n406_), .Y(u2_u1__abc_73914_new_n407_));
OAI21X1 OAI21X1_924 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n239_), .C(u2_u1__abc_73914_new_n407_), .Y(u2_u1__0bank2_open_0_0_));
OAI21X1 OAI21X1_925 ( .A(u2_u1__abc_73914_new_n404_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1__abc_73914_new_n410_), .Y(u2_u1__abc_73914_new_n411_));
OAI21X1 OAI21X1_926 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n137_), .C(u2_u1__abc_73914_new_n411_), .Y(u2_u1__0bank3_open_0_0_));
OAI21X1 OAI21X1_927 ( .A(u2_u1__abc_73914_new_n404_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1__abc_73914_new_n415_), .Y(u2_u1__abc_73914_new_n416_));
OAI21X1 OAI21X1_928 ( .A(u2_u1__abc_73914_new_n140_), .B(u2_u1__abc_73914_new_n209_), .C(u2_u1__abc_73914_new_n416_), .Y(u2_u1__0bank1_open_0_0_));
OAI21X1 OAI21X1_929 ( .A(u2_u1__abc_73914_new_n419_), .B(u2_u1__abc_73914_new_n418_), .C(u2_u1__abc_73914_new_n181_), .Y(u2_u1__0bank0_open_0_0_));
OAI21X1 OAI21X1_93 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_7_), .Y(_abc_81086_new_n389_));
OAI21X1 OAI21X1_930 ( .A(u3__abc_73372_new_n278_), .B(u3__abc_73372_new_n285_), .C(u3__abc_73372_new_n286_), .Y(u3__0mc_dp_o_3_0__0_));
OAI21X1 OAI21X1_931 ( .A(u3__abc_73372_new_n278_), .B(u3__abc_73372_new_n294_), .C(u3__abc_73372_new_n295_), .Y(u3__0mc_dp_o_3_0__1_));
OAI21X1 OAI21X1_932 ( .A(u3__abc_73372_new_n278_), .B(u3__abc_73372_new_n303_), .C(u3__abc_73372_new_n304_), .Y(u3__0mc_dp_o_3_0__2_));
OAI21X1 OAI21X1_933 ( .A(u3__abc_73372_new_n278_), .B(u3__abc_73372_new_n312_), .C(u3__abc_73372_new_n313_), .Y(u3__0mc_dp_o_3_0__3_));
OAI21X1 OAI21X1_934 ( .A(u3__abc_73372_new_n343_), .B(u3__abc_73372_new_n346_), .C(u3__abc_73372_new_n347_), .Y(u3__abc_73372_new_n348_));
OAI21X1 OAI21X1_935 ( .A(u3__abc_73372_new_n341_), .B(u3__abc_73372_new_n342_), .C(u3__abc_73372_new_n348_), .Y(u3__abc_73372_new_n349_));
OAI21X1 OAI21X1_936 ( .A(u3__abc_73372_new_n315_), .B(u3__abc_73372_new_n340_), .C(u3__abc_73372_new_n349_), .Y(u3__0byte1_7_0__0_));
OAI21X1 OAI21X1_937 ( .A(u3__abc_73372_new_n351_), .B(u3__abc_73372_new_n346_), .C(u3__abc_73372_new_n352_), .Y(u3__abc_73372_new_n353_));
OAI21X1 OAI21X1_938 ( .A(u3__abc_73372_new_n341_), .B(u3__abc_73372_new_n342_), .C(u3__abc_73372_new_n353_), .Y(u3__abc_73372_new_n354_));
OAI21X1 OAI21X1_939 ( .A(u3__abc_73372_new_n318_), .B(u3__abc_73372_new_n340_), .C(u3__abc_73372_new_n354_), .Y(u3__0byte1_7_0__1_));
OAI21X1 OAI21X1_94 ( .A(_abc_81086_new_n388_), .B(lmr_sel), .C(_abc_81086_new_n389_), .Y(csc_s_7_));
OAI21X1 OAI21X1_940 ( .A(u3__abc_73372_new_n356_), .B(u3__abc_73372_new_n346_), .C(u3__abc_73372_new_n357_), .Y(u3__abc_73372_new_n358_));
OAI21X1 OAI21X1_941 ( .A(u3__abc_73372_new_n341_), .B(u3__abc_73372_new_n342_), .C(u3__abc_73372_new_n358_), .Y(u3__abc_73372_new_n359_));
OAI21X1 OAI21X1_942 ( .A(u3__abc_73372_new_n321_), .B(u3__abc_73372_new_n340_), .C(u3__abc_73372_new_n359_), .Y(u3__0byte1_7_0__2_));
OAI21X1 OAI21X1_943 ( .A(u3__abc_73372_new_n361_), .B(u3__abc_73372_new_n346_), .C(u3__abc_73372_new_n362_), .Y(u3__abc_73372_new_n363_));
OAI21X1 OAI21X1_944 ( .A(u3__abc_73372_new_n341_), .B(u3__abc_73372_new_n342_), .C(u3__abc_73372_new_n363_), .Y(u3__abc_73372_new_n364_));
OAI21X1 OAI21X1_945 ( .A(u3__abc_73372_new_n324_), .B(u3__abc_73372_new_n340_), .C(u3__abc_73372_new_n364_), .Y(u3__0byte1_7_0__3_));
OAI21X1 OAI21X1_946 ( .A(u3__abc_73372_new_n366_), .B(u3__abc_73372_new_n346_), .C(u3__abc_73372_new_n367_), .Y(u3__abc_73372_new_n368_));
OAI21X1 OAI21X1_947 ( .A(u3__abc_73372_new_n341_), .B(u3__abc_73372_new_n342_), .C(u3__abc_73372_new_n368_), .Y(u3__abc_73372_new_n369_));
OAI21X1 OAI21X1_948 ( .A(u3__abc_73372_new_n327_), .B(u3__abc_73372_new_n340_), .C(u3__abc_73372_new_n369_), .Y(u3__0byte1_7_0__4_));
OAI21X1 OAI21X1_949 ( .A(u3__abc_73372_new_n371_), .B(u3__abc_73372_new_n346_), .C(u3__abc_73372_new_n372_), .Y(u3__abc_73372_new_n373_));
OAI21X1 OAI21X1_95 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_9_), .Y(_abc_81086_new_n395_));
OAI21X1 OAI21X1_950 ( .A(u3__abc_73372_new_n341_), .B(u3__abc_73372_new_n342_), .C(u3__abc_73372_new_n373_), .Y(u3__abc_73372_new_n374_));
OAI21X1 OAI21X1_951 ( .A(u3__abc_73372_new_n330_), .B(u3__abc_73372_new_n340_), .C(u3__abc_73372_new_n374_), .Y(u3__0byte1_7_0__5_));
OAI21X1 OAI21X1_952 ( .A(u3__abc_73372_new_n376_), .B(u3__abc_73372_new_n346_), .C(u3__abc_73372_new_n377_), .Y(u3__abc_73372_new_n378_));
OAI21X1 OAI21X1_953 ( .A(u3__abc_73372_new_n341_), .B(u3__abc_73372_new_n342_), .C(u3__abc_73372_new_n378_), .Y(u3__abc_73372_new_n379_));
OAI21X1 OAI21X1_954 ( .A(u3__abc_73372_new_n333_), .B(u3__abc_73372_new_n340_), .C(u3__abc_73372_new_n379_), .Y(u3__0byte1_7_0__6_));
OAI21X1 OAI21X1_955 ( .A(u3__abc_73372_new_n381_), .B(u3__abc_73372_new_n346_), .C(u3__abc_73372_new_n382_), .Y(u3__abc_73372_new_n383_));
OAI21X1 OAI21X1_956 ( .A(u3__abc_73372_new_n341_), .B(u3__abc_73372_new_n342_), .C(u3__abc_73372_new_n383_), .Y(u3__abc_73372_new_n384_));
OAI21X1 OAI21X1_957 ( .A(u3__abc_73372_new_n336_), .B(u3__abc_73372_new_n340_), .C(u3__abc_73372_new_n384_), .Y(u3__0byte1_7_0__7_));
OAI21X1 OAI21X1_958 ( .A(u3__abc_73372_new_n402_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n403_), .Y(u3__0mc_data_o_31_0__0_));
OAI21X1 OAI21X1_959 ( .A(u3__abc_73372_new_n405_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n406_), .Y(u3__0mc_data_o_31_0__1_));
OAI21X1 OAI21X1_96 ( .A(_abc_81086_new_n394_), .B(lmr_sel), .C(_abc_81086_new_n395_), .Y(u1_bas));
OAI21X1 OAI21X1_960 ( .A(u3__abc_73372_new_n408_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n409_), .Y(u3__0mc_data_o_31_0__2_));
OAI21X1 OAI21X1_961 ( .A(u3__abc_73372_new_n411_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n412_), .Y(u3__0mc_data_o_31_0__3_));
OAI21X1 OAI21X1_962 ( .A(u3__abc_73372_new_n414_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n415_), .Y(u3__0mc_data_o_31_0__4_));
OAI21X1 OAI21X1_963 ( .A(u3__abc_73372_new_n417_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n418_), .Y(u3__0mc_data_o_31_0__5_));
OAI21X1 OAI21X1_964 ( .A(u3__abc_73372_new_n420_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n421_), .Y(u3__0mc_data_o_31_0__6_));
OAI21X1 OAI21X1_965 ( .A(u3__abc_73372_new_n423_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n424_), .Y(u3__0mc_data_o_31_0__7_));
OAI21X1 OAI21X1_966 ( .A(u3__abc_73372_new_n426_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n427_), .Y(u3__0mc_data_o_31_0__8_));
OAI21X1 OAI21X1_967 ( .A(u3__abc_73372_new_n429_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n430_), .Y(u3__0mc_data_o_31_0__9_));
OAI21X1 OAI21X1_968 ( .A(u3__abc_73372_new_n432_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n433_), .Y(u3__0mc_data_o_31_0__10_));
OAI21X1 OAI21X1_969 ( .A(u3__abc_73372_new_n435_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n436_), .Y(u3__0mc_data_o_31_0__11_));
OAI21X1 OAI21X1_97 ( .A(init_ack), .B(lmr_ack), .C(sp_csc_10_), .Y(_abc_81086_new_n398_));
OAI21X1 OAI21X1_970 ( .A(u3__abc_73372_new_n438_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n439_), .Y(u3__0mc_data_o_31_0__12_));
OAI21X1 OAI21X1_971 ( .A(u3__abc_73372_new_n441_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n442_), .Y(u3__0mc_data_o_31_0__13_));
OAI21X1 OAI21X1_972 ( .A(u3__abc_73372_new_n444_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n445_), .Y(u3__0mc_data_o_31_0__14_));
OAI21X1 OAI21X1_973 ( .A(u3__abc_73372_new_n447_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n448_), .Y(u3__0mc_data_o_31_0__15_));
OAI21X1 OAI21X1_974 ( .A(u3__abc_73372_new_n450_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n451_), .Y(u3__0mc_data_o_31_0__16_));
OAI21X1 OAI21X1_975 ( .A(u3__abc_73372_new_n453_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n454_), .Y(u3__0mc_data_o_31_0__17_));
OAI21X1 OAI21X1_976 ( .A(u3__abc_73372_new_n456_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n457_), .Y(u3__0mc_data_o_31_0__18_));
OAI21X1 OAI21X1_977 ( .A(u3__abc_73372_new_n459_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n460_), .Y(u3__0mc_data_o_31_0__19_));
OAI21X1 OAI21X1_978 ( .A(u3__abc_73372_new_n462_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n463_), .Y(u3__0mc_data_o_31_0__20_));
OAI21X1 OAI21X1_979 ( .A(u3__abc_73372_new_n465_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n466_), .Y(u3__0mc_data_o_31_0__21_));
OAI21X1 OAI21X1_98 ( .A(_abc_81086_new_n397_), .B(lmr_sel), .C(_abc_81086_new_n398_), .Y(u5_kro));
OAI21X1 OAI21X1_980 ( .A(u3__abc_73372_new_n468_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n469_), .Y(u3__0mc_data_o_31_0__22_));
OAI21X1 OAI21X1_981 ( .A(u3__abc_73372_new_n471_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n472_), .Y(u3__0mc_data_o_31_0__23_));
OAI21X1 OAI21X1_982 ( .A(u3__abc_73372_new_n474_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n475_), .Y(u3__0mc_data_o_31_0__24_));
OAI21X1 OAI21X1_983 ( .A(u3__abc_73372_new_n477_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n478_), .Y(u3__0mc_data_o_31_0__25_));
OAI21X1 OAI21X1_984 ( .A(u3__abc_73372_new_n480_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n481_), .Y(u3__0mc_data_o_31_0__26_));
OAI21X1 OAI21X1_985 ( .A(u3__abc_73372_new_n483_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n484_), .Y(u3__0mc_data_o_31_0__27_));
OAI21X1 OAI21X1_986 ( .A(u3__abc_73372_new_n486_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n487_), .Y(u3__0mc_data_o_31_0__28_));
OAI21X1 OAI21X1_987 ( .A(u3__abc_73372_new_n489_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n490_), .Y(u3__0mc_data_o_31_0__29_));
OAI21X1 OAI21X1_988 ( .A(u3__abc_73372_new_n492_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n493_), .Y(u3__0mc_data_o_31_0__30_));
OAI21X1 OAI21X1_989 ( .A(u3__abc_73372_new_n495_), .B(u3__abc_73372_new_n277_), .C(u3__abc_73372_new_n496_), .Y(u3__0mc_data_o_31_0__31_));
OAI21X1 OAI21X1_99 ( .A(u0_init_req0), .B(u0__abc_74894_new_n1101_), .C(u0__abc_74894_new_n1103_), .Y(u0__abc_74894_new_n1104_));
OAI21X1 OAI21X1_990 ( .A(csc_5_), .B(u3_byte0_0_), .C(u3__abc_73372_new_n498_), .Y(u3__abc_73372_new_n499_));
OAI21X1 OAI21X1_991 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n499_), .C(u3__abc_73372_new_n500_), .Y(mem_dout_0_));
OAI21X1 OAI21X1_992 ( .A(csc_5_), .B(u3_byte0_1_), .C(u3__abc_73372_new_n502_), .Y(u3__abc_73372_new_n503_));
OAI21X1 OAI21X1_993 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n503_), .C(u3__abc_73372_new_n504_), .Y(mem_dout_1_));
OAI21X1 OAI21X1_994 ( .A(csc_5_), .B(u3_byte0_2_), .C(u3__abc_73372_new_n506_), .Y(u3__abc_73372_new_n507_));
OAI21X1 OAI21X1_995 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n507_), .C(u3__abc_73372_new_n508_), .Y(mem_dout_2_));
OAI21X1 OAI21X1_996 ( .A(csc_5_), .B(u3_byte0_3_), .C(u3__abc_73372_new_n510_), .Y(u3__abc_73372_new_n511_));
OAI21X1 OAI21X1_997 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n511_), .C(u3__abc_73372_new_n512_), .Y(mem_dout_3_));
OAI21X1 OAI21X1_998 ( .A(csc_5_), .B(u3_byte0_4_), .C(u3__abc_73372_new_n514_), .Y(u3__abc_73372_new_n515_));
OAI21X1 OAI21X1_999 ( .A(u3__abc_73372_new_n275_), .B(u3__abc_73372_new_n515_), .C(u3__abc_73372_new_n516_), .Y(mem_dout_4_));
OAI22X1 OAI22X1_1 ( .A(u0_sreq_cs_le), .B(u0__abc_74894_new_n1106_), .C(u0__abc_74894_new_n1110_), .D(u0__abc_74894_new_n1107_), .Y(u0__0spec_req_cs_7_0__1_));
OAI22X1 OAI22X1_10 ( .A(u0__abc_74894_new_n1299_), .B(u0__abc_74894_new_n3719_), .C(u0__abc_74894_new_n1297_), .D(u0__abc_74894_new_n3716_), .Y(u0__abc_74894_new_n3884_));
OAI22X1 OAI22X1_100 ( .A(u5__abc_78290_new_n763_), .B(u5_cmd_asserted), .C(u5__abc_78290_new_n2745_), .D(u5__abc_78290_new_n1412_), .Y(u5__abc_78290_new_n2746_));
OAI22X1 OAI22X1_101 ( .A(u5__abc_78290_new_n2615_), .B(u5__abc_78290_new_n2760_), .C(u5__abc_78290_new_n1229_), .D(u5__abc_78290_new_n2761_), .Y(u5__abc_78290_new_n2762_));
OAI22X1 OAI22X1_102 ( .A(u5_cmd_asserted), .B(u5__abc_78290_new_n553_), .C(u5__abc_78290_new_n2831_), .D(u5__abc_78290_new_n2830_), .Y(u5_next_state_27_));
OAI22X1 OAI22X1_103 ( .A(u5__abc_78290_new_n2873_), .B(u5__abc_78290_new_n2875_), .C(u5__abc_78290_new_n662_), .D(u5__abc_78290_new_n2584_), .Y(u5_next_state_38_));
OAI22X1 OAI22X1_104 ( .A(u5__abc_78290_new_n1335_), .B(u5__abc_78290_new_n2919_), .C(u5__abc_78290_new_n946_), .D(u5__abc_78290_new_n2591_), .Y(u5__abc_78290_new_n2920_));
OAI22X1 OAI22X1_105 ( .A(u5__abc_78290_new_n846_), .B(u5__abc_78290_new_n2591_), .C(u5__abc_78290_new_n1335_), .D(u5__abc_78290_new_n2967_), .Y(u5__abc_78290_new_n2968_));
OAI22X1 OAI22X1_106 ( .A(u5__abc_78290_new_n1363_), .B(u5__abc_78290_new_n3027_), .C(u5__abc_78290_new_n1186_), .D(u5__abc_78290_new_n3033_), .Y(mc_bg_d));
OAI22X1 OAI22X1_107 ( .A(u6__abc_81318_new_n142_), .B(u6__abc_81318_new_n144_), .C(u6__abc_81318_new_n135_), .D(u6__abc_81318_new_n141_), .Y(u6__0wb_ack_o_0_0_));
OAI22X1 OAI22X1_11 ( .A(u0__abc_74894_new_n1312_), .B(u0__abc_74894_new_n3736_), .C(u0__abc_74894_new_n1953_), .D(u0__abc_74894_new_n3733_), .Y(u0__abc_74894_new_n3890_));
OAI22X1 OAI22X1_12 ( .A(u0__abc_74894_new_n3517_), .B(u0__abc_74894_new_n3750_), .C(u0__abc_74894_new_n3619_), .D(u0__abc_74894_new_n3845_), .Y(u0__abc_74894_new_n3895_));
OAI22X1 OAI22X1_13 ( .A(u0__abc_74894_new_n1332_), .B(u0__abc_74894_new_n3736_), .C(u0__abc_74894_new_n1973_), .D(u0__abc_74894_new_n3733_), .Y(u0__abc_74894_new_n3913_));
OAI22X1 OAI22X1_14 ( .A(u0__abc_74894_new_n1430_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n2073_), .D(u0__abc_74894_new_n3733_), .Y(u0__abc_74894_new_n3999_));
OAI22X1 OAI22X1_15 ( .A(u0__abc_74894_new_n1439_), .B(u0__abc_74894_new_n3719_), .C(u0__abc_74894_new_n1450_), .D(u0__abc_74894_new_n3748_), .Y(u0__abc_74894_new_n4021_));
OAI22X1 OAI22X1_16 ( .A(u0__abc_74894_new_n1472_), .B(u0__abc_74894_new_n3736_), .C(u0__abc_74894_new_n2111_), .D(u0__abc_74894_new_n3732_), .Y(u0__abc_74894_new_n4042_));
OAI22X1 OAI22X1_17 ( .A(u0__abc_74894_new_n1512_), .B(u0__abc_74894_new_n3736_), .C(u0__abc_74894_new_n2151_), .D(u0__abc_74894_new_n3732_), .Y(u0__abc_74894_new_n4084_));
OAI22X1 OAI22X1_18 ( .A(u0__abc_74894_new_n1532_), .B(u0__abc_74894_new_n3736_), .C(u0__abc_74894_new_n2171_), .D(u0__abc_74894_new_n3732_), .Y(u0__abc_74894_new_n4106_));
OAI22X1 OAI22X1_19 ( .A(u0__abc_74894_new_n1550_), .B(u0__abc_74894_new_n3748_), .C(u0__abc_74894_new_n2193_), .D(u0__abc_74894_new_n3733_), .Y(u0__abc_74894_new_n4129_));
OAI22X1 OAI22X1_2 ( .A(u0_sreq_cs_le), .B(u0__abc_74894_new_n1112_), .C(u0__abc_74894_new_n1115_), .D(u0__abc_74894_new_n1117_), .Y(u0__0spec_req_cs_7_0__2_));
OAI22X1 OAI22X1_20 ( .A(u0_u0__abc_72207_new_n435_), .B(u0_u0__abc_72207_new_n436_), .C(u0_u0__abc_72207_new_n437_), .D(u0_u0__abc_72207_new_n438_), .Y(u0_u0__abc_72207_new_n439_));
OAI22X1 OAI22X1_21 ( .A(u0_u0__abc_72207_new_n443_), .B(u0_u0__abc_72207_new_n444_), .C(u0_u0__abc_72207_new_n445_), .D(u0_u0__abc_72207_new_n446_), .Y(u0_u0__abc_72207_new_n447_));
OAI22X1 OAI22X1_22 ( .A(u0_u0__abc_72207_new_n452_), .B(u0_u0__abc_72207_new_n453_), .C(u0_u0__abc_72207_new_n454_), .D(u0_u0__abc_72207_new_n455_), .Y(u0_u0__abc_72207_new_n456_));
OAI22X1 OAI22X1_23 ( .A(u0_init_ack0), .B(u0_u0__abc_72207_new_n462_), .C(u0_u0__abc_72207_new_n208_), .D(u0_u0__abc_72207_new_n464_), .Y(u0_u0__0init_req_0_0_));
OAI22X1 OAI22X1_24 ( .A(u0_u1__abc_72470_new_n412_), .B(u0_u1__abc_72470_new_n413_), .C(u0_u1__abc_72470_new_n414_), .D(u0_u1__abc_72470_new_n415_), .Y(u0_u1__abc_72470_new_n416_));
OAI22X1 OAI22X1_25 ( .A(u0_u1__abc_72470_new_n419_), .B(u0_u1__abc_72470_new_n420_), .C(u0_u1__abc_72470_new_n421_), .D(u0_u1__abc_72470_new_n422_), .Y(u0_u1__abc_72470_new_n423_));
OAI22X1 OAI22X1_26 ( .A(u0_u1__abc_72470_new_n428_), .B(u0_u1__abc_72470_new_n429_), .C(u0_u1__abc_72470_new_n430_), .D(u0_u1__abc_72470_new_n431_), .Y(u0_u1__abc_72470_new_n432_));
OAI22X1 OAI22X1_27 ( .A(u0_init_ack1), .B(u0_u1__abc_72470_new_n438_), .C(u0_u1__abc_72470_new_n440_), .D(u0_u1__abc_72470_new_n204_), .Y(u0_u1__0init_req_0_0_));
OAI22X1 OAI22X1_28 ( .A(u1__abc_72801_new_n258_), .B(u1__abc_72801_new_n259_), .C(u1__abc_72801_new_n261_), .D(u1__abc_72801_new_n263_), .Y(u1__abc_72801_new_n264_));
OAI22X1 OAI22X1_29 ( .A(u1__abc_72801_new_n259_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n263_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n299_));
OAI22X1 OAI22X1_3 ( .A(u0_sreq_cs_le), .B(u0__abc_74894_new_n1119_), .C(u0__abc_74894_new_n1123_), .D(u0__abc_74894_new_n1117_), .Y(u0__0spec_req_cs_7_0__3_));
OAI22X1 OAI22X1_30 ( .A(u1__abc_72801_new_n276_), .B(cs_le), .C(u1__abc_72801_new_n286_), .D(u1__abc_72801_new_n305_), .Y(u1__0bank_adr_1_0__0_));
OAI22X1 OAI22X1_31 ( .A(cs_le), .B(u1__abc_72801_new_n307_), .C(u1__abc_72801_new_n311_), .D(u1__abc_72801_new_n320_), .Y(u1__0bank_adr_1_0__1_));
OAI22X1 OAI22X1_32 ( .A(u1__abc_72801_new_n259_), .B(u1__abc_72801_new_n288_), .C(u1__abc_72801_new_n261_), .D(u1__abc_72801_new_n266_), .Y(u1__abc_72801_new_n350_));
OAI22X1 OAI22X1_33 ( .A(u1__abc_72801_new_n423_), .B(u1__abc_72801_new_n336_), .C(u1__abc_72801_new_n422_), .D(u1__abc_72801_new_n282_), .Y(u1__abc_72801_new_n424_));
OAI22X1 OAI22X1_34 ( .A(cs_le), .B(u1__abc_72801_new_n441_), .C(u1__abc_72801_new_n451_), .D(u1__abc_72801_new_n446_), .Y(u1__0row_adr_12_0__11_));
OAI22X1 OAI22X1_35 ( .A(u1__abc_72801_new_n464_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n467_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n507_));
OAI22X1 OAI22X1_36 ( .A(u1__abc_72801_new_n467_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n470_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n512_));
OAI22X1 OAI22X1_37 ( .A(u1__abc_72801_new_n470_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n473_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n517_));
OAI22X1 OAI22X1_38 ( .A(u1__abc_72801_new_n473_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n476_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n522_));
OAI22X1 OAI22X1_39 ( .A(u1__abc_72801_new_n476_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n479_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n527_));
OAI22X1 OAI22X1_4 ( .A(u0_sreq_cs_le), .B(u0__abc_74894_new_n1125_), .C(u0__abc_74894_new_n1129_), .D(u0__abc_74894_new_n1132_), .Y(u0__0spec_req_cs_7_0__4_));
OAI22X1 OAI22X1_40 ( .A(u1__abc_72801_new_n479_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n482_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n532_));
OAI22X1 OAI22X1_41 ( .A(u1__abc_72801_new_n537_), .B(u1__abc_72801_new_n288_), .C(u1__abc_72801_new_n482_), .D(u1__abc_72801_new_n261_), .Y(u1__abc_72801_new_n538_));
OAI22X1 OAI22X1_42 ( .A(u1__abc_72801_new_n543_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n277_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n550_));
OAI22X1 OAI22X1_43 ( .A(u1__abc_72801_new_n277_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n308_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n555_));
OAI22X1 OAI22X1_44 ( .A(u1__abc_72801_new_n308_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n324_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n560_));
OAI22X1 OAI22X1_45 ( .A(u1__abc_72801_new_n324_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n332_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n565_));
OAI22X1 OAI22X1_46 ( .A(u1__abc_72801_new_n399_), .B(u1__abc_72801_new_n261_), .C(u1__abc_72801_new_n408_), .D(u1__abc_72801_new_n288_), .Y(u1__abc_72801_new_n593_));
OAI22X1 OAI22X1_47 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n687_), .C(u1__abc_72801_new_n688_), .D(u1__abc_72801_new_n681_), .Y(mc_addr_d_0_));
OAI22X1 OAI22X1_48 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n695_), .C(u1__abc_72801_new_n696_), .D(u1__abc_72801_new_n692_), .Y(mc_addr_d_1_));
OAI22X1 OAI22X1_49 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n704_), .C(u1__abc_72801_new_n705_), .D(u1__abc_72801_new_n700_), .Y(mc_addr_d_2_));
OAI22X1 OAI22X1_5 ( .A(u0_sreq_cs_le), .B(u0__abc_74894_new_n1134_), .C(u0__abc_74894_new_n1138_), .D(u0__abc_74894_new_n1132_), .Y(u0__0spec_req_cs_7_0__5_));
OAI22X1 OAI22X1_50 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n712_), .C(u1__abc_72801_new_n713_), .D(u1__abc_72801_new_n709_), .Y(mc_addr_d_3_));
OAI22X1 OAI22X1_51 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n720_), .C(u1__abc_72801_new_n721_), .D(u1__abc_72801_new_n717_), .Y(mc_addr_d_4_));
OAI22X1 OAI22X1_52 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n728_), .C(u1__abc_72801_new_n729_), .D(u1__abc_72801_new_n725_), .Y(mc_addr_d_5_));
OAI22X1 OAI22X1_53 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n736_), .C(u1__abc_72801_new_n737_), .D(u1__abc_72801_new_n733_), .Y(mc_addr_d_6_));
OAI22X1 OAI22X1_54 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n744_), .C(u1__abc_72801_new_n745_), .D(u1__abc_72801_new_n741_), .Y(mc_addr_d_7_));
OAI22X1 OAI22X1_55 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n752_), .C(u1__abc_72801_new_n753_), .D(u1__abc_72801_new_n749_), .Y(mc_addr_d_8_));
OAI22X1 OAI22X1_56 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n761_), .C(u1__abc_72801_new_n762_), .D(u1__abc_72801_new_n757_), .Y(mc_addr_d_9_));
OAI22X1 OAI22X1_57 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n769_), .C(u1__abc_72801_new_n770_), .D(u1__abc_72801_new_n766_), .Y(mc_addr_d_11_));
OAI22X1 OAI22X1_58 ( .A(u1__abc_72801_new_n673_), .B(u1__abc_72801_new_n777_), .C(u1__abc_72801_new_n778_), .D(u1__abc_72801_new_n774_), .Y(mc_addr_d_12_));
OAI22X1 OAI22X1_59 ( .A(u1__abc_72801_new_n276_), .B(u1__abc_72801_new_n673_), .C(u1__abc_72801_new_n783_), .D(u1__abc_72801_new_n782_), .Y(mc_addr_d_13_));
OAI22X1 OAI22X1_6 ( .A(u0_sreq_cs_le), .B(u0__abc_74894_new_n1140_), .C(u0__abc_74894_new_n1145_), .D(u0__abc_74894_new_n1132_), .Y(u0__0spec_req_cs_7_0__6_));
OAI22X1 OAI22X1_60 ( .A(u1__abc_72801_new_n307_), .B(u1__abc_72801_new_n673_), .C(u1__abc_72801_new_n788_), .D(u1__abc_72801_new_n787_), .Y(mc_addr_d_14_));
OAI22X1 OAI22X1_61 ( .A(row_adr_8_), .B(u2_u0__abc_73914_new_n266_), .C(u2_u0__abc_73914_new_n267_), .D(row_adr_9_), .Y(u2_u0__abc_73914_new_n268_));
OAI22X1 OAI22X1_62 ( .A(u2_u0_b3_last_row_4_), .B(u2_u0__abc_73914_new_n152_), .C(u2_u0__abc_73914_new_n293_), .D(row_adr_6_), .Y(u2_u0__abc_73914_new_n294_));
OAI22X1 OAI22X1_63 ( .A(row_adr_2_), .B(u2_u0__abc_73914_new_n290_), .C(u2_u0_b3_last_row_6_), .D(u2_u0__abc_73914_new_n158_), .Y(u2_u0__abc_73914_new_n295_));
OAI22X1 OAI22X1_64 ( .A(u2_u0_b1_last_row_0_), .B(u2_u0__abc_73914_new_n136_), .C(u2_u0__abc_73914_new_n143_), .D(u2_u0_b1_last_row_1_), .Y(u2_u0__abc_73914_new_n298_));
OAI22X1 OAI22X1_65 ( .A(row_adr_3_), .B(u2_u0__abc_73914_new_n302_), .C(u2_u0__abc_73914_new_n155_), .D(u2_u0_b1_last_row_5_), .Y(u2_u0__abc_73914_new_n303_));
OAI22X1 OAI22X1_66 ( .A(u2_u0_b2_last_row_8_), .B(u2_u0__abc_73914_new_n164_), .C(u2_u0__abc_73914_new_n167_), .D(u2_u0_b2_last_row_9_), .Y(u2_u0__abc_73914_new_n365_));
OAI22X1 OAI22X1_67 ( .A(row_adr_6_), .B(u2_u0__abc_73914_new_n374_), .C(u2_u0__abc_73914_new_n146_), .D(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_73914_new_n375_));
OAI22X1 OAI22X1_68 ( .A(row_adr_2_), .B(u2_u0__abc_73914_new_n379_), .C(u2_u0__abc_73914_new_n143_), .D(u2_u0_b2_last_row_1_), .Y(u2_u0__abc_73914_new_n380_));
OAI22X1 OAI22X1_69 ( .A(row_adr_8_), .B(u2_u1__abc_73914_new_n266_), .C(u2_u1__abc_73914_new_n267_), .D(row_adr_9_), .Y(u2_u1__abc_73914_new_n268_));
OAI22X1 OAI22X1_7 ( .A(u0_sreq_cs_le), .B(u0__abc_74894_new_n1147_), .C(u0__abc_74894_new_n1152_), .D(u0__abc_74894_new_n1132_), .Y(u0__0spec_req_cs_7_0__7_));
OAI22X1 OAI22X1_70 ( .A(u2_u1_b3_last_row_4_), .B(u2_u1__abc_73914_new_n152_), .C(u2_u1__abc_73914_new_n293_), .D(row_adr_6_), .Y(u2_u1__abc_73914_new_n294_));
OAI22X1 OAI22X1_71 ( .A(row_adr_2_), .B(u2_u1__abc_73914_new_n290_), .C(u2_u1_b3_last_row_6_), .D(u2_u1__abc_73914_new_n158_), .Y(u2_u1__abc_73914_new_n295_));
OAI22X1 OAI22X1_72 ( .A(u2_u1_b1_last_row_0_), .B(u2_u1__abc_73914_new_n136_), .C(u2_u1__abc_73914_new_n143_), .D(u2_u1_b1_last_row_1_), .Y(u2_u1__abc_73914_new_n298_));
OAI22X1 OAI22X1_73 ( .A(row_adr_3_), .B(u2_u1__abc_73914_new_n302_), .C(u2_u1__abc_73914_new_n155_), .D(u2_u1_b1_last_row_5_), .Y(u2_u1__abc_73914_new_n303_));
OAI22X1 OAI22X1_74 ( .A(u2_u1_b2_last_row_8_), .B(u2_u1__abc_73914_new_n164_), .C(u2_u1__abc_73914_new_n167_), .D(u2_u1_b2_last_row_9_), .Y(u2_u1__abc_73914_new_n365_));
OAI22X1 OAI22X1_75 ( .A(row_adr_6_), .B(u2_u1__abc_73914_new_n374_), .C(u2_u1__abc_73914_new_n146_), .D(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_73914_new_n375_));
OAI22X1 OAI22X1_76 ( .A(row_adr_2_), .B(u2_u1__abc_73914_new_n379_), .C(u2_u1__abc_73914_new_n143_), .D(u2_u1_b2_last_row_1_), .Y(u2_u1__abc_73914_new_n380_));
OAI22X1 OAI22X1_77 ( .A(u3__abc_73372_new_n664_), .B(u3__abc_73372_new_n665_), .C(u3__abc_73372_new_n666_), .D(u3__abc_73372_new_n667_), .Y(u3__abc_73372_new_n668_));
OAI22X1 OAI22X1_78 ( .A(u3__abc_73372_new_n671_), .B(u3__abc_73372_new_n672_), .C(u3__abc_73372_new_n669_), .D(u3__abc_73372_new_n670_), .Y(u3__abc_73372_new_n673_));
OAI22X1 OAI22X1_79 ( .A(u3__abc_73372_new_n714_), .B(u3__abc_73372_new_n715_), .C(u3__abc_73372_new_n716_), .D(u3__abc_73372_new_n717_), .Y(u3__abc_73372_new_n718_));
OAI22X1 OAI22X1_8 ( .A(u0__abc_74894_new_n1177_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n1818_), .D(u0__abc_74894_new_n3707_), .Y(u0__abc_74894_new_n3763_));
OAI22X1 OAI22X1_80 ( .A(u3__abc_73372_new_n721_), .B(u3__abc_73372_new_n722_), .C(u3__abc_73372_new_n719_), .D(u3__abc_73372_new_n720_), .Y(u3__abc_73372_new_n723_));
OAI22X1 OAI22X1_81 ( .A(u4__abc_74770_new_n176_), .B(u4__abc_74770_new_n178_), .C(u4__abc_74770_new_n102_), .D(u4__abc_74770_new_n175_), .Y(u4__abc_74770_new_n179_));
OAI22X1 OAI22X1_82 ( .A(u5__abc_78290_new_n670_), .B(u5__abc_78290_new_n681_), .C(u5__abc_78290_new_n671_), .D(u5__abc_78290_new_n676_), .Y(u5__abc_78290_new_n682_));
OAI22X1 OAI22X1_83 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n691_), .C(u5__abc_78290_new_n671_), .D(u5__abc_78290_new_n696_), .Y(u5__abc_78290_new_n697_));
OAI22X1 OAI22X1_84 ( .A(u5__abc_78290_new_n448_), .B(u5__abc_78290_new_n804_), .C(u5__abc_78290_new_n808_), .D(u5__abc_78290_new_n670_), .Y(u5__abc_78290_new_n809_));
OAI22X1 OAI22X1_85 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n719_), .C(u5__abc_78290_new_n671_), .D(u5__abc_78290_new_n676_), .Y(u5__abc_78290_new_n993_));
OAI22X1 OAI22X1_86 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n519_), .C(u5__abc_78290_new_n551_), .D(u5__abc_78290_new_n552_), .Y(u5__abc_78290_new_n998_));
OAI22X1 OAI22X1_87 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n751_), .C(u5__abc_78290_new_n762_), .D(u5__abc_78290_new_n766_), .Y(u5__abc_78290_new_n1002_));
OAI22X1 OAI22X1_88 ( .A(u5__abc_78290_new_n756_), .B(u5__abc_78290_new_n759_), .C(u5__abc_78290_new_n454_), .D(u5__abc_78290_new_n893_), .Y(u5__abc_78290_new_n1005_));
OAI22X1 OAI22X1_89 ( .A(u5__abc_78290_new_n408_), .B(u5__abc_78290_new_n782_), .C(u5__abc_78290_new_n454_), .D(u5__abc_78290_new_n738_), .Y(u5__abc_78290_new_n1006_));
OAI22X1 OAI22X1_9 ( .A(u0__abc_74894_new_n1197_), .B(u0__abc_74894_new_n3716_), .C(u0__abc_74894_new_n1838_), .D(u0__abc_74894_new_n3707_), .Y(u0__abc_74894_new_n3788_));
OAI22X1 OAI22X1_90 ( .A(u5__abc_78290_new_n685_), .B(u5__abc_78290_new_n691_), .C(u5__abc_78290_new_n671_), .D(u5__abc_78290_new_n707_), .Y(u5__abc_78290_new_n2440_));
OAI22X1 OAI22X1_91 ( .A(u5__abc_78290_new_n2433_), .B(u5__abc_78290_new_n2425_), .C(u5__abc_78290_new_n2462_), .D(u5__abc_78290_new_n2460_), .Y(u5__0timer2_8_0__1_));
OAI22X1 OAI22X1_92 ( .A(u5__abc_78290_new_n2133_), .B(u5__abc_78290_new_n2425_), .C(u5__abc_78290_new_n2480_), .D(u5__abc_78290_new_n2508_), .Y(u5__0timer2_8_0__4_));
OAI22X1 OAI22X1_93 ( .A(u5__abc_78290_new_n2244_), .B(u5__abc_78290_new_n2425_), .C(u5__abc_78290_new_n2515_), .D(u5__abc_78290_new_n2518_), .Y(u5__0timer2_8_0__5_));
OAI22X1 OAI22X1_94 ( .A(u5__abc_78290_new_n2264_), .B(u5__abc_78290_new_n2425_), .C(u5__abc_78290_new_n2523_), .D(u5__abc_78290_new_n2524_), .Y(u5__0timer2_8_0__6_));
OAI22X1 OAI22X1_95 ( .A(u5__abc_78290_new_n2308_), .B(u5__abc_78290_new_n2425_), .C(u5__abc_78290_new_n2529_), .D(u5__abc_78290_new_n2524_), .Y(u5__0timer2_8_0__7_));
OAI22X1 OAI22X1_96 ( .A(u5__abc_78290_new_n2506_), .B(u5__abc_78290_new_n2425_), .C(u5__abc_78290_new_n2532_), .D(u5__abc_78290_new_n2524_), .Y(u5__0timer2_8_0__8_));
OAI22X1 OAI22X1_97 ( .A(u5_state_1_), .B(u5_tmr_done), .C(u5__abc_78290_new_n1058_), .D(u5__abc_78290_new_n1311_), .Y(u5__abc_78290_new_n2597_));
OAI22X1 OAI22X1_98 ( .A(u5__abc_78290_new_n1297_), .B(u5__abc_78290_new_n2661_), .C(u5__abc_78290_new_n771_), .D(u5__abc_78290_new_n2660_), .Y(u5_next_state_5_));
OAI22X1 OAI22X1_99 ( .A(u5__abc_78290_new_n732_), .B(u5__abc_78290_new_n2694_), .C(u5__abc_78290_new_n2692_), .D(u5__abc_78290_new_n2613_), .Y(u5_next_state_8_));
OR2X2 OR2X2_1 ( .A(u0__abc_74894_new_n1117_), .B(u0__abc_74894_new_n1131_), .Y(u0__abc_74894_new_n1132_));
OR2X2 OR2X2_10 ( .A(u0_u1_inited), .B(u0_init_ack1), .Y(u0_u1__0inited_0_0_));
OR2X2 OR2X2_100 ( .A(u5__abc_78290_new_n1307_), .B(u5__abc_78290_new_n1540_), .Y(u5__abc_78290_new_n1541_));
OR2X2 OR2X2_101 ( .A(u5__abc_78290_new_n1597_), .B(u5__abc_78290_new_n1604_), .Y(u5__abc_78290_new_n1605_));
OR2X2 OR2X2_102 ( .A(u5__abc_78290_new_n1823_), .B(u5__abc_78290_new_n454_), .Y(u5__abc_78290_new_n1824_));
OR2X2 OR2X2_103 ( .A(u5__abc_78290_new_n1928_), .B(u5__abc_78290_new_n477_), .Y(u5__abc_78290_new_n1929_));
OR2X2 OR2X2_104 ( .A(u5__abc_78290_new_n1932_), .B(u5__abc_78290_new_n477_), .Y(u5__abc_78290_new_n1933_));
OR2X2 OR2X2_105 ( .A(u5__abc_78290_new_n1235_), .B(u5__abc_78290_new_n1997_), .Y(u5__abc_78290_new_n1998_));
OR2X2 OR2X2_106 ( .A(u5__abc_78290_new_n1998_), .B(u5__abc_78290_new_n1999_), .Y(u5__abc_78290_new_n2000_));
OR2X2 OR2X2_107 ( .A(u5__abc_78290_new_n2002_), .B(u5__abc_78290_new_n969_), .Y(u5__abc_78290_new_n2004_));
OR2X2 OR2X2_108 ( .A(u5__abc_78290_new_n2003_), .B(u5_ir_cnt_1_), .Y(u5__abc_78290_new_n2015_));
OR2X2 OR2X2_109 ( .A(u5__abc_78290_new_n1556_), .B(u5__abc_78290_new_n2029_), .Y(u5__abc_78290_new_n2030_));
OR2X2 OR2X2_11 ( .A(csc_s_5_), .B(csc_s_4_), .Y(u1__abc_72801_new_n258_));
OR2X2 OR2X2_110 ( .A(u5__abc_78290_new_n2039_), .B(u5__abc_78290_new_n1186_), .Y(u5__abc_78290_new_n2040_));
OR2X2 OR2X2_111 ( .A(u5__abc_78290_new_n821_), .B(u5__abc_78290_new_n819_), .Y(u5__abc_78290_new_n2047_));
OR2X2 OR2X2_112 ( .A(u5__abc_78290_new_n670_), .B(u5__abc_78290_new_n808_), .Y(u5__abc_78290_new_n2050_));
OR2X2 OR2X2_113 ( .A(u5__abc_78290_new_n2054_), .B(u5__abc_78290_new_n2049_), .Y(u5__abc_78290_new_n2055_));
OR2X2 OR2X2_114 ( .A(u5__abc_78290_new_n2063_), .B(u5__abc_78290_new_n2062_), .Y(u5__abc_78290_new_n2064_));
OR2X2 OR2X2_115 ( .A(u5__abc_78290_new_n1008_), .B(u5__abc_78290_new_n1006_), .Y(u5__abc_78290_new_n2071_));
OR2X2 OR2X2_116 ( .A(u5__abc_78290_new_n2083_), .B(u5_timer_0_), .Y(u5__abc_78290_new_n2084_));
OR2X2 OR2X2_117 ( .A(u5__abc_78290_new_n2097_), .B(u5__abc_78290_new_n2103_), .Y(u5__abc_78290_new_n2104_));
OR2X2 OR2X2_118 ( .A(u5__abc_78290_new_n2158_), .B(u5__abc_78290_new_n923_), .Y(u5__abc_78290_new_n2159_));
OR2X2 OR2X2_119 ( .A(u5__abc_78290_new_n1294_), .B(u5__abc_78290_new_n2206_), .Y(u5__abc_78290_new_n2207_));
OR2X2 OR2X2_12 ( .A(csc_s_7_), .B(csc_s_6_), .Y(u1__abc_72801_new_n259_));
OR2X2 OR2X2_120 ( .A(u5__abc_78290_new_n2188_), .B(u5__abc_78290_new_n1687_), .Y(u5__abc_78290_new_n2263_));
OR2X2 OR2X2_121 ( .A(u5__abc_78290_new_n2317_), .B(u5__abc_78290_new_n2111_), .Y(u5__abc_78290_new_n2318_));
OR2X2 OR2X2_122 ( .A(u5__abc_78290_new_n1471_), .B(tms_s_11_), .Y(u5__abc_78290_new_n2326_));
OR2X2 OR2X2_123 ( .A(u5__abc_78290_new_n2176_), .B(u5__abc_78290_new_n1186_), .Y(u5__abc_78290_new_n2331_));
OR2X2 OR2X2_124 ( .A(u5__abc_78290_new_n1471_), .B(tms_s_6_), .Y(u5__abc_78290_new_n2360_));
OR2X2 OR2X2_125 ( .A(u5__abc_78290_new_n1471_), .B(tms_s_7_), .Y(u5__abc_78290_new_n2364_));
OR2X2 OR2X2_126 ( .A(u5__abc_78290_new_n631_), .B(u5__abc_78290_new_n454_), .Y(u5__abc_78290_new_n2374_));
OR2X2 OR2X2_127 ( .A(u5__abc_78290_new_n2409_), .B(u5__abc_78290_new_n1385_), .Y(u5__abc_78290_new_n2410_));
OR2X2 OR2X2_128 ( .A(u5__abc_78290_new_n2446_), .B(u5__abc_78290_new_n555_), .Y(u5__abc_78290_new_n2447_));
OR2X2 OR2X2_129 ( .A(u5__abc_78290_new_n2491_), .B(u5__abc_78290_new_n2379_), .Y(u5__abc_78290_new_n2492_));
OR2X2 OR2X2_13 ( .A(u1__abc_72801_new_n424_), .B(u1__abc_72801_new_n328_), .Y(u1__abc_72801_new_n445_));
OR2X2 OR2X2_130 ( .A(u5__abc_78290_new_n2593_), .B(u5__abc_78290_new_n1344_), .Y(u5__abc_78290_new_n2594_));
OR2X2 OR2X2_131 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1233_), .Y(u5__abc_78290_new_n2615_));
OR2X2 OR2X2_132 ( .A(u5__abc_78290_new_n2594_), .B(u5__abc_78290_new_n869_), .Y(u5__abc_78290_new_n2643_));
OR2X2 OR2X2_133 ( .A(u5__abc_78290_new_n2636_), .B(u5__abc_78290_new_n1990_), .Y(u5__abc_78290_new_n2731_));
OR2X2 OR2X2_134 ( .A(u5__abc_78290_new_n2790_), .B(u5__abc_78290_new_n2793_), .Y(u5_next_state_19_));
OR2X2 OR2X2_135 ( .A(u5__abc_78290_new_n2814_), .B(u5__abc_78290_new_n2818_), .Y(u5_next_state_24_));
OR2X2 OR2X2_136 ( .A(u5__abc_78290_new_n2834_), .B(u5__abc_78290_new_n2837_), .Y(u5_next_state_28_));
OR2X2 OR2X2_137 ( .A(u5__abc_78290_new_n1646_), .B(u5__abc_78290_new_n3094_), .Y(u5__abc_78290_new_n3095_));
OR2X2 OR2X2_138 ( .A(u5__abc_78290_new_n3097_), .B(u5__abc_78290_new_n3088_), .Y(u5__abc_78290_new_n3098_));
OR2X2 OR2X2_139 ( .A(u5__abc_78290_new_n3111_), .B(u5__abc_78290_new_n3110_), .Y(u5__abc_78290_new_n3112_));
OR2X2 OR2X2_14 ( .A(csc_s_3_), .B(csc_s_2_), .Y(u1__abc_72801_new_n671_));
OR2X2 OR2X2_140 ( .A(u5__abc_78290_new_n2000_), .B(u5__abc_78290_new_n3149_), .Y(u5__abc_78290_new_n3150_));
OR2X2 OR2X2_141 ( .A(par_err), .B(u0_wp_err), .Y(u6__abc_81318_new_n139_));
OR2X2 OR2X2_142 ( .A(u6__abc_81318_new_n133_), .B(\wb_addr_i[31] ), .Y(u6__abc_81318_new_n142_));
OR2X2 OR2X2_143 ( .A(u7__abc_73829_new_n76_), .B(u7_mc_dqm_r2_0_), .Y(u7__abc_73829_new_n77_));
OR2X2 OR2X2_144 ( .A(u7__abc_73829_new_n76_), .B(u7_mc_dqm_r2_1_), .Y(u7__abc_73829_new_n81_));
OR2X2 OR2X2_145 ( .A(u7__abc_73829_new_n76_), .B(u7_mc_dqm_r2_2_), .Y(u7__abc_73829_new_n83_));
OR2X2 OR2X2_146 ( .A(u7__abc_73829_new_n76_), .B(u7_mc_dqm_r2_3_), .Y(u7__abc_73829_new_n85_));
OR2X2 OR2X2_147 ( .A(susp_sel), .B(rfr_ack), .Y(u7__abc_73829_new_n107_));
OR2X2 OR2X2_148 ( .A(susp_sel), .B(oe_), .Y(u7__0mc_oe__0_0_));
OR2X2 OR2X2_15 ( .A(u1_u0__abc_72719_new_n71_), .B(u1_u0__abc_72719_new_n84_), .Y(u1_u0__abc_72719_new_n85_));
OR2X2 OR2X2_16 ( .A(bank_adr_0_), .B(bank_adr_1_), .Y(u2_u0__abc_73914_new_n179_));
OR2X2 OR2X2_17 ( .A(u2_u0__abc_73914_new_n209_), .B(u2_u0__abc_73914_new_n140_), .Y(u2_u0__abc_73914_new_n210_));
OR2X2 OR2X2_18 ( .A(u2_u0_b3_last_row_7_), .B(row_adr_7_), .Y(u2_u0__abc_73914_new_n278_));
OR2X2 OR2X2_19 ( .A(u2_u0_b3_last_row_5_), .B(row_adr_5_), .Y(u2_u0__abc_73914_new_n280_));
OR2X2 OR2X2_2 ( .A(1'h0), .B(u0_u1_wp_err), .Y(u0__abc_74894_new_n3471_));
OR2X2 OR2X2_20 ( .A(u2_u0__abc_73914_new_n294_), .B(u2_u0__abc_73914_new_n295_), .Y(u2_u0__abc_73914_new_n296_));
OR2X2 OR2X2_21 ( .A(row_adr_4_), .B(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_73914_new_n301_));
OR2X2 OR2X2_22 ( .A(row_adr_8_), .B(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_73914_new_n307_));
OR2X2 OR2X2_23 ( .A(row_adr_6_), .B(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_73914_new_n309_));
OR2X2 OR2X2_24 ( .A(u2_u0__abc_73914_new_n173_), .B(u2_u0_b1_last_row_11_), .Y(u2_u0__abc_73914_new_n320_));
OR2X2 OR2X2_25 ( .A(u2_u0__abc_73914_new_n161_), .B(u2_u0_b1_last_row_7_), .Y(u2_u0__abc_73914_new_n323_));
OR2X2 OR2X2_26 ( .A(u2_u0__abc_73914_new_n173_), .B(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_73914_new_n331_));
OR2X2 OR2X2_27 ( .A(u2_u0__abc_73914_new_n167_), .B(u2_u0_b0_last_row_9_), .Y(u2_u0__abc_73914_new_n332_));
OR2X2 OR2X2_28 ( .A(u2_u0__abc_73914_new_n164_), .B(u2_u0_b0_last_row_8_), .Y(u2_u0__abc_73914_new_n337_));
OR2X2 OR2X2_29 ( .A(row_adr_0_), .B(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_73914_new_n346_));
OR2X2 OR2X2_3 ( .A(u0__abc_74894_new_n3730_), .B(\wb_addr_i[6] ), .Y(u0__abc_74894_new_n3815_));
OR2X2 OR2X2_30 ( .A(row_adr_1_), .B(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_73914_new_n348_));
OR2X2 OR2X2_31 ( .A(row_adr_7_), .B(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_73914_new_n359_));
OR2X2 OR2X2_32 ( .A(row_adr_10_), .B(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_73914_new_n361_));
OR2X2 OR2X2_33 ( .A(row_adr_7_), .B(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_73914_new_n373_));
OR2X2 OR2X2_34 ( .A(row_adr_3_), .B(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_73914_new_n378_));
OR2X2 OR2X2_35 ( .A(u2_u0__abc_73914_new_n398_), .B(u2_bank_clr_all_0), .Y(u2_u0__abc_73914_new_n419_));
OR2X2 OR2X2_36 ( .A(bank_adr_0_), .B(bank_adr_1_), .Y(u2_u1__abc_73914_new_n179_));
OR2X2 OR2X2_37 ( .A(u2_u1__abc_73914_new_n209_), .B(u2_u1__abc_73914_new_n140_), .Y(u2_u1__abc_73914_new_n210_));
OR2X2 OR2X2_38 ( .A(u2_u1_b3_last_row_7_), .B(row_adr_7_), .Y(u2_u1__abc_73914_new_n278_));
OR2X2 OR2X2_39 ( .A(u2_u1_b3_last_row_5_), .B(row_adr_5_), .Y(u2_u1__abc_73914_new_n280_));
OR2X2 OR2X2_4 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n4449_));
OR2X2 OR2X2_40 ( .A(u2_u1__abc_73914_new_n294_), .B(u2_u1__abc_73914_new_n295_), .Y(u2_u1__abc_73914_new_n296_));
OR2X2 OR2X2_41 ( .A(row_adr_4_), .B(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_73914_new_n301_));
OR2X2 OR2X2_42 ( .A(row_adr_8_), .B(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_73914_new_n307_));
OR2X2 OR2X2_43 ( .A(row_adr_6_), .B(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_73914_new_n309_));
OR2X2 OR2X2_44 ( .A(u2_u1__abc_73914_new_n173_), .B(u2_u1_b1_last_row_11_), .Y(u2_u1__abc_73914_new_n320_));
OR2X2 OR2X2_45 ( .A(u2_u1__abc_73914_new_n161_), .B(u2_u1_b1_last_row_7_), .Y(u2_u1__abc_73914_new_n323_));
OR2X2 OR2X2_46 ( .A(u2_u1__abc_73914_new_n173_), .B(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_73914_new_n331_));
OR2X2 OR2X2_47 ( .A(u2_u1__abc_73914_new_n167_), .B(u2_u1_b0_last_row_9_), .Y(u2_u1__abc_73914_new_n332_));
OR2X2 OR2X2_48 ( .A(u2_u1__abc_73914_new_n164_), .B(u2_u1_b0_last_row_8_), .Y(u2_u1__abc_73914_new_n337_));
OR2X2 OR2X2_49 ( .A(row_adr_0_), .B(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_73914_new_n346_));
OR2X2 OR2X2_5 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n4455_));
OR2X2 OR2X2_50 ( .A(row_adr_1_), .B(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_73914_new_n348_));
OR2X2 OR2X2_51 ( .A(row_adr_7_), .B(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_73914_new_n359_));
OR2X2 OR2X2_52 ( .A(row_adr_10_), .B(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_73914_new_n361_));
OR2X2 OR2X2_53 ( .A(row_adr_7_), .B(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_73914_new_n373_));
OR2X2 OR2X2_54 ( .A(row_adr_3_), .B(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_73914_new_n378_));
OR2X2 OR2X2_55 ( .A(u2_u1__abc_73914_new_n398_), .B(u2_bank_clr_all_1), .Y(u2_u1__abc_73914_new_n419_));
OR2X2 OR2X2_56 ( .A(u3_rd_fifo_out_8_), .B(u3_rd_fifo_out_9_), .Y(u3__abc_73372_new_n631_));
OR2X2 OR2X2_57 ( .A(u3__abc_73372_new_n646_), .B(u3__abc_73372_new_n643_), .Y(u3__abc_73372_new_n647_));
OR2X2 OR2X2_58 ( .A(u3_rd_fifo_out_16_), .B(u3_rd_fifo_out_17_), .Y(u3__abc_73372_new_n653_));
OR2X2 OR2X2_59 ( .A(u3_rd_fifo_out_24_), .B(u3_rd_fifo_out_25_), .Y(u3__abc_73372_new_n703_));
OR2X2 OR2X2_6 ( .A(1'h0), .B(1'h0), .Y(u0__abc_74894_new_n4458_));
OR2X2 OR2X2_60 ( .A(u3_u0_rd_adr_0_), .B(u3_u0_rd_adr_3_), .Y(u3_u0__abc_74260_new_n734_));
OR2X2 OR2X2_61 ( .A(u3_u0__abc_74260_new_n735_), .B(u3_u0__abc_74260_new_n734_), .Y(u3_u0__abc_74260_new_n736_));
OR2X2 OR2X2_62 ( .A(u4_ps_cnt_3_), .B(rfr_ps_val_3_), .Y(u4__abc_74770_new_n71_));
OR2X2 OR2X2_63 ( .A(u4_ps_cnt_2_), .B(rfr_ps_val_2_), .Y(u4__abc_74770_new_n73_));
OR2X2 OR2X2_64 ( .A(u4_ps_cnt_7_), .B(rfr_ps_val_7_), .Y(u4__abc_74770_new_n76_));
OR2X2 OR2X2_65 ( .A(u4_ps_cnt_6_), .B(rfr_ps_val_6_), .Y(u4__abc_74770_new_n78_));
OR2X2 OR2X2_66 ( .A(u4_ps_cnt_0_), .B(rfr_ps_val_0_), .Y(u4__abc_74770_new_n84_));
OR2X2 OR2X2_67 ( .A(u4_ps_cnt_1_), .B(rfr_ps_val_1_), .Y(u4__abc_74770_new_n87_));
OR2X2 OR2X2_68 ( .A(u4__abc_74770_new_n112_), .B(rfr_ack), .Y(u4__abc_74770_new_n113_));
OR2X2 OR2X2_69 ( .A(u4__abc_74770_new_n139_), .B(u4_ps_cnt_2_), .Y(u4__abc_74770_new_n144_));
OR2X2 OR2X2_7 ( .A(init_req), .B(lmr_req), .Y(u0__abc_74894_new_n4465_));
OR2X2 OR2X2_70 ( .A(u4__abc_74770_new_n156_), .B(u4_ps_cnt_6_), .Y(u4__abc_74770_new_n162_));
OR2X2 OR2X2_71 ( .A(u5__abc_78290_new_n497_), .B(u5__abc_78290_new_n491_), .Y(u5__abc_78290_new_n498_));
OR2X2 OR2X2_72 ( .A(u5__abc_78290_new_n552_), .B(u5__abc_78290_new_n551_), .Y(u5__abc_78290_new_n553_));
OR2X2 OR2X2_73 ( .A(u5__abc_78290_new_n555_), .B(u5__abc_78290_new_n512_), .Y(u5__abc_78290_new_n556_));
OR2X2 OR2X2_74 ( .A(u5__abc_78290_new_n557_), .B(u5__abc_78290_new_n572_), .Y(u5__abc_78290_new_n573_));
OR2X2 OR2X2_75 ( .A(u5__abc_78290_new_n722_), .B(u5__abc_78290_new_n682_), .Y(u5__abc_78290_new_n723_));
OR2X2 OR2X2_76 ( .A(u5__abc_78290_new_n751_), .B(u5__abc_78290_new_n408_), .Y(u5__abc_78290_new_n752_));
OR2X2 OR2X2_77 ( .A(u5__abc_78290_new_n766_), .B(u5__abc_78290_new_n762_), .Y(u5__abc_78290_new_n767_));
OR2X2 OR2X2_78 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1127_), .Y(u5__abc_78290_new_n1128_));
OR2X2 OR2X2_79 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1228_), .Y(u5__abc_78290_new_n1229_));
OR2X2 OR2X2_8 ( .A(u0_u0_inited), .B(u0_init_ack0), .Y(u0_u0__0inited_0_0_));
OR2X2 OR2X2_80 ( .A(u5__abc_78290_new_n1234_), .B(u5__abc_78290_new_n1223_), .Y(u5__abc_78290_new_n1235_));
OR2X2 OR2X2_81 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1238_), .Y(u5__abc_78290_new_n1239_));
OR2X2 OR2X2_82 ( .A(u5__abc_78290_new_n1235_), .B(u5__abc_78290_new_n1251_), .Y(u5__abc_78290_new_n1252_));
OR2X2 OR2X2_83 ( .A(u5__abc_78290_new_n1258_), .B(u5__abc_78290_new_n1260_), .Y(u5__abc_78290_new_n1261_));
OR2X2 OR2X2_84 ( .A(u5__abc_78290_new_n1258_), .B(u5__abc_78290_new_n1265_), .Y(u5__abc_78290_new_n1266_));
OR2X2 OR2X2_85 ( .A(u5__abc_78290_new_n1053_), .B(u5__abc_78290_new_n1266_), .Y(u5__abc_78290_new_n1267_));
OR2X2 OR2X2_86 ( .A(u5__abc_78290_new_n1258_), .B(u5__abc_78290_new_n1276_), .Y(u5__abc_78290_new_n1277_));
OR2X2 OR2X2_87 ( .A(u5__abc_78290_new_n1284_), .B(u5__abc_78290_new_n1286_), .Y(u5__abc_78290_new_n1287_));
OR2X2 OR2X2_88 ( .A(u5__abc_78290_new_n1283_), .B(u5__abc_78290_new_n1292_), .Y(u5__abc_78290_new_n1293_));
OR2X2 OR2X2_89 ( .A(u5__abc_78290_new_n1275_), .B(u5__abc_78290_new_n1293_), .Y(u5__abc_78290_new_n1294_));
OR2X2 OR2X2_9 ( .A(u0_u1__abc_72470_new_n214_), .B(u0_u1__abc_72470_new_n212_), .Y(u0_u1__abc_72470_new_n215_));
OR2X2 OR2X2_90 ( .A(u5__abc_78290_new_n1307_), .B(u5__abc_78290_new_n1309_), .Y(u5__abc_78290_new_n1310_));
OR2X2 OR2X2_91 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1099_), .Y(u5__abc_78290_new_n1368_));
OR2X2 OR2X2_92 ( .A(u5__abc_78290_new_n1371_), .B(u5__abc_78290_new_n1360_), .Y(u5__abc_78290_new_n1372_));
OR2X2 OR2X2_93 ( .A(u5__abc_78290_new_n1038_), .B(u5__abc_78290_new_n1123_), .Y(u5__abc_78290_new_n1386_));
OR2X2 OR2X2_94 ( .A(u5__abc_78290_new_n1387_), .B(u5__abc_78290_new_n1388_), .Y(u5__abc_78290_new_n1389_));
OR2X2 OR2X2_95 ( .A(u5__abc_78290_new_n1410_), .B(u5_cnt), .Y(u5__abc_78290_new_n1415_));
OR2X2 OR2X2_96 ( .A(u5__abc_78290_new_n1435_), .B(u5__abc_78290_new_n1449_), .Y(u5_cmd_1_));
OR2X2 OR2X2_97 ( .A(u5__abc_78290_new_n1435_), .B(u5__abc_78290_new_n1463_), .Y(u5_cmd_2_));
OR2X2 OR2X2_98 ( .A(u5__abc_78290_new_n1471_), .B(tms_s_19_), .Y(u5__abc_78290_new_n1472_));
OR2X2 OR2X2_99 ( .A(u5__abc_78290_new_n1535_), .B(u5__abc_78290_new_n1536_), .Y(u5__abc_78290_new_n1537_));
XNOR2X1 XNOR2X1_1 ( .A(u1_u0__abc_72719_new_n52_), .B(u1_acs_addr_2_), .Y(u1_u0__0out_r_12_0__2_));
XNOR2X1 XNOR2X1_10 ( .A(u2_u0_b3_last_row_0_), .B(row_adr_0_), .Y(u2_u0__abc_73914_new_n274_));
XNOR2X1 XNOR2X1_11 ( .A(u2_u0_b3_last_row_12_), .B(row_adr_12_), .Y(u2_u0__abc_73914_new_n284_));
XNOR2X1 XNOR2X1_12 ( .A(row_adr_12_), .B(u2_u0_b1_last_row_12_), .Y(u2_u0__abc_73914_new_n311_));
XNOR2X1 XNOR2X1_13 ( .A(row_adr_2_), .B(u2_u0_b1_last_row_2_), .Y(u2_u0__abc_73914_new_n317_));
XNOR2X1 XNOR2X1_14 ( .A(row_adr_10_), .B(u2_u0_b1_last_row_10_), .Y(u2_u0__abc_73914_new_n321_));
XNOR2X1 XNOR2X1_15 ( .A(row_adr_5_), .B(u2_u0_b0_last_row_5_), .Y(u2_u0__abc_73914_new_n351_));
XNOR2X1 XNOR2X1_16 ( .A(row_adr_12_), .B(u2_u0_b2_last_row_12_), .Y(u2_u0__abc_73914_new_n384_));
XNOR2X1 XNOR2X1_17 ( .A(row_adr_0_), .B(u2_u0_b2_last_row_0_), .Y(u2_u0__abc_73914_new_n393_));
XNOR2X1 XNOR2X1_18 ( .A(u2_u1_b3_last_row_0_), .B(row_adr_0_), .Y(u2_u1__abc_73914_new_n274_));
XNOR2X1 XNOR2X1_19 ( .A(u2_u1_b3_last_row_12_), .B(row_adr_12_), .Y(u2_u1__abc_73914_new_n284_));
XNOR2X1 XNOR2X1_2 ( .A(u1_u0__abc_72719_new_n54_), .B(u1_acs_addr_3_), .Y(u1_u0__0out_r_12_0__3_));
XNOR2X1 XNOR2X1_20 ( .A(row_adr_12_), .B(u2_u1_b1_last_row_12_), .Y(u2_u1__abc_73914_new_n311_));
XNOR2X1 XNOR2X1_21 ( .A(row_adr_2_), .B(u2_u1_b1_last_row_2_), .Y(u2_u1__abc_73914_new_n317_));
XNOR2X1 XNOR2X1_22 ( .A(row_adr_10_), .B(u2_u1_b1_last_row_10_), .Y(u2_u1__abc_73914_new_n321_));
XNOR2X1 XNOR2X1_23 ( .A(row_adr_5_), .B(u2_u1_b0_last_row_5_), .Y(u2_u1__abc_73914_new_n351_));
XNOR2X1 XNOR2X1_24 ( .A(row_adr_12_), .B(u2_u1_b2_last_row_12_), .Y(u2_u1__abc_73914_new_n384_));
XNOR2X1 XNOR2X1_25 ( .A(row_adr_0_), .B(u2_u1_b2_last_row_0_), .Y(u2_u1__abc_73914_new_n393_));
XNOR2X1 XNOR2X1_26 ( .A(\wb_data_i[3] ), .B(\wb_data_i[2] ), .Y(u3__abc_73372_new_n279_));
XNOR2X1 XNOR2X1_27 ( .A(\wb_data_i[1] ), .B(\wb_data_i[0] ), .Y(u3__abc_73372_new_n280_));
XNOR2X1 XNOR2X1_28 ( .A(u3__abc_73372_new_n279_), .B(u3__abc_73372_new_n280_), .Y(u3__abc_73372_new_n281_));
XNOR2X1 XNOR2X1_29 ( .A(\wb_data_i[7] ), .B(\wb_data_i[6] ), .Y(u3__abc_73372_new_n282_));
XNOR2X1 XNOR2X1_3 ( .A(u1_u0__abc_72719_new_n58_), .B(u1_u0__abc_72719_new_n56_), .Y(u1_u0__0out_r_12_0__4_));
XNOR2X1 XNOR2X1_30 ( .A(\wb_data_i[5] ), .B(\wb_data_i[4] ), .Y(u3__abc_73372_new_n283_));
XNOR2X1 XNOR2X1_31 ( .A(u3__abc_73372_new_n282_), .B(u3__abc_73372_new_n283_), .Y(u3__abc_73372_new_n284_));
XNOR2X1 XNOR2X1_32 ( .A(u3__abc_73372_new_n281_), .B(u3__abc_73372_new_n284_), .Y(u3__abc_73372_new_n285_));
XNOR2X1 XNOR2X1_33 ( .A(\wb_data_i[9] ), .B(\wb_data_i[8] ), .Y(u3__abc_73372_new_n289_));
XNOR2X1 XNOR2X1_34 ( .A(u3__abc_73372_new_n288_), .B(u3__abc_73372_new_n289_), .Y(u3__abc_73372_new_n290_));
XNOR2X1 XNOR2X1_35 ( .A(\wb_data_i[13] ), .B(\wb_data_i[12] ), .Y(u3__abc_73372_new_n292_));
XNOR2X1 XNOR2X1_36 ( .A(u3__abc_73372_new_n291_), .B(u3__abc_73372_new_n292_), .Y(u3__abc_73372_new_n293_));
XNOR2X1 XNOR2X1_37 ( .A(u3__abc_73372_new_n290_), .B(u3__abc_73372_new_n293_), .Y(u3__abc_73372_new_n294_));
XNOR2X1 XNOR2X1_38 ( .A(\wb_data_i[17] ), .B(\wb_data_i[16] ), .Y(u3__abc_73372_new_n298_));
XNOR2X1 XNOR2X1_39 ( .A(u3__abc_73372_new_n297_), .B(u3__abc_73372_new_n298_), .Y(u3__abc_73372_new_n299_));
XNOR2X1 XNOR2X1_4 ( .A(u1_u0__abc_72719_new_n61_), .B(u1_acs_addr_6_), .Y(u1_u0__0out_r_12_0__6_));
XNOR2X1 XNOR2X1_40 ( .A(\wb_data_i[21] ), .B(\wb_data_i[20] ), .Y(u3__abc_73372_new_n301_));
XNOR2X1 XNOR2X1_41 ( .A(u3__abc_73372_new_n300_), .B(u3__abc_73372_new_n301_), .Y(u3__abc_73372_new_n302_));
XNOR2X1 XNOR2X1_42 ( .A(u3__abc_73372_new_n299_), .B(u3__abc_73372_new_n302_), .Y(u3__abc_73372_new_n303_));
XNOR2X1 XNOR2X1_43 ( .A(\wb_data_i[25] ), .B(\wb_data_i[24] ), .Y(u3__abc_73372_new_n307_));
XNOR2X1 XNOR2X1_44 ( .A(u3__abc_73372_new_n306_), .B(u3__abc_73372_new_n307_), .Y(u3__abc_73372_new_n308_));
XNOR2X1 XNOR2X1_45 ( .A(\wb_data_i[29] ), .B(\wb_data_i[28] ), .Y(u3__abc_73372_new_n310_));
XNOR2X1 XNOR2X1_46 ( .A(u3__abc_73372_new_n309_), .B(u3__abc_73372_new_n310_), .Y(u3__abc_73372_new_n311_));
XNOR2X1 XNOR2X1_47 ( .A(u3__abc_73372_new_n308_), .B(u3__abc_73372_new_n311_), .Y(u3__abc_73372_new_n312_));
XNOR2X1 XNOR2X1_48 ( .A(u3_rd_fifo_out_14_), .B(u3_rd_fifo_out_15_), .Y(u3__abc_73372_new_n639_));
XNOR2X1 XNOR2X1_49 ( .A(u3_rd_fifo_out_12_), .B(u3_rd_fifo_out_13_), .Y(u3__abc_73372_new_n644_));
XNOR2X1 XNOR2X1_5 ( .A(u1_u0__abc_72719_new_n71_), .B(u1_acs_addr_8_), .Y(u1_u0__0out_r_12_0__8_));
XNOR2X1 XNOR2X1_50 ( .A(u3_rd_fifo_out_10_), .B(u3_rd_fifo_out_11_), .Y(u3__abc_73372_new_n645_));
XNOR2X1 XNOR2X1_51 ( .A(u3__abc_73372_new_n644_), .B(u3__abc_73372_new_n645_), .Y(u3__abc_73372_new_n646_));
XNOR2X1 XNOR2X1_52 ( .A(u3_rd_fifo_out_22_), .B(u3_rd_fifo_out_23_), .Y(u3__abc_73372_new_n650_));
XNOR2X1 XNOR2X1_53 ( .A(u3_rd_fifo_out_6_), .B(u3_rd_fifo_out_7_), .Y(u3__abc_73372_new_n688_));
XNOR2X1 XNOR2X1_54 ( .A(u3_rd_fifo_out_4_), .B(u3_rd_fifo_out_5_), .Y(u3__abc_73372_new_n692_));
XNOR2X1 XNOR2X1_55 ( .A(u3_rd_fifo_out_2_), .B(u3_rd_fifo_out_3_), .Y(u3__abc_73372_new_n693_));
XNOR2X1 XNOR2X1_56 ( .A(u3__abc_73372_new_n692_), .B(u3__abc_73372_new_n693_), .Y(u3__abc_73372_new_n698_));
XNOR2X1 XNOR2X1_57 ( .A(u3_rd_fifo_out_30_), .B(u3_rd_fifo_out_31_), .Y(u3__abc_73372_new_n700_));
XNOR2X1 XNOR2X1_58 ( .A(u4_ps_cnt_4_), .B(rfr_ps_val_4_), .Y(u4__abc_74770_new_n82_));
XNOR2X1 XNOR2X1_59 ( .A(u4_ps_cnt_5_), .B(rfr_ps_val_5_), .Y(u4__abc_74770_new_n83_));
XNOR2X1 XNOR2X1_6 ( .A(u1_u0__abc_72719_new_n78_), .B(u1_acs_addr_10_), .Y(u1_u0__0out_r_12_0__10_));
XNOR2X1 XNOR2X1_60 ( .A(u4__abc_74770_new_n148_), .B(u4_ps_cnt_3_), .Y(u4__abc_74770_new_n149_));
XNOR2X1 XNOR2X1_61 ( .A(u5__abc_78290_new_n1953_), .B(u5_burst_cnt_7_), .Y(u5__abc_78290_new_n1954_));
XNOR2X1 XNOR2X1_62 ( .A(u5__abc_78290_new_n1969_), .B(u5_burst_cnt_9_), .Y(u5__abc_78290_new_n1970_));
XNOR2X1 XNOR2X1_63 ( .A(u5__abc_78290_new_n1975_), .B(u5_burst_cnt_10_), .Y(u5__abc_78290_new_n1976_));
XNOR2X1 XNOR2X1_64 ( .A(u5__abc_78290_new_n2234_), .B(u5_timer_2_), .Y(u5__abc_78290_new_n2294_));
XNOR2X1 XNOR2X1_65 ( .A(u5__abc_78290_new_n2554_), .B(u5_ack_cnt_3_), .Y(u5__abc_78290_new_n2555_));
XNOR2X1 XNOR2X1_7 ( .A(u1_u0__abc_72719_new_n91_), .B(u1_acs_addr_14_), .Y(u1_acs_addr_pl1_14_));
XNOR2X1 XNOR2X1_8 ( .A(u1_u0__abc_72719_new_n111_), .B(u1_acs_addr_21_), .Y(u1_acs_addr_pl1_21_));
XNOR2X1 XNOR2X1_9 ( .A(u1_u0__abc_72719_new_n121_), .B(u1_acs_addr_22_), .Y(u1_acs_addr_pl1_22_));
XOR2X1 XOR2X1_1 ( .A(u0_csc1_17_), .B(\wb_addr_i[22] ), .Y(u0_u1__abc_72470_new_n418_));
XOR2X1 XOR2X1_10 ( .A(\wb_data_i[27] ), .B(\wb_data_i[26] ), .Y(u3__abc_73372_new_n306_));
XOR2X1 XOR2X1_11 ( .A(\wb_data_i[31] ), .B(\wb_data_i[30] ), .Y(u3__abc_73372_new_n309_));
XOR2X1 XOR2X1_12 ( .A(u3_rd_fifo_out_14_), .B(u3_rd_fifo_out_15_), .Y(u3__abc_73372_new_n630_));
XOR2X1 XOR2X1_13 ( .A(u3_rd_fifo_out_6_), .B(u3_rd_fifo_out_7_), .Y(u3__abc_73372_new_n679_));
XOR2X1 XOR2X1_14 ( .A(u3__abc_73372_new_n692_), .B(u3__abc_73372_new_n693_), .Y(u3__abc_73372_new_n694_));
XOR2X1 XOR2X1_15 ( .A(u4__abc_74770_new_n151_), .B(u4_ps_cnt_4_), .Y(u4__abc_74770_new_n152_));
XOR2X1 XOR2X1_16 ( .A(u5__abc_78290_new_n2017_), .B(u5_ir_cnt_3_), .Y(u5__abc_78290_new_n2020_));
XOR2X1 XOR2X1_2 ( .A(u1_acs_addr_0_), .B(u1_acs_addr_1_), .Y(u1_u0__0out_r_12_0__1_));
XOR2X1 XOR2X1_3 ( .A(u1_u0__abc_72719_new_n89_), .B(u1_acs_addr_13_), .Y(u1_acs_addr_pl1_13_));
XOR2X1 XOR2X1_4 ( .A(u1_u0__abc_72719_new_n100_), .B(u1_acs_addr_16_), .Y(u1_acs_addr_pl1_16_));
XOR2X1 XOR2X1_5 ( .A(u1_u0__abc_72719_new_n104_), .B(u1_acs_addr_18_), .Y(u1_acs_addr_pl1_18_));
XOR2X1 XOR2X1_6 ( .A(\wb_data_i[11] ), .B(\wb_data_i[10] ), .Y(u3__abc_73372_new_n288_));
XOR2X1 XOR2X1_7 ( .A(\wb_data_i[15] ), .B(\wb_data_i[14] ), .Y(u3__abc_73372_new_n291_));
XOR2X1 XOR2X1_8 ( .A(\wb_data_i[19] ), .B(\wb_data_i[18] ), .Y(u3__abc_73372_new_n297_));
XOR2X1 XOR2X1_9 ( .A(\wb_data_i[23] ), .B(\wb_data_i[22] ), .Y(u3__abc_73372_new_n300_));


endmodule